magic
tech gf180mcuC
magscale 1 5
timestamp 1670224516
<< metal1 >>
rect 672 33333 24304 33350
rect 672 33307 2239 33333
rect 2265 33307 2291 33333
rect 2317 33307 2343 33333
rect 2369 33307 17599 33333
rect 17625 33307 17651 33333
rect 17677 33307 17703 33333
rect 17729 33307 24304 33333
rect 672 33290 24304 33307
rect 672 32941 24304 32958
rect 672 32915 9919 32941
rect 9945 32915 9971 32941
rect 9997 32915 10023 32941
rect 10049 32915 24304 32941
rect 672 32898 24304 32915
rect 672 32549 24304 32566
rect 672 32523 2239 32549
rect 2265 32523 2291 32549
rect 2317 32523 2343 32549
rect 2369 32523 17599 32549
rect 17625 32523 17651 32549
rect 17677 32523 17703 32549
rect 17729 32523 24304 32549
rect 672 32506 24304 32523
rect 672 32157 24304 32174
rect 672 32131 9919 32157
rect 9945 32131 9971 32157
rect 9997 32131 10023 32157
rect 10049 32131 24304 32157
rect 672 32114 24304 32131
rect 672 31765 24304 31782
rect 672 31739 2239 31765
rect 2265 31739 2291 31765
rect 2317 31739 2343 31765
rect 2369 31739 17599 31765
rect 17625 31739 17651 31765
rect 17677 31739 17703 31765
rect 17729 31739 24304 31765
rect 672 31722 24304 31739
rect 672 31373 24304 31390
rect 672 31347 9919 31373
rect 9945 31347 9971 31373
rect 9997 31347 10023 31373
rect 10049 31347 24304 31373
rect 672 31330 24304 31347
rect 672 30981 24304 30998
rect 672 30955 2239 30981
rect 2265 30955 2291 30981
rect 2317 30955 2343 30981
rect 2369 30955 17599 30981
rect 17625 30955 17651 30981
rect 17677 30955 17703 30981
rect 17729 30955 24304 30981
rect 672 30938 24304 30955
rect 672 30589 24304 30606
rect 672 30563 9919 30589
rect 9945 30563 9971 30589
rect 9997 30563 10023 30589
rect 10049 30563 24304 30589
rect 672 30546 24304 30563
rect 672 30197 24304 30214
rect 672 30171 2239 30197
rect 2265 30171 2291 30197
rect 2317 30171 2343 30197
rect 2369 30171 17599 30197
rect 17625 30171 17651 30197
rect 17677 30171 17703 30197
rect 17729 30171 24304 30197
rect 672 30154 24304 30171
rect 672 29805 24304 29822
rect 672 29779 9919 29805
rect 9945 29779 9971 29805
rect 9997 29779 10023 29805
rect 10049 29779 24304 29805
rect 672 29762 24304 29779
rect 23311 29609 23337 29615
rect 23311 29577 23337 29583
rect 23367 29609 23393 29615
rect 23367 29577 23393 29583
rect 23591 29609 23617 29615
rect 23591 29577 23617 29583
rect 672 29413 24304 29430
rect 672 29387 2239 29413
rect 2265 29387 2291 29413
rect 2317 29387 2343 29413
rect 2369 29387 17599 29413
rect 17625 29387 17651 29413
rect 17677 29387 17703 29413
rect 17729 29387 24304 29413
rect 672 29370 24304 29387
rect 23031 29217 23057 29223
rect 3929 29191 3935 29217
rect 3961 29191 3967 29217
rect 4377 29191 4383 29217
rect 4409 29191 4415 29217
rect 4601 29191 4607 29217
rect 4633 29191 4639 29217
rect 23031 29185 23057 29191
rect 23199 29217 23225 29223
rect 23199 29185 23225 29191
rect 23703 29217 23729 29223
rect 23703 29185 23729 29191
rect 23871 29217 23897 29223
rect 23871 29185 23897 29191
rect 23311 29161 23337 29167
rect 23311 29129 23337 29135
rect 23591 29161 23617 29167
rect 23591 29129 23617 29135
rect 672 29021 24304 29038
rect 672 28995 9919 29021
rect 9945 28995 9971 29021
rect 9997 28995 10023 29021
rect 10049 28995 24304 29021
rect 672 28978 24304 28995
rect 22415 28881 22441 28887
rect 4377 28855 4383 28881
rect 4409 28855 4415 28881
rect 5833 28855 5839 28881
rect 5865 28855 5871 28881
rect 22415 28849 22441 28855
rect 22695 28881 22721 28887
rect 22695 28849 22721 28855
rect 23087 28881 23113 28887
rect 23087 28849 23113 28855
rect 23255 28881 23281 28887
rect 23255 28849 23281 28855
rect 23535 28881 23561 28887
rect 23535 28849 23561 28855
rect 22583 28825 22609 28831
rect 3593 28799 3599 28825
rect 3625 28799 3631 28825
rect 4377 28799 4383 28825
rect 4409 28799 4415 28825
rect 5049 28799 5055 28825
rect 5081 28799 5087 28825
rect 5833 28799 5839 28825
rect 5865 28799 5871 28825
rect 22583 28793 22609 28799
rect 23031 28825 23057 28831
rect 23031 28793 23057 28799
rect 23647 28825 23673 28831
rect 23647 28793 23673 28799
rect 23815 28825 23841 28831
rect 23815 28793 23841 28799
rect 672 28629 24304 28646
rect 672 28603 2239 28629
rect 2265 28603 2291 28629
rect 2317 28603 2343 28629
rect 2369 28603 17599 28629
rect 17625 28603 17651 28629
rect 17677 28603 17703 28629
rect 17729 28603 24304 28629
rect 672 28586 24304 28603
rect 22135 28433 22161 28439
rect 3929 28407 3935 28433
rect 3961 28407 3967 28433
rect 4881 28407 4887 28433
rect 4913 28407 4919 28433
rect 22135 28401 22161 28407
rect 23031 28433 23057 28439
rect 23031 28401 23057 28407
rect 23591 28433 23617 28439
rect 23591 28401 23617 28407
rect 23759 28433 23785 28439
rect 23759 28401 23785 28407
rect 23871 28433 23897 28439
rect 23871 28401 23897 28407
rect 22191 28377 22217 28383
rect 4881 28351 4887 28377
rect 4913 28351 4919 28377
rect 22191 28345 22217 28351
rect 22359 28377 22385 28383
rect 22359 28345 22385 28351
rect 23143 28377 23169 28383
rect 23143 28345 23169 28351
rect 23311 28377 23337 28383
rect 23311 28345 23337 28351
rect 672 28237 24304 28254
rect 672 28211 9919 28237
rect 9945 28211 9971 28237
rect 9997 28211 10023 28237
rect 10049 28211 24304 28237
rect 672 28194 24304 28211
rect 22751 28097 22777 28103
rect 5833 28071 5839 28097
rect 5865 28071 5871 28097
rect 7513 28071 7519 28097
rect 7545 28071 7551 28097
rect 22751 28065 22777 28071
rect 23031 28097 23057 28103
rect 23031 28065 23057 28071
rect 23143 28097 23169 28103
rect 23143 28065 23169 28071
rect 23311 28097 23337 28103
rect 23311 28065 23337 28071
rect 23591 28097 23617 28103
rect 23591 28065 23617 28071
rect 23871 28097 23897 28103
rect 23871 28065 23897 28071
rect 21407 28041 21433 28047
rect 1857 28015 1863 28041
rect 1889 28015 1895 28041
rect 2305 28015 2311 28041
rect 2337 28015 2343 28041
rect 2529 28015 2535 28041
rect 2561 28015 2567 28041
rect 3593 28015 3599 28041
rect 3625 28015 3631 28041
rect 3873 28015 3879 28041
rect 3905 28015 3911 28041
rect 4041 28015 4047 28041
rect 4073 28015 4079 28041
rect 5049 28015 5055 28041
rect 5081 28015 5087 28041
rect 5833 28015 5839 28041
rect 5865 28015 5871 28041
rect 6617 28015 6623 28041
rect 6649 28015 6655 28041
rect 7513 28015 7519 28041
rect 7545 28015 7551 28041
rect 21407 28009 21433 28015
rect 21519 28041 21545 28047
rect 21519 28009 21545 28015
rect 21687 28041 21713 28047
rect 21687 28009 21713 28015
rect 21967 28041 21993 28047
rect 21967 28009 21993 28015
rect 22079 28041 22105 28047
rect 22079 28009 22105 28015
rect 22247 28041 22273 28047
rect 22247 28009 22273 28015
rect 22527 28041 22553 28047
rect 22527 28009 22553 28015
rect 22639 28041 22665 28047
rect 22639 28009 22665 28015
rect 23759 28041 23785 28047
rect 23759 28009 23785 28015
rect 672 27845 24304 27862
rect 672 27819 2239 27845
rect 2265 27819 2291 27845
rect 2317 27819 2343 27845
rect 2369 27819 17599 27845
rect 17625 27819 17651 27845
rect 17677 27819 17703 27845
rect 17729 27819 24304 27845
rect 672 27802 24304 27819
rect 21127 27649 21153 27655
rect 1353 27623 1359 27649
rect 1385 27623 1391 27649
rect 2473 27623 2479 27649
rect 2505 27623 2511 27649
rect 3313 27623 3319 27649
rect 3345 27623 3351 27649
rect 3985 27623 3991 27649
rect 4017 27623 4023 27649
rect 4769 27623 4775 27649
rect 4801 27623 4807 27649
rect 5441 27623 5447 27649
rect 5473 27623 5479 27649
rect 7121 27623 7127 27649
rect 7153 27623 7159 27649
rect 8017 27623 8023 27649
rect 8049 27623 8055 27649
rect 8409 27623 8415 27649
rect 8441 27623 8447 27649
rect 8857 27623 8863 27649
rect 8889 27623 8895 27649
rect 8969 27623 8975 27649
rect 9001 27623 9007 27649
rect 11041 27623 11047 27649
rect 11073 27623 11079 27649
rect 11377 27623 11383 27649
rect 11409 27623 11415 27649
rect 11489 27623 11495 27649
rect 11521 27623 11527 27649
rect 21127 27617 21153 27623
rect 21575 27649 21601 27655
rect 21575 27617 21601 27623
rect 21631 27649 21657 27655
rect 21631 27617 21657 27623
rect 21799 27649 21825 27655
rect 21799 27617 21825 27623
rect 22415 27649 22441 27655
rect 22415 27617 22441 27623
rect 20959 27593 20985 27599
rect 2473 27567 2479 27593
rect 2505 27567 2511 27593
rect 3985 27567 3991 27593
rect 4017 27567 4023 27593
rect 5441 27567 5447 27593
rect 5473 27567 5479 27593
rect 8017 27567 8023 27593
rect 8049 27567 8055 27593
rect 20959 27561 20985 27567
rect 21239 27593 21265 27599
rect 21239 27561 21265 27567
rect 22079 27593 22105 27599
rect 22079 27561 22105 27567
rect 22191 27593 22217 27599
rect 22191 27561 22217 27567
rect 22975 27593 23001 27599
rect 22975 27561 23001 27567
rect 23087 27593 23113 27599
rect 23087 27561 23113 27567
rect 23255 27593 23281 27599
rect 23255 27561 23281 27567
rect 23535 27593 23561 27599
rect 23535 27561 23561 27567
rect 23647 27593 23673 27599
rect 23647 27561 23673 27567
rect 23815 27593 23841 27599
rect 23815 27561 23841 27567
rect 672 27453 24304 27470
rect 672 27427 9919 27453
rect 9945 27427 9971 27453
rect 9997 27427 10023 27453
rect 10049 27427 24304 27453
rect 672 27410 24304 27427
rect 21071 27313 21097 27319
rect 7513 27287 7519 27313
rect 7545 27287 7551 27313
rect 10033 27287 10039 27313
rect 10065 27287 10071 27313
rect 11489 27287 11495 27313
rect 11521 27287 11527 27313
rect 21071 27281 21097 27287
rect 21631 27313 21657 27319
rect 21631 27281 21657 27287
rect 21183 27257 21209 27263
rect 1857 27231 1863 27257
rect 1889 27231 1895 27257
rect 2417 27231 2423 27257
rect 2449 27231 2455 27257
rect 2529 27231 2535 27257
rect 2561 27231 2567 27257
rect 3313 27231 3319 27257
rect 3345 27231 3351 27257
rect 3761 27231 3767 27257
rect 3793 27231 3799 27257
rect 3985 27231 3991 27257
rect 4017 27231 4023 27257
rect 5161 27231 5167 27257
rect 5193 27231 5199 27257
rect 5441 27231 5447 27257
rect 5473 27231 5479 27257
rect 5553 27231 5559 27257
rect 5585 27231 5591 27257
rect 6617 27231 6623 27257
rect 6649 27231 6655 27257
rect 7513 27231 7519 27257
rect 7545 27231 7551 27257
rect 8857 27231 8863 27257
rect 8889 27231 8895 27257
rect 10033 27231 10039 27257
rect 10065 27231 10071 27257
rect 10593 27231 10599 27257
rect 10625 27231 10631 27257
rect 11489 27231 11495 27257
rect 11521 27231 11527 27257
rect 21183 27225 21209 27231
rect 21351 27257 21377 27263
rect 21351 27225 21377 27231
rect 21743 27257 21769 27263
rect 21743 27225 21769 27231
rect 21967 27257 21993 27263
rect 21967 27225 21993 27231
rect 22191 27257 22217 27263
rect 22191 27225 22217 27231
rect 22359 27257 22385 27263
rect 22359 27225 22385 27231
rect 22527 27257 22553 27263
rect 22527 27225 22553 27231
rect 22751 27257 22777 27263
rect 22751 27225 22777 27231
rect 22919 27257 22945 27263
rect 22919 27225 22945 27231
rect 23031 27257 23057 27263
rect 23031 27225 23057 27231
rect 23311 27257 23337 27263
rect 23311 27225 23337 27231
rect 23423 27257 23449 27263
rect 23423 27225 23449 27231
rect 23647 27257 23673 27263
rect 23647 27225 23673 27231
rect 672 27061 24304 27078
rect 672 27035 2239 27061
rect 2265 27035 2291 27061
rect 2317 27035 2343 27061
rect 2369 27035 17599 27061
rect 17625 27035 17651 27061
rect 17677 27035 17703 27061
rect 17729 27035 24304 27061
rect 672 27018 24304 27035
rect 19783 26865 19809 26871
rect 1353 26839 1359 26865
rect 1385 26839 1391 26865
rect 2473 26839 2479 26865
rect 2505 26839 2511 26865
rect 3313 26839 3319 26865
rect 3345 26839 3351 26865
rect 3481 26839 3487 26865
rect 3513 26839 3519 26865
rect 3705 26839 3711 26865
rect 3737 26839 3743 26865
rect 4769 26839 4775 26865
rect 4801 26839 4807 26865
rect 5441 26839 5447 26865
rect 5473 26839 5479 26865
rect 7121 26839 7127 26865
rect 7153 26839 7159 26865
rect 8017 26839 8023 26865
rect 8049 26839 8055 26865
rect 8577 26839 8583 26865
rect 8609 26839 8615 26865
rect 8857 26839 8863 26865
rect 8889 26839 8895 26865
rect 8969 26839 8975 26865
rect 9001 26839 9007 26865
rect 11041 26839 11047 26865
rect 11073 26839 11079 26865
rect 11713 26839 11719 26865
rect 11745 26839 11751 26865
rect 19783 26833 19809 26839
rect 19951 26865 19977 26871
rect 19951 26833 19977 26839
rect 20343 26865 20369 26871
rect 20343 26833 20369 26839
rect 20511 26865 20537 26871
rect 20511 26833 20537 26839
rect 20679 26865 20705 26871
rect 20679 26833 20705 26839
rect 20959 26865 20985 26871
rect 20959 26833 20985 26839
rect 21127 26865 21153 26871
rect 21127 26833 21153 26839
rect 21239 26865 21265 26871
rect 21239 26833 21265 26839
rect 21631 26865 21657 26871
rect 21631 26833 21657 26839
rect 21799 26865 21825 26871
rect 21799 26833 21825 26839
rect 22135 26865 22161 26871
rect 22135 26833 22161 26839
rect 22247 26865 22273 26871
rect 22247 26833 22273 26839
rect 22415 26865 22441 26871
rect 22415 26833 22441 26839
rect 22751 26865 22777 26871
rect 22751 26833 22777 26839
rect 22919 26865 22945 26871
rect 22919 26833 22945 26839
rect 23087 26865 23113 26871
rect 23087 26833 23113 26839
rect 23423 26865 23449 26871
rect 23423 26833 23449 26839
rect 23647 26865 23673 26871
rect 23647 26833 23673 26839
rect 20119 26809 20145 26815
rect 2473 26783 2479 26809
rect 2505 26783 2511 26809
rect 5441 26783 5447 26809
rect 5473 26783 5479 26809
rect 8017 26783 8023 26809
rect 8049 26783 8055 26809
rect 11769 26783 11775 26809
rect 11801 26783 11807 26809
rect 20119 26777 20145 26783
rect 21519 26809 21545 26815
rect 21519 26777 21545 26783
rect 23311 26809 23337 26815
rect 23311 26777 23337 26783
rect 672 26669 24304 26686
rect 672 26643 9919 26669
rect 9945 26643 9971 26669
rect 9997 26643 10023 26669
rect 10049 26643 24304 26669
rect 672 26626 24304 26643
rect 21015 26529 21041 26535
rect 4265 26503 4271 26529
rect 4297 26503 4303 26529
rect 7513 26503 7519 26529
rect 7545 26503 7551 26529
rect 10033 26503 10039 26529
rect 10065 26503 10071 26529
rect 21015 26497 21041 26503
rect 21855 26529 21881 26535
rect 21855 26497 21881 26503
rect 22695 26529 22721 26535
rect 22695 26497 22721 26503
rect 22863 26529 22889 26535
rect 22863 26497 22889 26503
rect 21127 26473 21153 26479
rect 1857 26447 1863 26473
rect 1889 26447 1895 26473
rect 2417 26447 2423 26473
rect 2449 26447 2455 26473
rect 2529 26447 2535 26473
rect 2561 26447 2567 26473
rect 3313 26447 3319 26473
rect 3345 26447 3351 26473
rect 4209 26447 4215 26473
rect 4241 26447 4247 26473
rect 5161 26447 5167 26473
rect 5193 26447 5199 26473
rect 5329 26447 5335 26473
rect 5361 26447 5367 26473
rect 5553 26447 5559 26473
rect 5585 26447 5591 26473
rect 6337 26447 6343 26473
rect 6369 26447 6375 26473
rect 7513 26447 7519 26473
rect 7545 26447 7551 26473
rect 8913 26447 8919 26473
rect 8945 26447 8951 26473
rect 10033 26447 10039 26473
rect 10065 26447 10071 26473
rect 10593 26447 10599 26473
rect 10625 26447 10631 26473
rect 10873 26447 10879 26473
rect 10905 26447 10911 26473
rect 10985 26447 10991 26473
rect 11017 26447 11023 26473
rect 21127 26441 21153 26447
rect 21295 26473 21321 26479
rect 21295 26441 21321 26447
rect 21631 26473 21657 26479
rect 21631 26441 21657 26447
rect 21743 26473 21769 26479
rect 21743 26441 21769 26447
rect 22135 26473 22161 26479
rect 22135 26441 22161 26447
rect 22303 26473 22329 26479
rect 22303 26441 22329 26447
rect 22471 26473 22497 26479
rect 22471 26441 22497 26447
rect 22975 26473 23001 26479
rect 22975 26441 23001 26447
rect 23311 26473 23337 26479
rect 23311 26441 23337 26447
rect 23423 26473 23449 26479
rect 23423 26441 23449 26447
rect 23535 26473 23561 26479
rect 23535 26441 23561 26447
rect 672 26277 24304 26294
rect 672 26251 2239 26277
rect 2265 26251 2291 26277
rect 2317 26251 2343 26277
rect 2369 26251 17599 26277
rect 17625 26251 17651 26277
rect 17677 26251 17703 26277
rect 17729 26251 24304 26277
rect 672 26234 24304 26251
rect 21071 26081 21097 26087
rect 1353 26055 1359 26081
rect 1385 26055 1391 26081
rect 2473 26055 2479 26081
rect 2505 26055 2511 26081
rect 3313 26055 3319 26081
rect 3345 26055 3351 26081
rect 4209 26055 4215 26081
rect 4241 26055 4247 26081
rect 4769 26055 4775 26081
rect 4801 26055 4807 26081
rect 4937 26055 4943 26081
rect 4969 26055 4975 26081
rect 5161 26055 5167 26081
rect 5193 26055 5199 26081
rect 7121 26055 7127 26081
rect 7153 26055 7159 26081
rect 8017 26055 8023 26081
rect 8049 26055 8055 26081
rect 8577 26055 8583 26081
rect 8609 26055 8615 26081
rect 8857 26055 8863 26081
rect 8889 26055 8895 26081
rect 8969 26055 8975 26081
rect 9001 26055 9007 26081
rect 11097 26055 11103 26081
rect 11129 26055 11135 26081
rect 11713 26055 11719 26081
rect 11745 26055 11751 26081
rect 12553 26055 12559 26081
rect 12585 26055 12591 26081
rect 13337 26055 13343 26081
rect 13369 26055 13375 26081
rect 21071 26049 21097 26055
rect 21239 26081 21265 26087
rect 21239 26049 21265 26055
rect 21519 26081 21545 26087
rect 21519 26049 21545 26055
rect 21631 26081 21657 26087
rect 21631 26049 21657 26055
rect 21799 26081 21825 26087
rect 21799 26049 21825 26055
rect 22135 26081 22161 26087
rect 22135 26049 22161 26055
rect 22247 26081 22273 26087
rect 22247 26049 22273 26055
rect 22415 26081 22441 26087
rect 22415 26049 22441 26055
rect 23311 26081 23337 26087
rect 23311 26049 23337 26055
rect 23423 26081 23449 26087
rect 23423 26049 23449 26055
rect 20959 26025 20985 26031
rect 2473 25999 2479 26025
rect 2505 25999 2511 26025
rect 4209 25999 4215 26025
rect 4241 25999 4247 26025
rect 8017 25999 8023 26025
rect 8049 25999 8055 26025
rect 11769 25999 11775 26025
rect 11801 25999 11807 26025
rect 13337 25999 13343 26025
rect 13369 25999 13375 26025
rect 20959 25993 20985 25999
rect 23535 26025 23561 26031
rect 23535 25993 23561 25999
rect 672 25885 24304 25902
rect 672 25859 9919 25885
rect 9945 25859 9971 25885
rect 9997 25859 10023 25885
rect 10049 25859 24304 25885
rect 672 25842 24304 25859
rect 21575 25745 21601 25751
rect 3033 25719 3039 25745
rect 3065 25719 3071 25745
rect 4265 25719 4271 25745
rect 4297 25719 4303 25745
rect 7625 25719 7631 25745
rect 7657 25719 7663 25745
rect 10033 25719 10039 25745
rect 10065 25719 10071 25745
rect 11489 25719 11495 25745
rect 11521 25719 11527 25745
rect 21575 25713 21601 25719
rect 21855 25745 21881 25751
rect 21855 25713 21881 25719
rect 22135 25745 22161 25751
rect 22135 25713 22161 25719
rect 22695 25745 22721 25751
rect 22695 25713 22721 25719
rect 22863 25745 22889 25751
rect 22863 25713 22889 25719
rect 21743 25689 21769 25695
rect 2137 25663 2143 25689
rect 2169 25663 2175 25689
rect 3033 25663 3039 25689
rect 3065 25663 3071 25689
rect 3313 25663 3319 25689
rect 3345 25663 3351 25689
rect 4209 25663 4215 25689
rect 4241 25663 4247 25689
rect 5105 25663 5111 25689
rect 5137 25663 5143 25689
rect 5329 25663 5335 25689
rect 5361 25663 5367 25689
rect 5553 25663 5559 25689
rect 5585 25663 5591 25689
rect 6673 25663 6679 25689
rect 6705 25663 6711 25689
rect 7625 25663 7631 25689
rect 7657 25663 7663 25689
rect 9137 25663 9143 25689
rect 9169 25663 9175 25689
rect 10033 25663 10039 25689
rect 10065 25663 10071 25689
rect 10593 25663 10599 25689
rect 10625 25663 10631 25689
rect 11489 25663 11495 25689
rect 11521 25663 11527 25689
rect 13113 25663 13119 25689
rect 13145 25663 13151 25689
rect 13337 25663 13343 25689
rect 13369 25663 13375 25689
rect 13505 25663 13511 25689
rect 13537 25663 13543 25689
rect 21743 25657 21769 25663
rect 22303 25689 22329 25695
rect 22303 25657 22329 25663
rect 22471 25689 22497 25695
rect 22471 25657 22497 25663
rect 22975 25689 23001 25695
rect 22975 25657 23001 25663
rect 23311 25689 23337 25695
rect 23311 25657 23337 25663
rect 23423 25689 23449 25695
rect 23423 25657 23449 25663
rect 23535 25689 23561 25695
rect 23535 25657 23561 25663
rect 672 25493 24304 25510
rect 672 25467 2239 25493
rect 2265 25467 2291 25493
rect 2317 25467 2343 25493
rect 2369 25467 17599 25493
rect 17625 25467 17651 25493
rect 17677 25467 17703 25493
rect 17729 25467 24304 25493
rect 672 25450 24304 25467
rect 22135 25297 22161 25303
rect 1577 25271 1583 25297
rect 1609 25271 1615 25297
rect 2473 25271 2479 25297
rect 2505 25271 2511 25297
rect 3313 25271 3319 25297
rect 3345 25271 3351 25297
rect 4209 25271 4215 25297
rect 4241 25271 4247 25297
rect 4769 25271 4775 25297
rect 4801 25271 4807 25297
rect 4937 25271 4943 25297
rect 4969 25271 4975 25297
rect 5161 25271 5167 25297
rect 5193 25271 5199 25297
rect 7121 25271 7127 25297
rect 7153 25271 7159 25297
rect 8017 25271 8023 25297
rect 8049 25271 8055 25297
rect 8409 25271 8415 25297
rect 8441 25271 8447 25297
rect 8857 25271 8863 25297
rect 8889 25271 8895 25297
rect 8969 25271 8975 25297
rect 9001 25271 9007 25297
rect 11097 25271 11103 25297
rect 11129 25271 11135 25297
rect 11713 25271 11719 25297
rect 11745 25271 11751 25297
rect 12553 25271 12559 25297
rect 12585 25271 12591 25297
rect 12721 25271 12727 25297
rect 12753 25271 12759 25297
rect 12945 25271 12951 25297
rect 12977 25271 12983 25297
rect 22135 25265 22161 25271
rect 22247 25297 22273 25303
rect 22247 25265 22273 25271
rect 22359 25297 22385 25303
rect 22359 25265 22385 25271
rect 23311 25297 23337 25303
rect 23311 25265 23337 25271
rect 23423 25297 23449 25303
rect 23423 25265 23449 25271
rect 23591 25297 23617 25303
rect 23591 25265 23617 25271
rect 2473 25215 2479 25241
rect 2505 25215 2511 25241
rect 4209 25215 4215 25241
rect 4241 25215 4247 25241
rect 8017 25215 8023 25241
rect 8049 25215 8055 25241
rect 11769 25215 11775 25241
rect 11801 25215 11807 25241
rect 672 25101 24304 25118
rect 672 25075 9919 25101
rect 9945 25075 9971 25101
rect 9997 25075 10023 25101
rect 10049 25075 24304 25101
rect 672 25058 24304 25075
rect 22471 24961 22497 24967
rect 4489 24935 4495 24961
rect 4521 24935 4527 24961
rect 6169 24935 6175 24961
rect 6201 24935 6207 24961
rect 7625 24935 7631 24961
rect 7657 24935 7663 24961
rect 10033 24935 10039 24961
rect 10065 24935 10071 24961
rect 11489 24935 11495 24961
rect 11521 24935 11527 24961
rect 15241 24935 15247 24961
rect 15273 24935 15279 24961
rect 22471 24929 22497 24935
rect 22583 24961 22609 24967
rect 22583 24929 22609 24935
rect 22751 24961 22777 24967
rect 22751 24929 22777 24935
rect 23031 24961 23057 24967
rect 23031 24929 23057 24935
rect 23143 24961 23169 24967
rect 23143 24929 23169 24935
rect 23311 24961 23337 24967
rect 23311 24929 23337 24935
rect 23759 24905 23785 24911
rect 1857 24879 1863 24905
rect 1889 24879 1895 24905
rect 2417 24879 2423 24905
rect 2449 24879 2455 24905
rect 2529 24879 2535 24905
rect 2561 24879 2567 24905
rect 3369 24879 3375 24905
rect 3401 24879 3407 24905
rect 4489 24879 4495 24905
rect 4521 24879 4527 24905
rect 5049 24879 5055 24905
rect 5081 24879 5087 24905
rect 6169 24879 6175 24905
rect 6201 24879 6207 24905
rect 6673 24879 6679 24905
rect 6705 24879 6711 24905
rect 7625 24879 7631 24905
rect 7657 24879 7663 24905
rect 8913 24879 8919 24905
rect 8945 24879 8951 24905
rect 10033 24879 10039 24905
rect 10065 24879 10071 24905
rect 10313 24879 10319 24905
rect 10345 24879 10351 24905
rect 11489 24879 11495 24905
rect 11521 24879 11527 24905
rect 13113 24879 13119 24905
rect 13145 24879 13151 24905
rect 13393 24879 13399 24905
rect 13425 24879 13431 24905
rect 13505 24879 13511 24905
rect 13537 24879 13543 24905
rect 14513 24879 14519 24905
rect 14545 24879 14551 24905
rect 15129 24879 15135 24905
rect 15161 24879 15167 24905
rect 23759 24873 23785 24879
rect 23927 24905 23953 24911
rect 23927 24873 23953 24879
rect 24039 24905 24065 24911
rect 24039 24873 24065 24879
rect 672 24709 24304 24726
rect 672 24683 2239 24709
rect 2265 24683 2291 24709
rect 2317 24683 2343 24709
rect 2369 24683 17599 24709
rect 17625 24683 17651 24709
rect 17677 24683 17703 24709
rect 17729 24683 24304 24709
rect 672 24666 24304 24683
rect 23143 24513 23169 24519
rect 1353 24487 1359 24513
rect 1385 24487 1391 24513
rect 2473 24487 2479 24513
rect 2505 24487 2511 24513
rect 3817 24487 3823 24513
rect 3849 24487 3855 24513
rect 4377 24487 4383 24513
rect 4409 24487 4415 24513
rect 4489 24487 4495 24513
rect 4521 24487 4527 24513
rect 5273 24487 5279 24513
rect 5305 24487 5311 24513
rect 6449 24487 6455 24513
rect 6481 24487 6487 24513
rect 7121 24487 7127 24513
rect 7153 24487 7159 24513
rect 8017 24487 8023 24513
rect 8049 24487 8055 24513
rect 8577 24487 8583 24513
rect 8609 24487 8615 24513
rect 9473 24487 9479 24513
rect 9505 24487 9511 24513
rect 10817 24487 10823 24513
rect 10849 24487 10855 24513
rect 11377 24487 11383 24513
rect 11409 24487 11415 24513
rect 11489 24487 11495 24513
rect 11521 24487 11527 24513
rect 12553 24487 12559 24513
rect 12585 24487 12591 24513
rect 13337 24487 13343 24513
rect 13369 24487 13375 24513
rect 15073 24487 15079 24513
rect 15105 24487 15111 24513
rect 15241 24487 15247 24513
rect 15273 24487 15279 24513
rect 15465 24487 15471 24513
rect 15497 24487 15503 24513
rect 23143 24481 23169 24487
rect 23311 24513 23337 24519
rect 23311 24481 23337 24487
rect 23759 24513 23785 24519
rect 23759 24481 23785 24487
rect 23871 24513 23897 24519
rect 23871 24481 23897 24487
rect 23479 24457 23505 24463
rect 2473 24431 2479 24457
rect 2505 24431 2511 24457
rect 6449 24431 6455 24457
rect 6481 24431 6487 24457
rect 8017 24431 8023 24457
rect 8049 24431 8055 24457
rect 9473 24431 9479 24457
rect 9505 24431 9511 24457
rect 13337 24431 13343 24457
rect 13369 24431 13375 24457
rect 23479 24425 23505 24431
rect 24039 24457 24065 24463
rect 24039 24425 24065 24431
rect 672 24317 24304 24334
rect 672 24291 9919 24317
rect 9945 24291 9971 24317
rect 9997 24291 10023 24317
rect 10049 24291 24304 24317
rect 672 24274 24304 24291
rect 23927 24177 23953 24183
rect 3033 24151 3039 24177
rect 3065 24151 3071 24177
rect 4489 24151 4495 24177
rect 4521 24151 4527 24177
rect 6169 24151 6175 24177
rect 6201 24151 6207 24177
rect 7625 24151 7631 24177
rect 7657 24151 7663 24177
rect 10033 24151 10039 24177
rect 10065 24151 10071 24177
rect 11489 24151 11495 24177
rect 11521 24151 11527 24177
rect 15241 24151 15247 24177
rect 15273 24151 15279 24177
rect 23927 24145 23953 24151
rect 23759 24121 23785 24127
rect 1857 24095 1863 24121
rect 1889 24095 1895 24121
rect 3033 24095 3039 24121
rect 3065 24095 3071 24121
rect 3369 24095 3375 24121
rect 3401 24095 3407 24121
rect 4489 24095 4495 24121
rect 4521 24095 4527 24121
rect 5049 24095 5055 24121
rect 5081 24095 5087 24121
rect 6169 24095 6175 24121
rect 6201 24095 6207 24121
rect 6673 24095 6679 24121
rect 6705 24095 6711 24121
rect 7625 24095 7631 24121
rect 7657 24095 7663 24121
rect 9081 24095 9087 24121
rect 9113 24095 9119 24121
rect 10033 24095 10039 24121
rect 10065 24095 10071 24121
rect 10593 24095 10599 24121
rect 10625 24095 10631 24121
rect 11489 24095 11495 24121
rect 11521 24095 11527 24121
rect 13113 24095 13119 24121
rect 13145 24095 13151 24121
rect 13337 24095 13343 24121
rect 13369 24095 13375 24121
rect 13505 24095 13511 24121
rect 13537 24095 13543 24121
rect 14513 24095 14519 24121
rect 14545 24095 14551 24121
rect 15129 24095 15135 24121
rect 15161 24095 15167 24121
rect 23759 24089 23785 24095
rect 24039 24121 24065 24127
rect 24039 24089 24065 24095
rect 672 23925 24304 23942
rect 672 23899 2239 23925
rect 2265 23899 2291 23925
rect 2317 23899 2343 23925
rect 2369 23899 17599 23925
rect 17625 23899 17651 23925
rect 17677 23899 17703 23925
rect 17729 23899 24304 23925
rect 672 23882 24304 23899
rect 1353 23703 1359 23729
rect 1385 23703 1391 23729
rect 2473 23703 2479 23729
rect 2505 23703 2511 23729
rect 4097 23703 4103 23729
rect 4129 23703 4135 23729
rect 4993 23703 4999 23729
rect 5025 23703 5031 23729
rect 5553 23703 5559 23729
rect 5585 23703 5591 23729
rect 6449 23703 6455 23729
rect 6481 23703 6487 23729
rect 7121 23703 7127 23729
rect 7153 23703 7159 23729
rect 8017 23703 8023 23729
rect 8049 23703 8055 23729
rect 8577 23703 8583 23729
rect 8609 23703 8615 23729
rect 9473 23703 9479 23729
rect 9505 23703 9511 23729
rect 11097 23703 11103 23729
rect 11129 23703 11135 23729
rect 11713 23703 11719 23729
rect 11745 23703 11751 23729
rect 12273 23703 12279 23729
rect 12305 23703 12311 23729
rect 13449 23703 13455 23729
rect 13481 23703 13487 23729
rect 15073 23703 15079 23729
rect 15105 23703 15111 23729
rect 15241 23703 15247 23729
rect 15273 23703 15279 23729
rect 15465 23703 15471 23729
rect 15497 23703 15503 23729
rect 2473 23647 2479 23673
rect 2505 23647 2511 23673
rect 4993 23647 4999 23673
rect 5025 23647 5031 23673
rect 6449 23647 6455 23673
rect 6481 23647 6487 23673
rect 8017 23647 8023 23673
rect 8049 23647 8055 23673
rect 9473 23647 9479 23673
rect 9505 23647 9511 23673
rect 11769 23647 11775 23673
rect 11801 23647 11807 23673
rect 13449 23647 13455 23673
rect 13481 23647 13487 23673
rect 672 23533 24304 23550
rect 672 23507 9919 23533
rect 9945 23507 9971 23533
rect 9997 23507 10023 23533
rect 10049 23507 24304 23533
rect 672 23490 24304 23507
rect 3033 23367 3039 23393
rect 3065 23367 3071 23393
rect 4489 23367 4495 23393
rect 4521 23367 4527 23393
rect 6169 23367 6175 23393
rect 6201 23367 6207 23393
rect 7513 23367 7519 23393
rect 7545 23367 7551 23393
rect 13953 23367 13959 23393
rect 13985 23367 13991 23393
rect 15297 23367 15303 23393
rect 15329 23367 15335 23393
rect 23703 23337 23729 23343
rect 1857 23311 1863 23337
rect 1889 23311 1895 23337
rect 3033 23311 3039 23337
rect 3065 23311 3071 23337
rect 3369 23311 3375 23337
rect 3401 23311 3407 23337
rect 4489 23311 4495 23337
rect 4521 23311 4527 23337
rect 5049 23311 5055 23337
rect 5081 23311 5087 23337
rect 6169 23311 6175 23337
rect 6201 23311 6207 23337
rect 6673 23311 6679 23337
rect 6705 23311 6711 23337
rect 7513 23311 7519 23337
rect 7545 23311 7551 23337
rect 9081 23311 9087 23337
rect 9113 23311 9119 23337
rect 9305 23311 9311 23337
rect 9337 23311 9343 23337
rect 9529 23311 9535 23337
rect 9561 23311 9567 23337
rect 10313 23311 10319 23337
rect 10345 23311 10351 23337
rect 10873 23311 10879 23337
rect 10905 23311 10911 23337
rect 10985 23311 10991 23337
rect 11017 23311 11023 23337
rect 12833 23311 12839 23337
rect 12865 23311 12871 23337
rect 13953 23311 13959 23337
rect 13985 23311 13991 23337
rect 14569 23311 14575 23337
rect 14601 23311 14607 23337
rect 15297 23311 15303 23337
rect 15329 23311 15335 23337
rect 23703 23305 23729 23311
rect 23871 23337 23897 23343
rect 23871 23305 23897 23311
rect 23983 23337 24009 23343
rect 23983 23305 24009 23311
rect 672 23141 24304 23158
rect 672 23115 2239 23141
rect 2265 23115 2291 23141
rect 2317 23115 2343 23141
rect 2369 23115 17599 23141
rect 17625 23115 17651 23141
rect 17677 23115 17703 23141
rect 17729 23115 24304 23141
rect 672 23098 24304 23115
rect 23871 22945 23897 22951
rect 1353 22919 1359 22945
rect 1385 22919 1391 22945
rect 2473 22919 2479 22945
rect 2505 22919 2511 22945
rect 4097 22919 4103 22945
rect 4129 22919 4135 22945
rect 4993 22919 4999 22945
rect 5025 22919 5031 22945
rect 5273 22919 5279 22945
rect 5305 22919 5311 22945
rect 6169 22919 6175 22945
rect 6201 22919 6207 22945
rect 8129 22919 8135 22945
rect 8161 22919 8167 22945
rect 9025 22919 9031 22945
rect 9057 22919 9063 22945
rect 10817 22919 10823 22945
rect 10849 22919 10855 22945
rect 11265 22919 11271 22945
rect 11297 22919 11303 22945
rect 11489 22919 11495 22945
rect 11521 22919 11527 22945
rect 12273 22919 12279 22945
rect 12305 22919 12311 22945
rect 13449 22919 13455 22945
rect 13481 22919 13487 22945
rect 14793 22919 14799 22945
rect 14825 22919 14831 22945
rect 15297 22919 15303 22945
rect 15329 22919 15335 22945
rect 15465 22919 15471 22945
rect 15497 22919 15503 22945
rect 16249 22919 16255 22945
rect 16281 22919 16287 22945
rect 16809 22919 16815 22945
rect 16841 22919 16847 22945
rect 16921 22919 16927 22945
rect 16953 22919 16959 22945
rect 23871 22913 23897 22919
rect 23983 22945 24009 22951
rect 23983 22913 24009 22919
rect 23199 22889 23225 22895
rect 2473 22863 2479 22889
rect 2505 22863 2511 22889
rect 4993 22863 4999 22889
rect 5025 22863 5031 22889
rect 6225 22863 6231 22889
rect 6257 22863 6263 22889
rect 9025 22863 9031 22889
rect 9057 22863 9063 22889
rect 13449 22863 13455 22889
rect 13481 22863 13487 22889
rect 23199 22857 23225 22863
rect 23367 22889 23393 22895
rect 23367 22857 23393 22863
rect 23479 22889 23505 22895
rect 23479 22857 23505 22863
rect 23759 22889 23785 22895
rect 23759 22857 23785 22863
rect 672 22749 24304 22766
rect 672 22723 9919 22749
rect 9945 22723 9971 22749
rect 9997 22723 10023 22749
rect 10049 22723 24304 22749
rect 672 22706 24304 22723
rect 2977 22583 2983 22609
rect 3009 22583 3015 22609
rect 4489 22583 4495 22609
rect 4521 22583 4527 22609
rect 7009 22583 7015 22609
rect 7041 22583 7047 22609
rect 8241 22583 8247 22609
rect 8273 22583 8279 22609
rect 11265 22583 11271 22609
rect 11297 22583 11303 22609
rect 13953 22583 13959 22609
rect 13985 22583 13991 22609
rect 15297 22583 15303 22609
rect 15329 22583 15335 22609
rect 23759 22553 23785 22559
rect 1857 22527 1863 22553
rect 1889 22527 1895 22553
rect 2977 22527 2983 22553
rect 3009 22527 3015 22553
rect 3369 22527 3375 22553
rect 3401 22527 3407 22553
rect 4489 22527 4495 22553
rect 4521 22527 4527 22553
rect 5833 22527 5839 22553
rect 5865 22527 5871 22553
rect 7009 22527 7015 22553
rect 7041 22527 7047 22553
rect 7569 22527 7575 22553
rect 7601 22527 7607 22553
rect 8241 22527 8247 22553
rect 8273 22527 8279 22553
rect 9081 22527 9087 22553
rect 9113 22527 9119 22553
rect 9305 22527 9311 22553
rect 9337 22527 9343 22553
rect 9529 22527 9535 22553
rect 9561 22527 9567 22553
rect 10313 22527 10319 22553
rect 10345 22527 10351 22553
rect 11265 22527 11271 22553
rect 11297 22527 11303 22553
rect 12833 22527 12839 22553
rect 12865 22527 12871 22553
rect 13953 22527 13959 22553
rect 13985 22527 13991 22553
rect 14569 22527 14575 22553
rect 14601 22527 14607 22553
rect 15297 22527 15303 22553
rect 15329 22527 15335 22553
rect 16809 22527 16815 22553
rect 16841 22527 16847 22553
rect 17257 22527 17263 22553
rect 17289 22527 17295 22553
rect 17481 22527 17487 22553
rect 17513 22527 17519 22553
rect 23759 22521 23785 22527
rect 23871 22553 23897 22559
rect 23871 22521 23897 22527
rect 23983 22553 24009 22559
rect 23983 22521 24009 22527
rect 672 22357 24304 22374
rect 672 22331 2239 22357
rect 2265 22331 2291 22357
rect 2317 22331 2343 22357
rect 2369 22331 17599 22357
rect 17625 22331 17651 22357
rect 17677 22331 17703 22357
rect 17729 22331 24304 22357
rect 672 22314 24304 22331
rect 1353 22135 1359 22161
rect 1385 22135 1391 22161
rect 2473 22135 2479 22161
rect 2505 22135 2511 22161
rect 4097 22135 4103 22161
rect 4129 22135 4135 22161
rect 4993 22135 4999 22161
rect 5025 22135 5031 22161
rect 5273 22135 5279 22161
rect 5305 22135 5311 22161
rect 6225 22135 6231 22161
rect 6257 22135 6263 22161
rect 8129 22135 8135 22161
rect 8161 22135 8167 22161
rect 9025 22135 9031 22161
rect 9057 22135 9063 22161
rect 10817 22135 10823 22161
rect 10849 22135 10855 22161
rect 11265 22135 11271 22161
rect 11297 22135 11303 22161
rect 11489 22135 11495 22161
rect 11521 22135 11527 22161
rect 12273 22135 12279 22161
rect 12305 22135 12311 22161
rect 13225 22135 13231 22161
rect 13257 22135 13263 22161
rect 14793 22135 14799 22161
rect 14825 22135 14831 22161
rect 15297 22135 15303 22161
rect 15329 22135 15335 22161
rect 15465 22135 15471 22161
rect 15497 22135 15503 22161
rect 16249 22135 16255 22161
rect 16281 22135 16287 22161
rect 16753 22135 16759 22161
rect 16785 22135 16791 22161
rect 16921 22135 16927 22161
rect 16953 22135 16959 22161
rect 2473 22079 2479 22105
rect 2505 22079 2511 22105
rect 4993 22079 4999 22105
rect 5025 22079 5031 22105
rect 6225 22079 6231 22105
rect 6257 22079 6263 22105
rect 9025 22079 9031 22105
rect 9057 22079 9063 22105
rect 13225 22079 13231 22105
rect 13257 22079 13263 22105
rect 672 21965 24304 21982
rect 672 21939 9919 21965
rect 9945 21939 9971 21965
rect 9997 21939 10023 21965
rect 10049 21939 24304 21965
rect 672 21922 24304 21939
rect 4377 21799 4383 21825
rect 4409 21799 4415 21825
rect 8241 21799 8247 21825
rect 8273 21799 8279 21825
rect 11265 21799 11271 21825
rect 11297 21799 11303 21825
rect 15353 21799 15359 21825
rect 15385 21799 15391 21825
rect 17985 21799 17991 21825
rect 18017 21799 18023 21825
rect 19273 21799 19279 21825
rect 19305 21799 19311 21825
rect 2137 21743 2143 21769
rect 2169 21743 2175 21769
rect 2417 21743 2423 21769
rect 2449 21743 2455 21769
rect 2529 21743 2535 21769
rect 2561 21743 2567 21769
rect 3593 21743 3599 21769
rect 3625 21743 3631 21769
rect 4377 21743 4383 21769
rect 4409 21743 4415 21769
rect 5833 21743 5839 21769
rect 5865 21743 5871 21769
rect 6393 21743 6399 21769
rect 6425 21743 6431 21769
rect 6505 21743 6511 21769
rect 6537 21743 6543 21769
rect 7289 21743 7295 21769
rect 7321 21743 7327 21769
rect 8241 21743 8247 21769
rect 8273 21743 8279 21769
rect 9081 21743 9087 21769
rect 9113 21743 9119 21769
rect 9305 21743 9311 21769
rect 9337 21743 9343 21769
rect 9529 21743 9535 21769
rect 9561 21743 9567 21769
rect 10313 21743 10319 21769
rect 10345 21743 10351 21769
rect 11265 21743 11271 21769
rect 11297 21743 11303 21769
rect 12833 21743 12839 21769
rect 12865 21743 12871 21769
rect 13393 21743 13399 21769
rect 13425 21743 13431 21769
rect 13505 21743 13511 21769
rect 13537 21743 13543 21769
rect 14569 21743 14575 21769
rect 14601 21743 14607 21769
rect 15353 21743 15359 21769
rect 15385 21743 15391 21769
rect 17089 21743 17095 21769
rect 17121 21743 17127 21769
rect 17985 21743 17991 21769
rect 18017 21743 18023 21769
rect 18545 21743 18551 21769
rect 18577 21743 18583 21769
rect 19273 21743 19279 21769
rect 19305 21743 19311 21769
rect 672 21573 24304 21590
rect 672 21547 2239 21573
rect 2265 21547 2291 21573
rect 2317 21547 2343 21573
rect 2369 21547 17599 21573
rect 17625 21547 17651 21573
rect 17677 21547 17703 21573
rect 17729 21547 24304 21573
rect 672 21530 24304 21547
rect 1577 21351 1583 21377
rect 1609 21351 1615 21377
rect 2473 21351 2479 21377
rect 2505 21351 2511 21377
rect 3817 21351 3823 21377
rect 3849 21351 3855 21377
rect 4377 21351 4383 21377
rect 4409 21351 4415 21377
rect 4489 21351 4495 21377
rect 4521 21351 4527 21377
rect 5273 21351 5279 21377
rect 5305 21351 5311 21377
rect 6393 21351 6399 21377
rect 6425 21351 6431 21377
rect 8129 21351 8135 21377
rect 8161 21351 8167 21377
rect 9025 21351 9031 21377
rect 9057 21351 9063 21377
rect 10817 21351 10823 21377
rect 10849 21351 10855 21377
rect 11265 21351 11271 21377
rect 11297 21351 11303 21377
rect 11489 21351 11495 21377
rect 11521 21351 11527 21377
rect 12273 21351 12279 21377
rect 12305 21351 12311 21377
rect 13449 21351 13455 21377
rect 13481 21351 13487 21377
rect 14793 21351 14799 21377
rect 14825 21351 14831 21377
rect 15353 21351 15359 21377
rect 15385 21351 15391 21377
rect 15465 21351 15471 21377
rect 15497 21351 15503 21377
rect 16249 21351 16255 21377
rect 16281 21351 16287 21377
rect 17425 21351 17431 21377
rect 17457 21351 17463 21377
rect 19049 21351 19055 21377
rect 19081 21351 19087 21377
rect 19273 21351 19279 21377
rect 19305 21351 19311 21377
rect 19441 21351 19447 21377
rect 19473 21351 19479 21377
rect 2473 21295 2479 21321
rect 2505 21295 2511 21321
rect 6393 21295 6399 21321
rect 6425 21295 6431 21321
rect 9025 21295 9031 21321
rect 9057 21295 9063 21321
rect 13449 21295 13455 21321
rect 13481 21295 13487 21321
rect 17425 21295 17431 21321
rect 17457 21295 17463 21321
rect 672 21181 24304 21198
rect 672 21155 9919 21181
rect 9945 21155 9971 21181
rect 9997 21155 10023 21181
rect 10049 21155 24304 21181
rect 672 21138 24304 21155
rect 4377 21015 4383 21041
rect 4409 21015 4415 21041
rect 7009 21015 7015 21041
rect 7041 21015 7047 21041
rect 8241 21015 8247 21041
rect 8273 21015 8279 21041
rect 9809 21015 9815 21041
rect 9841 21015 9847 21041
rect 11265 21015 11271 21041
rect 11297 21015 11303 21041
rect 14009 21015 14015 21041
rect 14041 21015 14047 21041
rect 15353 21015 15359 21041
rect 15385 21015 15391 21041
rect 17929 21015 17935 21041
rect 17961 21015 17967 21041
rect 19441 21015 19447 21041
rect 19473 21015 19479 21041
rect 2137 20959 2143 20985
rect 2169 20959 2175 20985
rect 2417 20959 2423 20985
rect 2449 20959 2455 20985
rect 2529 20959 2535 20985
rect 2561 20959 2567 20985
rect 3593 20959 3599 20985
rect 3625 20959 3631 20985
rect 4377 20959 4383 20985
rect 4409 20959 4415 20985
rect 5833 20959 5839 20985
rect 5865 20959 5871 20985
rect 7009 20959 7015 20985
rect 7041 20959 7047 20985
rect 7289 20959 7295 20985
rect 7321 20959 7327 20985
rect 8241 20959 8247 20985
rect 8273 20959 8279 20985
rect 9137 20959 9143 20985
rect 9169 20959 9175 20985
rect 9809 20959 9815 20985
rect 9841 20959 9847 20985
rect 10313 20959 10319 20985
rect 10345 20959 10351 20985
rect 11265 20959 11271 20985
rect 11297 20959 11303 20985
rect 12945 20959 12951 20985
rect 12977 20959 12983 20985
rect 14009 20959 14015 20985
rect 14041 20959 14047 20985
rect 14569 20959 14575 20985
rect 14601 20959 14607 20985
rect 15353 20959 15359 20985
rect 15385 20959 15391 20985
rect 16809 20959 16815 20985
rect 16841 20959 16847 20985
rect 17929 20959 17935 20985
rect 17961 20959 17967 20985
rect 18545 20959 18551 20985
rect 18577 20959 18583 20985
rect 19441 20959 19447 20985
rect 19473 20959 19479 20985
rect 672 20789 24304 20806
rect 672 20763 2239 20789
rect 2265 20763 2291 20789
rect 2317 20763 2343 20789
rect 2369 20763 17599 20789
rect 17625 20763 17651 20789
rect 17677 20763 17703 20789
rect 17729 20763 24304 20789
rect 672 20746 24304 20763
rect 1577 20567 1583 20593
rect 1609 20567 1615 20593
rect 2473 20567 2479 20593
rect 2505 20567 2511 20593
rect 3817 20567 3823 20593
rect 3849 20567 3855 20593
rect 4265 20567 4271 20593
rect 4297 20567 4303 20593
rect 4489 20567 4495 20593
rect 4521 20567 4527 20593
rect 5273 20567 5279 20593
rect 5305 20567 5311 20593
rect 6449 20567 6455 20593
rect 6481 20567 6487 20593
rect 8129 20567 8135 20593
rect 8161 20567 8167 20593
rect 9025 20567 9031 20593
rect 9057 20567 9063 20593
rect 10817 20567 10823 20593
rect 10849 20567 10855 20593
rect 11265 20567 11271 20593
rect 11297 20567 11303 20593
rect 11489 20567 11495 20593
rect 11521 20567 11527 20593
rect 12273 20567 12279 20593
rect 12305 20567 12311 20593
rect 13449 20567 13455 20593
rect 13481 20567 13487 20593
rect 14905 20567 14911 20593
rect 14937 20567 14943 20593
rect 15353 20567 15359 20593
rect 15385 20567 15391 20593
rect 15465 20567 15471 20593
rect 15497 20567 15503 20593
rect 16529 20567 16535 20593
rect 16561 20567 16567 20593
rect 17425 20567 17431 20593
rect 17457 20567 17463 20593
rect 19049 20567 19055 20593
rect 19081 20567 19087 20593
rect 19945 20567 19951 20593
rect 19977 20567 19983 20593
rect 20505 20567 20511 20593
rect 20537 20567 20543 20593
rect 21233 20567 21239 20593
rect 21265 20567 21271 20593
rect 2473 20511 2479 20537
rect 2505 20511 2511 20537
rect 6449 20511 6455 20537
rect 6481 20511 6487 20537
rect 9025 20511 9031 20537
rect 9057 20511 9063 20537
rect 13449 20511 13455 20537
rect 13481 20511 13487 20537
rect 17425 20511 17431 20537
rect 17457 20511 17463 20537
rect 19945 20511 19951 20537
rect 19977 20511 19983 20537
rect 21233 20511 21239 20537
rect 21265 20511 21271 20537
rect 672 20397 24304 20414
rect 672 20371 9919 20397
rect 9945 20371 9971 20397
rect 9997 20371 10023 20397
rect 10049 20371 24304 20397
rect 672 20354 24304 20371
rect 4265 20231 4271 20257
rect 4297 20231 4303 20257
rect 7009 20231 7015 20257
rect 7041 20231 7047 20257
rect 8241 20231 8247 20257
rect 8273 20231 8279 20257
rect 9809 20231 9815 20257
rect 9841 20231 9847 20257
rect 11265 20231 11271 20257
rect 11297 20231 11303 20257
rect 14009 20231 14015 20257
rect 14041 20231 14047 20257
rect 15353 20231 15359 20257
rect 15385 20231 15391 20257
rect 17985 20231 17991 20257
rect 18017 20231 18023 20257
rect 19273 20231 19279 20257
rect 19305 20231 19311 20257
rect 2137 20175 2143 20201
rect 2169 20175 2175 20201
rect 2417 20175 2423 20201
rect 2449 20175 2455 20201
rect 2529 20175 2535 20201
rect 2561 20175 2567 20201
rect 3593 20175 3599 20201
rect 3625 20175 3631 20201
rect 4209 20175 4215 20201
rect 4241 20175 4247 20201
rect 5833 20175 5839 20201
rect 5865 20175 5871 20201
rect 7009 20175 7015 20201
rect 7041 20175 7047 20201
rect 7289 20175 7295 20201
rect 7321 20175 7327 20201
rect 8241 20175 8247 20201
rect 8273 20175 8279 20201
rect 9137 20175 9143 20201
rect 9169 20175 9175 20201
rect 9809 20175 9815 20201
rect 9841 20175 9847 20201
rect 10313 20175 10319 20201
rect 10345 20175 10351 20201
rect 11265 20175 11271 20201
rect 11297 20175 11303 20201
rect 12945 20175 12951 20201
rect 12977 20175 12983 20201
rect 14009 20175 14015 20201
rect 14041 20175 14047 20201
rect 14289 20175 14295 20201
rect 14321 20175 14327 20201
rect 15353 20175 15359 20201
rect 15385 20175 15391 20201
rect 16809 20175 16815 20201
rect 16841 20175 16847 20201
rect 17985 20175 17991 20201
rect 18017 20175 18023 20201
rect 18545 20175 18551 20201
rect 18577 20175 18583 20201
rect 19273 20175 19279 20201
rect 19305 20175 19311 20201
rect 20953 20175 20959 20201
rect 20985 20175 20991 20201
rect 21233 20175 21239 20201
rect 21265 20175 21271 20201
rect 21457 20175 21463 20201
rect 21489 20175 21495 20201
rect 672 20005 24304 20022
rect 672 19979 2239 20005
rect 2265 19979 2291 20005
rect 2317 19979 2343 20005
rect 2369 19979 17599 20005
rect 17625 19979 17651 20005
rect 17677 19979 17703 20005
rect 17729 19979 24304 20005
rect 672 19962 24304 19979
rect 23759 19809 23785 19815
rect 1577 19783 1583 19809
rect 1609 19783 1615 19809
rect 2473 19783 2479 19809
rect 2505 19783 2511 19809
rect 3817 19783 3823 19809
rect 3849 19783 3855 19809
rect 4377 19783 4383 19809
rect 4409 19783 4415 19809
rect 4545 19783 4551 19809
rect 4577 19783 4583 19809
rect 5273 19783 5279 19809
rect 5305 19783 5311 19809
rect 6449 19783 6455 19809
rect 6481 19783 6487 19809
rect 8129 19783 8135 19809
rect 8161 19783 8167 19809
rect 9025 19783 9031 19809
rect 9057 19783 9063 19809
rect 10817 19783 10823 19809
rect 10849 19783 10855 19809
rect 11265 19783 11271 19809
rect 11297 19783 11303 19809
rect 11489 19783 11495 19809
rect 11521 19783 11527 19809
rect 12273 19783 12279 19809
rect 12305 19783 12311 19809
rect 13449 19783 13455 19809
rect 13481 19783 13487 19809
rect 14793 19783 14799 19809
rect 14825 19783 14831 19809
rect 15913 19783 15919 19809
rect 15945 19783 15951 19809
rect 16249 19783 16255 19809
rect 16281 19783 16287 19809
rect 17425 19783 17431 19809
rect 17457 19783 17463 19809
rect 19049 19783 19055 19809
rect 19081 19783 19087 19809
rect 19329 19783 19335 19809
rect 19361 19783 19367 19809
rect 19441 19783 19447 19809
rect 19473 19783 19479 19809
rect 20505 19783 20511 19809
rect 20537 19783 20543 19809
rect 21177 19783 21183 19809
rect 21209 19783 21215 19809
rect 23759 19777 23785 19783
rect 23871 19809 23897 19815
rect 23871 19777 23897 19783
rect 24039 19753 24065 19759
rect 2473 19727 2479 19753
rect 2505 19727 2511 19753
rect 6449 19727 6455 19753
rect 6481 19727 6487 19753
rect 9025 19727 9031 19753
rect 9057 19727 9063 19753
rect 13449 19727 13455 19753
rect 13481 19727 13487 19753
rect 15913 19727 15919 19753
rect 15945 19727 15951 19753
rect 17425 19727 17431 19753
rect 17457 19727 17463 19753
rect 21177 19727 21183 19753
rect 21209 19727 21215 19753
rect 24039 19721 24065 19727
rect 672 19613 24304 19630
rect 672 19587 9919 19613
rect 9945 19587 9971 19613
rect 9997 19587 10023 19613
rect 10049 19587 24304 19613
rect 672 19570 24304 19587
rect 4433 19447 4439 19473
rect 4465 19447 4471 19473
rect 7009 19447 7015 19473
rect 7041 19447 7047 19473
rect 8241 19447 8247 19473
rect 8273 19447 8279 19473
rect 9809 19447 9815 19473
rect 9841 19447 9847 19473
rect 11265 19447 11271 19473
rect 11297 19447 11303 19473
rect 14009 19447 14015 19473
rect 14041 19447 14047 19473
rect 15465 19447 15471 19473
rect 15497 19447 15503 19473
rect 17985 19447 17991 19473
rect 18017 19447 18023 19473
rect 19329 19447 19335 19473
rect 19361 19447 19367 19473
rect 21793 19447 21799 19473
rect 21825 19447 21831 19473
rect 23249 19447 23255 19473
rect 23281 19447 23287 19473
rect 23703 19417 23729 19423
rect 2137 19391 2143 19417
rect 2169 19391 2175 19417
rect 2417 19391 2423 19417
rect 2449 19391 2455 19417
rect 2529 19391 2535 19417
rect 2561 19391 2567 19417
rect 3593 19391 3599 19417
rect 3625 19391 3631 19417
rect 4433 19391 4439 19417
rect 4465 19391 4471 19417
rect 5833 19391 5839 19417
rect 5865 19391 5871 19417
rect 7009 19391 7015 19417
rect 7041 19391 7047 19417
rect 7289 19391 7295 19417
rect 7321 19391 7327 19417
rect 8241 19391 8247 19417
rect 8273 19391 8279 19417
rect 9137 19391 9143 19417
rect 9169 19391 9175 19417
rect 9809 19391 9815 19417
rect 9841 19391 9847 19417
rect 10313 19391 10319 19417
rect 10345 19391 10351 19417
rect 11265 19391 11271 19417
rect 11297 19391 11303 19417
rect 12945 19391 12951 19417
rect 12977 19391 12983 19417
rect 14009 19391 14015 19417
rect 14041 19391 14047 19417
rect 14289 19391 14295 19417
rect 14321 19391 14327 19417
rect 15465 19391 15471 19417
rect 15497 19391 15503 19417
rect 16865 19391 16871 19417
rect 16897 19391 16903 19417
rect 17985 19391 17991 19417
rect 18017 19391 18023 19417
rect 18545 19391 18551 19417
rect 18577 19391 18583 19417
rect 19329 19391 19335 19417
rect 19361 19391 19367 19417
rect 20953 19391 20959 19417
rect 20985 19391 20991 19417
rect 21793 19391 21799 19417
rect 21825 19391 21831 19417
rect 22521 19391 22527 19417
rect 22553 19391 22559 19417
rect 23249 19391 23255 19417
rect 23281 19391 23287 19417
rect 23703 19385 23729 19391
rect 23871 19417 23897 19423
rect 23871 19385 23897 19391
rect 24039 19417 24065 19423
rect 24039 19385 24065 19391
rect 672 19221 24304 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 24304 19221
rect 672 19178 24304 19195
rect 1577 18999 1583 19025
rect 1609 18999 1615 19025
rect 2473 18999 2479 19025
rect 2505 18999 2511 19025
rect 3817 18999 3823 19025
rect 3849 18999 3855 19025
rect 4377 18999 4383 19025
rect 4409 18999 4415 19025
rect 4489 18999 4495 19025
rect 4521 18999 4527 19025
rect 5273 18999 5279 19025
rect 5305 18999 5311 19025
rect 6449 18999 6455 19025
rect 6481 18999 6487 19025
rect 8129 18999 8135 19025
rect 8161 18999 8167 19025
rect 9025 18999 9031 19025
rect 9057 18999 9063 19025
rect 10817 18999 10823 19025
rect 10849 18999 10855 19025
rect 11265 18999 11271 19025
rect 11297 18999 11303 19025
rect 11489 18999 11495 19025
rect 11521 18999 11527 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 13449 18999 13455 19025
rect 13481 18999 13487 19025
rect 14905 18999 14911 19025
rect 14937 18999 14943 19025
rect 15353 18999 15359 19025
rect 15385 18999 15391 19025
rect 15465 18999 15471 19025
rect 15497 18999 15503 19025
rect 16249 18999 16255 19025
rect 16281 18999 16287 19025
rect 17425 18999 17431 19025
rect 17457 18999 17463 19025
rect 19049 18999 19055 19025
rect 19081 18999 19087 19025
rect 19329 18999 19335 19025
rect 19361 18999 19367 19025
rect 19441 18999 19447 19025
rect 19473 18999 19479 19025
rect 20225 18999 20231 19025
rect 20257 18999 20263 19025
rect 21233 18999 21239 19025
rect 21265 18999 21271 19025
rect 22745 18999 22751 19025
rect 22777 18999 22783 19025
rect 23249 18999 23255 19025
rect 23281 18999 23287 19025
rect 23417 18999 23423 19025
rect 23449 18999 23455 19025
rect 2473 18943 2479 18969
rect 2505 18943 2511 18969
rect 6449 18943 6455 18969
rect 6481 18943 6487 18969
rect 9025 18943 9031 18969
rect 9057 18943 9063 18969
rect 13449 18943 13455 18969
rect 13481 18943 13487 18969
rect 17425 18943 17431 18969
rect 17457 18943 17463 18969
rect 21233 18943 21239 18969
rect 21265 18943 21271 18969
rect 672 18829 24304 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 24304 18829
rect 672 18786 24304 18803
rect 4433 18663 4439 18689
rect 4465 18663 4471 18689
rect 7009 18663 7015 18689
rect 7041 18663 7047 18689
rect 8409 18663 8415 18689
rect 8441 18663 8447 18689
rect 10033 18663 10039 18689
rect 10065 18663 10071 18689
rect 11265 18663 11271 18689
rect 11297 18663 11303 18689
rect 15465 18663 15471 18689
rect 15497 18663 15503 18689
rect 17985 18663 17991 18689
rect 18017 18663 18023 18689
rect 19329 18663 19335 18689
rect 19361 18663 19367 18689
rect 23417 18663 23423 18689
rect 23449 18663 23455 18689
rect 2137 18607 2143 18633
rect 2169 18607 2175 18633
rect 2417 18607 2423 18633
rect 2449 18607 2455 18633
rect 2529 18607 2535 18633
rect 2561 18607 2567 18633
rect 3593 18607 3599 18633
rect 3625 18607 3631 18633
rect 4433 18607 4439 18633
rect 4465 18607 4471 18633
rect 5833 18607 5839 18633
rect 5865 18607 5871 18633
rect 7009 18607 7015 18633
rect 7041 18607 7047 18633
rect 7289 18607 7295 18633
rect 7321 18607 7327 18633
rect 8409 18607 8415 18633
rect 8441 18607 8447 18633
rect 9137 18607 9143 18633
rect 9169 18607 9175 18633
rect 10033 18607 10039 18633
rect 10065 18607 10071 18633
rect 10313 18607 10319 18633
rect 10345 18607 10351 18633
rect 11265 18607 11271 18633
rect 11297 18607 11303 18633
rect 12833 18607 12839 18633
rect 12865 18607 12871 18633
rect 13393 18607 13399 18633
rect 13425 18607 13431 18633
rect 13505 18607 13511 18633
rect 13537 18607 13543 18633
rect 14569 18607 14575 18633
rect 14601 18607 14607 18633
rect 15465 18607 15471 18633
rect 15497 18607 15503 18633
rect 16865 18607 16871 18633
rect 16897 18607 16903 18633
rect 17985 18607 17991 18633
rect 18017 18607 18023 18633
rect 18545 18607 18551 18633
rect 18577 18607 18583 18633
rect 19329 18607 19335 18633
rect 19361 18607 19367 18633
rect 20953 18607 20959 18633
rect 20985 18607 20991 18633
rect 21233 18607 21239 18633
rect 21265 18607 21271 18633
rect 21457 18607 21463 18633
rect 21489 18607 21495 18633
rect 22521 18607 22527 18633
rect 22553 18607 22559 18633
rect 23417 18607 23423 18633
rect 23449 18607 23455 18633
rect 672 18437 24304 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 24304 18437
rect 672 18394 24304 18411
rect 1577 18215 1583 18241
rect 1609 18215 1615 18241
rect 2473 18215 2479 18241
rect 2505 18215 2511 18241
rect 3817 18215 3823 18241
rect 3849 18215 3855 18241
rect 4377 18215 4383 18241
rect 4409 18215 4415 18241
rect 4489 18215 4495 18241
rect 4521 18215 4527 18241
rect 5273 18215 5279 18241
rect 5305 18215 5311 18241
rect 6449 18215 6455 18241
rect 6481 18215 6487 18241
rect 8129 18215 8135 18241
rect 8161 18215 8167 18241
rect 9025 18215 9031 18241
rect 9057 18215 9063 18241
rect 10817 18215 10823 18241
rect 10849 18215 10855 18241
rect 11265 18215 11271 18241
rect 11297 18215 11303 18241
rect 11489 18215 11495 18241
rect 11521 18215 11527 18241
rect 12273 18215 12279 18241
rect 12305 18215 12311 18241
rect 13449 18215 13455 18241
rect 13481 18215 13487 18241
rect 14793 18215 14799 18241
rect 14825 18215 14831 18241
rect 15913 18215 15919 18241
rect 15945 18215 15951 18241
rect 16249 18215 16255 18241
rect 16281 18215 16287 18241
rect 17425 18215 17431 18241
rect 17457 18215 17463 18241
rect 19049 18215 19055 18241
rect 19081 18215 19087 18241
rect 19329 18215 19335 18241
rect 19361 18215 19367 18241
rect 19441 18215 19447 18241
rect 19473 18215 19479 18241
rect 20225 18215 20231 18241
rect 20257 18215 20263 18241
rect 21233 18215 21239 18241
rect 21265 18215 21271 18241
rect 22745 18215 22751 18241
rect 22777 18215 22783 18241
rect 23249 18215 23255 18241
rect 23281 18215 23287 18241
rect 23417 18215 23423 18241
rect 23449 18215 23455 18241
rect 2473 18159 2479 18185
rect 2505 18159 2511 18185
rect 6449 18159 6455 18185
rect 6481 18159 6487 18185
rect 9025 18159 9031 18185
rect 9057 18159 9063 18185
rect 13449 18159 13455 18185
rect 13481 18159 13487 18185
rect 15913 18159 15919 18185
rect 15945 18159 15951 18185
rect 17425 18159 17431 18185
rect 17457 18159 17463 18185
rect 21233 18159 21239 18185
rect 21265 18159 21271 18185
rect 672 18045 24304 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 24304 18045
rect 672 18002 24304 18019
rect 3033 17879 3039 17905
rect 3065 17879 3071 17905
rect 7009 17879 7015 17905
rect 7041 17879 7047 17905
rect 8409 17879 8415 17905
rect 8441 17879 8447 17905
rect 9809 17879 9815 17905
rect 9841 17879 9847 17905
rect 11265 17879 11271 17905
rect 11297 17879 11303 17905
rect 15465 17879 15471 17905
rect 15497 17879 15503 17905
rect 17985 17879 17991 17905
rect 18017 17879 18023 17905
rect 19329 17879 19335 17905
rect 19361 17879 19367 17905
rect 23417 17879 23423 17905
rect 23449 17879 23455 17905
rect 2137 17823 2143 17849
rect 2169 17823 2175 17849
rect 3033 17823 3039 17849
rect 3065 17823 3071 17849
rect 3593 17823 3599 17849
rect 3625 17823 3631 17849
rect 3873 17823 3879 17849
rect 3905 17823 3911 17849
rect 4153 17823 4159 17849
rect 4185 17823 4191 17849
rect 5833 17823 5839 17849
rect 5865 17823 5871 17849
rect 7009 17823 7015 17849
rect 7041 17823 7047 17849
rect 7289 17823 7295 17849
rect 7321 17823 7327 17849
rect 8409 17823 8415 17849
rect 8441 17823 8447 17849
rect 9137 17823 9143 17849
rect 9169 17823 9175 17849
rect 9809 17823 9815 17849
rect 9841 17823 9847 17849
rect 10313 17823 10319 17849
rect 10345 17823 10351 17849
rect 11265 17823 11271 17849
rect 11297 17823 11303 17849
rect 13113 17823 13119 17849
rect 13145 17823 13151 17849
rect 13393 17823 13399 17849
rect 13425 17823 13431 17849
rect 13505 17823 13511 17849
rect 13537 17823 13543 17849
rect 14569 17823 14575 17849
rect 14601 17823 14607 17849
rect 15465 17823 15471 17849
rect 15497 17823 15503 17849
rect 16865 17823 16871 17849
rect 16897 17823 16903 17849
rect 17985 17823 17991 17849
rect 18017 17823 18023 17849
rect 18545 17823 18551 17849
rect 18577 17823 18583 17849
rect 19329 17823 19335 17849
rect 19361 17823 19367 17849
rect 20953 17823 20959 17849
rect 20985 17823 20991 17849
rect 21233 17823 21239 17849
rect 21265 17823 21271 17849
rect 21457 17823 21463 17849
rect 21489 17823 21495 17849
rect 22521 17823 22527 17849
rect 22553 17823 22559 17849
rect 23417 17823 23423 17849
rect 23449 17823 23455 17849
rect 672 17653 24304 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 24304 17653
rect 672 17610 24304 17627
rect 1577 17431 1583 17457
rect 1609 17431 1615 17457
rect 2473 17431 2479 17457
rect 2505 17431 2511 17457
rect 4097 17431 4103 17457
rect 4129 17431 4135 17457
rect 4377 17431 4383 17457
rect 4409 17431 4415 17457
rect 4489 17431 4495 17457
rect 4521 17431 4527 17457
rect 5273 17431 5279 17457
rect 5305 17431 5311 17457
rect 6449 17431 6455 17457
rect 6481 17431 6487 17457
rect 8129 17431 8135 17457
rect 8161 17431 8167 17457
rect 8409 17431 8415 17457
rect 8441 17431 8447 17457
rect 8521 17431 8527 17457
rect 8553 17431 8559 17457
rect 10817 17431 10823 17457
rect 10849 17431 10855 17457
rect 11265 17431 11271 17457
rect 11297 17431 11303 17457
rect 11489 17431 11495 17457
rect 11521 17431 11527 17457
rect 12553 17431 12559 17457
rect 12585 17431 12591 17457
rect 13449 17431 13455 17457
rect 13481 17431 13487 17457
rect 14793 17431 14799 17457
rect 14825 17431 14831 17457
rect 15913 17431 15919 17457
rect 15945 17431 15951 17457
rect 16249 17431 16255 17457
rect 16281 17431 16287 17457
rect 16809 17431 16815 17457
rect 16841 17431 16847 17457
rect 16921 17431 16927 17457
rect 16953 17431 16959 17457
rect 19049 17431 19055 17457
rect 19081 17431 19087 17457
rect 19329 17431 19335 17457
rect 19361 17431 19367 17457
rect 19441 17431 19447 17457
rect 19473 17431 19479 17457
rect 20225 17431 20231 17457
rect 20257 17431 20263 17457
rect 21233 17431 21239 17457
rect 21265 17431 21271 17457
rect 22745 17431 22751 17457
rect 22777 17431 22783 17457
rect 23249 17431 23255 17457
rect 23281 17431 23287 17457
rect 23417 17431 23423 17457
rect 23449 17431 23455 17457
rect 2473 17375 2479 17401
rect 2505 17375 2511 17401
rect 6449 17375 6455 17401
rect 6481 17375 6487 17401
rect 13449 17375 13455 17401
rect 13481 17375 13487 17401
rect 15913 17375 15919 17401
rect 15945 17375 15951 17401
rect 21233 17375 21239 17401
rect 21265 17375 21271 17401
rect 672 17261 24304 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 24304 17261
rect 672 17218 24304 17235
rect 3033 17095 3039 17121
rect 3065 17095 3071 17121
rect 4433 17095 4439 17121
rect 4465 17095 4471 17121
rect 7009 17095 7015 17121
rect 7041 17095 7047 17121
rect 8409 17095 8415 17121
rect 8441 17095 8447 17121
rect 9809 17095 9815 17121
rect 9841 17095 9847 17121
rect 11265 17095 11271 17121
rect 11297 17095 11303 17121
rect 15241 17095 15247 17121
rect 15273 17095 15279 17121
rect 17985 17095 17991 17121
rect 18017 17095 18023 17121
rect 19329 17095 19335 17121
rect 19361 17095 19367 17121
rect 23249 17095 23255 17121
rect 23281 17095 23287 17121
rect 1857 17039 1863 17065
rect 1889 17039 1895 17065
rect 3033 17039 3039 17065
rect 3065 17039 3071 17065
rect 3593 17039 3599 17065
rect 3625 17039 3631 17065
rect 4433 17039 4439 17065
rect 4465 17039 4471 17065
rect 5833 17039 5839 17065
rect 5865 17039 5871 17065
rect 7009 17039 7015 17065
rect 7041 17039 7047 17065
rect 7289 17039 7295 17065
rect 7321 17039 7327 17065
rect 8409 17039 8415 17065
rect 8441 17039 8447 17065
rect 9137 17039 9143 17065
rect 9169 17039 9175 17065
rect 9809 17039 9815 17065
rect 9841 17039 9847 17065
rect 10313 17039 10319 17065
rect 10345 17039 10351 17065
rect 11265 17039 11271 17065
rect 11297 17039 11303 17065
rect 12889 17039 12895 17065
rect 12921 17039 12927 17065
rect 13393 17039 13399 17065
rect 13425 17039 13431 17065
rect 13505 17039 13511 17065
rect 13537 17039 13543 17065
rect 14401 17039 14407 17065
rect 14433 17039 14439 17065
rect 15241 17039 15247 17065
rect 15273 17039 15279 17065
rect 16977 17039 16983 17065
rect 17009 17039 17015 17065
rect 17985 17039 17991 17065
rect 18017 17039 18023 17065
rect 18545 17039 18551 17065
rect 18577 17039 18583 17065
rect 19329 17039 19335 17065
rect 19361 17039 19367 17065
rect 20953 17039 20959 17065
rect 20985 17039 20991 17065
rect 21233 17039 21239 17065
rect 21265 17039 21271 17065
rect 21457 17039 21463 17065
rect 21489 17039 21495 17065
rect 22241 17039 22247 17065
rect 22273 17039 22279 17065
rect 23249 17039 23255 17065
rect 23281 17039 23287 17065
rect 672 16869 24304 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 24304 16869
rect 672 16826 24304 16843
rect 1577 16647 1583 16673
rect 1609 16647 1615 16673
rect 2473 16647 2479 16673
rect 2505 16647 2511 16673
rect 4097 16647 4103 16673
rect 4129 16647 4135 16673
rect 4377 16647 4383 16673
rect 4409 16647 4415 16673
rect 4545 16647 4551 16673
rect 4577 16647 4583 16673
rect 5273 16647 5279 16673
rect 5305 16647 5311 16673
rect 6449 16647 6455 16673
rect 6481 16647 6487 16673
rect 8129 16647 8135 16673
rect 8161 16647 8167 16673
rect 8409 16647 8415 16673
rect 8441 16647 8447 16673
rect 8521 16647 8527 16673
rect 8553 16647 8559 16673
rect 10817 16647 10823 16673
rect 10849 16647 10855 16673
rect 11265 16647 11271 16673
rect 11297 16647 11303 16673
rect 11489 16647 11495 16673
rect 11521 16647 11527 16673
rect 12553 16647 12559 16673
rect 12585 16647 12591 16673
rect 13449 16647 13455 16673
rect 13481 16647 13487 16673
rect 14793 16647 14799 16673
rect 14825 16647 14831 16673
rect 15241 16647 15247 16673
rect 15273 16647 15279 16673
rect 15465 16647 15471 16673
rect 15497 16647 15503 16673
rect 16249 16647 16255 16673
rect 16281 16647 16287 16673
rect 16921 16647 16927 16673
rect 16953 16647 16959 16673
rect 19049 16647 19055 16673
rect 19081 16647 19087 16673
rect 19329 16647 19335 16673
rect 19361 16647 19367 16673
rect 19441 16647 19447 16673
rect 19473 16647 19479 16673
rect 20225 16647 20231 16673
rect 20257 16647 20263 16673
rect 21233 16647 21239 16673
rect 21265 16647 21271 16673
rect 22745 16647 22751 16673
rect 22777 16647 22783 16673
rect 23249 16647 23255 16673
rect 23281 16647 23287 16673
rect 23417 16647 23423 16673
rect 23449 16647 23455 16673
rect 2473 16591 2479 16617
rect 2505 16591 2511 16617
rect 6449 16591 6455 16617
rect 6481 16591 6487 16617
rect 13449 16591 13455 16617
rect 13481 16591 13487 16617
rect 17313 16591 17319 16617
rect 17345 16591 17351 16617
rect 21233 16591 21239 16617
rect 21265 16591 21271 16617
rect 672 16477 24304 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 24304 16477
rect 672 16434 24304 16451
rect 2977 16311 2983 16337
rect 3009 16311 3015 16337
rect 4321 16311 4327 16337
rect 4353 16311 4359 16337
rect 7009 16311 7015 16337
rect 7041 16311 7047 16337
rect 8409 16311 8415 16337
rect 8441 16311 8447 16337
rect 9809 16311 9815 16337
rect 9841 16311 9847 16337
rect 11265 16311 11271 16337
rect 11297 16311 11303 16337
rect 15241 16311 15247 16337
rect 15273 16311 15279 16337
rect 19217 16311 19223 16337
rect 19249 16311 19255 16337
rect 23249 16311 23255 16337
rect 23281 16311 23287 16337
rect 1857 16255 1863 16281
rect 1889 16255 1895 16281
rect 2977 16255 2983 16281
rect 3009 16255 3015 16281
rect 3593 16255 3599 16281
rect 3625 16255 3631 16281
rect 4321 16255 4327 16281
rect 4353 16255 4359 16281
rect 5833 16255 5839 16281
rect 5865 16255 5871 16281
rect 7009 16255 7015 16281
rect 7041 16255 7047 16281
rect 7289 16255 7295 16281
rect 7321 16255 7327 16281
rect 8409 16255 8415 16281
rect 8441 16255 8447 16281
rect 9137 16255 9143 16281
rect 9169 16255 9175 16281
rect 9809 16255 9815 16281
rect 9841 16255 9847 16281
rect 10593 16255 10599 16281
rect 10625 16255 10631 16281
rect 11265 16255 11271 16281
rect 11297 16255 11303 16281
rect 12889 16255 12895 16281
rect 12921 16255 12927 16281
rect 13393 16255 13399 16281
rect 13425 16255 13431 16281
rect 13505 16255 13511 16281
rect 13537 16255 13543 16281
rect 14401 16255 14407 16281
rect 14433 16255 14439 16281
rect 15241 16255 15247 16281
rect 15273 16255 15279 16281
rect 16977 16255 16983 16281
rect 17009 16255 17015 16281
rect 17313 16255 17319 16281
rect 17345 16255 17351 16281
rect 17481 16255 17487 16281
rect 17513 16255 17519 16281
rect 18545 16255 18551 16281
rect 18577 16255 18583 16281
rect 19217 16255 19223 16281
rect 19249 16255 19255 16281
rect 20953 16255 20959 16281
rect 20985 16255 20991 16281
rect 21233 16255 21239 16281
rect 21265 16255 21271 16281
rect 21457 16255 21463 16281
rect 21489 16255 21495 16281
rect 22241 16255 22247 16281
rect 22273 16255 22279 16281
rect 23249 16255 23255 16281
rect 23281 16255 23287 16281
rect 672 16085 24304 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 24304 16085
rect 672 16042 24304 16059
rect 1577 15863 1583 15889
rect 1609 15863 1615 15889
rect 2417 15863 2423 15889
rect 2449 15863 2455 15889
rect 3817 15863 3823 15889
rect 3849 15863 3855 15889
rect 4937 15863 4943 15889
rect 4969 15863 4975 15889
rect 5553 15863 5559 15889
rect 5585 15863 5591 15889
rect 5945 15863 5951 15889
rect 5977 15863 5983 15889
rect 7905 15863 7911 15889
rect 7937 15863 7943 15889
rect 9025 15863 9031 15889
rect 9057 15863 9063 15889
rect 11097 15863 11103 15889
rect 11129 15863 11135 15889
rect 11377 15863 11383 15889
rect 11409 15863 11415 15889
rect 11489 15863 11495 15889
rect 11521 15863 11527 15889
rect 12553 15863 12559 15889
rect 12585 15863 12591 15889
rect 12721 15863 12727 15889
rect 12753 15863 12759 15889
rect 12945 15863 12951 15889
rect 12977 15863 12983 15889
rect 14793 15863 14799 15889
rect 14825 15863 14831 15889
rect 15241 15863 15247 15889
rect 15273 15863 15279 15889
rect 15465 15863 15471 15889
rect 15497 15863 15503 15889
rect 16249 15863 16255 15889
rect 16281 15863 16287 15889
rect 17425 15863 17431 15889
rect 17457 15863 17463 15889
rect 19049 15863 19055 15889
rect 19081 15863 19087 15889
rect 19945 15863 19951 15889
rect 19977 15863 19983 15889
rect 20225 15863 20231 15889
rect 20257 15863 20263 15889
rect 21009 15863 21015 15889
rect 21041 15863 21047 15889
rect 22745 15863 22751 15889
rect 22777 15863 22783 15889
rect 23193 15863 23199 15889
rect 23225 15863 23231 15889
rect 23417 15863 23423 15889
rect 23449 15863 23455 15889
rect 2417 15807 2423 15833
rect 2449 15807 2455 15833
rect 4937 15807 4943 15833
rect 4969 15807 4975 15833
rect 6225 15807 6231 15833
rect 6257 15807 6263 15833
rect 9025 15807 9031 15833
rect 9057 15807 9063 15833
rect 17425 15807 17431 15833
rect 17457 15807 17463 15833
rect 19945 15807 19951 15833
rect 19977 15807 19983 15833
rect 21177 15807 21183 15833
rect 21209 15807 21215 15833
rect 672 15693 24304 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 24304 15693
rect 672 15650 24304 15667
rect 4489 15527 4495 15553
rect 4521 15527 4527 15553
rect 8465 15527 8471 15553
rect 8497 15527 8503 15553
rect 11489 15527 11495 15553
rect 11521 15527 11527 15553
rect 15241 15527 15247 15553
rect 15273 15527 15279 15553
rect 17985 15527 17991 15553
rect 18017 15527 18023 15553
rect 19273 15527 19279 15553
rect 19305 15527 19311 15553
rect 1857 15471 1863 15497
rect 1889 15471 1895 15497
rect 2417 15471 2423 15497
rect 2449 15471 2455 15497
rect 2529 15471 2535 15497
rect 2561 15471 2567 15497
rect 3593 15471 3599 15497
rect 3625 15471 3631 15497
rect 4489 15471 4495 15497
rect 4521 15471 4527 15497
rect 6113 15471 6119 15497
rect 6145 15471 6151 15497
rect 6281 15471 6287 15497
rect 6313 15471 6319 15497
rect 6505 15471 6511 15497
rect 6537 15471 6543 15497
rect 7289 15471 7295 15497
rect 7321 15471 7327 15497
rect 8465 15471 8471 15497
rect 8497 15471 8503 15497
rect 8857 15471 8863 15497
rect 8889 15471 8895 15497
rect 9305 15471 9311 15497
rect 9337 15471 9343 15497
rect 9529 15471 9535 15497
rect 9561 15471 9567 15497
rect 10593 15471 10599 15497
rect 10625 15471 10631 15497
rect 11489 15471 11495 15497
rect 11521 15471 11527 15497
rect 13113 15471 13119 15497
rect 13145 15471 13151 15497
rect 13281 15471 13287 15497
rect 13313 15471 13319 15497
rect 13505 15471 13511 15497
rect 13537 15471 13543 15497
rect 14569 15471 14575 15497
rect 14601 15471 14607 15497
rect 15241 15471 15247 15497
rect 15273 15471 15279 15497
rect 17089 15471 17095 15497
rect 17121 15471 17127 15497
rect 17985 15471 17991 15497
rect 18017 15471 18023 15497
rect 18265 15471 18271 15497
rect 18297 15471 18303 15497
rect 19273 15471 19279 15497
rect 19305 15471 19311 15497
rect 20785 15471 20791 15497
rect 20817 15471 20823 15497
rect 21233 15471 21239 15497
rect 21265 15471 21271 15497
rect 21457 15471 21463 15497
rect 21489 15471 21495 15497
rect 22241 15471 22247 15497
rect 22273 15471 22279 15497
rect 22689 15471 22695 15497
rect 22721 15471 22727 15497
rect 22913 15471 22919 15497
rect 22945 15471 22951 15497
rect 672 15301 24304 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 24304 15301
rect 672 15258 24304 15275
rect 1353 15079 1359 15105
rect 1385 15079 1391 15105
rect 2361 15079 2367 15105
rect 2393 15079 2399 15105
rect 3817 15079 3823 15105
rect 3849 15079 3855 15105
rect 4937 15079 4943 15105
rect 4969 15079 4975 15105
rect 5273 15079 5279 15105
rect 5305 15079 5311 15105
rect 6449 15079 6455 15105
rect 6481 15079 6487 15105
rect 7905 15079 7911 15105
rect 7937 15079 7943 15105
rect 9025 15079 9031 15105
rect 9057 15079 9063 15105
rect 11097 15079 11103 15105
rect 11129 15079 11135 15105
rect 11377 15079 11383 15105
rect 11409 15079 11415 15105
rect 11489 15079 11495 15105
rect 11521 15079 11527 15105
rect 12553 15079 12559 15105
rect 12585 15079 12591 15105
rect 12721 15079 12727 15105
rect 12753 15079 12759 15105
rect 12945 15079 12951 15105
rect 12977 15079 12983 15105
rect 14793 15079 14799 15105
rect 14825 15079 14831 15105
rect 15241 15079 15247 15105
rect 15273 15079 15279 15105
rect 15465 15079 15471 15105
rect 15497 15079 15503 15105
rect 16249 15079 16255 15105
rect 16281 15079 16287 15105
rect 17425 15079 17431 15105
rect 17457 15079 17463 15105
rect 19049 15079 19055 15105
rect 19081 15079 19087 15105
rect 19329 15079 19335 15105
rect 19361 15079 19367 15105
rect 19441 15079 19447 15105
rect 19473 15079 19479 15105
rect 20225 15079 20231 15105
rect 20257 15079 20263 15105
rect 21009 15079 21015 15105
rect 21041 15079 21047 15105
rect 22745 15079 22751 15105
rect 22777 15079 22783 15105
rect 23193 15079 23199 15105
rect 23225 15079 23231 15105
rect 23417 15079 23423 15105
rect 23449 15079 23455 15105
rect 2361 15023 2367 15049
rect 2393 15023 2399 15049
rect 4937 15023 4943 15049
rect 4969 15023 4975 15049
rect 6449 15023 6455 15049
rect 6481 15023 6487 15049
rect 9025 15023 9031 15049
rect 9057 15023 9063 15049
rect 17425 15023 17431 15049
rect 17457 15023 17463 15049
rect 21177 15023 21183 15049
rect 21209 15023 21215 15049
rect 672 14909 24304 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 24304 14909
rect 672 14866 24304 14883
rect 4489 14743 4495 14769
rect 4521 14743 4527 14769
rect 6169 14743 6175 14769
rect 6201 14743 6207 14769
rect 11489 14743 11495 14769
rect 11521 14743 11527 14769
rect 15241 14743 15247 14769
rect 15273 14743 15279 14769
rect 19441 14743 19447 14769
rect 19473 14743 19479 14769
rect 1857 14687 1863 14713
rect 1889 14687 1895 14713
rect 2361 14687 2367 14713
rect 2393 14687 2399 14713
rect 2585 14687 2591 14713
rect 2617 14687 2623 14713
rect 3593 14687 3599 14713
rect 3625 14687 3631 14713
rect 4489 14687 4495 14713
rect 4521 14687 4527 14713
rect 5273 14687 5279 14713
rect 5305 14687 5311 14713
rect 6169 14687 6175 14713
rect 6201 14687 6207 14713
rect 6729 14687 6735 14713
rect 6761 14687 6767 14713
rect 6897 14687 6903 14713
rect 6929 14687 6935 14713
rect 7121 14687 7127 14713
rect 7153 14687 7159 14713
rect 8857 14687 8863 14713
rect 8889 14687 8895 14713
rect 9417 14687 9423 14713
rect 9449 14687 9455 14713
rect 9529 14687 9535 14713
rect 9561 14687 9567 14713
rect 10593 14687 10599 14713
rect 10625 14687 10631 14713
rect 11489 14687 11495 14713
rect 11521 14687 11527 14713
rect 13113 14687 13119 14713
rect 13145 14687 13151 14713
rect 13281 14687 13287 14713
rect 13313 14687 13319 14713
rect 13505 14687 13511 14713
rect 13537 14687 13543 14713
rect 14569 14687 14575 14713
rect 14601 14687 14607 14713
rect 15241 14687 15247 14713
rect 15273 14687 15279 14713
rect 17089 14687 17095 14713
rect 17121 14687 17127 14713
rect 17369 14687 17375 14713
rect 17401 14687 17407 14713
rect 17481 14687 17487 14713
rect 17513 14687 17519 14713
rect 18265 14687 18271 14713
rect 18297 14687 18303 14713
rect 19441 14687 19447 14713
rect 19473 14687 19479 14713
rect 20785 14687 20791 14713
rect 20817 14687 20823 14713
rect 21233 14687 21239 14713
rect 21265 14687 21271 14713
rect 21457 14687 21463 14713
rect 21489 14687 21495 14713
rect 22241 14687 22247 14713
rect 22273 14687 22279 14713
rect 22745 14687 22751 14713
rect 22777 14687 22783 14713
rect 22913 14687 22919 14713
rect 22945 14687 22951 14713
rect 672 14517 24304 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 24304 14517
rect 672 14474 24304 14491
rect 1577 14295 1583 14321
rect 1609 14295 1615 14321
rect 2137 14295 2143 14321
rect 2169 14295 2175 14321
rect 3817 14295 3823 14321
rect 3849 14295 3855 14321
rect 4993 14295 4999 14321
rect 5025 14295 5031 14321
rect 5553 14295 5559 14321
rect 5585 14295 5591 14321
rect 6169 14295 6175 14321
rect 6201 14295 6207 14321
rect 6841 14295 6847 14321
rect 6873 14295 6879 14321
rect 7289 14295 7295 14321
rect 7321 14295 7327 14321
rect 7513 14295 7519 14321
rect 7545 14295 7551 14321
rect 8409 14295 8415 14321
rect 8441 14295 8447 14321
rect 9417 14295 9423 14321
rect 9449 14295 9455 14321
rect 11097 14295 11103 14321
rect 11129 14295 11135 14321
rect 11377 14295 11383 14321
rect 11409 14295 11415 14321
rect 11489 14295 11495 14321
rect 11521 14295 11527 14321
rect 12553 14295 12559 14321
rect 12585 14295 12591 14321
rect 12721 14295 12727 14321
rect 12753 14295 12759 14321
rect 12945 14295 12951 14321
rect 12977 14295 12983 14321
rect 14793 14295 14799 14321
rect 14825 14295 14831 14321
rect 15241 14295 15247 14321
rect 15273 14295 15279 14321
rect 15465 14295 15471 14321
rect 15497 14295 15503 14321
rect 16249 14295 16255 14321
rect 16281 14295 16287 14321
rect 17425 14295 17431 14321
rect 17457 14295 17463 14321
rect 19049 14295 19055 14321
rect 19081 14295 19087 14321
rect 19329 14295 19335 14321
rect 19361 14295 19367 14321
rect 19441 14295 19447 14321
rect 19473 14295 19479 14321
rect 20225 14295 20231 14321
rect 20257 14295 20263 14321
rect 21009 14295 21015 14321
rect 21041 14295 21047 14321
rect 22857 14295 22863 14321
rect 22889 14295 22895 14321
rect 24033 14295 24039 14321
rect 24065 14295 24071 14321
rect 2249 14239 2255 14265
rect 2281 14239 2287 14265
rect 4993 14239 4999 14265
rect 5025 14239 5031 14265
rect 6225 14239 6231 14265
rect 6257 14239 6263 14265
rect 9417 14239 9423 14265
rect 9449 14239 9455 14265
rect 17425 14239 17431 14265
rect 17457 14239 17463 14265
rect 21177 14239 21183 14265
rect 21209 14239 21215 14265
rect 22857 14239 22863 14265
rect 22889 14239 22895 14265
rect 672 14125 24304 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 24304 14125
rect 672 14082 24304 14099
rect 4489 13959 4495 13985
rect 4521 13959 4527 13985
rect 8185 13959 8191 13985
rect 8217 13959 8223 13985
rect 11489 13959 11495 13985
rect 11521 13959 11527 13985
rect 15241 13959 15247 13985
rect 15273 13959 15279 13985
rect 19441 13959 19447 13985
rect 19473 13959 19479 13985
rect 22857 13959 22863 13985
rect 22889 13959 22895 13985
rect 2137 13903 2143 13929
rect 2169 13903 2175 13929
rect 2305 13903 2311 13929
rect 2337 13903 2343 13929
rect 2529 13903 2535 13929
rect 2561 13903 2567 13929
rect 3369 13903 3375 13929
rect 3401 13903 3407 13929
rect 4489 13903 4495 13929
rect 4521 13903 4527 13929
rect 5553 13903 5559 13929
rect 5585 13903 5591 13929
rect 6113 13903 6119 13929
rect 6145 13903 6151 13929
rect 6225 13903 6231 13929
rect 6257 13903 6263 13929
rect 7009 13903 7015 13929
rect 7041 13903 7047 13929
rect 8185 13903 8191 13929
rect 8217 13903 8223 13929
rect 8857 13903 8863 13929
rect 8889 13903 8895 13929
rect 9417 13903 9423 13929
rect 9449 13903 9455 13929
rect 9529 13903 9535 13929
rect 9561 13903 9567 13929
rect 10593 13903 10599 13929
rect 10625 13903 10631 13929
rect 11489 13903 11495 13929
rect 11521 13903 11527 13929
rect 13113 13903 13119 13929
rect 13145 13903 13151 13929
rect 13281 13903 13287 13929
rect 13313 13903 13319 13929
rect 13505 13903 13511 13929
rect 13537 13903 13543 13929
rect 14569 13903 14575 13929
rect 14601 13903 14607 13929
rect 15241 13903 15247 13929
rect 15273 13903 15279 13929
rect 17089 13903 17095 13929
rect 17121 13903 17127 13929
rect 17369 13903 17375 13929
rect 17401 13903 17407 13929
rect 17481 13903 17487 13929
rect 17513 13903 17519 13929
rect 18265 13903 18271 13929
rect 18297 13903 18303 13929
rect 19441 13903 19447 13929
rect 19473 13903 19479 13929
rect 20953 13903 20959 13929
rect 20985 13903 20991 13929
rect 21233 13903 21239 13929
rect 21265 13903 21271 13929
rect 21457 13903 21463 13929
rect 21489 13903 21495 13929
rect 22857 13903 22863 13929
rect 22889 13903 22895 13929
rect 24033 13903 24039 13929
rect 24065 13903 24071 13929
rect 672 13733 24304 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 24304 13733
rect 672 13690 24304 13707
rect 1577 13511 1583 13537
rect 1609 13511 1615 13537
rect 2473 13511 2479 13537
rect 2505 13511 2511 13537
rect 3817 13511 3823 13537
rect 3849 13511 3855 13537
rect 4993 13511 4999 13537
rect 5025 13511 5031 13537
rect 5497 13511 5503 13537
rect 5529 13511 5535 13537
rect 6113 13511 6119 13537
rect 6145 13511 6151 13537
rect 7009 13511 7015 13537
rect 7041 13511 7047 13537
rect 8185 13511 8191 13537
rect 8217 13511 8223 13537
rect 8465 13511 8471 13537
rect 8497 13511 8503 13537
rect 9417 13511 9423 13537
rect 9449 13511 9455 13537
rect 11097 13511 11103 13537
rect 11129 13511 11135 13537
rect 11377 13511 11383 13537
rect 11409 13511 11415 13537
rect 11489 13511 11495 13537
rect 11521 13511 11527 13537
rect 12553 13511 12559 13537
rect 12585 13511 12591 13537
rect 12721 13511 12727 13537
rect 12753 13511 12759 13537
rect 12945 13511 12951 13537
rect 12977 13511 12983 13537
rect 14793 13511 14799 13537
rect 14825 13511 14831 13537
rect 15241 13511 15247 13537
rect 15273 13511 15279 13537
rect 15465 13511 15471 13537
rect 15497 13511 15503 13537
rect 16249 13511 16255 13537
rect 16281 13511 16287 13537
rect 17425 13511 17431 13537
rect 17457 13511 17463 13537
rect 19049 13511 19055 13537
rect 19081 13511 19087 13537
rect 19329 13511 19335 13537
rect 19361 13511 19367 13537
rect 19441 13511 19447 13537
rect 19473 13511 19479 13537
rect 20505 13511 20511 13537
rect 20537 13511 20543 13537
rect 21401 13511 21407 13537
rect 21433 13511 21439 13537
rect 22857 13511 22863 13537
rect 22889 13511 22895 13537
rect 24033 13511 24039 13537
rect 24065 13511 24071 13537
rect 2473 13455 2479 13481
rect 2505 13455 2511 13481
rect 4993 13455 4999 13481
rect 5025 13455 5031 13481
rect 6225 13455 6231 13481
rect 6257 13455 6263 13481
rect 8185 13455 8191 13481
rect 8217 13455 8223 13481
rect 9417 13455 9423 13481
rect 9449 13455 9455 13481
rect 17425 13455 17431 13481
rect 17457 13455 17463 13481
rect 21401 13455 21407 13481
rect 21433 13455 21439 13481
rect 22857 13455 22863 13481
rect 22889 13455 22895 13481
rect 672 13341 24304 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 24304 13341
rect 672 13298 24304 13315
rect 4489 13175 4495 13201
rect 4521 13175 4527 13201
rect 8129 13175 8135 13201
rect 8161 13175 8167 13201
rect 11489 13175 11495 13201
rect 11521 13175 11527 13201
rect 15241 13175 15247 13201
rect 15273 13175 15279 13201
rect 22857 13175 22863 13201
rect 22889 13175 22895 13201
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 2417 13119 2423 13145
rect 2449 13119 2455 13145
rect 2529 13119 2535 13145
rect 2561 13119 2567 13145
rect 3369 13119 3375 13145
rect 3401 13119 3407 13145
rect 4489 13119 4495 13145
rect 4521 13119 4527 13145
rect 5497 13119 5503 13145
rect 5529 13119 5535 13145
rect 6057 13119 6063 13145
rect 6089 13119 6095 13145
rect 6225 13119 6231 13145
rect 6257 13119 6263 13145
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 8129 13119 8135 13145
rect 8161 13119 8167 13145
rect 8857 13119 8863 13145
rect 8889 13119 8895 13145
rect 9417 13119 9423 13145
rect 9449 13119 9455 13145
rect 9529 13119 9535 13145
rect 9561 13119 9567 13145
rect 10593 13119 10599 13145
rect 10625 13119 10631 13145
rect 11489 13119 11495 13145
rect 11521 13119 11527 13145
rect 13113 13119 13119 13145
rect 13145 13119 13151 13145
rect 13281 13119 13287 13145
rect 13313 13119 13319 13145
rect 13505 13119 13511 13145
rect 13537 13119 13543 13145
rect 14569 13119 14575 13145
rect 14601 13119 14607 13145
rect 15241 13119 15247 13145
rect 15273 13119 15279 13145
rect 17089 13119 17095 13145
rect 17121 13119 17127 13145
rect 17257 13119 17263 13145
rect 17289 13119 17295 13145
rect 17481 13119 17487 13145
rect 17513 13119 17519 13145
rect 18265 13119 18271 13145
rect 18297 13119 18303 13145
rect 18713 13119 18719 13145
rect 18745 13119 18751 13145
rect 18937 13119 18943 13145
rect 18969 13119 18975 13145
rect 20953 13119 20959 13145
rect 20985 13119 20991 13145
rect 21233 13119 21239 13145
rect 21265 13119 21271 13145
rect 21457 13119 21463 13145
rect 21489 13119 21495 13145
rect 22857 13119 22863 13145
rect 22889 13119 22895 13145
rect 24033 13119 24039 13145
rect 24065 13119 24071 13145
rect 672 12949 24304 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 24304 12949
rect 672 12906 24304 12923
rect 1577 12727 1583 12753
rect 1609 12727 1615 12753
rect 2361 12727 2367 12753
rect 2393 12727 2399 12753
rect 3817 12727 3823 12753
rect 3849 12727 3855 12753
rect 4993 12727 4999 12753
rect 5025 12727 5031 12753
rect 5497 12727 5503 12753
rect 5529 12727 5535 12753
rect 6057 12727 6063 12753
rect 6089 12727 6095 12753
rect 7009 12727 7015 12753
rect 7041 12727 7047 12753
rect 8185 12727 8191 12753
rect 8217 12727 8223 12753
rect 8465 12727 8471 12753
rect 8497 12727 8503 12753
rect 9417 12727 9423 12753
rect 9449 12727 9455 12753
rect 11097 12727 11103 12753
rect 11129 12727 11135 12753
rect 11377 12727 11383 12753
rect 11409 12727 11415 12753
rect 11489 12727 11495 12753
rect 11521 12727 11527 12753
rect 12553 12727 12559 12753
rect 12585 12727 12591 12753
rect 12721 12727 12727 12753
rect 12753 12727 12759 12753
rect 12945 12727 12951 12753
rect 12977 12727 12983 12753
rect 14793 12727 14799 12753
rect 14825 12727 14831 12753
rect 15241 12727 15247 12753
rect 15273 12727 15279 12753
rect 15465 12727 15471 12753
rect 15497 12727 15503 12753
rect 16249 12727 16255 12753
rect 16281 12727 16287 12753
rect 17257 12727 17263 12753
rect 17289 12727 17295 12753
rect 19049 12727 19055 12753
rect 19081 12727 19087 12753
rect 19329 12727 19335 12753
rect 19361 12727 19367 12753
rect 19441 12727 19447 12753
rect 19473 12727 19479 12753
rect 20505 12727 20511 12753
rect 20537 12727 20543 12753
rect 21233 12727 21239 12753
rect 21265 12727 21271 12753
rect 22857 12727 22863 12753
rect 22889 12727 22895 12753
rect 24033 12727 24039 12753
rect 24065 12727 24071 12753
rect 2361 12671 2367 12697
rect 2393 12671 2399 12697
rect 4993 12671 4999 12697
rect 5025 12671 5031 12697
rect 6225 12671 6231 12697
rect 6257 12671 6263 12697
rect 8185 12671 8191 12697
rect 8217 12671 8223 12697
rect 9417 12671 9423 12697
rect 9449 12671 9455 12697
rect 17257 12671 17263 12697
rect 17289 12671 17295 12697
rect 21233 12671 21239 12697
rect 21265 12671 21271 12697
rect 22857 12671 22863 12697
rect 22889 12671 22895 12697
rect 672 12557 24304 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 24304 12557
rect 672 12514 24304 12531
rect 8129 12391 8135 12417
rect 8161 12391 8167 12417
rect 11489 12391 11495 12417
rect 11521 12391 11527 12417
rect 15241 12391 15247 12417
rect 15273 12391 15279 12417
rect 19273 12391 19279 12417
rect 19305 12391 19311 12417
rect 22857 12391 22863 12417
rect 22889 12391 22895 12417
rect 2137 12335 2143 12361
rect 2169 12335 2175 12361
rect 2417 12335 2423 12361
rect 2449 12335 2455 12361
rect 2529 12335 2535 12361
rect 2561 12335 2567 12361
rect 3593 12335 3599 12361
rect 3625 12335 3631 12361
rect 3761 12335 3767 12361
rect 3793 12335 3799 12361
rect 3985 12335 3991 12361
rect 4017 12335 4023 12361
rect 5497 12335 5503 12361
rect 5529 12335 5535 12361
rect 6057 12335 6063 12361
rect 6089 12335 6095 12361
rect 6225 12335 6231 12361
rect 6257 12335 6263 12361
rect 6953 12335 6959 12361
rect 6985 12335 6991 12361
rect 8129 12335 8135 12361
rect 8161 12335 8167 12361
rect 8857 12335 8863 12361
rect 8889 12335 8895 12361
rect 9417 12335 9423 12361
rect 9449 12335 9455 12361
rect 9529 12335 9535 12361
rect 9561 12335 9567 12361
rect 10593 12335 10599 12361
rect 10625 12335 10631 12361
rect 11489 12335 11495 12361
rect 11521 12335 11527 12361
rect 13113 12335 13119 12361
rect 13145 12335 13151 12361
rect 13281 12335 13287 12361
rect 13313 12335 13319 12361
rect 13505 12335 13511 12361
rect 13537 12335 13543 12361
rect 14569 12335 14575 12361
rect 14601 12335 14607 12361
rect 15129 12335 15135 12361
rect 15161 12335 15167 12361
rect 17089 12335 17095 12361
rect 17121 12335 17127 12361
rect 17257 12335 17263 12361
rect 17289 12335 17295 12361
rect 17481 12335 17487 12361
rect 17513 12335 17519 12361
rect 18545 12335 18551 12361
rect 18577 12335 18583 12361
rect 19273 12335 19279 12361
rect 19305 12335 19311 12361
rect 21625 12335 21631 12361
rect 21657 12335 21663 12361
rect 22129 12335 22135 12361
rect 22161 12335 22167 12361
rect 22577 12335 22583 12361
rect 22609 12335 22615 12361
rect 22857 12335 22863 12361
rect 22889 12335 22895 12361
rect 24033 12335 24039 12361
rect 24065 12335 24071 12361
rect 672 12165 24304 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 24304 12165
rect 672 12122 24304 12139
rect 1577 11943 1583 11969
rect 1609 11943 1615 11969
rect 2473 11943 2479 11969
rect 2505 11943 2511 11969
rect 3313 11943 3319 11969
rect 3345 11943 3351 11969
rect 3761 11943 3767 11969
rect 3793 11943 3799 11969
rect 4489 11943 4495 11969
rect 4521 11943 4527 11969
rect 5665 11943 5671 11969
rect 5697 11943 5703 11969
rect 7009 11943 7015 11969
rect 7041 11943 7047 11969
rect 8185 11943 8191 11969
rect 8217 11943 8223 11969
rect 8465 11943 8471 11969
rect 8497 11943 8503 11969
rect 9417 11943 9423 11969
rect 9449 11943 9455 11969
rect 11097 11943 11103 11969
rect 11129 11943 11135 11969
rect 11377 11943 11383 11969
rect 11409 11943 11415 11969
rect 11489 11943 11495 11969
rect 11521 11943 11527 11969
rect 12553 11943 12559 11969
rect 12585 11943 12591 11969
rect 12721 11943 12727 11969
rect 12753 11943 12759 11969
rect 12945 11943 12951 11969
rect 12977 11943 12983 11969
rect 14793 11943 14799 11969
rect 14825 11943 14831 11969
rect 15913 11943 15919 11969
rect 15945 11943 15951 11969
rect 16249 11943 16255 11969
rect 16281 11943 16287 11969
rect 17425 11943 17431 11969
rect 17457 11943 17463 11969
rect 19049 11943 19055 11969
rect 19081 11943 19087 11969
rect 19217 11943 19223 11969
rect 19249 11943 19255 11969
rect 19441 11943 19447 11969
rect 19473 11943 19479 11969
rect 21625 11943 21631 11969
rect 21657 11943 21663 11969
rect 21793 11943 21799 11969
rect 21825 11943 21831 11969
rect 22353 11943 22359 11969
rect 22385 11943 22391 11969
rect 22857 11943 22863 11969
rect 22889 11943 22895 11969
rect 24033 11943 24039 11969
rect 24065 11943 24071 11969
rect 2473 11887 2479 11913
rect 2505 11887 2511 11913
rect 3985 11887 3991 11913
rect 4017 11887 4023 11913
rect 5665 11887 5671 11913
rect 5697 11887 5703 11913
rect 8185 11887 8191 11913
rect 8217 11887 8223 11913
rect 9417 11887 9423 11913
rect 9449 11887 9455 11913
rect 15913 11887 15919 11913
rect 15945 11887 15951 11913
rect 17425 11887 17431 11913
rect 17457 11887 17463 11913
rect 22857 11887 22863 11913
rect 22889 11887 22895 11913
rect 672 11773 24304 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 24304 11773
rect 672 11730 24304 11747
rect 2865 11607 2871 11633
rect 2897 11607 2903 11633
rect 4489 11607 4495 11633
rect 4521 11607 4527 11633
rect 5833 11607 5839 11633
rect 5865 11607 5871 11633
rect 8185 11607 8191 11633
rect 8217 11607 8223 11633
rect 10033 11607 10039 11633
rect 10065 11607 10071 11633
rect 11489 11607 11495 11633
rect 11521 11607 11527 11633
rect 15465 11607 15471 11633
rect 15497 11607 15503 11633
rect 17817 11607 17823 11633
rect 17849 11607 17855 11633
rect 21625 11607 21631 11633
rect 21657 11607 21663 11633
rect 22857 11607 22863 11633
rect 22889 11607 22895 11633
rect 2137 11551 2143 11577
rect 2169 11551 2175 11577
rect 2865 11551 2871 11577
rect 2897 11551 2903 11577
rect 3425 11551 3431 11577
rect 3457 11551 3463 11577
rect 4489 11551 4495 11577
rect 4521 11551 4527 11577
rect 5049 11551 5055 11577
rect 5081 11551 5087 11577
rect 5833 11551 5839 11577
rect 5865 11551 5871 11577
rect 7289 11551 7295 11577
rect 7321 11551 7327 11577
rect 8185 11551 8191 11577
rect 8217 11551 8223 11577
rect 8857 11551 8863 11577
rect 8889 11551 8895 11577
rect 10033 11551 10039 11577
rect 10065 11551 10071 11577
rect 10593 11551 10599 11577
rect 10625 11551 10631 11577
rect 11489 11551 11495 11577
rect 11521 11551 11527 11577
rect 13113 11551 13119 11577
rect 13145 11551 13151 11577
rect 13281 11551 13287 11577
rect 13313 11551 13319 11577
rect 13505 11551 13511 11577
rect 13537 11551 13543 11577
rect 14569 11551 14575 11577
rect 14601 11551 14607 11577
rect 15465 11551 15471 11577
rect 15497 11551 15503 11577
rect 17089 11551 17095 11577
rect 17121 11551 17127 11577
rect 17817 11551 17823 11577
rect 17849 11551 17855 11577
rect 18433 11551 18439 11577
rect 18465 11551 18471 11577
rect 18713 11551 18719 11577
rect 18745 11551 18751 11577
rect 18937 11551 18943 11577
rect 18969 11551 18975 11577
rect 21681 11551 21687 11577
rect 21713 11551 21719 11577
rect 22577 11551 22583 11577
rect 22609 11551 22615 11577
rect 22857 11551 22863 11577
rect 22889 11551 22895 11577
rect 24033 11551 24039 11577
rect 24065 11551 24071 11577
rect 672 11381 24304 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 24304 11381
rect 672 11338 24304 11355
rect 1577 11159 1583 11185
rect 1609 11159 1615 11185
rect 2473 11159 2479 11185
rect 2505 11159 2511 11185
rect 3425 11159 3431 11185
rect 3457 11159 3463 11185
rect 4601 11159 4607 11185
rect 4633 11159 4639 11185
rect 5049 11159 5055 11185
rect 5081 11159 5087 11185
rect 5833 11159 5839 11185
rect 5865 11159 5871 11185
rect 7233 11159 7239 11185
rect 7265 11159 7271 11185
rect 8073 11159 8079 11185
rect 8105 11159 8111 11185
rect 8409 11159 8415 11185
rect 8441 11159 8447 11185
rect 9417 11159 9423 11185
rect 9449 11159 9455 11185
rect 11097 11159 11103 11185
rect 11129 11159 11135 11185
rect 11377 11159 11383 11185
rect 11409 11159 11415 11185
rect 11489 11159 11495 11185
rect 11521 11159 11527 11185
rect 12553 11159 12559 11185
rect 12585 11159 12591 11185
rect 12721 11159 12727 11185
rect 12753 11159 12759 11185
rect 12945 11159 12951 11185
rect 12977 11159 12983 11185
rect 14793 11159 14799 11185
rect 14825 11159 14831 11185
rect 15353 11159 15359 11185
rect 15385 11159 15391 11185
rect 15465 11159 15471 11185
rect 15497 11159 15503 11185
rect 16529 11159 16535 11185
rect 16561 11159 16567 11185
rect 16809 11159 16815 11185
rect 16841 11159 16847 11185
rect 16921 11159 16927 11185
rect 16953 11159 16959 11185
rect 20225 11159 20231 11185
rect 20257 11159 20263 11185
rect 20393 11159 20399 11185
rect 20425 11159 20431 11185
rect 20897 11159 20903 11185
rect 20929 11159 20935 11185
rect 21681 11159 21687 11185
rect 21713 11159 21719 11185
rect 21793 11159 21799 11185
rect 21825 11159 21831 11185
rect 22353 11159 22359 11185
rect 22385 11159 22391 11185
rect 22969 11159 22975 11185
rect 23001 11159 23007 11185
rect 24033 11159 24039 11185
rect 24065 11159 24071 11185
rect 2473 11103 2479 11129
rect 2505 11103 2511 11129
rect 4601 11103 4607 11129
rect 4633 11103 4639 11129
rect 5833 11103 5839 11129
rect 5865 11103 5871 11129
rect 8073 11103 8079 11129
rect 8105 11103 8111 11129
rect 9417 11103 9423 11129
rect 9449 11103 9455 11129
rect 22969 11103 22975 11129
rect 23001 11103 23007 11129
rect 672 10989 24304 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 24304 10989
rect 672 10946 24304 10963
rect 2809 10823 2815 10849
rect 2841 10823 2847 10849
rect 4489 10823 4495 10849
rect 4521 10823 4527 10849
rect 5833 10823 5839 10849
rect 5865 10823 5871 10849
rect 8073 10823 8079 10849
rect 8105 10823 8111 10849
rect 11489 10823 11495 10849
rect 11521 10823 11527 10849
rect 13785 10823 13791 10849
rect 13817 10823 13823 10849
rect 15353 10823 15359 10849
rect 15385 10823 15391 10849
rect 17761 10823 17767 10849
rect 17793 10823 17799 10849
rect 20393 10823 20399 10849
rect 20425 10823 20431 10849
rect 22969 10823 22975 10849
rect 23001 10823 23007 10849
rect 2137 10767 2143 10793
rect 2169 10767 2175 10793
rect 2809 10767 2815 10793
rect 2841 10767 2847 10793
rect 3425 10767 3431 10793
rect 3457 10767 3463 10793
rect 4489 10767 4495 10793
rect 4521 10767 4527 10793
rect 5049 10767 5055 10793
rect 5081 10767 5087 10793
rect 5833 10767 5839 10793
rect 5865 10767 5871 10793
rect 7233 10767 7239 10793
rect 7265 10767 7271 10793
rect 8073 10767 8079 10793
rect 8105 10767 8111 10793
rect 8857 10767 8863 10793
rect 8889 10767 8895 10793
rect 9417 10767 9423 10793
rect 9449 10767 9455 10793
rect 9585 10767 9591 10793
rect 9617 10767 9623 10793
rect 10593 10767 10599 10793
rect 10625 10767 10631 10793
rect 11489 10767 11495 10793
rect 11521 10767 11527 10793
rect 13113 10767 13119 10793
rect 13145 10767 13151 10793
rect 13785 10767 13791 10793
rect 13817 10767 13823 10793
rect 14569 10767 14575 10793
rect 14601 10767 14607 10793
rect 15353 10767 15359 10793
rect 15385 10767 15391 10793
rect 17089 10767 17095 10793
rect 17121 10767 17127 10793
rect 17761 10767 17767 10793
rect 17793 10767 17799 10793
rect 19441 10767 19447 10793
rect 19473 10767 19479 10793
rect 20393 10767 20399 10793
rect 20425 10767 20431 10793
rect 21625 10767 21631 10793
rect 21657 10767 21663 10793
rect 21849 10767 21855 10793
rect 21881 10767 21887 10793
rect 22073 10767 22079 10793
rect 22105 10767 22111 10793
rect 22969 10767 22975 10793
rect 23001 10767 23007 10793
rect 24033 10767 24039 10793
rect 24065 10767 24071 10793
rect 672 10597 24304 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 24304 10597
rect 672 10554 24304 10571
rect 1577 10375 1583 10401
rect 1609 10375 1615 10401
rect 2473 10375 2479 10401
rect 2505 10375 2511 10401
rect 3425 10375 3431 10401
rect 3457 10375 3463 10401
rect 4601 10375 4607 10401
rect 4633 10375 4639 10401
rect 5049 10375 5055 10401
rect 5081 10375 5087 10401
rect 5833 10375 5839 10401
rect 5865 10375 5871 10401
rect 7233 10375 7239 10401
rect 7265 10375 7271 10401
rect 8073 10375 8079 10401
rect 8105 10375 8111 10401
rect 8409 10375 8415 10401
rect 8441 10375 8447 10401
rect 9585 10375 9591 10401
rect 9617 10375 9623 10401
rect 11097 10375 11103 10401
rect 11129 10375 11135 10401
rect 11377 10375 11383 10401
rect 11409 10375 11415 10401
rect 11489 10375 11495 10401
rect 11521 10375 11527 10401
rect 12553 10375 12559 10401
rect 12585 10375 12591 10401
rect 13449 10375 13455 10401
rect 13481 10375 13487 10401
rect 14793 10375 14799 10401
rect 14825 10375 14831 10401
rect 15353 10375 15359 10401
rect 15385 10375 15391 10401
rect 15465 10375 15471 10401
rect 15497 10375 15503 10401
rect 16473 10375 16479 10401
rect 16505 10375 16511 10401
rect 16809 10375 16815 10401
rect 16841 10375 16847 10401
rect 16921 10375 16927 10401
rect 16953 10375 16959 10401
rect 20001 10375 20007 10401
rect 20033 10375 20039 10401
rect 20897 10375 20903 10401
rect 20929 10375 20935 10401
rect 21457 10375 21463 10401
rect 21489 10375 21495 10401
rect 22073 10375 22079 10401
rect 22105 10375 22111 10401
rect 22969 10375 22975 10401
rect 23001 10375 23007 10401
rect 24033 10375 24039 10401
rect 24065 10375 24071 10401
rect 2473 10319 2479 10345
rect 2505 10319 2511 10345
rect 4601 10319 4607 10345
rect 4633 10319 4639 10345
rect 5833 10319 5839 10345
rect 5865 10319 5871 10345
rect 8073 10319 8079 10345
rect 8105 10319 8111 10345
rect 9585 10319 9591 10345
rect 9617 10319 9623 10345
rect 13449 10319 13455 10345
rect 13481 10319 13487 10345
rect 20897 10319 20903 10345
rect 20929 10319 20935 10345
rect 22129 10319 22135 10345
rect 22161 10319 22167 10345
rect 22969 10319 22975 10345
rect 23001 10319 23007 10345
rect 672 10205 24304 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 24304 10205
rect 672 10162 24304 10179
rect 4489 10039 4495 10065
rect 4521 10039 4527 10065
rect 6673 10039 6679 10065
rect 6705 10039 6711 10065
rect 8129 10039 8135 10065
rect 8161 10039 8167 10065
rect 9809 10039 9815 10065
rect 9841 10039 9847 10065
rect 14009 10039 14015 10065
rect 14041 10039 14047 10065
rect 15353 10039 15359 10065
rect 15385 10039 15391 10065
rect 17985 10039 17991 10065
rect 18017 10039 18023 10065
rect 22577 10039 22583 10065
rect 22609 10039 22615 10065
rect 22913 10039 22919 10065
rect 22945 10039 22951 10065
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 2417 9983 2423 10009
rect 2449 9983 2455 10009
rect 2529 9983 2535 10009
rect 2561 9983 2567 10009
rect 3593 9983 3599 10009
rect 3625 9983 3631 10009
rect 4489 9983 4495 10009
rect 4521 9983 4527 10009
rect 5497 9983 5503 10009
rect 5529 9983 5535 10009
rect 6673 9983 6679 10009
rect 6705 9983 6711 10009
rect 7233 9983 7239 10009
rect 7265 9983 7271 10009
rect 8129 9983 8135 10009
rect 8161 9983 8167 10009
rect 9137 9983 9143 10009
rect 9169 9983 9175 10009
rect 9809 9983 9815 10009
rect 9841 9983 9847 10009
rect 10313 9983 10319 10009
rect 10345 9983 10351 10009
rect 10873 9983 10879 10009
rect 10905 9983 10911 10009
rect 10985 9983 10991 10009
rect 11017 9983 11023 10009
rect 12833 9983 12839 10009
rect 12865 9983 12871 10009
rect 14009 9983 14015 10009
rect 14041 9983 14047 10009
rect 14289 9983 14295 10009
rect 14321 9983 14327 10009
rect 15353 9983 15359 10009
rect 15385 9983 15391 10009
rect 17089 9983 17095 10009
rect 17121 9983 17127 10009
rect 17985 9983 17991 10009
rect 18017 9983 18023 10009
rect 21681 9983 21687 10009
rect 21713 9983 21719 10009
rect 22577 9983 22583 10009
rect 22609 9983 22615 10009
rect 22913 9983 22919 10009
rect 22945 9983 22951 10009
rect 23753 9983 23759 10009
rect 23785 9983 23791 10009
rect 672 9813 24304 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 24304 9813
rect 672 9770 24304 9787
rect 1353 9591 1359 9617
rect 1385 9591 1391 9617
rect 2473 9591 2479 9617
rect 2505 9591 2511 9617
rect 3817 9591 3823 9617
rect 3849 9591 3855 9617
rect 4377 9591 4383 9617
rect 4409 9591 4415 9617
rect 4489 9591 4495 9617
rect 4521 9591 4527 9617
rect 5441 9591 5447 9617
rect 5473 9591 5479 9617
rect 6449 9591 6455 9617
rect 6481 9591 6487 9617
rect 7177 9591 7183 9617
rect 7209 9591 7215 9617
rect 8073 9591 8079 9617
rect 8105 9591 8111 9617
rect 8633 9591 8639 9617
rect 8665 9591 8671 9617
rect 9529 9591 9535 9617
rect 9561 9591 9567 9617
rect 11097 9591 11103 9617
rect 11129 9591 11135 9617
rect 11377 9591 11383 9617
rect 11409 9591 11415 9617
rect 11489 9591 11495 9617
rect 11521 9591 11527 9617
rect 12273 9591 12279 9617
rect 12305 9591 12311 9617
rect 13449 9591 13455 9617
rect 13481 9591 13487 9617
rect 14793 9591 14799 9617
rect 14825 9591 14831 9617
rect 15745 9591 15751 9617
rect 15777 9591 15783 9617
rect 16529 9591 16535 9617
rect 16561 9591 16567 9617
rect 17425 9591 17431 9617
rect 17457 9591 17463 9617
rect 21177 9591 21183 9617
rect 21209 9591 21215 9617
rect 22353 9591 22359 9617
rect 22385 9591 22391 9617
rect 22913 9591 22919 9617
rect 22945 9591 22951 9617
rect 23753 9591 23759 9617
rect 23785 9591 23791 9617
rect 2473 9535 2479 9561
rect 2505 9535 2511 9561
rect 6449 9535 6455 9561
rect 6481 9535 6487 9561
rect 8073 9535 8079 9561
rect 8105 9535 8111 9561
rect 9529 9535 9535 9561
rect 9561 9535 9567 9561
rect 13449 9535 13455 9561
rect 13481 9535 13487 9561
rect 15745 9535 15751 9561
rect 15777 9535 15783 9561
rect 17425 9535 17431 9561
rect 17457 9535 17463 9561
rect 22353 9535 22359 9561
rect 22385 9535 22391 9561
rect 22913 9535 22919 9561
rect 22945 9535 22951 9561
rect 672 9421 24304 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 24304 9421
rect 672 9378 24304 9395
rect 4489 9255 4495 9281
rect 4521 9255 4527 9281
rect 6673 9255 6679 9281
rect 6705 9255 6711 9281
rect 8129 9255 8135 9281
rect 8161 9255 8167 9281
rect 10033 9255 10039 9281
rect 10065 9255 10071 9281
rect 11489 9255 11495 9281
rect 11521 9255 11527 9281
rect 15465 9255 15471 9281
rect 15497 9255 15503 9281
rect 17985 9255 17991 9281
rect 18017 9255 18023 9281
rect 19217 9255 19223 9281
rect 19249 9255 19255 9281
rect 22577 9255 22583 9281
rect 22609 9255 22615 9281
rect 22913 9255 22919 9281
rect 22945 9255 22951 9281
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 2417 9199 2423 9225
rect 2449 9199 2455 9225
rect 2529 9199 2535 9225
rect 2561 9199 2567 9225
rect 3593 9199 3599 9225
rect 3625 9199 3631 9225
rect 4489 9199 4495 9225
rect 4521 9199 4527 9225
rect 5497 9199 5503 9225
rect 5529 9199 5535 9225
rect 6673 9199 6679 9225
rect 6705 9199 6711 9225
rect 7233 9199 7239 9225
rect 7265 9199 7271 9225
rect 8129 9199 8135 9225
rect 8161 9199 8167 9225
rect 9137 9199 9143 9225
rect 9169 9199 9175 9225
rect 10033 9199 10039 9225
rect 10065 9199 10071 9225
rect 10313 9199 10319 9225
rect 10345 9199 10351 9225
rect 11489 9199 11495 9225
rect 11521 9199 11527 9225
rect 12833 9199 12839 9225
rect 12865 9199 12871 9225
rect 13393 9199 13399 9225
rect 13425 9199 13431 9225
rect 13505 9199 13511 9225
rect 13537 9199 13543 9225
rect 14569 9199 14575 9225
rect 14601 9199 14607 9225
rect 15465 9199 15471 9225
rect 15497 9199 15503 9225
rect 17089 9199 17095 9225
rect 17121 9199 17127 9225
rect 17985 9199 17991 9225
rect 18017 9199 18023 9225
rect 18545 9199 18551 9225
rect 18577 9199 18583 9225
rect 19217 9199 19223 9225
rect 19249 9199 19255 9225
rect 21401 9199 21407 9225
rect 21433 9199 21439 9225
rect 22577 9199 22583 9225
rect 22609 9199 22615 9225
rect 22913 9199 22919 9225
rect 22945 9199 22951 9225
rect 23753 9199 23759 9225
rect 23785 9199 23791 9225
rect 672 9029 24304 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 24304 9029
rect 672 8986 24304 9003
rect 1353 8807 1359 8833
rect 1385 8807 1391 8833
rect 2473 8807 2479 8833
rect 2505 8807 2511 8833
rect 3817 8807 3823 8833
rect 3849 8807 3855 8833
rect 4377 8807 4383 8833
rect 4409 8807 4415 8833
rect 4489 8807 4495 8833
rect 4521 8807 4527 8833
rect 5273 8807 5279 8833
rect 5305 8807 5311 8833
rect 6449 8807 6455 8833
rect 6481 8807 6487 8833
rect 7177 8807 7183 8833
rect 7209 8807 7215 8833
rect 8073 8807 8079 8833
rect 8105 8807 8111 8833
rect 8633 8807 8639 8833
rect 8665 8807 8671 8833
rect 9529 8807 9535 8833
rect 9561 8807 9567 8833
rect 11097 8807 11103 8833
rect 11129 8807 11135 8833
rect 11713 8807 11719 8833
rect 11745 8807 11751 8833
rect 12273 8807 12279 8833
rect 12305 8807 12311 8833
rect 13393 8807 13399 8833
rect 13425 8807 13431 8833
rect 14793 8807 14799 8833
rect 14825 8807 14831 8833
rect 15353 8807 15359 8833
rect 15385 8807 15391 8833
rect 15465 8807 15471 8833
rect 15497 8807 15503 8833
rect 16529 8807 16535 8833
rect 16561 8807 16567 8833
rect 17145 8807 17151 8833
rect 17177 8807 17183 8833
rect 19049 8807 19055 8833
rect 19081 8807 19087 8833
rect 19217 8807 19223 8833
rect 19249 8807 19255 8833
rect 19441 8807 19447 8833
rect 19473 8807 19479 8833
rect 22857 8807 22863 8833
rect 22889 8807 22895 8833
rect 23753 8807 23759 8833
rect 23785 8807 23791 8833
rect 2473 8751 2479 8777
rect 2505 8751 2511 8777
rect 6449 8751 6455 8777
rect 6481 8751 6487 8777
rect 8073 8751 8079 8777
rect 8105 8751 8111 8777
rect 9529 8751 9535 8777
rect 9561 8751 9567 8777
rect 11769 8751 11775 8777
rect 11801 8751 11807 8777
rect 13393 8751 13399 8777
rect 13425 8751 13431 8777
rect 17201 8751 17207 8777
rect 17233 8751 17239 8777
rect 22857 8751 22863 8777
rect 22889 8751 22895 8777
rect 672 8637 24304 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 24304 8637
rect 672 8594 24304 8611
rect 6617 8471 6623 8497
rect 6649 8471 6655 8497
rect 8073 8471 8079 8497
rect 8105 8471 8111 8497
rect 11489 8471 11495 8497
rect 11521 8471 11527 8497
rect 14009 8471 14015 8497
rect 14041 8471 14047 8497
rect 15353 8471 15359 8497
rect 15385 8471 15391 8497
rect 19217 8471 19223 8497
rect 19249 8471 19255 8497
rect 22857 8471 22863 8497
rect 22889 8471 22895 8497
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 2417 8415 2423 8441
rect 2449 8415 2455 8441
rect 2529 8415 2535 8441
rect 2561 8415 2567 8441
rect 3593 8415 3599 8441
rect 3625 8415 3631 8441
rect 3761 8415 3767 8441
rect 3793 8415 3799 8441
rect 4489 8415 4495 8441
rect 4521 8415 4527 8441
rect 5441 8415 5447 8441
rect 5473 8415 5479 8441
rect 6617 8415 6623 8441
rect 6649 8415 6655 8441
rect 7177 8415 7183 8441
rect 7209 8415 7215 8441
rect 8073 8415 8079 8441
rect 8105 8415 8111 8441
rect 9137 8415 9143 8441
rect 9169 8415 9175 8441
rect 9417 8415 9423 8441
rect 9449 8415 9455 8441
rect 9529 8415 9535 8441
rect 9561 8415 9567 8441
rect 10313 8415 10319 8441
rect 10345 8415 10351 8441
rect 11489 8415 11495 8441
rect 11521 8415 11527 8441
rect 13113 8415 13119 8441
rect 13145 8415 13151 8441
rect 14009 8415 14015 8441
rect 14041 8415 14047 8441
rect 14569 8415 14575 8441
rect 14601 8415 14607 8441
rect 15353 8415 15359 8441
rect 15385 8415 15391 8441
rect 17089 8415 17095 8441
rect 17121 8415 17127 8441
rect 17257 8415 17263 8441
rect 17289 8415 17295 8441
rect 17481 8415 17487 8441
rect 17513 8415 17519 8441
rect 18545 8415 18551 8441
rect 18577 8415 18583 8441
rect 19217 8415 19223 8441
rect 19249 8415 19255 8441
rect 22857 8415 22863 8441
rect 22889 8415 22895 8441
rect 23753 8415 23759 8441
rect 23785 8415 23791 8441
rect 672 8245 24304 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 24304 8245
rect 672 8202 24304 8219
rect 1353 8023 1359 8049
rect 1385 8023 1391 8049
rect 2473 8023 2479 8049
rect 2505 8023 2511 8049
rect 3817 8023 3823 8049
rect 3849 8023 3855 8049
rect 4993 8023 4999 8049
rect 5025 8023 5031 8049
rect 5273 8023 5279 8049
rect 5305 8023 5311 8049
rect 6449 8023 6455 8049
rect 6481 8023 6487 8049
rect 7233 8023 7239 8049
rect 7265 8023 7271 8049
rect 8129 8023 8135 8049
rect 8161 8023 8167 8049
rect 8689 8023 8695 8049
rect 8721 8023 8727 8049
rect 9417 8023 9423 8049
rect 9449 8023 9455 8049
rect 11097 8023 11103 8049
rect 11129 8023 11135 8049
rect 11377 8023 11383 8049
rect 11409 8023 11415 8049
rect 11489 8023 11495 8049
rect 11521 8023 11527 8049
rect 12553 8023 12559 8049
rect 12585 8023 12591 8049
rect 13449 8023 13455 8049
rect 13481 8023 13487 8049
rect 14793 8023 14799 8049
rect 14825 8023 14831 8049
rect 15353 8023 15359 8049
rect 15385 8023 15391 8049
rect 15465 8023 15471 8049
rect 15497 8023 15503 8049
rect 16529 8023 16535 8049
rect 16561 8023 16567 8049
rect 17425 8023 17431 8049
rect 17457 8023 17463 8049
rect 19049 8023 19055 8049
rect 19081 8023 19087 8049
rect 19217 8023 19223 8049
rect 19249 8023 19255 8049
rect 19441 8023 19447 8049
rect 19473 8023 19479 8049
rect 20225 8023 20231 8049
rect 20257 8023 20263 8049
rect 21009 8023 21015 8049
rect 21041 8023 21047 8049
rect 22913 8023 22919 8049
rect 22945 8023 22951 8049
rect 24033 8023 24039 8049
rect 24065 8023 24071 8049
rect 2473 7967 2479 7993
rect 2505 7967 2511 7993
rect 4993 7967 4999 7993
rect 5025 7967 5031 7993
rect 6449 7967 6455 7993
rect 6481 7967 6487 7993
rect 8129 7967 8135 7993
rect 8161 7967 8167 7993
rect 9417 7967 9423 7993
rect 9449 7967 9455 7993
rect 13449 7967 13455 7993
rect 13481 7967 13487 7993
rect 17425 7967 17431 7993
rect 17457 7967 17463 7993
rect 21177 7967 21183 7993
rect 21209 7967 21215 7993
rect 22913 7967 22919 7993
rect 22945 7967 22951 7993
rect 672 7853 24304 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 24304 7853
rect 672 7810 24304 7827
rect 4489 7687 4495 7713
rect 4521 7687 4527 7713
rect 5833 7687 5839 7713
rect 5865 7687 5871 7713
rect 8129 7687 8135 7713
rect 8161 7687 8167 7713
rect 10033 7687 10039 7713
rect 10065 7687 10071 7713
rect 11489 7687 11495 7713
rect 11521 7687 11527 7713
rect 14009 7687 14015 7713
rect 14041 7687 14047 7713
rect 15465 7687 15471 7713
rect 15497 7687 15503 7713
rect 22857 7687 22863 7713
rect 22889 7687 22895 7713
rect 2137 7631 2143 7657
rect 2169 7631 2175 7657
rect 2417 7631 2423 7657
rect 2449 7631 2455 7657
rect 2529 7631 2535 7657
rect 2561 7631 2567 7657
rect 3593 7631 3599 7657
rect 3625 7631 3631 7657
rect 4489 7631 4495 7657
rect 4521 7631 4527 7657
rect 5161 7631 5167 7657
rect 5193 7631 5199 7657
rect 5833 7631 5839 7657
rect 5865 7631 5871 7657
rect 7233 7631 7239 7657
rect 7265 7631 7271 7657
rect 8129 7631 8135 7657
rect 8161 7631 8167 7657
rect 9137 7631 9143 7657
rect 9169 7631 9175 7657
rect 10033 7631 10039 7657
rect 10065 7631 10071 7657
rect 10313 7631 10319 7657
rect 10345 7631 10351 7657
rect 11489 7631 11495 7657
rect 11521 7631 11527 7657
rect 13113 7631 13119 7657
rect 13145 7631 13151 7657
rect 14009 7631 14015 7657
rect 14041 7631 14047 7657
rect 14569 7631 14575 7657
rect 14601 7631 14607 7657
rect 15465 7631 15471 7657
rect 15497 7631 15503 7657
rect 17089 7631 17095 7657
rect 17121 7631 17127 7657
rect 17369 7631 17375 7657
rect 17401 7631 17407 7657
rect 17481 7631 17487 7657
rect 17513 7631 17519 7657
rect 18545 7631 18551 7657
rect 18577 7631 18583 7657
rect 18713 7631 18719 7657
rect 18745 7631 18751 7657
rect 18937 7631 18943 7657
rect 18969 7631 18975 7657
rect 20785 7631 20791 7657
rect 20817 7631 20823 7657
rect 21233 7631 21239 7657
rect 21265 7631 21271 7657
rect 21457 7631 21463 7657
rect 21489 7631 21495 7657
rect 22857 7631 22863 7657
rect 22889 7631 22895 7657
rect 24033 7631 24039 7657
rect 24065 7631 24071 7657
rect 672 7461 24304 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 24304 7461
rect 672 7418 24304 7435
rect 1353 7239 1359 7265
rect 1385 7239 1391 7265
rect 2025 7239 2031 7265
rect 2057 7239 2063 7265
rect 3593 7239 3599 7265
rect 3625 7239 3631 7265
rect 4489 7239 4495 7265
rect 4521 7239 4527 7265
rect 4881 7239 4887 7265
rect 4913 7239 4919 7265
rect 5833 7239 5839 7265
rect 5865 7239 5871 7265
rect 7233 7239 7239 7265
rect 7265 7239 7271 7265
rect 8129 7239 8135 7265
rect 8161 7239 8167 7265
rect 8689 7239 8695 7265
rect 8721 7239 8727 7265
rect 9585 7239 9591 7265
rect 9617 7239 9623 7265
rect 11097 7239 11103 7265
rect 11129 7239 11135 7265
rect 11377 7239 11383 7265
rect 11409 7239 11415 7265
rect 11489 7239 11495 7265
rect 11521 7239 11527 7265
rect 12553 7239 12559 7265
rect 12585 7239 12591 7265
rect 13449 7239 13455 7265
rect 13481 7239 13487 7265
rect 14793 7239 14799 7265
rect 14825 7239 14831 7265
rect 15353 7239 15359 7265
rect 15385 7239 15391 7265
rect 15465 7239 15471 7265
rect 15497 7239 15503 7265
rect 16529 7239 16535 7265
rect 16561 7239 16567 7265
rect 17425 7239 17431 7265
rect 17457 7239 17463 7265
rect 18769 7239 18775 7265
rect 18801 7239 18807 7265
rect 19217 7239 19223 7265
rect 19249 7239 19255 7265
rect 19441 7239 19447 7265
rect 19473 7239 19479 7265
rect 20225 7239 20231 7265
rect 20257 7239 20263 7265
rect 21009 7239 21015 7265
rect 21041 7239 21047 7265
rect 22913 7239 22919 7265
rect 22945 7239 22951 7265
rect 23809 7239 23815 7265
rect 23841 7239 23847 7265
rect 2249 7183 2255 7209
rect 2281 7183 2287 7209
rect 4489 7183 4495 7209
rect 4521 7183 4527 7209
rect 5833 7183 5839 7209
rect 5865 7183 5871 7209
rect 8129 7183 8135 7209
rect 8161 7183 8167 7209
rect 9585 7183 9591 7209
rect 9617 7183 9623 7209
rect 13449 7183 13455 7209
rect 13481 7183 13487 7209
rect 17425 7183 17431 7209
rect 17457 7183 17463 7209
rect 21177 7183 21183 7209
rect 21209 7183 21215 7209
rect 22913 7183 22919 7209
rect 22945 7183 22951 7209
rect 672 7069 24304 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 24304 7069
rect 672 7026 24304 7043
rect 2865 6903 2871 6929
rect 2897 6903 2903 6929
rect 4489 6903 4495 6929
rect 4521 6903 4527 6929
rect 5833 6903 5839 6929
rect 5865 6903 5871 6929
rect 8073 6903 8079 6929
rect 8105 6903 8111 6929
rect 10873 6903 10879 6929
rect 10905 6903 10911 6929
rect 12441 6903 12447 6929
rect 12473 6903 12479 6929
rect 14009 6903 14015 6929
rect 14041 6903 14047 6929
rect 15353 6903 15359 6929
rect 15385 6903 15391 6929
rect 22857 6903 22863 6929
rect 22889 6903 22895 6929
rect 1913 6847 1919 6873
rect 1945 6847 1951 6873
rect 2865 6847 2871 6873
rect 2897 6847 2903 6873
rect 3593 6847 3599 6873
rect 3625 6847 3631 6873
rect 4489 6847 4495 6873
rect 4521 6847 4527 6873
rect 4881 6847 4887 6873
rect 4913 6847 4919 6873
rect 5833 6847 5839 6873
rect 5865 6847 5871 6873
rect 7177 6847 7183 6873
rect 7209 6847 7215 6873
rect 8073 6847 8079 6873
rect 8105 6847 8111 6873
rect 9809 6847 9815 6873
rect 9841 6847 9847 6873
rect 10873 6847 10879 6873
rect 10905 6847 10911 6873
rect 11545 6847 11551 6873
rect 11577 6847 11583 6873
rect 12441 6847 12447 6873
rect 12473 6847 12479 6873
rect 13113 6847 13119 6873
rect 13145 6847 13151 6873
rect 14009 6847 14015 6873
rect 14041 6847 14047 6873
rect 14569 6847 14575 6873
rect 14601 6847 14607 6873
rect 15353 6847 15359 6873
rect 15385 6847 15391 6873
rect 17089 6847 17095 6873
rect 17121 6847 17127 6873
rect 17257 6847 17263 6873
rect 17289 6847 17295 6873
rect 17481 6847 17487 6873
rect 17513 6847 17519 6873
rect 18265 6847 18271 6873
rect 18297 6847 18303 6873
rect 18713 6847 18719 6873
rect 18745 6847 18751 6873
rect 18937 6847 18943 6873
rect 18969 6847 18975 6873
rect 22857 6847 22863 6873
rect 22889 6847 22895 6873
rect 23753 6847 23759 6873
rect 23785 6847 23791 6873
rect 672 6677 24304 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 24304 6677
rect 672 6634 24304 6651
rect 1577 6455 1583 6481
rect 1609 6455 1615 6481
rect 2473 6455 2479 6481
rect 2505 6455 2511 6481
rect 4153 6455 4159 6481
rect 4185 6455 4191 6481
rect 4993 6455 4999 6481
rect 5025 6455 5031 6481
rect 5273 6455 5279 6481
rect 5305 6455 5311 6481
rect 6449 6455 6455 6481
rect 6481 6455 6487 6481
rect 7793 6455 7799 6481
rect 7825 6455 7831 6481
rect 8969 6455 8975 6481
rect 9001 6455 9007 6481
rect 9529 6455 9535 6481
rect 9561 6455 9567 6481
rect 10425 6455 10431 6481
rect 10457 6455 10463 6481
rect 12049 6455 12055 6481
rect 12081 6455 12087 6481
rect 12945 6455 12951 6481
rect 12977 6455 12983 6481
rect 13393 6455 13399 6481
rect 13425 6455 13431 6481
rect 14233 6455 14239 6481
rect 14265 6455 14271 6481
rect 14793 6455 14799 6481
rect 14825 6455 14831 6481
rect 15353 6455 15359 6481
rect 15385 6455 15391 6481
rect 15465 6455 15471 6481
rect 15497 6455 15503 6481
rect 16529 6455 16535 6481
rect 16561 6455 16567 6481
rect 17201 6455 17207 6481
rect 17233 6455 17239 6481
rect 18769 6455 18775 6481
rect 18801 6455 18807 6481
rect 19217 6455 19223 6481
rect 19249 6455 19255 6481
rect 19441 6455 19447 6481
rect 19473 6455 19479 6481
rect 20225 6455 20231 6481
rect 20257 6455 20263 6481
rect 20673 6455 20679 6481
rect 20705 6455 20711 6481
rect 21009 6455 21015 6481
rect 21041 6455 21047 6481
rect 22857 6455 22863 6481
rect 22889 6455 22895 6481
rect 23809 6455 23815 6481
rect 23841 6455 23847 6481
rect 2473 6399 2479 6425
rect 2505 6399 2511 6425
rect 4041 6399 4047 6425
rect 4073 6399 4079 6425
rect 5273 6399 5279 6425
rect 5305 6399 5311 6425
rect 7793 6399 7799 6425
rect 7825 6399 7831 6425
rect 10425 6399 10431 6425
rect 10457 6399 10463 6425
rect 12945 6399 12951 6425
rect 12977 6399 12983 6425
rect 14233 6399 14239 6425
rect 14265 6399 14271 6425
rect 17201 6399 17207 6425
rect 17233 6399 17239 6425
rect 22857 6399 22863 6425
rect 22889 6399 22895 6425
rect 672 6285 24304 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 24304 6285
rect 672 6242 24304 6259
rect 2081 6119 2087 6145
rect 2113 6119 2119 6145
rect 5833 6119 5839 6145
rect 5865 6119 5871 6145
rect 7513 6119 7519 6145
rect 7545 6119 7551 6145
rect 10873 6119 10879 6145
rect 10905 6119 10911 6145
rect 12441 6119 12447 6145
rect 12473 6119 12479 6145
rect 14009 6119 14015 6145
rect 14041 6119 14047 6145
rect 15353 6119 15359 6145
rect 15385 6119 15391 6145
rect 17761 6119 17767 6145
rect 17793 6119 17799 6145
rect 1185 6063 1191 6089
rect 1217 6063 1223 6089
rect 2081 6063 2087 6089
rect 2113 6063 2119 6089
rect 2529 6063 2535 6089
rect 2561 6063 2567 6089
rect 2809 6063 2815 6089
rect 2841 6063 2847 6089
rect 3033 6063 3039 6089
rect 3065 6063 3071 6089
rect 5833 6063 5839 6089
rect 5865 6063 5871 6089
rect 7009 6063 7015 6089
rect 7041 6063 7047 6089
rect 7569 6063 7575 6089
rect 7601 6063 7607 6089
rect 8465 6063 8471 6089
rect 8497 6063 8503 6089
rect 9809 6063 9815 6089
rect 9841 6063 9847 6089
rect 10873 6063 10879 6089
rect 10905 6063 10911 6089
rect 11545 6063 11551 6089
rect 11577 6063 11583 6089
rect 12441 6063 12447 6089
rect 12473 6063 12479 6089
rect 13113 6063 13119 6089
rect 13145 6063 13151 6089
rect 14009 6063 14015 6089
rect 14041 6063 14047 6089
rect 14569 6063 14575 6089
rect 14601 6063 14607 6089
rect 15353 6063 15359 6089
rect 15385 6063 15391 6089
rect 16809 6063 16815 6089
rect 16841 6063 16847 6089
rect 17761 6063 17767 6089
rect 17793 6063 17799 6089
rect 18265 6063 18271 6089
rect 18297 6063 18303 6089
rect 18825 6063 18831 6089
rect 18857 6063 18863 6089
rect 18937 6063 18943 6089
rect 18969 6063 18975 6089
rect 672 5893 24304 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 24304 5893
rect 672 5850 24304 5867
rect 1185 5671 1191 5697
rect 1217 5671 1223 5697
rect 2081 5671 2087 5697
rect 2113 5671 2119 5697
rect 2865 5671 2871 5697
rect 2897 5671 2903 5697
rect 3313 5671 3319 5697
rect 3345 5671 3351 5697
rect 3537 5671 3543 5697
rect 3569 5671 3575 5697
rect 5553 5671 5559 5697
rect 5585 5671 5591 5697
rect 6449 5671 6455 5697
rect 6481 5671 6487 5697
rect 7793 5671 7799 5697
rect 7825 5671 7831 5697
rect 8969 5671 8975 5697
rect 9001 5671 9007 5697
rect 9529 5671 9535 5697
rect 9561 5671 9567 5697
rect 10425 5671 10431 5697
rect 10457 5671 10463 5697
rect 12049 5671 12055 5697
rect 12081 5671 12087 5697
rect 12889 5671 12895 5697
rect 12921 5671 12927 5697
rect 13393 5671 13399 5697
rect 13425 5671 13431 5697
rect 14009 5671 14015 5697
rect 14041 5671 14047 5697
rect 14793 5671 14799 5697
rect 14825 5671 14831 5697
rect 15913 5671 15919 5697
rect 15945 5671 15951 5697
rect 16529 5671 16535 5697
rect 16561 5671 16567 5697
rect 17425 5671 17431 5697
rect 17457 5671 17463 5697
rect 19049 5671 19055 5697
rect 19081 5671 19087 5697
rect 19217 5671 19223 5697
rect 19249 5671 19255 5697
rect 19441 5671 19447 5697
rect 19473 5671 19479 5697
rect 2081 5615 2087 5641
rect 2113 5615 2119 5641
rect 6449 5615 6455 5641
rect 6481 5615 6487 5641
rect 7793 5615 7799 5641
rect 7825 5615 7831 5641
rect 10425 5615 10431 5641
rect 10457 5615 10463 5641
rect 12889 5615 12895 5641
rect 12921 5615 12927 5641
rect 14177 5615 14183 5641
rect 14209 5615 14215 5641
rect 15913 5615 15919 5641
rect 15945 5615 15951 5641
rect 17425 5615 17431 5641
rect 17457 5615 17463 5641
rect 672 5501 24304 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 24304 5501
rect 672 5458 24304 5475
rect 2081 5335 2087 5361
rect 2113 5335 2119 5361
rect 12441 5335 12447 5361
rect 12473 5335 12479 5361
rect 14009 5335 14015 5361
rect 14041 5335 14047 5361
rect 15465 5335 15471 5361
rect 15497 5335 15503 5361
rect 17761 5335 17767 5361
rect 17793 5335 17799 5361
rect 1185 5279 1191 5305
rect 1217 5279 1223 5305
rect 2081 5279 2087 5305
rect 2113 5279 2119 5305
rect 2529 5279 2535 5305
rect 2561 5279 2567 5305
rect 2809 5279 2815 5305
rect 2841 5279 2847 5305
rect 3033 5279 3039 5305
rect 3065 5279 3071 5305
rect 6113 5279 6119 5305
rect 6145 5279 6151 5305
rect 6393 5279 6399 5305
rect 6425 5279 6431 5305
rect 6505 5279 6511 5305
rect 6537 5279 6543 5305
rect 7513 5279 7519 5305
rect 7545 5279 7551 5305
rect 7793 5279 7799 5305
rect 7825 5279 7831 5305
rect 7961 5279 7967 5305
rect 7993 5279 7999 5305
rect 9809 5279 9815 5305
rect 9841 5279 9847 5305
rect 10369 5279 10375 5305
rect 10401 5279 10407 5305
rect 10481 5279 10487 5305
rect 10513 5279 10519 5305
rect 11545 5279 11551 5305
rect 11577 5279 11583 5305
rect 12441 5279 12447 5305
rect 12473 5279 12479 5305
rect 13113 5279 13119 5305
rect 13145 5279 13151 5305
rect 14009 5279 14015 5305
rect 14041 5279 14047 5305
rect 14569 5279 14575 5305
rect 14601 5279 14607 5305
rect 15465 5279 15471 5305
rect 15497 5279 15503 5305
rect 16809 5279 16815 5305
rect 16841 5279 16847 5305
rect 17761 5279 17767 5305
rect 17793 5279 17799 5305
rect 18545 5279 18551 5305
rect 18577 5279 18583 5305
rect 18713 5279 18719 5305
rect 18745 5279 18751 5305
rect 18937 5279 18943 5305
rect 18969 5279 18975 5305
rect 672 5109 24304 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 24304 5109
rect 672 5066 24304 5083
rect 1185 4887 1191 4913
rect 1217 4887 1223 4913
rect 2025 4887 2031 4913
rect 2057 4887 2063 4913
rect 2865 4887 2871 4913
rect 2897 4887 2903 4913
rect 3313 4887 3319 4913
rect 3345 4887 3351 4913
rect 3537 4887 3543 4913
rect 3569 4887 3575 4913
rect 8073 4887 8079 4913
rect 8105 4887 8111 4913
rect 8241 4887 8247 4913
rect 8273 4887 8279 4913
rect 8465 4887 8471 4913
rect 8497 4887 8503 4913
rect 9529 4887 9535 4913
rect 9561 4887 9567 4913
rect 10425 4887 10431 4913
rect 10457 4887 10463 4913
rect 12049 4887 12055 4913
rect 12081 4887 12087 4913
rect 12889 4887 12895 4913
rect 12921 4887 12927 4913
rect 13393 4887 13399 4913
rect 13425 4887 13431 4913
rect 14233 4887 14239 4913
rect 14265 4887 14271 4913
rect 14793 4887 14799 4913
rect 14825 4887 14831 4913
rect 15913 4887 15919 4913
rect 15945 4887 15951 4913
rect 16529 4887 16535 4913
rect 16561 4887 16567 4913
rect 17425 4887 17431 4913
rect 17457 4887 17463 4913
rect 2025 4831 2031 4857
rect 2057 4831 2063 4857
rect 10425 4831 10431 4857
rect 10457 4831 10463 4857
rect 12889 4831 12895 4857
rect 12921 4831 12927 4857
rect 14233 4831 14239 4857
rect 14265 4831 14271 4857
rect 15913 4831 15919 4857
rect 15945 4831 15951 4857
rect 17425 4831 17431 4857
rect 17457 4831 17463 4857
rect 672 4717 24304 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 24304 4717
rect 672 4674 24304 4691
rect 2025 4551 2031 4577
rect 2057 4551 2063 4577
rect 3313 4551 3319 4577
rect 3345 4551 3351 4577
rect 10873 4551 10879 4577
rect 10905 4551 10911 4577
rect 12385 4551 12391 4577
rect 12417 4551 12423 4577
rect 13953 4551 13959 4577
rect 13985 4551 13991 4577
rect 15465 4551 15471 4577
rect 15497 4551 15503 4577
rect 1185 4495 1191 4521
rect 1217 4495 1223 4521
rect 2025 4495 2031 4521
rect 2057 4495 2063 4521
rect 2529 4495 2535 4521
rect 2561 4495 2567 4521
rect 3313 4495 3319 4521
rect 3345 4495 3351 4521
rect 6337 4495 6343 4521
rect 6369 4495 6375 4521
rect 6505 4495 6511 4521
rect 6537 4495 6543 4521
rect 7009 4495 7015 4521
rect 7041 4495 7047 4521
rect 7513 4495 7519 4521
rect 7545 4495 7551 4521
rect 7737 4495 7743 4521
rect 7769 4495 7775 4521
rect 7961 4495 7967 4521
rect 7993 4495 7999 4521
rect 10033 4495 10039 4521
rect 10065 4495 10071 4521
rect 10873 4495 10879 4521
rect 10905 4495 10911 4521
rect 11545 4495 11551 4521
rect 11577 4495 11583 4521
rect 12385 4495 12391 4521
rect 12417 4495 12423 4521
rect 13113 4495 13119 4521
rect 13145 4495 13151 4521
rect 13953 4495 13959 4521
rect 13985 4495 13991 4521
rect 14569 4495 14575 4521
rect 14601 4495 14607 4521
rect 15465 4495 15471 4521
rect 15497 4495 15503 4521
rect 17089 4495 17095 4521
rect 17121 4495 17127 4521
rect 17369 4495 17375 4521
rect 17401 4495 17407 4521
rect 17481 4495 17487 4521
rect 17513 4495 17519 4521
rect 672 4325 24304 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 24304 4325
rect 672 4282 24304 4299
rect 1017 4103 1023 4129
rect 1049 4103 1055 4129
rect 1857 4103 1863 4129
rect 1889 4103 1895 4129
rect 5777 4103 5783 4129
rect 5809 4103 5815 4129
rect 5889 4103 5895 4129
rect 5921 4103 5927 4129
rect 6449 4103 6455 4129
rect 6481 4103 6487 4129
rect 7793 4103 7799 4129
rect 7825 4103 7831 4129
rect 8241 4103 8247 4129
rect 8273 4103 8279 4129
rect 8465 4103 8471 4129
rect 8497 4103 8503 4129
rect 9529 4103 9535 4129
rect 9561 4103 9567 4129
rect 10369 4103 10375 4129
rect 10401 4103 10407 4129
rect 11769 4103 11775 4129
rect 11801 4103 11807 4129
rect 12945 4103 12951 4129
rect 12977 4103 12983 4129
rect 13225 4103 13231 4129
rect 13257 4103 13263 4129
rect 14177 4103 14183 4129
rect 14209 4103 14215 4129
rect 15073 4103 15079 4129
rect 15105 4103 15111 4129
rect 15913 4103 15919 4129
rect 15945 4103 15951 4129
rect 16249 4103 16255 4129
rect 16281 4103 16287 4129
rect 17201 4103 17207 4129
rect 17233 4103 17239 4129
rect 22913 4103 22919 4129
rect 22945 4103 22951 4129
rect 24033 4103 24039 4129
rect 24065 4103 24071 4129
rect 1857 4047 1863 4073
rect 1889 4047 1895 4073
rect 10369 4047 10375 4073
rect 10401 4047 10407 4073
rect 12945 4047 12951 4073
rect 12977 4047 12983 4073
rect 14177 4047 14183 4073
rect 14209 4047 14215 4073
rect 15913 4047 15919 4073
rect 15945 4047 15951 4073
rect 17201 4047 17207 4073
rect 17233 4047 17239 4073
rect 22913 4047 22919 4073
rect 22945 4047 22951 4073
rect 672 3933 24304 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 24304 3933
rect 672 3890 24304 3907
rect 1857 3767 1863 3793
rect 1889 3767 1895 3793
rect 5833 3767 5839 3793
rect 5865 3767 5871 3793
rect 10873 3767 10879 3793
rect 10905 3767 10911 3793
rect 12441 3767 12447 3793
rect 12473 3767 12479 3793
rect 13953 3767 13959 3793
rect 13985 3767 13991 3793
rect 15465 3767 15471 3793
rect 15497 3767 15503 3793
rect 1017 3711 1023 3737
rect 1049 3711 1055 3737
rect 1857 3711 1863 3737
rect 1889 3711 1895 3737
rect 5833 3711 5839 3737
rect 5865 3711 5871 3737
rect 7009 3711 7015 3737
rect 7041 3711 7047 3737
rect 7513 3711 7519 3737
rect 7545 3711 7551 3737
rect 7793 3711 7799 3737
rect 7825 3711 7831 3737
rect 7961 3711 7967 3737
rect 7993 3711 7999 3737
rect 9809 3711 9815 3737
rect 9841 3711 9847 3737
rect 10873 3711 10879 3737
rect 10905 3711 10911 3737
rect 11265 3711 11271 3737
rect 11297 3711 11303 3737
rect 12441 3711 12447 3737
rect 12473 3711 12479 3737
rect 12833 3711 12839 3737
rect 12865 3711 12871 3737
rect 13953 3711 13959 3737
rect 13985 3711 13991 3737
rect 14569 3711 14575 3737
rect 14601 3711 14607 3737
rect 15465 3711 15471 3737
rect 15497 3711 15503 3737
rect 16809 3711 16815 3737
rect 16841 3711 16847 3737
rect 17257 3711 17263 3737
rect 17289 3711 17295 3737
rect 17481 3711 17487 3737
rect 17513 3711 17519 3737
rect 672 3541 24304 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 24304 3541
rect 672 3498 24304 3515
rect 8073 3319 8079 3345
rect 8105 3319 8111 3345
rect 8241 3319 8247 3345
rect 8273 3319 8279 3345
rect 8465 3319 8471 3345
rect 8497 3319 8503 3345
rect 9529 3319 9535 3345
rect 9561 3319 9567 3345
rect 10425 3319 10431 3345
rect 10457 3319 10463 3345
rect 11769 3319 11775 3345
rect 11801 3319 11807 3345
rect 12889 3319 12895 3345
rect 12921 3319 12927 3345
rect 13393 3319 13399 3345
rect 13425 3319 13431 3345
rect 14121 3319 14127 3345
rect 14153 3319 14159 3345
rect 15073 3319 15079 3345
rect 15105 3319 15111 3345
rect 15577 3319 15583 3345
rect 15609 3319 15615 3345
rect 16249 3319 16255 3345
rect 16281 3319 16287 3345
rect 17201 3319 17207 3345
rect 17233 3319 17239 3345
rect 10425 3263 10431 3289
rect 10457 3263 10463 3289
rect 12889 3263 12895 3289
rect 12921 3263 12927 3289
rect 14121 3263 14127 3289
rect 14153 3263 14159 3289
rect 15745 3263 15751 3289
rect 15777 3263 15783 3289
rect 17201 3263 17207 3289
rect 17233 3263 17239 3289
rect 672 3149 24304 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 24304 3149
rect 672 3106 24304 3123
rect 1857 2983 1863 3009
rect 1889 2983 1895 3009
rect 5833 2983 5839 3009
rect 5865 2983 5871 3009
rect 8465 2983 8471 3009
rect 8497 2983 8503 3009
rect 10761 2983 10767 3009
rect 10793 2983 10799 3009
rect 12329 2983 12335 3009
rect 12361 2983 12367 3009
rect 14009 2983 14015 3009
rect 14041 2983 14047 3009
rect 15465 2983 15471 3009
rect 15497 2983 15503 3009
rect 905 2927 911 2953
rect 937 2927 943 2953
rect 1857 2927 1863 2953
rect 1889 2927 1895 2953
rect 5833 2927 5839 2953
rect 5865 2927 5871 2953
rect 7009 2927 7015 2953
rect 7041 2927 7047 2953
rect 7569 2927 7575 2953
rect 7601 2927 7607 2953
rect 8465 2927 8471 2953
rect 8497 2927 8503 2953
rect 10033 2927 10039 2953
rect 10065 2927 10071 2953
rect 10761 2927 10767 2953
rect 10793 2927 10799 2953
rect 11545 2927 11551 2953
rect 11577 2927 11583 2953
rect 12329 2927 12335 2953
rect 12361 2927 12367 2953
rect 13113 2927 13119 2953
rect 13145 2927 13151 2953
rect 14009 2927 14015 2953
rect 14041 2927 14047 2953
rect 14569 2927 14575 2953
rect 14601 2927 14607 2953
rect 15465 2927 15471 2953
rect 15497 2927 15503 2953
rect 672 2757 24304 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 24304 2757
rect 672 2714 24304 2731
rect 905 2535 911 2561
rect 937 2535 943 2561
rect 2081 2535 2087 2561
rect 2113 2535 2119 2561
rect 5273 2535 5279 2561
rect 5305 2535 5311 2561
rect 6225 2535 6231 2561
rect 6257 2535 6263 2561
rect 8073 2535 8079 2561
rect 8105 2535 8111 2561
rect 8969 2535 8975 2561
rect 9001 2535 9007 2561
rect 9249 2535 9255 2561
rect 9281 2535 9287 2561
rect 10425 2535 10431 2561
rect 10457 2535 10463 2561
rect 11769 2535 11775 2561
rect 11801 2535 11807 2561
rect 12889 2535 12895 2561
rect 12921 2535 12927 2561
rect 13169 2535 13175 2561
rect 13201 2535 13207 2561
rect 14009 2535 14015 2561
rect 14041 2535 14047 2561
rect 14793 2535 14799 2561
rect 14825 2535 14831 2561
rect 15353 2535 15359 2561
rect 15385 2535 15391 2561
rect 15465 2535 15471 2561
rect 15497 2535 15503 2561
rect 2081 2479 2087 2505
rect 2113 2479 2119 2505
rect 5273 2479 5279 2505
rect 5305 2479 5311 2505
rect 8969 2479 8975 2505
rect 9001 2479 9007 2505
rect 10425 2479 10431 2505
rect 10457 2479 10463 2505
rect 12889 2479 12895 2505
rect 12921 2479 12927 2505
rect 14121 2479 14127 2505
rect 14153 2479 14159 2505
rect 672 2365 24304 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 24304 2365
rect 672 2322 24304 2339
rect 3761 2199 3767 2225
rect 3793 2199 3799 2225
rect 10761 2199 10767 2225
rect 10793 2199 10799 2225
rect 12441 2199 12447 2225
rect 12473 2199 12479 2225
rect 14009 2199 14015 2225
rect 14041 2199 14047 2225
rect 15353 2199 15359 2225
rect 15385 2199 15391 2225
rect 2865 2143 2871 2169
rect 2897 2143 2903 2169
rect 3761 2143 3767 2169
rect 3793 2143 3799 2169
rect 7009 2143 7015 2169
rect 7041 2143 7047 2169
rect 7569 2143 7575 2169
rect 7601 2143 7607 2169
rect 7681 2143 7687 2169
rect 7713 2143 7719 2169
rect 9809 2143 9815 2169
rect 9841 2143 9847 2169
rect 10761 2143 10767 2169
rect 10793 2143 10799 2169
rect 11545 2143 11551 2169
rect 11577 2143 11583 2169
rect 12441 2143 12447 2169
rect 12473 2143 12479 2169
rect 13113 2143 13119 2169
rect 13145 2143 13151 2169
rect 14009 2143 14015 2169
rect 14041 2143 14047 2169
rect 14289 2143 14295 2169
rect 14321 2143 14327 2169
rect 15353 2143 15359 2169
rect 15385 2143 15391 2169
rect 672 1973 24304 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 24304 1973
rect 672 1930 24304 1947
rect 2865 1751 2871 1777
rect 2897 1751 2903 1777
rect 3817 1751 3823 1777
rect 3849 1751 3855 1777
rect 7009 1751 7015 1777
rect 7041 1751 7047 1777
rect 7569 1751 7575 1777
rect 7601 1751 7607 1777
rect 7681 1751 7687 1777
rect 7713 1751 7719 1777
rect 9417 1751 9423 1777
rect 9449 1751 9455 1777
rect 9585 1751 9591 1777
rect 9617 1751 9623 1777
rect 9809 1751 9815 1777
rect 9841 1751 9847 1777
rect 11097 1751 11103 1777
rect 11129 1751 11135 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 12945 1751 12951 1777
rect 12977 1751 12983 1777
rect 13841 1751 13847 1777
rect 13873 1751 13879 1777
rect 3817 1695 3823 1721
rect 3849 1695 3855 1721
rect 12273 1695 12279 1721
rect 12305 1695 12311 1721
rect 13841 1695 13847 1721
rect 13873 1695 13879 1721
rect 672 1581 24304 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 24304 1581
rect 672 1538 24304 1555
<< via1 >>
rect 2239 33307 2265 33333
rect 2291 33307 2317 33333
rect 2343 33307 2369 33333
rect 17599 33307 17625 33333
rect 17651 33307 17677 33333
rect 17703 33307 17729 33333
rect 9919 32915 9945 32941
rect 9971 32915 9997 32941
rect 10023 32915 10049 32941
rect 2239 32523 2265 32549
rect 2291 32523 2317 32549
rect 2343 32523 2369 32549
rect 17599 32523 17625 32549
rect 17651 32523 17677 32549
rect 17703 32523 17729 32549
rect 9919 32131 9945 32157
rect 9971 32131 9997 32157
rect 10023 32131 10049 32157
rect 2239 31739 2265 31765
rect 2291 31739 2317 31765
rect 2343 31739 2369 31765
rect 17599 31739 17625 31765
rect 17651 31739 17677 31765
rect 17703 31739 17729 31765
rect 9919 31347 9945 31373
rect 9971 31347 9997 31373
rect 10023 31347 10049 31373
rect 2239 30955 2265 30981
rect 2291 30955 2317 30981
rect 2343 30955 2369 30981
rect 17599 30955 17625 30981
rect 17651 30955 17677 30981
rect 17703 30955 17729 30981
rect 9919 30563 9945 30589
rect 9971 30563 9997 30589
rect 10023 30563 10049 30589
rect 2239 30171 2265 30197
rect 2291 30171 2317 30197
rect 2343 30171 2369 30197
rect 17599 30171 17625 30197
rect 17651 30171 17677 30197
rect 17703 30171 17729 30197
rect 9919 29779 9945 29805
rect 9971 29779 9997 29805
rect 10023 29779 10049 29805
rect 23311 29583 23337 29609
rect 23367 29583 23393 29609
rect 23591 29583 23617 29609
rect 2239 29387 2265 29413
rect 2291 29387 2317 29413
rect 2343 29387 2369 29413
rect 17599 29387 17625 29413
rect 17651 29387 17677 29413
rect 17703 29387 17729 29413
rect 3935 29191 3961 29217
rect 4383 29191 4409 29217
rect 4607 29191 4633 29217
rect 23031 29191 23057 29217
rect 23199 29191 23225 29217
rect 23703 29191 23729 29217
rect 23871 29191 23897 29217
rect 23311 29135 23337 29161
rect 23591 29135 23617 29161
rect 9919 28995 9945 29021
rect 9971 28995 9997 29021
rect 10023 28995 10049 29021
rect 4383 28855 4409 28881
rect 5839 28855 5865 28881
rect 22415 28855 22441 28881
rect 22695 28855 22721 28881
rect 23087 28855 23113 28881
rect 23255 28855 23281 28881
rect 23535 28855 23561 28881
rect 3599 28799 3625 28825
rect 4383 28799 4409 28825
rect 5055 28799 5081 28825
rect 5839 28799 5865 28825
rect 22583 28799 22609 28825
rect 23031 28799 23057 28825
rect 23647 28799 23673 28825
rect 23815 28799 23841 28825
rect 2239 28603 2265 28629
rect 2291 28603 2317 28629
rect 2343 28603 2369 28629
rect 17599 28603 17625 28629
rect 17651 28603 17677 28629
rect 17703 28603 17729 28629
rect 3935 28407 3961 28433
rect 4887 28407 4913 28433
rect 22135 28407 22161 28433
rect 23031 28407 23057 28433
rect 23591 28407 23617 28433
rect 23759 28407 23785 28433
rect 23871 28407 23897 28433
rect 4887 28351 4913 28377
rect 22191 28351 22217 28377
rect 22359 28351 22385 28377
rect 23143 28351 23169 28377
rect 23311 28351 23337 28377
rect 9919 28211 9945 28237
rect 9971 28211 9997 28237
rect 10023 28211 10049 28237
rect 5839 28071 5865 28097
rect 7519 28071 7545 28097
rect 22751 28071 22777 28097
rect 23031 28071 23057 28097
rect 23143 28071 23169 28097
rect 23311 28071 23337 28097
rect 23591 28071 23617 28097
rect 23871 28071 23897 28097
rect 1863 28015 1889 28041
rect 2311 28015 2337 28041
rect 2535 28015 2561 28041
rect 3599 28015 3625 28041
rect 3879 28015 3905 28041
rect 4047 28015 4073 28041
rect 5055 28015 5081 28041
rect 5839 28015 5865 28041
rect 6623 28015 6649 28041
rect 7519 28015 7545 28041
rect 21407 28015 21433 28041
rect 21519 28015 21545 28041
rect 21687 28015 21713 28041
rect 21967 28015 21993 28041
rect 22079 28015 22105 28041
rect 22247 28015 22273 28041
rect 22527 28015 22553 28041
rect 22639 28015 22665 28041
rect 23759 28015 23785 28041
rect 2239 27819 2265 27845
rect 2291 27819 2317 27845
rect 2343 27819 2369 27845
rect 17599 27819 17625 27845
rect 17651 27819 17677 27845
rect 17703 27819 17729 27845
rect 1359 27623 1385 27649
rect 2479 27623 2505 27649
rect 3319 27623 3345 27649
rect 3991 27623 4017 27649
rect 4775 27623 4801 27649
rect 5447 27623 5473 27649
rect 7127 27623 7153 27649
rect 8023 27623 8049 27649
rect 8415 27623 8441 27649
rect 8863 27623 8889 27649
rect 8975 27623 9001 27649
rect 11047 27623 11073 27649
rect 11383 27623 11409 27649
rect 11495 27623 11521 27649
rect 21127 27623 21153 27649
rect 21575 27623 21601 27649
rect 21631 27623 21657 27649
rect 21799 27623 21825 27649
rect 22415 27623 22441 27649
rect 2479 27567 2505 27593
rect 3991 27567 4017 27593
rect 5447 27567 5473 27593
rect 8023 27567 8049 27593
rect 20959 27567 20985 27593
rect 21239 27567 21265 27593
rect 22079 27567 22105 27593
rect 22191 27567 22217 27593
rect 22975 27567 23001 27593
rect 23087 27567 23113 27593
rect 23255 27567 23281 27593
rect 23535 27567 23561 27593
rect 23647 27567 23673 27593
rect 23815 27567 23841 27593
rect 9919 27427 9945 27453
rect 9971 27427 9997 27453
rect 10023 27427 10049 27453
rect 7519 27287 7545 27313
rect 10039 27287 10065 27313
rect 11495 27287 11521 27313
rect 21071 27287 21097 27313
rect 21631 27287 21657 27313
rect 1863 27231 1889 27257
rect 2423 27231 2449 27257
rect 2535 27231 2561 27257
rect 3319 27231 3345 27257
rect 3767 27231 3793 27257
rect 3991 27231 4017 27257
rect 5167 27231 5193 27257
rect 5447 27231 5473 27257
rect 5559 27231 5585 27257
rect 6623 27231 6649 27257
rect 7519 27231 7545 27257
rect 8863 27231 8889 27257
rect 10039 27231 10065 27257
rect 10599 27231 10625 27257
rect 11495 27231 11521 27257
rect 21183 27231 21209 27257
rect 21351 27231 21377 27257
rect 21743 27231 21769 27257
rect 21967 27231 21993 27257
rect 22191 27231 22217 27257
rect 22359 27231 22385 27257
rect 22527 27231 22553 27257
rect 22751 27231 22777 27257
rect 22919 27231 22945 27257
rect 23031 27231 23057 27257
rect 23311 27231 23337 27257
rect 23423 27231 23449 27257
rect 23647 27231 23673 27257
rect 2239 27035 2265 27061
rect 2291 27035 2317 27061
rect 2343 27035 2369 27061
rect 17599 27035 17625 27061
rect 17651 27035 17677 27061
rect 17703 27035 17729 27061
rect 1359 26839 1385 26865
rect 2479 26839 2505 26865
rect 3319 26839 3345 26865
rect 3487 26839 3513 26865
rect 3711 26839 3737 26865
rect 4775 26839 4801 26865
rect 5447 26839 5473 26865
rect 7127 26839 7153 26865
rect 8023 26839 8049 26865
rect 8583 26839 8609 26865
rect 8863 26839 8889 26865
rect 8975 26839 9001 26865
rect 11047 26839 11073 26865
rect 11719 26839 11745 26865
rect 19783 26839 19809 26865
rect 19951 26839 19977 26865
rect 20343 26839 20369 26865
rect 20511 26839 20537 26865
rect 20679 26839 20705 26865
rect 20959 26839 20985 26865
rect 21127 26839 21153 26865
rect 21239 26839 21265 26865
rect 21631 26839 21657 26865
rect 21799 26839 21825 26865
rect 22135 26839 22161 26865
rect 22247 26839 22273 26865
rect 22415 26839 22441 26865
rect 22751 26839 22777 26865
rect 22919 26839 22945 26865
rect 23087 26839 23113 26865
rect 23423 26839 23449 26865
rect 23647 26839 23673 26865
rect 2479 26783 2505 26809
rect 5447 26783 5473 26809
rect 8023 26783 8049 26809
rect 11775 26783 11801 26809
rect 20119 26783 20145 26809
rect 21519 26783 21545 26809
rect 23311 26783 23337 26809
rect 9919 26643 9945 26669
rect 9971 26643 9997 26669
rect 10023 26643 10049 26669
rect 4271 26503 4297 26529
rect 7519 26503 7545 26529
rect 10039 26503 10065 26529
rect 21015 26503 21041 26529
rect 21855 26503 21881 26529
rect 22695 26503 22721 26529
rect 22863 26503 22889 26529
rect 1863 26447 1889 26473
rect 2423 26447 2449 26473
rect 2535 26447 2561 26473
rect 3319 26447 3345 26473
rect 4215 26447 4241 26473
rect 5167 26447 5193 26473
rect 5335 26447 5361 26473
rect 5559 26447 5585 26473
rect 6343 26447 6369 26473
rect 7519 26447 7545 26473
rect 8919 26447 8945 26473
rect 10039 26447 10065 26473
rect 10599 26447 10625 26473
rect 10879 26447 10905 26473
rect 10991 26447 11017 26473
rect 21127 26447 21153 26473
rect 21295 26447 21321 26473
rect 21631 26447 21657 26473
rect 21743 26447 21769 26473
rect 22135 26447 22161 26473
rect 22303 26447 22329 26473
rect 22471 26447 22497 26473
rect 22975 26447 23001 26473
rect 23311 26447 23337 26473
rect 23423 26447 23449 26473
rect 23535 26447 23561 26473
rect 2239 26251 2265 26277
rect 2291 26251 2317 26277
rect 2343 26251 2369 26277
rect 17599 26251 17625 26277
rect 17651 26251 17677 26277
rect 17703 26251 17729 26277
rect 1359 26055 1385 26081
rect 2479 26055 2505 26081
rect 3319 26055 3345 26081
rect 4215 26055 4241 26081
rect 4775 26055 4801 26081
rect 4943 26055 4969 26081
rect 5167 26055 5193 26081
rect 7127 26055 7153 26081
rect 8023 26055 8049 26081
rect 8583 26055 8609 26081
rect 8863 26055 8889 26081
rect 8975 26055 9001 26081
rect 11103 26055 11129 26081
rect 11719 26055 11745 26081
rect 12559 26055 12585 26081
rect 13343 26055 13369 26081
rect 21071 26055 21097 26081
rect 21239 26055 21265 26081
rect 21519 26055 21545 26081
rect 21631 26055 21657 26081
rect 21799 26055 21825 26081
rect 22135 26055 22161 26081
rect 22247 26055 22273 26081
rect 22415 26055 22441 26081
rect 23311 26055 23337 26081
rect 23423 26055 23449 26081
rect 2479 25999 2505 26025
rect 4215 25999 4241 26025
rect 8023 25999 8049 26025
rect 11775 25999 11801 26025
rect 13343 25999 13369 26025
rect 20959 25999 20985 26025
rect 23535 25999 23561 26025
rect 9919 25859 9945 25885
rect 9971 25859 9997 25885
rect 10023 25859 10049 25885
rect 3039 25719 3065 25745
rect 4271 25719 4297 25745
rect 7631 25719 7657 25745
rect 10039 25719 10065 25745
rect 11495 25719 11521 25745
rect 21575 25719 21601 25745
rect 21855 25719 21881 25745
rect 22135 25719 22161 25745
rect 22695 25719 22721 25745
rect 22863 25719 22889 25745
rect 2143 25663 2169 25689
rect 3039 25663 3065 25689
rect 3319 25663 3345 25689
rect 4215 25663 4241 25689
rect 5111 25663 5137 25689
rect 5335 25663 5361 25689
rect 5559 25663 5585 25689
rect 6679 25663 6705 25689
rect 7631 25663 7657 25689
rect 9143 25663 9169 25689
rect 10039 25663 10065 25689
rect 10599 25663 10625 25689
rect 11495 25663 11521 25689
rect 13119 25663 13145 25689
rect 13343 25663 13369 25689
rect 13511 25663 13537 25689
rect 21743 25663 21769 25689
rect 22303 25663 22329 25689
rect 22471 25663 22497 25689
rect 22975 25663 23001 25689
rect 23311 25663 23337 25689
rect 23423 25663 23449 25689
rect 23535 25663 23561 25689
rect 2239 25467 2265 25493
rect 2291 25467 2317 25493
rect 2343 25467 2369 25493
rect 17599 25467 17625 25493
rect 17651 25467 17677 25493
rect 17703 25467 17729 25493
rect 1583 25271 1609 25297
rect 2479 25271 2505 25297
rect 3319 25271 3345 25297
rect 4215 25271 4241 25297
rect 4775 25271 4801 25297
rect 4943 25271 4969 25297
rect 5167 25271 5193 25297
rect 7127 25271 7153 25297
rect 8023 25271 8049 25297
rect 8415 25271 8441 25297
rect 8863 25271 8889 25297
rect 8975 25271 9001 25297
rect 11103 25271 11129 25297
rect 11719 25271 11745 25297
rect 12559 25271 12585 25297
rect 12727 25271 12753 25297
rect 12951 25271 12977 25297
rect 22135 25271 22161 25297
rect 22247 25271 22273 25297
rect 22359 25271 22385 25297
rect 23311 25271 23337 25297
rect 23423 25271 23449 25297
rect 23591 25271 23617 25297
rect 2479 25215 2505 25241
rect 4215 25215 4241 25241
rect 8023 25215 8049 25241
rect 11775 25215 11801 25241
rect 9919 25075 9945 25101
rect 9971 25075 9997 25101
rect 10023 25075 10049 25101
rect 4495 24935 4521 24961
rect 6175 24935 6201 24961
rect 7631 24935 7657 24961
rect 10039 24935 10065 24961
rect 11495 24935 11521 24961
rect 15247 24935 15273 24961
rect 22471 24935 22497 24961
rect 22583 24935 22609 24961
rect 22751 24935 22777 24961
rect 23031 24935 23057 24961
rect 23143 24935 23169 24961
rect 23311 24935 23337 24961
rect 1863 24879 1889 24905
rect 2423 24879 2449 24905
rect 2535 24879 2561 24905
rect 3375 24879 3401 24905
rect 4495 24879 4521 24905
rect 5055 24879 5081 24905
rect 6175 24879 6201 24905
rect 6679 24879 6705 24905
rect 7631 24879 7657 24905
rect 8919 24879 8945 24905
rect 10039 24879 10065 24905
rect 10319 24879 10345 24905
rect 11495 24879 11521 24905
rect 13119 24879 13145 24905
rect 13399 24879 13425 24905
rect 13511 24879 13537 24905
rect 14519 24879 14545 24905
rect 15135 24879 15161 24905
rect 23759 24879 23785 24905
rect 23927 24879 23953 24905
rect 24039 24879 24065 24905
rect 2239 24683 2265 24709
rect 2291 24683 2317 24709
rect 2343 24683 2369 24709
rect 17599 24683 17625 24709
rect 17651 24683 17677 24709
rect 17703 24683 17729 24709
rect 1359 24487 1385 24513
rect 2479 24487 2505 24513
rect 3823 24487 3849 24513
rect 4383 24487 4409 24513
rect 4495 24487 4521 24513
rect 5279 24487 5305 24513
rect 6455 24487 6481 24513
rect 7127 24487 7153 24513
rect 8023 24487 8049 24513
rect 8583 24487 8609 24513
rect 9479 24487 9505 24513
rect 10823 24487 10849 24513
rect 11383 24487 11409 24513
rect 11495 24487 11521 24513
rect 12559 24487 12585 24513
rect 13343 24487 13369 24513
rect 15079 24487 15105 24513
rect 15247 24487 15273 24513
rect 15471 24487 15497 24513
rect 23143 24487 23169 24513
rect 23311 24487 23337 24513
rect 23759 24487 23785 24513
rect 23871 24487 23897 24513
rect 2479 24431 2505 24457
rect 6455 24431 6481 24457
rect 8023 24431 8049 24457
rect 9479 24431 9505 24457
rect 13343 24431 13369 24457
rect 23479 24431 23505 24457
rect 24039 24431 24065 24457
rect 9919 24291 9945 24317
rect 9971 24291 9997 24317
rect 10023 24291 10049 24317
rect 3039 24151 3065 24177
rect 4495 24151 4521 24177
rect 6175 24151 6201 24177
rect 7631 24151 7657 24177
rect 10039 24151 10065 24177
rect 11495 24151 11521 24177
rect 15247 24151 15273 24177
rect 23927 24151 23953 24177
rect 1863 24095 1889 24121
rect 3039 24095 3065 24121
rect 3375 24095 3401 24121
rect 4495 24095 4521 24121
rect 5055 24095 5081 24121
rect 6175 24095 6201 24121
rect 6679 24095 6705 24121
rect 7631 24095 7657 24121
rect 9087 24095 9113 24121
rect 10039 24095 10065 24121
rect 10599 24095 10625 24121
rect 11495 24095 11521 24121
rect 13119 24095 13145 24121
rect 13343 24095 13369 24121
rect 13511 24095 13537 24121
rect 14519 24095 14545 24121
rect 15135 24095 15161 24121
rect 23759 24095 23785 24121
rect 24039 24095 24065 24121
rect 2239 23899 2265 23925
rect 2291 23899 2317 23925
rect 2343 23899 2369 23925
rect 17599 23899 17625 23925
rect 17651 23899 17677 23925
rect 17703 23899 17729 23925
rect 1359 23703 1385 23729
rect 2479 23703 2505 23729
rect 4103 23703 4129 23729
rect 4999 23703 5025 23729
rect 5559 23703 5585 23729
rect 6455 23703 6481 23729
rect 7127 23703 7153 23729
rect 8023 23703 8049 23729
rect 8583 23703 8609 23729
rect 9479 23703 9505 23729
rect 11103 23703 11129 23729
rect 11719 23703 11745 23729
rect 12279 23703 12305 23729
rect 13455 23703 13481 23729
rect 15079 23703 15105 23729
rect 15247 23703 15273 23729
rect 15471 23703 15497 23729
rect 2479 23647 2505 23673
rect 4999 23647 5025 23673
rect 6455 23647 6481 23673
rect 8023 23647 8049 23673
rect 9479 23647 9505 23673
rect 11775 23647 11801 23673
rect 13455 23647 13481 23673
rect 9919 23507 9945 23533
rect 9971 23507 9997 23533
rect 10023 23507 10049 23533
rect 3039 23367 3065 23393
rect 4495 23367 4521 23393
rect 6175 23367 6201 23393
rect 7519 23367 7545 23393
rect 13959 23367 13985 23393
rect 15303 23367 15329 23393
rect 1863 23311 1889 23337
rect 3039 23311 3065 23337
rect 3375 23311 3401 23337
rect 4495 23311 4521 23337
rect 5055 23311 5081 23337
rect 6175 23311 6201 23337
rect 6679 23311 6705 23337
rect 7519 23311 7545 23337
rect 9087 23311 9113 23337
rect 9311 23311 9337 23337
rect 9535 23311 9561 23337
rect 10319 23311 10345 23337
rect 10879 23311 10905 23337
rect 10991 23311 11017 23337
rect 12839 23311 12865 23337
rect 13959 23311 13985 23337
rect 14575 23311 14601 23337
rect 15303 23311 15329 23337
rect 23703 23311 23729 23337
rect 23871 23311 23897 23337
rect 23983 23311 24009 23337
rect 2239 23115 2265 23141
rect 2291 23115 2317 23141
rect 2343 23115 2369 23141
rect 17599 23115 17625 23141
rect 17651 23115 17677 23141
rect 17703 23115 17729 23141
rect 1359 22919 1385 22945
rect 2479 22919 2505 22945
rect 4103 22919 4129 22945
rect 4999 22919 5025 22945
rect 5279 22919 5305 22945
rect 6175 22919 6201 22945
rect 8135 22919 8161 22945
rect 9031 22919 9057 22945
rect 10823 22919 10849 22945
rect 11271 22919 11297 22945
rect 11495 22919 11521 22945
rect 12279 22919 12305 22945
rect 13455 22919 13481 22945
rect 14799 22919 14825 22945
rect 15303 22919 15329 22945
rect 15471 22919 15497 22945
rect 16255 22919 16281 22945
rect 16815 22919 16841 22945
rect 16927 22919 16953 22945
rect 23871 22919 23897 22945
rect 23983 22919 24009 22945
rect 2479 22863 2505 22889
rect 4999 22863 5025 22889
rect 6231 22863 6257 22889
rect 9031 22863 9057 22889
rect 13455 22863 13481 22889
rect 23199 22863 23225 22889
rect 23367 22863 23393 22889
rect 23479 22863 23505 22889
rect 23759 22863 23785 22889
rect 9919 22723 9945 22749
rect 9971 22723 9997 22749
rect 10023 22723 10049 22749
rect 2983 22583 3009 22609
rect 4495 22583 4521 22609
rect 7015 22583 7041 22609
rect 8247 22583 8273 22609
rect 11271 22583 11297 22609
rect 13959 22583 13985 22609
rect 15303 22583 15329 22609
rect 1863 22527 1889 22553
rect 2983 22527 3009 22553
rect 3375 22527 3401 22553
rect 4495 22527 4521 22553
rect 5839 22527 5865 22553
rect 7015 22527 7041 22553
rect 7575 22527 7601 22553
rect 8247 22527 8273 22553
rect 9087 22527 9113 22553
rect 9311 22527 9337 22553
rect 9535 22527 9561 22553
rect 10319 22527 10345 22553
rect 11271 22527 11297 22553
rect 12839 22527 12865 22553
rect 13959 22527 13985 22553
rect 14575 22527 14601 22553
rect 15303 22527 15329 22553
rect 16815 22527 16841 22553
rect 17263 22527 17289 22553
rect 17487 22527 17513 22553
rect 23759 22527 23785 22553
rect 23871 22527 23897 22553
rect 23983 22527 24009 22553
rect 2239 22331 2265 22357
rect 2291 22331 2317 22357
rect 2343 22331 2369 22357
rect 17599 22331 17625 22357
rect 17651 22331 17677 22357
rect 17703 22331 17729 22357
rect 1359 22135 1385 22161
rect 2479 22135 2505 22161
rect 4103 22135 4129 22161
rect 4999 22135 5025 22161
rect 5279 22135 5305 22161
rect 6231 22135 6257 22161
rect 8135 22135 8161 22161
rect 9031 22135 9057 22161
rect 10823 22135 10849 22161
rect 11271 22135 11297 22161
rect 11495 22135 11521 22161
rect 12279 22135 12305 22161
rect 13231 22135 13257 22161
rect 14799 22135 14825 22161
rect 15303 22135 15329 22161
rect 15471 22135 15497 22161
rect 16255 22135 16281 22161
rect 16759 22135 16785 22161
rect 16927 22135 16953 22161
rect 2479 22079 2505 22105
rect 4999 22079 5025 22105
rect 6231 22079 6257 22105
rect 9031 22079 9057 22105
rect 13231 22079 13257 22105
rect 9919 21939 9945 21965
rect 9971 21939 9997 21965
rect 10023 21939 10049 21965
rect 4383 21799 4409 21825
rect 8247 21799 8273 21825
rect 11271 21799 11297 21825
rect 15359 21799 15385 21825
rect 17991 21799 18017 21825
rect 19279 21799 19305 21825
rect 2143 21743 2169 21769
rect 2423 21743 2449 21769
rect 2535 21743 2561 21769
rect 3599 21743 3625 21769
rect 4383 21743 4409 21769
rect 5839 21743 5865 21769
rect 6399 21743 6425 21769
rect 6511 21743 6537 21769
rect 7295 21743 7321 21769
rect 8247 21743 8273 21769
rect 9087 21743 9113 21769
rect 9311 21743 9337 21769
rect 9535 21743 9561 21769
rect 10319 21743 10345 21769
rect 11271 21743 11297 21769
rect 12839 21743 12865 21769
rect 13399 21743 13425 21769
rect 13511 21743 13537 21769
rect 14575 21743 14601 21769
rect 15359 21743 15385 21769
rect 17095 21743 17121 21769
rect 17991 21743 18017 21769
rect 18551 21743 18577 21769
rect 19279 21743 19305 21769
rect 2239 21547 2265 21573
rect 2291 21547 2317 21573
rect 2343 21547 2369 21573
rect 17599 21547 17625 21573
rect 17651 21547 17677 21573
rect 17703 21547 17729 21573
rect 1583 21351 1609 21377
rect 2479 21351 2505 21377
rect 3823 21351 3849 21377
rect 4383 21351 4409 21377
rect 4495 21351 4521 21377
rect 5279 21351 5305 21377
rect 6399 21351 6425 21377
rect 8135 21351 8161 21377
rect 9031 21351 9057 21377
rect 10823 21351 10849 21377
rect 11271 21351 11297 21377
rect 11495 21351 11521 21377
rect 12279 21351 12305 21377
rect 13455 21351 13481 21377
rect 14799 21351 14825 21377
rect 15359 21351 15385 21377
rect 15471 21351 15497 21377
rect 16255 21351 16281 21377
rect 17431 21351 17457 21377
rect 19055 21351 19081 21377
rect 19279 21351 19305 21377
rect 19447 21351 19473 21377
rect 2479 21295 2505 21321
rect 6399 21295 6425 21321
rect 9031 21295 9057 21321
rect 13455 21295 13481 21321
rect 17431 21295 17457 21321
rect 9919 21155 9945 21181
rect 9971 21155 9997 21181
rect 10023 21155 10049 21181
rect 4383 21015 4409 21041
rect 7015 21015 7041 21041
rect 8247 21015 8273 21041
rect 9815 21015 9841 21041
rect 11271 21015 11297 21041
rect 14015 21015 14041 21041
rect 15359 21015 15385 21041
rect 17935 21015 17961 21041
rect 19447 21015 19473 21041
rect 2143 20959 2169 20985
rect 2423 20959 2449 20985
rect 2535 20959 2561 20985
rect 3599 20959 3625 20985
rect 4383 20959 4409 20985
rect 5839 20959 5865 20985
rect 7015 20959 7041 20985
rect 7295 20959 7321 20985
rect 8247 20959 8273 20985
rect 9143 20959 9169 20985
rect 9815 20959 9841 20985
rect 10319 20959 10345 20985
rect 11271 20959 11297 20985
rect 12951 20959 12977 20985
rect 14015 20959 14041 20985
rect 14575 20959 14601 20985
rect 15359 20959 15385 20985
rect 16815 20959 16841 20985
rect 17935 20959 17961 20985
rect 18551 20959 18577 20985
rect 19447 20959 19473 20985
rect 2239 20763 2265 20789
rect 2291 20763 2317 20789
rect 2343 20763 2369 20789
rect 17599 20763 17625 20789
rect 17651 20763 17677 20789
rect 17703 20763 17729 20789
rect 1583 20567 1609 20593
rect 2479 20567 2505 20593
rect 3823 20567 3849 20593
rect 4271 20567 4297 20593
rect 4495 20567 4521 20593
rect 5279 20567 5305 20593
rect 6455 20567 6481 20593
rect 8135 20567 8161 20593
rect 9031 20567 9057 20593
rect 10823 20567 10849 20593
rect 11271 20567 11297 20593
rect 11495 20567 11521 20593
rect 12279 20567 12305 20593
rect 13455 20567 13481 20593
rect 14911 20567 14937 20593
rect 15359 20567 15385 20593
rect 15471 20567 15497 20593
rect 16535 20567 16561 20593
rect 17431 20567 17457 20593
rect 19055 20567 19081 20593
rect 19951 20567 19977 20593
rect 20511 20567 20537 20593
rect 21239 20567 21265 20593
rect 2479 20511 2505 20537
rect 6455 20511 6481 20537
rect 9031 20511 9057 20537
rect 13455 20511 13481 20537
rect 17431 20511 17457 20537
rect 19951 20511 19977 20537
rect 21239 20511 21265 20537
rect 9919 20371 9945 20397
rect 9971 20371 9997 20397
rect 10023 20371 10049 20397
rect 4271 20231 4297 20257
rect 7015 20231 7041 20257
rect 8247 20231 8273 20257
rect 9815 20231 9841 20257
rect 11271 20231 11297 20257
rect 14015 20231 14041 20257
rect 15359 20231 15385 20257
rect 17991 20231 18017 20257
rect 19279 20231 19305 20257
rect 2143 20175 2169 20201
rect 2423 20175 2449 20201
rect 2535 20175 2561 20201
rect 3599 20175 3625 20201
rect 4215 20175 4241 20201
rect 5839 20175 5865 20201
rect 7015 20175 7041 20201
rect 7295 20175 7321 20201
rect 8247 20175 8273 20201
rect 9143 20175 9169 20201
rect 9815 20175 9841 20201
rect 10319 20175 10345 20201
rect 11271 20175 11297 20201
rect 12951 20175 12977 20201
rect 14015 20175 14041 20201
rect 14295 20175 14321 20201
rect 15359 20175 15385 20201
rect 16815 20175 16841 20201
rect 17991 20175 18017 20201
rect 18551 20175 18577 20201
rect 19279 20175 19305 20201
rect 20959 20175 20985 20201
rect 21239 20175 21265 20201
rect 21463 20175 21489 20201
rect 2239 19979 2265 20005
rect 2291 19979 2317 20005
rect 2343 19979 2369 20005
rect 17599 19979 17625 20005
rect 17651 19979 17677 20005
rect 17703 19979 17729 20005
rect 1583 19783 1609 19809
rect 2479 19783 2505 19809
rect 3823 19783 3849 19809
rect 4383 19783 4409 19809
rect 4551 19783 4577 19809
rect 5279 19783 5305 19809
rect 6455 19783 6481 19809
rect 8135 19783 8161 19809
rect 9031 19783 9057 19809
rect 10823 19783 10849 19809
rect 11271 19783 11297 19809
rect 11495 19783 11521 19809
rect 12279 19783 12305 19809
rect 13455 19783 13481 19809
rect 14799 19783 14825 19809
rect 15919 19783 15945 19809
rect 16255 19783 16281 19809
rect 17431 19783 17457 19809
rect 19055 19783 19081 19809
rect 19335 19783 19361 19809
rect 19447 19783 19473 19809
rect 20511 19783 20537 19809
rect 21183 19783 21209 19809
rect 23759 19783 23785 19809
rect 23871 19783 23897 19809
rect 2479 19727 2505 19753
rect 6455 19727 6481 19753
rect 9031 19727 9057 19753
rect 13455 19727 13481 19753
rect 15919 19727 15945 19753
rect 17431 19727 17457 19753
rect 21183 19727 21209 19753
rect 24039 19727 24065 19753
rect 9919 19587 9945 19613
rect 9971 19587 9997 19613
rect 10023 19587 10049 19613
rect 4439 19447 4465 19473
rect 7015 19447 7041 19473
rect 8247 19447 8273 19473
rect 9815 19447 9841 19473
rect 11271 19447 11297 19473
rect 14015 19447 14041 19473
rect 15471 19447 15497 19473
rect 17991 19447 18017 19473
rect 19335 19447 19361 19473
rect 21799 19447 21825 19473
rect 23255 19447 23281 19473
rect 2143 19391 2169 19417
rect 2423 19391 2449 19417
rect 2535 19391 2561 19417
rect 3599 19391 3625 19417
rect 4439 19391 4465 19417
rect 5839 19391 5865 19417
rect 7015 19391 7041 19417
rect 7295 19391 7321 19417
rect 8247 19391 8273 19417
rect 9143 19391 9169 19417
rect 9815 19391 9841 19417
rect 10319 19391 10345 19417
rect 11271 19391 11297 19417
rect 12951 19391 12977 19417
rect 14015 19391 14041 19417
rect 14295 19391 14321 19417
rect 15471 19391 15497 19417
rect 16871 19391 16897 19417
rect 17991 19391 18017 19417
rect 18551 19391 18577 19417
rect 19335 19391 19361 19417
rect 20959 19391 20985 19417
rect 21799 19391 21825 19417
rect 22527 19391 22553 19417
rect 23255 19391 23281 19417
rect 23703 19391 23729 19417
rect 23871 19391 23897 19417
rect 24039 19391 24065 19417
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 1583 18999 1609 19025
rect 2479 18999 2505 19025
rect 3823 18999 3849 19025
rect 4383 18999 4409 19025
rect 4495 18999 4521 19025
rect 5279 18999 5305 19025
rect 6455 18999 6481 19025
rect 8135 18999 8161 19025
rect 9031 18999 9057 19025
rect 10823 18999 10849 19025
rect 11271 18999 11297 19025
rect 11495 18999 11521 19025
rect 12279 18999 12305 19025
rect 13455 18999 13481 19025
rect 14911 18999 14937 19025
rect 15359 18999 15385 19025
rect 15471 18999 15497 19025
rect 16255 18999 16281 19025
rect 17431 18999 17457 19025
rect 19055 18999 19081 19025
rect 19335 18999 19361 19025
rect 19447 18999 19473 19025
rect 20231 18999 20257 19025
rect 21239 18999 21265 19025
rect 22751 18999 22777 19025
rect 23255 18999 23281 19025
rect 23423 18999 23449 19025
rect 2479 18943 2505 18969
rect 6455 18943 6481 18969
rect 9031 18943 9057 18969
rect 13455 18943 13481 18969
rect 17431 18943 17457 18969
rect 21239 18943 21265 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 4439 18663 4465 18689
rect 7015 18663 7041 18689
rect 8415 18663 8441 18689
rect 10039 18663 10065 18689
rect 11271 18663 11297 18689
rect 15471 18663 15497 18689
rect 17991 18663 18017 18689
rect 19335 18663 19361 18689
rect 23423 18663 23449 18689
rect 2143 18607 2169 18633
rect 2423 18607 2449 18633
rect 2535 18607 2561 18633
rect 3599 18607 3625 18633
rect 4439 18607 4465 18633
rect 5839 18607 5865 18633
rect 7015 18607 7041 18633
rect 7295 18607 7321 18633
rect 8415 18607 8441 18633
rect 9143 18607 9169 18633
rect 10039 18607 10065 18633
rect 10319 18607 10345 18633
rect 11271 18607 11297 18633
rect 12839 18607 12865 18633
rect 13399 18607 13425 18633
rect 13511 18607 13537 18633
rect 14575 18607 14601 18633
rect 15471 18607 15497 18633
rect 16871 18607 16897 18633
rect 17991 18607 18017 18633
rect 18551 18607 18577 18633
rect 19335 18607 19361 18633
rect 20959 18607 20985 18633
rect 21239 18607 21265 18633
rect 21463 18607 21489 18633
rect 22527 18607 22553 18633
rect 23423 18607 23449 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 1583 18215 1609 18241
rect 2479 18215 2505 18241
rect 3823 18215 3849 18241
rect 4383 18215 4409 18241
rect 4495 18215 4521 18241
rect 5279 18215 5305 18241
rect 6455 18215 6481 18241
rect 8135 18215 8161 18241
rect 9031 18215 9057 18241
rect 10823 18215 10849 18241
rect 11271 18215 11297 18241
rect 11495 18215 11521 18241
rect 12279 18215 12305 18241
rect 13455 18215 13481 18241
rect 14799 18215 14825 18241
rect 15919 18215 15945 18241
rect 16255 18215 16281 18241
rect 17431 18215 17457 18241
rect 19055 18215 19081 18241
rect 19335 18215 19361 18241
rect 19447 18215 19473 18241
rect 20231 18215 20257 18241
rect 21239 18215 21265 18241
rect 22751 18215 22777 18241
rect 23255 18215 23281 18241
rect 23423 18215 23449 18241
rect 2479 18159 2505 18185
rect 6455 18159 6481 18185
rect 9031 18159 9057 18185
rect 13455 18159 13481 18185
rect 15919 18159 15945 18185
rect 17431 18159 17457 18185
rect 21239 18159 21265 18185
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 3039 17879 3065 17905
rect 7015 17879 7041 17905
rect 8415 17879 8441 17905
rect 9815 17879 9841 17905
rect 11271 17879 11297 17905
rect 15471 17879 15497 17905
rect 17991 17879 18017 17905
rect 19335 17879 19361 17905
rect 23423 17879 23449 17905
rect 2143 17823 2169 17849
rect 3039 17823 3065 17849
rect 3599 17823 3625 17849
rect 3879 17823 3905 17849
rect 4159 17823 4185 17849
rect 5839 17823 5865 17849
rect 7015 17823 7041 17849
rect 7295 17823 7321 17849
rect 8415 17823 8441 17849
rect 9143 17823 9169 17849
rect 9815 17823 9841 17849
rect 10319 17823 10345 17849
rect 11271 17823 11297 17849
rect 13119 17823 13145 17849
rect 13399 17823 13425 17849
rect 13511 17823 13537 17849
rect 14575 17823 14601 17849
rect 15471 17823 15497 17849
rect 16871 17823 16897 17849
rect 17991 17823 18017 17849
rect 18551 17823 18577 17849
rect 19335 17823 19361 17849
rect 20959 17823 20985 17849
rect 21239 17823 21265 17849
rect 21463 17823 21489 17849
rect 22527 17823 22553 17849
rect 23423 17823 23449 17849
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 1583 17431 1609 17457
rect 2479 17431 2505 17457
rect 4103 17431 4129 17457
rect 4383 17431 4409 17457
rect 4495 17431 4521 17457
rect 5279 17431 5305 17457
rect 6455 17431 6481 17457
rect 8135 17431 8161 17457
rect 8415 17431 8441 17457
rect 8527 17431 8553 17457
rect 10823 17431 10849 17457
rect 11271 17431 11297 17457
rect 11495 17431 11521 17457
rect 12559 17431 12585 17457
rect 13455 17431 13481 17457
rect 14799 17431 14825 17457
rect 15919 17431 15945 17457
rect 16255 17431 16281 17457
rect 16815 17431 16841 17457
rect 16927 17431 16953 17457
rect 19055 17431 19081 17457
rect 19335 17431 19361 17457
rect 19447 17431 19473 17457
rect 20231 17431 20257 17457
rect 21239 17431 21265 17457
rect 22751 17431 22777 17457
rect 23255 17431 23281 17457
rect 23423 17431 23449 17457
rect 2479 17375 2505 17401
rect 6455 17375 6481 17401
rect 13455 17375 13481 17401
rect 15919 17375 15945 17401
rect 21239 17375 21265 17401
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 3039 17095 3065 17121
rect 4439 17095 4465 17121
rect 7015 17095 7041 17121
rect 8415 17095 8441 17121
rect 9815 17095 9841 17121
rect 11271 17095 11297 17121
rect 15247 17095 15273 17121
rect 17991 17095 18017 17121
rect 19335 17095 19361 17121
rect 23255 17095 23281 17121
rect 1863 17039 1889 17065
rect 3039 17039 3065 17065
rect 3599 17039 3625 17065
rect 4439 17039 4465 17065
rect 5839 17039 5865 17065
rect 7015 17039 7041 17065
rect 7295 17039 7321 17065
rect 8415 17039 8441 17065
rect 9143 17039 9169 17065
rect 9815 17039 9841 17065
rect 10319 17039 10345 17065
rect 11271 17039 11297 17065
rect 12895 17039 12921 17065
rect 13399 17039 13425 17065
rect 13511 17039 13537 17065
rect 14407 17039 14433 17065
rect 15247 17039 15273 17065
rect 16983 17039 17009 17065
rect 17991 17039 18017 17065
rect 18551 17039 18577 17065
rect 19335 17039 19361 17065
rect 20959 17039 20985 17065
rect 21239 17039 21265 17065
rect 21463 17039 21489 17065
rect 22247 17039 22273 17065
rect 23255 17039 23281 17065
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 1583 16647 1609 16673
rect 2479 16647 2505 16673
rect 4103 16647 4129 16673
rect 4383 16647 4409 16673
rect 4551 16647 4577 16673
rect 5279 16647 5305 16673
rect 6455 16647 6481 16673
rect 8135 16647 8161 16673
rect 8415 16647 8441 16673
rect 8527 16647 8553 16673
rect 10823 16647 10849 16673
rect 11271 16647 11297 16673
rect 11495 16647 11521 16673
rect 12559 16647 12585 16673
rect 13455 16647 13481 16673
rect 14799 16647 14825 16673
rect 15247 16647 15273 16673
rect 15471 16647 15497 16673
rect 16255 16647 16281 16673
rect 16927 16647 16953 16673
rect 19055 16647 19081 16673
rect 19335 16647 19361 16673
rect 19447 16647 19473 16673
rect 20231 16647 20257 16673
rect 21239 16647 21265 16673
rect 22751 16647 22777 16673
rect 23255 16647 23281 16673
rect 23423 16647 23449 16673
rect 2479 16591 2505 16617
rect 6455 16591 6481 16617
rect 13455 16591 13481 16617
rect 17319 16591 17345 16617
rect 21239 16591 21265 16617
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2983 16311 3009 16337
rect 4327 16311 4353 16337
rect 7015 16311 7041 16337
rect 8415 16311 8441 16337
rect 9815 16311 9841 16337
rect 11271 16311 11297 16337
rect 15247 16311 15273 16337
rect 19223 16311 19249 16337
rect 23255 16311 23281 16337
rect 1863 16255 1889 16281
rect 2983 16255 3009 16281
rect 3599 16255 3625 16281
rect 4327 16255 4353 16281
rect 5839 16255 5865 16281
rect 7015 16255 7041 16281
rect 7295 16255 7321 16281
rect 8415 16255 8441 16281
rect 9143 16255 9169 16281
rect 9815 16255 9841 16281
rect 10599 16255 10625 16281
rect 11271 16255 11297 16281
rect 12895 16255 12921 16281
rect 13399 16255 13425 16281
rect 13511 16255 13537 16281
rect 14407 16255 14433 16281
rect 15247 16255 15273 16281
rect 16983 16255 17009 16281
rect 17319 16255 17345 16281
rect 17487 16255 17513 16281
rect 18551 16255 18577 16281
rect 19223 16255 19249 16281
rect 20959 16255 20985 16281
rect 21239 16255 21265 16281
rect 21463 16255 21489 16281
rect 22247 16255 22273 16281
rect 23255 16255 23281 16281
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 1583 15863 1609 15889
rect 2423 15863 2449 15889
rect 3823 15863 3849 15889
rect 4943 15863 4969 15889
rect 5559 15863 5585 15889
rect 5951 15863 5977 15889
rect 7911 15863 7937 15889
rect 9031 15863 9057 15889
rect 11103 15863 11129 15889
rect 11383 15863 11409 15889
rect 11495 15863 11521 15889
rect 12559 15863 12585 15889
rect 12727 15863 12753 15889
rect 12951 15863 12977 15889
rect 14799 15863 14825 15889
rect 15247 15863 15273 15889
rect 15471 15863 15497 15889
rect 16255 15863 16281 15889
rect 17431 15863 17457 15889
rect 19055 15863 19081 15889
rect 19951 15863 19977 15889
rect 20231 15863 20257 15889
rect 21015 15863 21041 15889
rect 22751 15863 22777 15889
rect 23199 15863 23225 15889
rect 23423 15863 23449 15889
rect 2423 15807 2449 15833
rect 4943 15807 4969 15833
rect 6231 15807 6257 15833
rect 9031 15807 9057 15833
rect 17431 15807 17457 15833
rect 19951 15807 19977 15833
rect 21183 15807 21209 15833
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 4495 15527 4521 15553
rect 8471 15527 8497 15553
rect 11495 15527 11521 15553
rect 15247 15527 15273 15553
rect 17991 15527 18017 15553
rect 19279 15527 19305 15553
rect 1863 15471 1889 15497
rect 2423 15471 2449 15497
rect 2535 15471 2561 15497
rect 3599 15471 3625 15497
rect 4495 15471 4521 15497
rect 6119 15471 6145 15497
rect 6287 15471 6313 15497
rect 6511 15471 6537 15497
rect 7295 15471 7321 15497
rect 8471 15471 8497 15497
rect 8863 15471 8889 15497
rect 9311 15471 9337 15497
rect 9535 15471 9561 15497
rect 10599 15471 10625 15497
rect 11495 15471 11521 15497
rect 13119 15471 13145 15497
rect 13287 15471 13313 15497
rect 13511 15471 13537 15497
rect 14575 15471 14601 15497
rect 15247 15471 15273 15497
rect 17095 15471 17121 15497
rect 17991 15471 18017 15497
rect 18271 15471 18297 15497
rect 19279 15471 19305 15497
rect 20791 15471 20817 15497
rect 21239 15471 21265 15497
rect 21463 15471 21489 15497
rect 22247 15471 22273 15497
rect 22695 15471 22721 15497
rect 22919 15471 22945 15497
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 1359 15079 1385 15105
rect 2367 15079 2393 15105
rect 3823 15079 3849 15105
rect 4943 15079 4969 15105
rect 5279 15079 5305 15105
rect 6455 15079 6481 15105
rect 7911 15079 7937 15105
rect 9031 15079 9057 15105
rect 11103 15079 11129 15105
rect 11383 15079 11409 15105
rect 11495 15079 11521 15105
rect 12559 15079 12585 15105
rect 12727 15079 12753 15105
rect 12951 15079 12977 15105
rect 14799 15079 14825 15105
rect 15247 15079 15273 15105
rect 15471 15079 15497 15105
rect 16255 15079 16281 15105
rect 17431 15079 17457 15105
rect 19055 15079 19081 15105
rect 19335 15079 19361 15105
rect 19447 15079 19473 15105
rect 20231 15079 20257 15105
rect 21015 15079 21041 15105
rect 22751 15079 22777 15105
rect 23199 15079 23225 15105
rect 23423 15079 23449 15105
rect 2367 15023 2393 15049
rect 4943 15023 4969 15049
rect 6455 15023 6481 15049
rect 9031 15023 9057 15049
rect 17431 15023 17457 15049
rect 21183 15023 21209 15049
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 4495 14743 4521 14769
rect 6175 14743 6201 14769
rect 11495 14743 11521 14769
rect 15247 14743 15273 14769
rect 19447 14743 19473 14769
rect 1863 14687 1889 14713
rect 2367 14687 2393 14713
rect 2591 14687 2617 14713
rect 3599 14687 3625 14713
rect 4495 14687 4521 14713
rect 5279 14687 5305 14713
rect 6175 14687 6201 14713
rect 6735 14687 6761 14713
rect 6903 14687 6929 14713
rect 7127 14687 7153 14713
rect 8863 14687 8889 14713
rect 9423 14687 9449 14713
rect 9535 14687 9561 14713
rect 10599 14687 10625 14713
rect 11495 14687 11521 14713
rect 13119 14687 13145 14713
rect 13287 14687 13313 14713
rect 13511 14687 13537 14713
rect 14575 14687 14601 14713
rect 15247 14687 15273 14713
rect 17095 14687 17121 14713
rect 17375 14687 17401 14713
rect 17487 14687 17513 14713
rect 18271 14687 18297 14713
rect 19447 14687 19473 14713
rect 20791 14687 20817 14713
rect 21239 14687 21265 14713
rect 21463 14687 21489 14713
rect 22247 14687 22273 14713
rect 22751 14687 22777 14713
rect 22919 14687 22945 14713
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 1583 14295 1609 14321
rect 2143 14295 2169 14321
rect 3823 14295 3849 14321
rect 4999 14295 5025 14321
rect 5559 14295 5585 14321
rect 6175 14295 6201 14321
rect 6847 14295 6873 14321
rect 7295 14295 7321 14321
rect 7519 14295 7545 14321
rect 8415 14295 8441 14321
rect 9423 14295 9449 14321
rect 11103 14295 11129 14321
rect 11383 14295 11409 14321
rect 11495 14295 11521 14321
rect 12559 14295 12585 14321
rect 12727 14295 12753 14321
rect 12951 14295 12977 14321
rect 14799 14295 14825 14321
rect 15247 14295 15273 14321
rect 15471 14295 15497 14321
rect 16255 14295 16281 14321
rect 17431 14295 17457 14321
rect 19055 14295 19081 14321
rect 19335 14295 19361 14321
rect 19447 14295 19473 14321
rect 20231 14295 20257 14321
rect 21015 14295 21041 14321
rect 22863 14295 22889 14321
rect 24039 14295 24065 14321
rect 2255 14239 2281 14265
rect 4999 14239 5025 14265
rect 6231 14239 6257 14265
rect 9423 14239 9449 14265
rect 17431 14239 17457 14265
rect 21183 14239 21209 14265
rect 22863 14239 22889 14265
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 4495 13959 4521 13985
rect 8191 13959 8217 13985
rect 11495 13959 11521 13985
rect 15247 13959 15273 13985
rect 19447 13959 19473 13985
rect 22863 13959 22889 13985
rect 2143 13903 2169 13929
rect 2311 13903 2337 13929
rect 2535 13903 2561 13929
rect 3375 13903 3401 13929
rect 4495 13903 4521 13929
rect 5559 13903 5585 13929
rect 6119 13903 6145 13929
rect 6231 13903 6257 13929
rect 7015 13903 7041 13929
rect 8191 13903 8217 13929
rect 8863 13903 8889 13929
rect 9423 13903 9449 13929
rect 9535 13903 9561 13929
rect 10599 13903 10625 13929
rect 11495 13903 11521 13929
rect 13119 13903 13145 13929
rect 13287 13903 13313 13929
rect 13511 13903 13537 13929
rect 14575 13903 14601 13929
rect 15247 13903 15273 13929
rect 17095 13903 17121 13929
rect 17375 13903 17401 13929
rect 17487 13903 17513 13929
rect 18271 13903 18297 13929
rect 19447 13903 19473 13929
rect 20959 13903 20985 13929
rect 21239 13903 21265 13929
rect 21463 13903 21489 13929
rect 22863 13903 22889 13929
rect 24039 13903 24065 13929
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 1583 13511 1609 13537
rect 2479 13511 2505 13537
rect 3823 13511 3849 13537
rect 4999 13511 5025 13537
rect 5503 13511 5529 13537
rect 6119 13511 6145 13537
rect 7015 13511 7041 13537
rect 8191 13511 8217 13537
rect 8471 13511 8497 13537
rect 9423 13511 9449 13537
rect 11103 13511 11129 13537
rect 11383 13511 11409 13537
rect 11495 13511 11521 13537
rect 12559 13511 12585 13537
rect 12727 13511 12753 13537
rect 12951 13511 12977 13537
rect 14799 13511 14825 13537
rect 15247 13511 15273 13537
rect 15471 13511 15497 13537
rect 16255 13511 16281 13537
rect 17431 13511 17457 13537
rect 19055 13511 19081 13537
rect 19335 13511 19361 13537
rect 19447 13511 19473 13537
rect 20511 13511 20537 13537
rect 21407 13511 21433 13537
rect 22863 13511 22889 13537
rect 24039 13511 24065 13537
rect 2479 13455 2505 13481
rect 4999 13455 5025 13481
rect 6231 13455 6257 13481
rect 8191 13455 8217 13481
rect 9423 13455 9449 13481
rect 17431 13455 17457 13481
rect 21407 13455 21433 13481
rect 22863 13455 22889 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 4495 13175 4521 13201
rect 8135 13175 8161 13201
rect 11495 13175 11521 13201
rect 15247 13175 15273 13201
rect 22863 13175 22889 13201
rect 2143 13119 2169 13145
rect 2423 13119 2449 13145
rect 2535 13119 2561 13145
rect 3375 13119 3401 13145
rect 4495 13119 4521 13145
rect 5503 13119 5529 13145
rect 6063 13119 6089 13145
rect 6231 13119 6257 13145
rect 6959 13119 6985 13145
rect 8135 13119 8161 13145
rect 8863 13119 8889 13145
rect 9423 13119 9449 13145
rect 9535 13119 9561 13145
rect 10599 13119 10625 13145
rect 11495 13119 11521 13145
rect 13119 13119 13145 13145
rect 13287 13119 13313 13145
rect 13511 13119 13537 13145
rect 14575 13119 14601 13145
rect 15247 13119 15273 13145
rect 17095 13119 17121 13145
rect 17263 13119 17289 13145
rect 17487 13119 17513 13145
rect 18271 13119 18297 13145
rect 18719 13119 18745 13145
rect 18943 13119 18969 13145
rect 20959 13119 20985 13145
rect 21239 13119 21265 13145
rect 21463 13119 21489 13145
rect 22863 13119 22889 13145
rect 24039 13119 24065 13145
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 1583 12727 1609 12753
rect 2367 12727 2393 12753
rect 3823 12727 3849 12753
rect 4999 12727 5025 12753
rect 5503 12727 5529 12753
rect 6063 12727 6089 12753
rect 7015 12727 7041 12753
rect 8191 12727 8217 12753
rect 8471 12727 8497 12753
rect 9423 12727 9449 12753
rect 11103 12727 11129 12753
rect 11383 12727 11409 12753
rect 11495 12727 11521 12753
rect 12559 12727 12585 12753
rect 12727 12727 12753 12753
rect 12951 12727 12977 12753
rect 14799 12727 14825 12753
rect 15247 12727 15273 12753
rect 15471 12727 15497 12753
rect 16255 12727 16281 12753
rect 17263 12727 17289 12753
rect 19055 12727 19081 12753
rect 19335 12727 19361 12753
rect 19447 12727 19473 12753
rect 20511 12727 20537 12753
rect 21239 12727 21265 12753
rect 22863 12727 22889 12753
rect 24039 12727 24065 12753
rect 2367 12671 2393 12697
rect 4999 12671 5025 12697
rect 6231 12671 6257 12697
rect 8191 12671 8217 12697
rect 9423 12671 9449 12697
rect 17263 12671 17289 12697
rect 21239 12671 21265 12697
rect 22863 12671 22889 12697
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8135 12391 8161 12417
rect 11495 12391 11521 12417
rect 15247 12391 15273 12417
rect 19279 12391 19305 12417
rect 22863 12391 22889 12417
rect 2143 12335 2169 12361
rect 2423 12335 2449 12361
rect 2535 12335 2561 12361
rect 3599 12335 3625 12361
rect 3767 12335 3793 12361
rect 3991 12335 4017 12361
rect 5503 12335 5529 12361
rect 6063 12335 6089 12361
rect 6231 12335 6257 12361
rect 6959 12335 6985 12361
rect 8135 12335 8161 12361
rect 8863 12335 8889 12361
rect 9423 12335 9449 12361
rect 9535 12335 9561 12361
rect 10599 12335 10625 12361
rect 11495 12335 11521 12361
rect 13119 12335 13145 12361
rect 13287 12335 13313 12361
rect 13511 12335 13537 12361
rect 14575 12335 14601 12361
rect 15135 12335 15161 12361
rect 17095 12335 17121 12361
rect 17263 12335 17289 12361
rect 17487 12335 17513 12361
rect 18551 12335 18577 12361
rect 19279 12335 19305 12361
rect 21631 12335 21657 12361
rect 22135 12335 22161 12361
rect 22583 12335 22609 12361
rect 22863 12335 22889 12361
rect 24039 12335 24065 12361
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 1583 11943 1609 11969
rect 2479 11943 2505 11969
rect 3319 11943 3345 11969
rect 3767 11943 3793 11969
rect 4495 11943 4521 11969
rect 5671 11943 5697 11969
rect 7015 11943 7041 11969
rect 8191 11943 8217 11969
rect 8471 11943 8497 11969
rect 9423 11943 9449 11969
rect 11103 11943 11129 11969
rect 11383 11943 11409 11969
rect 11495 11943 11521 11969
rect 12559 11943 12585 11969
rect 12727 11943 12753 11969
rect 12951 11943 12977 11969
rect 14799 11943 14825 11969
rect 15919 11943 15945 11969
rect 16255 11943 16281 11969
rect 17431 11943 17457 11969
rect 19055 11943 19081 11969
rect 19223 11943 19249 11969
rect 19447 11943 19473 11969
rect 21631 11943 21657 11969
rect 21799 11943 21825 11969
rect 22359 11943 22385 11969
rect 22863 11943 22889 11969
rect 24039 11943 24065 11969
rect 2479 11887 2505 11913
rect 3991 11887 4017 11913
rect 5671 11887 5697 11913
rect 8191 11887 8217 11913
rect 9423 11887 9449 11913
rect 15919 11887 15945 11913
rect 17431 11887 17457 11913
rect 22863 11887 22889 11913
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 2871 11607 2897 11633
rect 4495 11607 4521 11633
rect 5839 11607 5865 11633
rect 8191 11607 8217 11633
rect 10039 11607 10065 11633
rect 11495 11607 11521 11633
rect 15471 11607 15497 11633
rect 17823 11607 17849 11633
rect 21631 11607 21657 11633
rect 22863 11607 22889 11633
rect 2143 11551 2169 11577
rect 2871 11551 2897 11577
rect 3431 11551 3457 11577
rect 4495 11551 4521 11577
rect 5055 11551 5081 11577
rect 5839 11551 5865 11577
rect 7295 11551 7321 11577
rect 8191 11551 8217 11577
rect 8863 11551 8889 11577
rect 10039 11551 10065 11577
rect 10599 11551 10625 11577
rect 11495 11551 11521 11577
rect 13119 11551 13145 11577
rect 13287 11551 13313 11577
rect 13511 11551 13537 11577
rect 14575 11551 14601 11577
rect 15471 11551 15497 11577
rect 17095 11551 17121 11577
rect 17823 11551 17849 11577
rect 18439 11551 18465 11577
rect 18719 11551 18745 11577
rect 18943 11551 18969 11577
rect 21687 11551 21713 11577
rect 22583 11551 22609 11577
rect 22863 11551 22889 11577
rect 24039 11551 24065 11577
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 1583 11159 1609 11185
rect 2479 11159 2505 11185
rect 3431 11159 3457 11185
rect 4607 11159 4633 11185
rect 5055 11159 5081 11185
rect 5839 11159 5865 11185
rect 7239 11159 7265 11185
rect 8079 11159 8105 11185
rect 8415 11159 8441 11185
rect 9423 11159 9449 11185
rect 11103 11159 11129 11185
rect 11383 11159 11409 11185
rect 11495 11159 11521 11185
rect 12559 11159 12585 11185
rect 12727 11159 12753 11185
rect 12951 11159 12977 11185
rect 14799 11159 14825 11185
rect 15359 11159 15385 11185
rect 15471 11159 15497 11185
rect 16535 11159 16561 11185
rect 16815 11159 16841 11185
rect 16927 11159 16953 11185
rect 20231 11159 20257 11185
rect 20399 11159 20425 11185
rect 20903 11159 20929 11185
rect 21687 11159 21713 11185
rect 21799 11159 21825 11185
rect 22359 11159 22385 11185
rect 22975 11159 23001 11185
rect 24039 11159 24065 11185
rect 2479 11103 2505 11129
rect 4607 11103 4633 11129
rect 5839 11103 5865 11129
rect 8079 11103 8105 11129
rect 9423 11103 9449 11129
rect 22975 11103 23001 11129
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 2815 10823 2841 10849
rect 4495 10823 4521 10849
rect 5839 10823 5865 10849
rect 8079 10823 8105 10849
rect 11495 10823 11521 10849
rect 13791 10823 13817 10849
rect 15359 10823 15385 10849
rect 17767 10823 17793 10849
rect 20399 10823 20425 10849
rect 22975 10823 23001 10849
rect 2143 10767 2169 10793
rect 2815 10767 2841 10793
rect 3431 10767 3457 10793
rect 4495 10767 4521 10793
rect 5055 10767 5081 10793
rect 5839 10767 5865 10793
rect 7239 10767 7265 10793
rect 8079 10767 8105 10793
rect 8863 10767 8889 10793
rect 9423 10767 9449 10793
rect 9591 10767 9617 10793
rect 10599 10767 10625 10793
rect 11495 10767 11521 10793
rect 13119 10767 13145 10793
rect 13791 10767 13817 10793
rect 14575 10767 14601 10793
rect 15359 10767 15385 10793
rect 17095 10767 17121 10793
rect 17767 10767 17793 10793
rect 19447 10767 19473 10793
rect 20399 10767 20425 10793
rect 21631 10767 21657 10793
rect 21855 10767 21881 10793
rect 22079 10767 22105 10793
rect 22975 10767 23001 10793
rect 24039 10767 24065 10793
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 1583 10375 1609 10401
rect 2479 10375 2505 10401
rect 3431 10375 3457 10401
rect 4607 10375 4633 10401
rect 5055 10375 5081 10401
rect 5839 10375 5865 10401
rect 7239 10375 7265 10401
rect 8079 10375 8105 10401
rect 8415 10375 8441 10401
rect 9591 10375 9617 10401
rect 11103 10375 11129 10401
rect 11383 10375 11409 10401
rect 11495 10375 11521 10401
rect 12559 10375 12585 10401
rect 13455 10375 13481 10401
rect 14799 10375 14825 10401
rect 15359 10375 15385 10401
rect 15471 10375 15497 10401
rect 16479 10375 16505 10401
rect 16815 10375 16841 10401
rect 16927 10375 16953 10401
rect 20007 10375 20033 10401
rect 20903 10375 20929 10401
rect 21463 10375 21489 10401
rect 22079 10375 22105 10401
rect 22975 10375 23001 10401
rect 24039 10375 24065 10401
rect 2479 10319 2505 10345
rect 4607 10319 4633 10345
rect 5839 10319 5865 10345
rect 8079 10319 8105 10345
rect 9591 10319 9617 10345
rect 13455 10319 13481 10345
rect 20903 10319 20929 10345
rect 22135 10319 22161 10345
rect 22975 10319 23001 10345
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 4495 10039 4521 10065
rect 6679 10039 6705 10065
rect 8135 10039 8161 10065
rect 9815 10039 9841 10065
rect 14015 10039 14041 10065
rect 15359 10039 15385 10065
rect 17991 10039 18017 10065
rect 22583 10039 22609 10065
rect 22919 10039 22945 10065
rect 2143 9983 2169 10009
rect 2423 9983 2449 10009
rect 2535 9983 2561 10009
rect 3599 9983 3625 10009
rect 4495 9983 4521 10009
rect 5503 9983 5529 10009
rect 6679 9983 6705 10009
rect 7239 9983 7265 10009
rect 8135 9983 8161 10009
rect 9143 9983 9169 10009
rect 9815 9983 9841 10009
rect 10319 9983 10345 10009
rect 10879 9983 10905 10009
rect 10991 9983 11017 10009
rect 12839 9983 12865 10009
rect 14015 9983 14041 10009
rect 14295 9983 14321 10009
rect 15359 9983 15385 10009
rect 17095 9983 17121 10009
rect 17991 9983 18017 10009
rect 21687 9983 21713 10009
rect 22583 9983 22609 10009
rect 22919 9983 22945 10009
rect 23759 9983 23785 10009
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 1359 9591 1385 9617
rect 2479 9591 2505 9617
rect 3823 9591 3849 9617
rect 4383 9591 4409 9617
rect 4495 9591 4521 9617
rect 5447 9591 5473 9617
rect 6455 9591 6481 9617
rect 7183 9591 7209 9617
rect 8079 9591 8105 9617
rect 8639 9591 8665 9617
rect 9535 9591 9561 9617
rect 11103 9591 11129 9617
rect 11383 9591 11409 9617
rect 11495 9591 11521 9617
rect 12279 9591 12305 9617
rect 13455 9591 13481 9617
rect 14799 9591 14825 9617
rect 15751 9591 15777 9617
rect 16535 9591 16561 9617
rect 17431 9591 17457 9617
rect 21183 9591 21209 9617
rect 22359 9591 22385 9617
rect 22919 9591 22945 9617
rect 23759 9591 23785 9617
rect 2479 9535 2505 9561
rect 6455 9535 6481 9561
rect 8079 9535 8105 9561
rect 9535 9535 9561 9561
rect 13455 9535 13481 9561
rect 15751 9535 15777 9561
rect 17431 9535 17457 9561
rect 22359 9535 22385 9561
rect 22919 9535 22945 9561
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 4495 9255 4521 9281
rect 6679 9255 6705 9281
rect 8135 9255 8161 9281
rect 10039 9255 10065 9281
rect 11495 9255 11521 9281
rect 15471 9255 15497 9281
rect 17991 9255 18017 9281
rect 19223 9255 19249 9281
rect 22583 9255 22609 9281
rect 22919 9255 22945 9281
rect 2143 9199 2169 9225
rect 2423 9199 2449 9225
rect 2535 9199 2561 9225
rect 3599 9199 3625 9225
rect 4495 9199 4521 9225
rect 5503 9199 5529 9225
rect 6679 9199 6705 9225
rect 7239 9199 7265 9225
rect 8135 9199 8161 9225
rect 9143 9199 9169 9225
rect 10039 9199 10065 9225
rect 10319 9199 10345 9225
rect 11495 9199 11521 9225
rect 12839 9199 12865 9225
rect 13399 9199 13425 9225
rect 13511 9199 13537 9225
rect 14575 9199 14601 9225
rect 15471 9199 15497 9225
rect 17095 9199 17121 9225
rect 17991 9199 18017 9225
rect 18551 9199 18577 9225
rect 19223 9199 19249 9225
rect 21407 9199 21433 9225
rect 22583 9199 22609 9225
rect 22919 9199 22945 9225
rect 23759 9199 23785 9225
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 1359 8807 1385 8833
rect 2479 8807 2505 8833
rect 3823 8807 3849 8833
rect 4383 8807 4409 8833
rect 4495 8807 4521 8833
rect 5279 8807 5305 8833
rect 6455 8807 6481 8833
rect 7183 8807 7209 8833
rect 8079 8807 8105 8833
rect 8639 8807 8665 8833
rect 9535 8807 9561 8833
rect 11103 8807 11129 8833
rect 11719 8807 11745 8833
rect 12279 8807 12305 8833
rect 13399 8807 13425 8833
rect 14799 8807 14825 8833
rect 15359 8807 15385 8833
rect 15471 8807 15497 8833
rect 16535 8807 16561 8833
rect 17151 8807 17177 8833
rect 19055 8807 19081 8833
rect 19223 8807 19249 8833
rect 19447 8807 19473 8833
rect 22863 8807 22889 8833
rect 23759 8807 23785 8833
rect 2479 8751 2505 8777
rect 6455 8751 6481 8777
rect 8079 8751 8105 8777
rect 9535 8751 9561 8777
rect 11775 8751 11801 8777
rect 13399 8751 13425 8777
rect 17207 8751 17233 8777
rect 22863 8751 22889 8777
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 6623 8471 6649 8497
rect 8079 8471 8105 8497
rect 11495 8471 11521 8497
rect 14015 8471 14041 8497
rect 15359 8471 15385 8497
rect 19223 8471 19249 8497
rect 22863 8471 22889 8497
rect 2143 8415 2169 8441
rect 2423 8415 2449 8441
rect 2535 8415 2561 8441
rect 3599 8415 3625 8441
rect 3767 8415 3793 8441
rect 4495 8415 4521 8441
rect 5447 8415 5473 8441
rect 6623 8415 6649 8441
rect 7183 8415 7209 8441
rect 8079 8415 8105 8441
rect 9143 8415 9169 8441
rect 9423 8415 9449 8441
rect 9535 8415 9561 8441
rect 10319 8415 10345 8441
rect 11495 8415 11521 8441
rect 13119 8415 13145 8441
rect 14015 8415 14041 8441
rect 14575 8415 14601 8441
rect 15359 8415 15385 8441
rect 17095 8415 17121 8441
rect 17263 8415 17289 8441
rect 17487 8415 17513 8441
rect 18551 8415 18577 8441
rect 19223 8415 19249 8441
rect 22863 8415 22889 8441
rect 23759 8415 23785 8441
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 1359 8023 1385 8049
rect 2479 8023 2505 8049
rect 3823 8023 3849 8049
rect 4999 8023 5025 8049
rect 5279 8023 5305 8049
rect 6455 8023 6481 8049
rect 7239 8023 7265 8049
rect 8135 8023 8161 8049
rect 8695 8023 8721 8049
rect 9423 8023 9449 8049
rect 11103 8023 11129 8049
rect 11383 8023 11409 8049
rect 11495 8023 11521 8049
rect 12559 8023 12585 8049
rect 13455 8023 13481 8049
rect 14799 8023 14825 8049
rect 15359 8023 15385 8049
rect 15471 8023 15497 8049
rect 16535 8023 16561 8049
rect 17431 8023 17457 8049
rect 19055 8023 19081 8049
rect 19223 8023 19249 8049
rect 19447 8023 19473 8049
rect 20231 8023 20257 8049
rect 21015 8023 21041 8049
rect 22919 8023 22945 8049
rect 24039 8023 24065 8049
rect 2479 7967 2505 7993
rect 4999 7967 5025 7993
rect 6455 7967 6481 7993
rect 8135 7967 8161 7993
rect 9423 7967 9449 7993
rect 13455 7967 13481 7993
rect 17431 7967 17457 7993
rect 21183 7967 21209 7993
rect 22919 7967 22945 7993
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 4495 7687 4521 7713
rect 5839 7687 5865 7713
rect 8135 7687 8161 7713
rect 10039 7687 10065 7713
rect 11495 7687 11521 7713
rect 14015 7687 14041 7713
rect 15471 7687 15497 7713
rect 22863 7687 22889 7713
rect 2143 7631 2169 7657
rect 2423 7631 2449 7657
rect 2535 7631 2561 7657
rect 3599 7631 3625 7657
rect 4495 7631 4521 7657
rect 5167 7631 5193 7657
rect 5839 7631 5865 7657
rect 7239 7631 7265 7657
rect 8135 7631 8161 7657
rect 9143 7631 9169 7657
rect 10039 7631 10065 7657
rect 10319 7631 10345 7657
rect 11495 7631 11521 7657
rect 13119 7631 13145 7657
rect 14015 7631 14041 7657
rect 14575 7631 14601 7657
rect 15471 7631 15497 7657
rect 17095 7631 17121 7657
rect 17375 7631 17401 7657
rect 17487 7631 17513 7657
rect 18551 7631 18577 7657
rect 18719 7631 18745 7657
rect 18943 7631 18969 7657
rect 20791 7631 20817 7657
rect 21239 7631 21265 7657
rect 21463 7631 21489 7657
rect 22863 7631 22889 7657
rect 24039 7631 24065 7657
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 1359 7239 1385 7265
rect 2031 7239 2057 7265
rect 3599 7239 3625 7265
rect 4495 7239 4521 7265
rect 4887 7239 4913 7265
rect 5839 7239 5865 7265
rect 7239 7239 7265 7265
rect 8135 7239 8161 7265
rect 8695 7239 8721 7265
rect 9591 7239 9617 7265
rect 11103 7239 11129 7265
rect 11383 7239 11409 7265
rect 11495 7239 11521 7265
rect 12559 7239 12585 7265
rect 13455 7239 13481 7265
rect 14799 7239 14825 7265
rect 15359 7239 15385 7265
rect 15471 7239 15497 7265
rect 16535 7239 16561 7265
rect 17431 7239 17457 7265
rect 18775 7239 18801 7265
rect 19223 7239 19249 7265
rect 19447 7239 19473 7265
rect 20231 7239 20257 7265
rect 21015 7239 21041 7265
rect 22919 7239 22945 7265
rect 23815 7239 23841 7265
rect 2255 7183 2281 7209
rect 4495 7183 4521 7209
rect 5839 7183 5865 7209
rect 8135 7183 8161 7209
rect 9591 7183 9617 7209
rect 13455 7183 13481 7209
rect 17431 7183 17457 7209
rect 21183 7183 21209 7209
rect 22919 7183 22945 7209
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 2871 6903 2897 6929
rect 4495 6903 4521 6929
rect 5839 6903 5865 6929
rect 8079 6903 8105 6929
rect 10879 6903 10905 6929
rect 12447 6903 12473 6929
rect 14015 6903 14041 6929
rect 15359 6903 15385 6929
rect 22863 6903 22889 6929
rect 1919 6847 1945 6873
rect 2871 6847 2897 6873
rect 3599 6847 3625 6873
rect 4495 6847 4521 6873
rect 4887 6847 4913 6873
rect 5839 6847 5865 6873
rect 7183 6847 7209 6873
rect 8079 6847 8105 6873
rect 9815 6847 9841 6873
rect 10879 6847 10905 6873
rect 11551 6847 11577 6873
rect 12447 6847 12473 6873
rect 13119 6847 13145 6873
rect 14015 6847 14041 6873
rect 14575 6847 14601 6873
rect 15359 6847 15385 6873
rect 17095 6847 17121 6873
rect 17263 6847 17289 6873
rect 17487 6847 17513 6873
rect 18271 6847 18297 6873
rect 18719 6847 18745 6873
rect 18943 6847 18969 6873
rect 22863 6847 22889 6873
rect 23759 6847 23785 6873
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 1583 6455 1609 6481
rect 2479 6455 2505 6481
rect 4159 6455 4185 6481
rect 4999 6455 5025 6481
rect 5279 6455 5305 6481
rect 6455 6455 6481 6481
rect 7799 6455 7825 6481
rect 8975 6455 9001 6481
rect 9535 6455 9561 6481
rect 10431 6455 10457 6481
rect 12055 6455 12081 6481
rect 12951 6455 12977 6481
rect 13399 6455 13425 6481
rect 14239 6455 14265 6481
rect 14799 6455 14825 6481
rect 15359 6455 15385 6481
rect 15471 6455 15497 6481
rect 16535 6455 16561 6481
rect 17207 6455 17233 6481
rect 18775 6455 18801 6481
rect 19223 6455 19249 6481
rect 19447 6455 19473 6481
rect 20231 6455 20257 6481
rect 20679 6455 20705 6481
rect 21015 6455 21041 6481
rect 22863 6455 22889 6481
rect 23815 6455 23841 6481
rect 2479 6399 2505 6425
rect 4047 6399 4073 6425
rect 5279 6399 5305 6425
rect 7799 6399 7825 6425
rect 10431 6399 10457 6425
rect 12951 6399 12977 6425
rect 14239 6399 14265 6425
rect 17207 6399 17233 6425
rect 22863 6399 22889 6425
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2087 6119 2113 6145
rect 5839 6119 5865 6145
rect 7519 6119 7545 6145
rect 10879 6119 10905 6145
rect 12447 6119 12473 6145
rect 14015 6119 14041 6145
rect 15359 6119 15385 6145
rect 17767 6119 17793 6145
rect 1191 6063 1217 6089
rect 2087 6063 2113 6089
rect 2535 6063 2561 6089
rect 2815 6063 2841 6089
rect 3039 6063 3065 6089
rect 5839 6063 5865 6089
rect 7015 6063 7041 6089
rect 7575 6063 7601 6089
rect 8471 6063 8497 6089
rect 9815 6063 9841 6089
rect 10879 6063 10905 6089
rect 11551 6063 11577 6089
rect 12447 6063 12473 6089
rect 13119 6063 13145 6089
rect 14015 6063 14041 6089
rect 14575 6063 14601 6089
rect 15359 6063 15385 6089
rect 16815 6063 16841 6089
rect 17767 6063 17793 6089
rect 18271 6063 18297 6089
rect 18831 6063 18857 6089
rect 18943 6063 18969 6089
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 1191 5671 1217 5697
rect 2087 5671 2113 5697
rect 2871 5671 2897 5697
rect 3319 5671 3345 5697
rect 3543 5671 3569 5697
rect 5559 5671 5585 5697
rect 6455 5671 6481 5697
rect 7799 5671 7825 5697
rect 8975 5671 9001 5697
rect 9535 5671 9561 5697
rect 10431 5671 10457 5697
rect 12055 5671 12081 5697
rect 12895 5671 12921 5697
rect 13399 5671 13425 5697
rect 14015 5671 14041 5697
rect 14799 5671 14825 5697
rect 15919 5671 15945 5697
rect 16535 5671 16561 5697
rect 17431 5671 17457 5697
rect 19055 5671 19081 5697
rect 19223 5671 19249 5697
rect 19447 5671 19473 5697
rect 2087 5615 2113 5641
rect 6455 5615 6481 5641
rect 7799 5615 7825 5641
rect 10431 5615 10457 5641
rect 12895 5615 12921 5641
rect 14183 5615 14209 5641
rect 15919 5615 15945 5641
rect 17431 5615 17457 5641
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2087 5335 2113 5361
rect 12447 5335 12473 5361
rect 14015 5335 14041 5361
rect 15471 5335 15497 5361
rect 17767 5335 17793 5361
rect 1191 5279 1217 5305
rect 2087 5279 2113 5305
rect 2535 5279 2561 5305
rect 2815 5279 2841 5305
rect 3039 5279 3065 5305
rect 6119 5279 6145 5305
rect 6399 5279 6425 5305
rect 6511 5279 6537 5305
rect 7519 5279 7545 5305
rect 7799 5279 7825 5305
rect 7967 5279 7993 5305
rect 9815 5279 9841 5305
rect 10375 5279 10401 5305
rect 10487 5279 10513 5305
rect 11551 5279 11577 5305
rect 12447 5279 12473 5305
rect 13119 5279 13145 5305
rect 14015 5279 14041 5305
rect 14575 5279 14601 5305
rect 15471 5279 15497 5305
rect 16815 5279 16841 5305
rect 17767 5279 17793 5305
rect 18551 5279 18577 5305
rect 18719 5279 18745 5305
rect 18943 5279 18969 5305
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 1191 4887 1217 4913
rect 2031 4887 2057 4913
rect 2871 4887 2897 4913
rect 3319 4887 3345 4913
rect 3543 4887 3569 4913
rect 8079 4887 8105 4913
rect 8247 4887 8273 4913
rect 8471 4887 8497 4913
rect 9535 4887 9561 4913
rect 10431 4887 10457 4913
rect 12055 4887 12081 4913
rect 12895 4887 12921 4913
rect 13399 4887 13425 4913
rect 14239 4887 14265 4913
rect 14799 4887 14825 4913
rect 15919 4887 15945 4913
rect 16535 4887 16561 4913
rect 17431 4887 17457 4913
rect 2031 4831 2057 4857
rect 10431 4831 10457 4857
rect 12895 4831 12921 4857
rect 14239 4831 14265 4857
rect 15919 4831 15945 4857
rect 17431 4831 17457 4857
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2031 4551 2057 4577
rect 3319 4551 3345 4577
rect 10879 4551 10905 4577
rect 12391 4551 12417 4577
rect 13959 4551 13985 4577
rect 15471 4551 15497 4577
rect 1191 4495 1217 4521
rect 2031 4495 2057 4521
rect 2535 4495 2561 4521
rect 3319 4495 3345 4521
rect 6343 4495 6369 4521
rect 6511 4495 6537 4521
rect 7015 4495 7041 4521
rect 7519 4495 7545 4521
rect 7743 4495 7769 4521
rect 7967 4495 7993 4521
rect 10039 4495 10065 4521
rect 10879 4495 10905 4521
rect 11551 4495 11577 4521
rect 12391 4495 12417 4521
rect 13119 4495 13145 4521
rect 13959 4495 13985 4521
rect 14575 4495 14601 4521
rect 15471 4495 15497 4521
rect 17095 4495 17121 4521
rect 17375 4495 17401 4521
rect 17487 4495 17513 4521
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 1023 4103 1049 4129
rect 1863 4103 1889 4129
rect 5783 4103 5809 4129
rect 5895 4103 5921 4129
rect 6455 4103 6481 4129
rect 7799 4103 7825 4129
rect 8247 4103 8273 4129
rect 8471 4103 8497 4129
rect 9535 4103 9561 4129
rect 10375 4103 10401 4129
rect 11775 4103 11801 4129
rect 12951 4103 12977 4129
rect 13231 4103 13257 4129
rect 14183 4103 14209 4129
rect 15079 4103 15105 4129
rect 15919 4103 15945 4129
rect 16255 4103 16281 4129
rect 17207 4103 17233 4129
rect 22919 4103 22945 4129
rect 24039 4103 24065 4129
rect 1863 4047 1889 4073
rect 10375 4047 10401 4073
rect 12951 4047 12977 4073
rect 14183 4047 14209 4073
rect 15919 4047 15945 4073
rect 17207 4047 17233 4073
rect 22919 4047 22945 4073
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 1863 3767 1889 3793
rect 5839 3767 5865 3793
rect 10879 3767 10905 3793
rect 12447 3767 12473 3793
rect 13959 3767 13985 3793
rect 15471 3767 15497 3793
rect 1023 3711 1049 3737
rect 1863 3711 1889 3737
rect 5839 3711 5865 3737
rect 7015 3711 7041 3737
rect 7519 3711 7545 3737
rect 7799 3711 7825 3737
rect 7967 3711 7993 3737
rect 9815 3711 9841 3737
rect 10879 3711 10905 3737
rect 11271 3711 11297 3737
rect 12447 3711 12473 3737
rect 12839 3711 12865 3737
rect 13959 3711 13985 3737
rect 14575 3711 14601 3737
rect 15471 3711 15497 3737
rect 16815 3711 16841 3737
rect 17263 3711 17289 3737
rect 17487 3711 17513 3737
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 8079 3319 8105 3345
rect 8247 3319 8273 3345
rect 8471 3319 8497 3345
rect 9535 3319 9561 3345
rect 10431 3319 10457 3345
rect 11775 3319 11801 3345
rect 12895 3319 12921 3345
rect 13399 3319 13425 3345
rect 14127 3319 14153 3345
rect 15079 3319 15105 3345
rect 15583 3319 15609 3345
rect 16255 3319 16281 3345
rect 17207 3319 17233 3345
rect 10431 3263 10457 3289
rect 12895 3263 12921 3289
rect 14127 3263 14153 3289
rect 15751 3263 15777 3289
rect 17207 3263 17233 3289
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 1863 2983 1889 3009
rect 5839 2983 5865 3009
rect 8471 2983 8497 3009
rect 10767 2983 10793 3009
rect 12335 2983 12361 3009
rect 14015 2983 14041 3009
rect 15471 2983 15497 3009
rect 911 2927 937 2953
rect 1863 2927 1889 2953
rect 5839 2927 5865 2953
rect 7015 2927 7041 2953
rect 7575 2927 7601 2953
rect 8471 2927 8497 2953
rect 10039 2927 10065 2953
rect 10767 2927 10793 2953
rect 11551 2927 11577 2953
rect 12335 2927 12361 2953
rect 13119 2927 13145 2953
rect 14015 2927 14041 2953
rect 14575 2927 14601 2953
rect 15471 2927 15497 2953
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 911 2535 937 2561
rect 2087 2535 2113 2561
rect 5279 2535 5305 2561
rect 6231 2535 6257 2561
rect 8079 2535 8105 2561
rect 8975 2535 9001 2561
rect 9255 2535 9281 2561
rect 10431 2535 10457 2561
rect 11775 2535 11801 2561
rect 12895 2535 12921 2561
rect 13175 2535 13201 2561
rect 14015 2535 14041 2561
rect 14799 2535 14825 2561
rect 15359 2535 15385 2561
rect 15471 2535 15497 2561
rect 2087 2479 2113 2505
rect 5279 2479 5305 2505
rect 8975 2479 9001 2505
rect 10431 2479 10457 2505
rect 12895 2479 12921 2505
rect 14127 2479 14153 2505
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 3767 2199 3793 2225
rect 10767 2199 10793 2225
rect 12447 2199 12473 2225
rect 14015 2199 14041 2225
rect 15359 2199 15385 2225
rect 2871 2143 2897 2169
rect 3767 2143 3793 2169
rect 7015 2143 7041 2169
rect 7575 2143 7601 2169
rect 7687 2143 7713 2169
rect 9815 2143 9841 2169
rect 10767 2143 10793 2169
rect 11551 2143 11577 2169
rect 12447 2143 12473 2169
rect 13119 2143 13145 2169
rect 14015 2143 14041 2169
rect 14295 2143 14321 2169
rect 15359 2143 15385 2169
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 2871 1751 2897 1777
rect 3823 1751 3849 1777
rect 7015 1751 7041 1777
rect 7575 1751 7601 1777
rect 7687 1751 7713 1777
rect 9423 1751 9449 1777
rect 9591 1751 9617 1777
rect 9815 1751 9841 1777
rect 11103 1751 11129 1777
rect 12279 1751 12305 1777
rect 12951 1751 12977 1777
rect 13847 1751 13873 1777
rect 3823 1695 3849 1721
rect 12279 1695 12305 1721
rect 13847 1695 13873 1721
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 1680 34600 1736 35000
rect 4214 34622 4634 34650
rect 1694 33614 1722 34600
rect 4214 33614 4242 34622
rect 4606 34538 4634 34622
rect 4760 34600 4816 35000
rect 7840 34600 7896 35000
rect 10920 34600 10976 35000
rect 14000 34600 14056 35000
rect 17080 34600 17136 35000
rect 20160 34600 20216 35000
rect 22694 34622 23114 34650
rect 4774 34538 4802 34600
rect 4606 34510 4802 34538
rect 1694 33586 2170 33614
rect 4214 33586 4354 33614
rect 1750 32802 1778 32807
rect 1358 27649 1386 27655
rect 1358 27623 1359 27649
rect 1385 27623 1386 27649
rect 1358 26922 1386 27623
rect 1358 26865 1386 26894
rect 1358 26839 1359 26865
rect 1385 26839 1386 26865
rect 1358 26081 1386 26839
rect 1358 26055 1359 26081
rect 1385 26055 1386 26081
rect 1358 24513 1386 26055
rect 1582 25690 1610 25695
rect 1582 25297 1610 25662
rect 1750 25690 1778 32774
rect 1750 25657 1778 25662
rect 1806 28434 1834 28439
rect 1582 25271 1583 25297
rect 1609 25271 1610 25297
rect 1582 25265 1610 25271
rect 1358 24487 1359 24513
rect 1385 24487 1386 24513
rect 1358 24066 1386 24487
rect 1358 23729 1386 24038
rect 1358 23703 1359 23729
rect 1385 23703 1386 23729
rect 1358 23562 1386 23703
rect 1358 22945 1386 23534
rect 1358 22919 1359 22945
rect 1385 22919 1386 22945
rect 1358 22161 1386 22919
rect 1806 22554 1834 28406
rect 1862 28041 1890 28047
rect 1862 28015 1863 28041
rect 1889 28015 1890 28041
rect 1862 27257 1890 28015
rect 2142 28042 2170 33586
rect 2238 33334 2370 33339
rect 2266 33306 2290 33334
rect 2318 33306 2342 33334
rect 2238 33301 2370 33306
rect 2238 32550 2370 32555
rect 2266 32522 2290 32550
rect 2318 32522 2342 32550
rect 2238 32517 2370 32522
rect 2238 31766 2370 31771
rect 2266 31738 2290 31766
rect 2318 31738 2342 31766
rect 2238 31733 2370 31738
rect 2238 30982 2370 30987
rect 2266 30954 2290 30982
rect 2318 30954 2342 30982
rect 2238 30949 2370 30954
rect 2238 30198 2370 30203
rect 2266 30170 2290 30198
rect 2318 30170 2342 30198
rect 2238 30165 2370 30170
rect 2238 29414 2370 29419
rect 2266 29386 2290 29414
rect 2318 29386 2342 29414
rect 2238 29381 2370 29386
rect 3934 29217 3962 29223
rect 3934 29191 3935 29217
rect 3961 29191 3962 29217
rect 3598 28826 3626 28831
rect 3934 28826 3962 29191
rect 3598 28825 3962 28826
rect 3598 28799 3599 28825
rect 3625 28799 3962 28825
rect 3598 28798 3962 28799
rect 2238 28630 2370 28635
rect 2266 28602 2290 28630
rect 2318 28602 2342 28630
rect 2238 28597 2370 28602
rect 2310 28042 2338 28047
rect 2534 28042 2562 28047
rect 2142 28041 2562 28042
rect 2142 28015 2311 28041
rect 2337 28015 2535 28041
rect 2561 28015 2562 28041
rect 2142 28014 2562 28015
rect 2310 28009 2338 28014
rect 2238 27846 2370 27851
rect 2266 27818 2290 27846
rect 2318 27818 2342 27846
rect 2238 27813 2370 27818
rect 2478 27649 2506 28014
rect 2534 28009 2562 28014
rect 3598 28041 3626 28798
rect 3934 28433 3962 28798
rect 4326 28714 4354 33586
rect 7854 29610 7882 34600
rect 9918 32942 10050 32947
rect 9946 32914 9970 32942
rect 9998 32914 10022 32942
rect 9918 32909 10050 32914
rect 9918 32158 10050 32163
rect 9946 32130 9970 32158
rect 9998 32130 10022 32158
rect 9918 32125 10050 32130
rect 9918 31374 10050 31379
rect 9946 31346 9970 31374
rect 9998 31346 10022 31374
rect 9918 31341 10050 31346
rect 9918 30590 10050 30595
rect 9946 30562 9970 30590
rect 9998 30562 10022 30590
rect 9918 30557 10050 30562
rect 9918 29806 10050 29811
rect 9946 29778 9970 29806
rect 9998 29778 10022 29806
rect 9918 29773 10050 29778
rect 7854 29577 7882 29582
rect 3934 28407 3935 28433
rect 3961 28407 3962 28433
rect 3934 28401 3962 28407
rect 4214 28686 4354 28714
rect 4382 29218 4410 29223
rect 4606 29218 4634 29223
rect 4382 29217 4634 29218
rect 4382 29191 4383 29217
rect 4409 29191 4607 29217
rect 4633 29191 4634 29217
rect 4382 29190 4634 29191
rect 4382 28881 4410 29190
rect 4606 29185 4634 29190
rect 9918 29022 10050 29027
rect 9946 28994 9970 29022
rect 9998 28994 10022 29022
rect 9918 28989 10050 28994
rect 4382 28855 4383 28881
rect 4409 28855 4410 28881
rect 4382 28825 4410 28855
rect 5838 28881 5866 28887
rect 5838 28855 5839 28881
rect 5865 28855 5866 28881
rect 4382 28799 4383 28825
rect 4409 28799 4410 28825
rect 3598 28015 3599 28041
rect 3625 28015 3626 28041
rect 3598 27734 3626 28015
rect 3878 28042 3906 28047
rect 4046 28042 4074 28047
rect 3878 28041 4074 28042
rect 3878 28015 3879 28041
rect 3905 28015 4047 28041
rect 4073 28015 4074 28041
rect 3878 28014 4074 28015
rect 3878 28009 3906 28014
rect 4046 27734 4074 28014
rect 2478 27623 2479 27649
rect 2505 27623 2506 27649
rect 2478 27593 2506 27623
rect 2478 27567 2479 27593
rect 2505 27567 2506 27593
rect 1862 27231 1863 27257
rect 1889 27231 1890 27257
rect 1862 26922 1890 27231
rect 2422 27258 2450 27263
rect 2478 27258 2506 27567
rect 3318 27706 3626 27734
rect 3990 27706 4074 27734
rect 3318 27649 3346 27706
rect 3318 27623 3319 27649
rect 3345 27623 3346 27649
rect 2534 27258 2562 27263
rect 2422 27257 2562 27258
rect 2422 27231 2423 27257
rect 2449 27231 2535 27257
rect 2561 27231 2562 27257
rect 2422 27230 2562 27231
rect 2422 27225 2450 27230
rect 1862 26473 1890 26894
rect 1862 26447 1863 26473
rect 1889 26447 1890 26473
rect 1862 26441 1890 26447
rect 2086 27202 2114 27207
rect 1862 24905 1890 24911
rect 1862 24879 1863 24905
rect 1889 24879 1890 24905
rect 1862 24346 1890 24879
rect 1862 24121 1890 24318
rect 1862 24095 1863 24121
rect 1889 24095 1890 24121
rect 1862 23562 1890 24095
rect 1862 23337 1890 23534
rect 1862 23311 1863 23337
rect 1889 23311 1890 23337
rect 1862 23305 1890 23311
rect 1862 22554 1890 22559
rect 1806 22553 1890 22554
rect 1806 22527 1863 22553
rect 1889 22527 1890 22553
rect 1806 22526 1890 22527
rect 1358 22135 1359 22161
rect 1385 22135 1386 22161
rect 1358 15105 1386 22135
rect 1862 21770 1890 22526
rect 1862 21737 1890 21742
rect 1582 21377 1610 21383
rect 1582 21351 1583 21377
rect 1609 21351 1610 21377
rect 1582 20593 1610 21351
rect 1582 20567 1583 20593
rect 1609 20567 1610 20593
rect 1582 19809 1610 20567
rect 1582 19783 1583 19809
rect 1609 19783 1610 19809
rect 1582 19025 1610 19783
rect 2086 19698 2114 27174
rect 2238 27062 2370 27067
rect 2266 27034 2290 27062
rect 2318 27034 2342 27062
rect 2238 27029 2370 27034
rect 2534 26922 2562 27230
rect 2478 26894 2534 26922
rect 2478 26865 2506 26894
rect 2534 26889 2562 26894
rect 3318 27257 3346 27623
rect 3990 27649 4018 27678
rect 3990 27623 3991 27649
rect 4017 27623 4018 27649
rect 3990 27593 4018 27623
rect 3990 27567 3991 27593
rect 4017 27567 4018 27593
rect 3766 27258 3794 27263
rect 3990 27258 4018 27567
rect 3318 27231 3319 27257
rect 3345 27231 3346 27257
rect 2478 26839 2479 26865
rect 2505 26839 2506 26865
rect 2478 26809 2506 26839
rect 2478 26783 2479 26809
rect 2505 26783 2506 26809
rect 2422 26474 2450 26479
rect 2478 26474 2506 26783
rect 3318 26865 3346 27231
rect 3710 27257 4018 27258
rect 3710 27231 3767 27257
rect 3793 27231 3991 27257
rect 4017 27231 4018 27257
rect 3710 27230 4018 27231
rect 3318 26839 3319 26865
rect 3345 26839 3346 26865
rect 2534 26474 2562 26479
rect 2422 26473 2562 26474
rect 2422 26447 2423 26473
rect 2449 26447 2535 26473
rect 2561 26447 2562 26473
rect 2422 26446 2562 26447
rect 2422 26441 2450 26446
rect 2238 26278 2370 26283
rect 2266 26250 2290 26278
rect 2318 26250 2342 26278
rect 2238 26245 2370 26250
rect 2478 26081 2506 26446
rect 2534 26441 2562 26446
rect 3318 26473 3346 26839
rect 3486 26922 3514 26927
rect 3486 26865 3514 26894
rect 3486 26839 3487 26865
rect 3513 26839 3514 26865
rect 3486 26833 3514 26839
rect 3710 26922 3738 27230
rect 3766 27225 3794 27230
rect 3990 27225 4018 27230
rect 3710 26865 3738 26894
rect 3710 26839 3711 26865
rect 3737 26839 3738 26865
rect 3710 26833 3738 26839
rect 3318 26447 3319 26473
rect 3345 26447 3346 26473
rect 2478 26055 2479 26081
rect 2505 26055 2506 26081
rect 2478 26025 2506 26055
rect 2478 25999 2479 26025
rect 2505 25999 2506 26025
rect 2142 25690 2170 25695
rect 2142 25643 2170 25662
rect 2238 25494 2370 25499
rect 2266 25466 2290 25494
rect 2318 25466 2342 25494
rect 2238 25461 2370 25466
rect 2478 25298 2506 25999
rect 3318 26081 3346 26447
rect 3318 26055 3319 26081
rect 3345 26055 3346 26081
rect 3038 25745 3066 25751
rect 3038 25719 3039 25745
rect 3065 25719 3066 25745
rect 3038 25690 3066 25719
rect 3038 25689 3178 25690
rect 3038 25663 3039 25689
rect 3065 25663 3178 25689
rect 3038 25662 3178 25663
rect 3038 25657 3066 25662
rect 2478 25241 2506 25270
rect 2478 25215 2479 25241
rect 2505 25215 2506 25241
rect 2478 25209 2506 25215
rect 3150 25298 3178 25662
rect 2422 24906 2450 24911
rect 2534 24906 2562 24911
rect 2422 24905 2562 24906
rect 2422 24879 2423 24905
rect 2449 24879 2535 24905
rect 2561 24879 2562 24905
rect 2422 24878 2562 24879
rect 2422 24873 2450 24878
rect 2238 24710 2370 24715
rect 2266 24682 2290 24710
rect 2318 24682 2342 24710
rect 2238 24677 2370 24682
rect 2478 24513 2506 24878
rect 2534 24873 2562 24878
rect 2478 24487 2479 24513
rect 2505 24487 2506 24513
rect 2478 24457 2506 24487
rect 2478 24431 2479 24457
rect 2505 24431 2506 24457
rect 2238 23926 2370 23931
rect 2266 23898 2290 23926
rect 2318 23898 2342 23926
rect 2238 23893 2370 23898
rect 2478 23729 2506 24431
rect 2478 23703 2479 23729
rect 2505 23703 2506 23729
rect 2478 23674 2506 23703
rect 2238 23142 2370 23147
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2238 23109 2370 23114
rect 2478 22945 2506 23646
rect 3038 24177 3066 24183
rect 3038 24151 3039 24177
rect 3065 24151 3066 24177
rect 3038 24122 3066 24151
rect 3038 23674 3066 24094
rect 3038 23393 3066 23646
rect 3150 23674 3178 25270
rect 3318 25689 3346 26055
rect 3318 25663 3319 25689
rect 3345 25663 3346 25689
rect 3318 25298 3346 25663
rect 4214 26530 4242 28686
rect 4382 27734 4410 28799
rect 5054 28825 5082 28831
rect 5054 28799 5055 28825
rect 5081 28799 5082 28825
rect 4886 28433 4914 28439
rect 4886 28407 4887 28433
rect 4913 28407 4914 28433
rect 4886 28378 4914 28407
rect 4886 28377 5026 28378
rect 4886 28351 4887 28377
rect 4913 28351 5026 28377
rect 4886 28350 5026 28351
rect 4886 28345 4914 28350
rect 4270 27706 4410 27734
rect 4998 27706 5026 28350
rect 5054 28041 5082 28799
rect 5054 28015 5055 28041
rect 5081 28015 5082 28041
rect 5054 27734 5082 28015
rect 5838 28825 5866 28855
rect 5838 28799 5839 28825
rect 5865 28799 5866 28825
rect 5838 28097 5866 28799
rect 9918 28238 10050 28243
rect 9946 28210 9970 28238
rect 9998 28210 10022 28238
rect 9918 28205 10050 28210
rect 5838 28071 5839 28097
rect 5865 28071 5866 28097
rect 5838 28041 5866 28071
rect 7518 28097 7546 28103
rect 7518 28071 7519 28097
rect 7545 28071 7546 28097
rect 5838 28015 5839 28041
rect 5865 28015 5866 28041
rect 5838 27762 5866 28015
rect 5054 27706 5194 27734
rect 5838 27729 5866 27734
rect 6622 28041 6650 28047
rect 6622 28015 6623 28041
rect 6649 28015 6650 28041
rect 4270 27673 4298 27678
rect 4998 27673 5026 27678
rect 4774 27649 4802 27655
rect 4774 27623 4775 27649
rect 4801 27623 4802 27649
rect 4774 26865 4802 27623
rect 4774 26839 4775 26865
rect 4801 26839 4802 26865
rect 4270 26530 4298 26535
rect 4214 26529 4298 26530
rect 4214 26503 4271 26529
rect 4297 26503 4298 26529
rect 4214 26502 4298 26503
rect 4214 26473 4242 26502
rect 4270 26497 4298 26502
rect 4214 26447 4215 26473
rect 4241 26447 4242 26473
rect 4214 26081 4242 26447
rect 4214 26055 4215 26081
rect 4241 26055 4242 26081
rect 4214 26025 4242 26055
rect 4214 25999 4215 26025
rect 4241 25999 4242 26025
rect 4214 25746 4242 25999
rect 4774 26081 4802 26839
rect 5166 27258 5194 27706
rect 5166 26474 5194 27230
rect 5446 27649 5474 27655
rect 5446 27623 5447 27649
rect 5473 27623 5474 27649
rect 5446 27593 5474 27623
rect 5446 27567 5447 27593
rect 5473 27567 5474 27593
rect 5446 27258 5474 27567
rect 5558 27258 5586 27263
rect 5446 27257 5586 27258
rect 5446 27231 5447 27257
rect 5473 27231 5559 27257
rect 5585 27231 5586 27257
rect 5446 27230 5586 27231
rect 5446 26865 5474 27230
rect 5558 27225 5586 27230
rect 6622 27258 6650 28015
rect 7518 28041 7546 28071
rect 7518 28015 7519 28041
rect 7545 28015 7546 28041
rect 6622 27211 6650 27230
rect 7126 27649 7154 27655
rect 7126 27623 7127 27649
rect 7153 27623 7154 27649
rect 7126 27258 7154 27623
rect 5446 26839 5447 26865
rect 5473 26839 5474 26865
rect 5446 26809 5474 26839
rect 7126 26922 7154 27230
rect 7126 26865 7154 26894
rect 7126 26839 7127 26865
rect 7153 26839 7154 26865
rect 7126 26833 7154 26839
rect 7518 27313 7546 28015
rect 10934 27986 10962 34600
rect 14014 33614 14042 34600
rect 17094 33614 17122 34600
rect 14014 33586 14210 33614
rect 17094 33586 17178 33614
rect 10934 27953 10962 27958
rect 7518 27287 7519 27313
rect 7545 27287 7546 27313
rect 7518 27257 7546 27287
rect 7518 27231 7519 27257
rect 7545 27231 7546 27257
rect 5446 26783 5447 26809
rect 5473 26783 5474 26809
rect 5110 26473 5194 26474
rect 5110 26447 5167 26473
rect 5193 26447 5194 26473
rect 5110 26446 5194 26447
rect 4774 26055 4775 26081
rect 4801 26055 4802 26081
rect 4270 25746 4298 25751
rect 4214 25745 4298 25746
rect 4214 25719 4271 25745
rect 4297 25719 4298 25745
rect 4214 25718 4298 25719
rect 4214 25689 4242 25718
rect 4270 25713 4298 25718
rect 4214 25663 4215 25689
rect 4241 25663 4242 25689
rect 3822 25298 3850 25303
rect 3318 25297 3402 25298
rect 3318 25271 3319 25297
rect 3345 25271 3402 25297
rect 3318 25270 3402 25271
rect 3318 25265 3346 25270
rect 3374 24905 3402 25270
rect 3374 24879 3375 24905
rect 3401 24879 3402 24905
rect 3374 24346 3402 24879
rect 3374 24121 3402 24318
rect 3822 24513 3850 25270
rect 4214 25297 4242 25663
rect 4214 25271 4215 25297
rect 4241 25271 4242 25297
rect 4214 25242 4242 25271
rect 4774 25578 4802 26055
rect 4774 25298 4802 25550
rect 4214 25241 4522 25242
rect 4214 25215 4215 25241
rect 4241 25215 4522 25241
rect 4774 25232 4802 25270
rect 4942 26082 4970 26087
rect 4942 25298 4970 26054
rect 5110 25689 5138 26446
rect 5166 26441 5194 26446
rect 5334 26474 5362 26479
rect 5446 26474 5474 26783
rect 7518 26529 7546 27231
rect 7518 26503 7519 26529
rect 7545 26503 7546 26529
rect 5558 26474 5586 26479
rect 5334 26473 5586 26474
rect 5334 26447 5335 26473
rect 5361 26447 5559 26473
rect 5585 26447 5586 26473
rect 5334 26446 5586 26447
rect 5166 26082 5194 26087
rect 5166 26035 5194 26054
rect 5334 26082 5362 26446
rect 5558 26441 5586 26446
rect 6342 26473 6370 26479
rect 6342 26447 6343 26473
rect 6369 26447 6370 26473
rect 5110 25663 5111 25689
rect 5137 25663 5138 25689
rect 5110 25578 5138 25663
rect 5334 25690 5362 26054
rect 5558 25690 5586 25695
rect 5334 25689 5586 25690
rect 5334 25663 5335 25689
rect 5361 25663 5559 25689
rect 5585 25663 5586 25689
rect 5334 25662 5586 25663
rect 5334 25657 5362 25662
rect 5558 25657 5586 25662
rect 6342 25690 6370 26447
rect 7518 26473 7546 26503
rect 7518 26447 7519 26473
rect 7545 26447 7546 26473
rect 7126 26081 7154 26087
rect 7126 26055 7127 26081
rect 7153 26055 7154 26081
rect 6342 25657 6370 25662
rect 6678 25689 6706 25695
rect 6678 25663 6679 25689
rect 6705 25663 6706 25689
rect 5110 25545 5138 25550
rect 5166 25298 5194 25303
rect 4942 25297 5194 25298
rect 4942 25271 4943 25297
rect 4969 25271 5167 25297
rect 5193 25271 5194 25297
rect 4942 25270 5194 25271
rect 4214 25214 4522 25215
rect 4214 25209 4242 25214
rect 4494 25186 4522 25214
rect 4942 25186 4970 25270
rect 5166 25265 5194 25270
rect 4494 25158 4970 25186
rect 4494 24961 4522 25158
rect 4494 24935 4495 24961
rect 4521 24935 4522 24961
rect 4494 24905 4522 24935
rect 6174 24961 6202 24967
rect 6174 24935 6175 24961
rect 6201 24935 6202 24961
rect 4494 24879 4495 24905
rect 4521 24879 4522 24905
rect 3822 24487 3823 24513
rect 3849 24487 3850 24513
rect 3822 24346 3850 24487
rect 4382 24514 4410 24519
rect 4494 24514 4522 24879
rect 4382 24513 4522 24514
rect 4382 24487 4383 24513
rect 4409 24487 4495 24513
rect 4521 24487 4522 24513
rect 4382 24486 4522 24487
rect 4382 24481 4410 24486
rect 3822 24313 3850 24318
rect 3374 24095 3375 24121
rect 3401 24095 3402 24121
rect 3374 24089 3402 24095
rect 4494 24177 4522 24486
rect 4494 24151 4495 24177
rect 4521 24151 4522 24177
rect 4494 24122 4522 24151
rect 5054 24905 5082 24911
rect 5054 24879 5055 24905
rect 5081 24879 5082 24905
rect 5054 24514 5082 24879
rect 6174 24905 6202 24935
rect 6174 24879 6175 24905
rect 6201 24879 6202 24905
rect 5278 24514 5306 24519
rect 5054 24513 5306 24514
rect 5054 24487 5279 24513
rect 5305 24487 5306 24513
rect 5054 24486 5306 24487
rect 4522 24094 4578 24122
rect 4494 24056 4522 24094
rect 3150 23641 3178 23646
rect 4102 23729 4130 23735
rect 4102 23703 4103 23729
rect 4129 23703 4130 23729
rect 4102 23618 4130 23703
rect 4102 23585 4130 23590
rect 4494 23674 4522 23679
rect 3038 23367 3039 23393
rect 3065 23367 3066 23393
rect 3038 23337 3066 23367
rect 4494 23393 4522 23646
rect 4494 23367 4495 23393
rect 4521 23367 4522 23393
rect 3038 23311 3039 23337
rect 3065 23311 3066 23337
rect 3038 23305 3066 23311
rect 3374 23337 3402 23343
rect 3374 23311 3375 23337
rect 3401 23311 3402 23337
rect 2478 22919 2479 22945
rect 2505 22919 2506 22945
rect 2478 22889 2506 22919
rect 2478 22863 2479 22889
rect 2505 22863 2506 22889
rect 2238 22358 2370 22363
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2238 22325 2370 22330
rect 2478 22161 2506 22863
rect 2478 22135 2479 22161
rect 2505 22135 2506 22161
rect 2478 22105 2506 22135
rect 2478 22079 2479 22105
rect 2505 22079 2506 22105
rect 2478 22073 2506 22079
rect 2982 22609 3010 22615
rect 2982 22583 2983 22609
rect 3009 22583 3010 22609
rect 2982 22553 3010 22583
rect 2982 22527 2983 22553
rect 3009 22527 3010 22553
rect 2982 21854 3010 22527
rect 2534 21826 3010 21854
rect 3374 22553 3402 23311
rect 4494 23337 4522 23367
rect 4494 23311 4495 23337
rect 4521 23311 4522 23337
rect 3374 22527 3375 22553
rect 3401 22527 3402 22553
rect 2086 19665 2114 19670
rect 2142 21770 2170 21775
rect 2142 20985 2170 21742
rect 2422 21770 2450 21775
rect 2534 21770 2562 21826
rect 2422 21769 2562 21770
rect 2422 21743 2423 21769
rect 2449 21743 2535 21769
rect 2561 21743 2562 21769
rect 2422 21742 2562 21743
rect 3374 21770 3402 22527
rect 4102 22946 4130 22951
rect 4102 22161 4130 22918
rect 4494 22609 4522 23311
rect 4494 22583 4495 22609
rect 4521 22583 4522 22609
rect 4494 22554 4522 22583
rect 4102 22135 4103 22161
rect 4129 22135 4130 22161
rect 4102 21854 4130 22135
rect 3822 21826 4130 21854
rect 4382 22526 4494 22554
rect 3598 21770 3626 21775
rect 3374 21769 3626 21770
rect 3374 21743 3599 21769
rect 3625 21743 3626 21769
rect 3374 21742 3626 21743
rect 2422 21737 2450 21742
rect 2238 21574 2370 21579
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2238 21541 2370 21546
rect 2478 21377 2506 21742
rect 2534 21737 2562 21742
rect 2478 21351 2479 21377
rect 2505 21351 2506 21377
rect 2478 21321 2506 21351
rect 2478 21295 2479 21321
rect 2505 21295 2506 21321
rect 2142 20959 2143 20985
rect 2169 20959 2170 20985
rect 2142 20201 2170 20959
rect 2422 20986 2450 20991
rect 2478 20986 2506 21295
rect 2534 20986 2562 20991
rect 2422 20985 2562 20986
rect 2422 20959 2423 20985
rect 2449 20959 2535 20985
rect 2561 20959 2562 20985
rect 2422 20958 2562 20959
rect 2238 20790 2370 20795
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2238 20757 2370 20762
rect 2422 20594 2450 20958
rect 2534 20953 2562 20958
rect 3598 20985 3626 21742
rect 3598 20959 3599 20985
rect 3625 20959 3626 20985
rect 2478 20594 2506 20599
rect 2422 20593 2506 20594
rect 2422 20567 2479 20593
rect 2505 20567 2506 20593
rect 2422 20566 2506 20567
rect 2478 20537 2506 20566
rect 2478 20511 2479 20537
rect 2505 20511 2506 20537
rect 2142 20175 2143 20201
rect 2169 20175 2170 20201
rect 1582 18999 1583 19025
rect 1609 18999 1610 19025
rect 1582 18242 1610 18999
rect 2142 19417 2170 20175
rect 2422 20202 2450 20207
rect 2478 20202 2506 20511
rect 2534 20202 2562 20207
rect 2422 20201 2534 20202
rect 2422 20175 2423 20201
rect 2449 20175 2534 20201
rect 2422 20174 2534 20175
rect 2238 20006 2370 20011
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2238 19973 2370 19978
rect 2422 19810 2450 20174
rect 2534 20136 2562 20174
rect 3598 20201 3626 20959
rect 3598 20175 3599 20201
rect 3625 20175 3626 20201
rect 2478 19810 2506 19815
rect 2422 19809 2506 19810
rect 2422 19783 2479 19809
rect 2505 19783 2506 19809
rect 2422 19782 2506 19783
rect 2478 19753 2506 19782
rect 2478 19727 2479 19753
rect 2505 19727 2506 19753
rect 2142 19391 2143 19417
rect 2169 19391 2170 19417
rect 2142 18633 2170 19391
rect 2422 19418 2450 19423
rect 2478 19418 2506 19727
rect 2534 19418 2562 19423
rect 2422 19417 2562 19418
rect 2422 19391 2423 19417
rect 2449 19391 2535 19417
rect 2561 19391 2562 19417
rect 2422 19390 2562 19391
rect 2422 19385 2450 19390
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2478 19025 2506 19390
rect 2534 19385 2562 19390
rect 3598 19417 3626 20175
rect 3598 19391 3599 19417
rect 3625 19391 3626 19417
rect 2478 18999 2479 19025
rect 2505 18999 2506 19025
rect 2478 18969 2506 18999
rect 2478 18943 2479 18969
rect 2505 18943 2506 18969
rect 2142 18607 2143 18633
rect 2169 18607 2170 18633
rect 2142 18242 2170 18607
rect 2422 18634 2450 18639
rect 2478 18634 2506 18943
rect 2534 18634 2562 18639
rect 2422 18633 2562 18634
rect 2422 18607 2423 18633
rect 2449 18607 2535 18633
rect 2561 18607 2562 18633
rect 2422 18606 2562 18607
rect 2422 18601 2450 18606
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 1582 18241 2170 18242
rect 1582 18215 1583 18241
rect 1609 18215 2170 18241
rect 1582 18214 2170 18215
rect 1582 18209 1610 18214
rect 2142 17850 2170 18214
rect 2142 17803 2170 17822
rect 2478 18241 2506 18606
rect 2534 18601 2562 18606
rect 3598 18633 3626 19391
rect 3598 18607 3599 18633
rect 3625 18607 3626 18633
rect 2478 18215 2479 18241
rect 2505 18215 2506 18241
rect 2478 18185 2506 18215
rect 2478 18159 2479 18185
rect 2505 18159 2506 18185
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 1358 15079 1359 15105
rect 1385 15079 1386 15105
rect 1358 14714 1386 15079
rect 1358 14681 1386 14686
rect 1582 17457 1610 17463
rect 1582 17431 1583 17457
rect 1609 17431 1610 17457
rect 1582 17066 1610 17431
rect 2142 17458 2170 17463
rect 1862 17066 1890 17071
rect 1582 17065 1890 17066
rect 1582 17039 1863 17065
rect 1889 17039 1890 17065
rect 1582 17038 1890 17039
rect 1582 16673 1610 17038
rect 1582 16647 1583 16673
rect 1609 16647 1610 16673
rect 1582 15889 1610 16647
rect 1582 15863 1583 15889
rect 1609 15863 1610 15889
rect 1582 14321 1610 15863
rect 1862 16281 1890 17038
rect 1862 16255 1863 16281
rect 1889 16255 1890 16281
rect 1862 15497 1890 16255
rect 1862 15471 1863 15497
rect 1889 15471 1890 15497
rect 1862 15465 1890 15471
rect 1918 15330 1946 15335
rect 1862 14714 1890 14719
rect 1862 14667 1890 14686
rect 1582 14295 1583 14321
rect 1609 14295 1610 14321
rect 1582 13537 1610 14295
rect 1582 13511 1583 13537
rect 1609 13511 1610 13537
rect 1582 12753 1610 13511
rect 1582 12727 1583 12753
rect 1609 12727 1610 12753
rect 1582 11970 1610 12727
rect 1582 11185 1610 11942
rect 1582 11159 1583 11185
rect 1609 11159 1610 11185
rect 1582 10401 1610 11159
rect 1918 11858 1946 15302
rect 2142 14322 2170 17430
rect 2478 17458 2506 18159
rect 3598 18242 3626 18607
rect 3822 21377 3850 21826
rect 3822 21351 3823 21377
rect 3849 21351 3850 21377
rect 3822 20593 3850 21351
rect 4382 21825 4410 22526
rect 4494 22507 4522 22526
rect 4382 21799 4383 21825
rect 4409 21799 4410 21825
rect 4382 21769 4410 21799
rect 4382 21743 4383 21769
rect 4409 21743 4410 21769
rect 4382 21378 4410 21743
rect 4494 21378 4522 21383
rect 4382 21377 4522 21378
rect 4382 21351 4383 21377
rect 4409 21351 4495 21377
rect 4521 21351 4522 21377
rect 4382 21350 4522 21351
rect 4382 21041 4410 21350
rect 4494 21345 4522 21350
rect 4382 21015 4383 21041
rect 4409 21015 4410 21041
rect 4382 20985 4410 21015
rect 4382 20959 4383 20985
rect 4409 20959 4410 20985
rect 3822 20567 3823 20593
rect 3849 20567 3850 20593
rect 3822 19809 3850 20567
rect 4270 20594 4298 20599
rect 4382 20594 4410 20959
rect 4494 20594 4522 20599
rect 4270 20593 4522 20594
rect 4270 20567 4271 20593
rect 4297 20567 4495 20593
rect 4521 20567 4522 20593
rect 4270 20566 4522 20567
rect 4270 20258 4298 20566
rect 4494 20561 4522 20566
rect 4214 20257 4298 20258
rect 4214 20231 4271 20257
rect 4297 20231 4298 20257
rect 4214 20230 4298 20231
rect 4214 20202 4242 20230
rect 4270 20225 4298 20230
rect 4214 20155 4242 20174
rect 3822 19783 3823 19809
rect 3849 19783 3850 19809
rect 3822 19025 3850 19783
rect 4382 19810 4410 19815
rect 4550 19810 4578 24094
rect 5054 24121 5082 24486
rect 5278 24481 5306 24486
rect 5054 24095 5055 24121
rect 5081 24095 5082 24121
rect 4998 23729 5026 23735
rect 4998 23703 4999 23729
rect 5025 23703 5026 23729
rect 4998 23673 5026 23703
rect 4998 23647 4999 23673
rect 5025 23647 5026 23673
rect 4998 23562 5026 23647
rect 4998 22945 5026 23534
rect 5054 23618 5082 24095
rect 6174 24177 6202 24879
rect 6678 24905 6706 25663
rect 6678 24879 6679 24905
rect 6705 24879 6706 24905
rect 6174 24151 6175 24177
rect 6201 24151 6202 24177
rect 6174 24122 6202 24151
rect 5558 23730 5586 23735
rect 5558 23683 5586 23702
rect 5054 23338 5082 23590
rect 6174 23562 6202 24094
rect 6454 24513 6482 24519
rect 6454 24487 6455 24513
rect 6481 24487 6482 24513
rect 6454 24457 6482 24487
rect 6454 24431 6455 24457
rect 6481 24431 6482 24457
rect 6454 24122 6482 24431
rect 6454 23729 6482 24094
rect 6454 23703 6455 23729
rect 6481 23703 6482 23729
rect 6454 23674 6482 23703
rect 6454 23627 6482 23646
rect 6678 24121 6706 24879
rect 6678 24095 6679 24121
rect 6705 24095 6706 24121
rect 6678 23730 6706 24095
rect 6174 23393 6202 23534
rect 6174 23367 6175 23393
rect 6201 23367 6202 23393
rect 5054 23337 5306 23338
rect 5054 23311 5055 23337
rect 5081 23311 5306 23337
rect 5054 23310 5306 23311
rect 5054 23305 5082 23310
rect 4998 22919 4999 22945
rect 5025 22919 5026 22945
rect 4998 22889 5026 22919
rect 5278 22945 5306 23310
rect 5278 22919 5279 22945
rect 5305 22919 5306 22945
rect 5278 22913 5306 22919
rect 6174 23337 6202 23367
rect 6174 23311 6175 23337
rect 6201 23311 6202 23337
rect 6174 22946 6202 23311
rect 6678 23337 6706 23702
rect 7126 25297 7154 26055
rect 7518 25746 7546 26447
rect 8022 27649 8050 27655
rect 8022 27623 8023 27649
rect 8049 27623 8050 27649
rect 8022 27593 8050 27623
rect 8022 27567 8023 27593
rect 8049 27567 8050 27593
rect 8022 26865 8050 27567
rect 8414 27649 8442 27655
rect 8414 27623 8415 27649
rect 8441 27623 8442 27649
rect 8414 27202 8442 27623
rect 8862 27650 8890 27655
rect 8974 27650 9002 27655
rect 8862 27649 9002 27650
rect 8862 27623 8863 27649
rect 8889 27623 8975 27649
rect 9001 27623 9002 27649
rect 8862 27622 9002 27623
rect 8862 27617 8890 27622
rect 8414 27169 8442 27174
rect 8862 27257 8890 27263
rect 8862 27231 8863 27257
rect 8889 27231 8890 27257
rect 8862 27202 8890 27231
rect 8862 27169 8890 27174
rect 8022 26839 8023 26865
rect 8049 26839 8050 26865
rect 8022 26809 8050 26839
rect 8022 26783 8023 26809
rect 8049 26783 8050 26809
rect 8022 26081 8050 26783
rect 8022 26055 8023 26081
rect 8049 26055 8050 26081
rect 8022 26025 8050 26055
rect 8022 25999 8023 26025
rect 8049 25999 8050 26025
rect 7630 25746 7658 25751
rect 7518 25745 7658 25746
rect 7518 25719 7631 25745
rect 7657 25719 7658 25745
rect 7518 25718 7658 25719
rect 7126 25271 7127 25297
rect 7153 25271 7154 25297
rect 7126 24513 7154 25271
rect 7126 24487 7127 24513
rect 7153 24487 7154 24513
rect 7126 23730 7154 24487
rect 7630 25689 7658 25718
rect 7630 25663 7631 25689
rect 7657 25663 7658 25689
rect 7630 24961 7658 25663
rect 7630 24935 7631 24961
rect 7657 24935 7658 24961
rect 7630 24905 7658 24935
rect 7630 24879 7631 24905
rect 7657 24879 7658 24905
rect 7630 24234 7658 24879
rect 7630 24177 7658 24206
rect 7630 24151 7631 24177
rect 7657 24151 7658 24177
rect 7630 24121 7658 24151
rect 7630 24095 7631 24121
rect 7657 24095 7658 24121
rect 7630 24089 7658 24095
rect 8022 25297 8050 25999
rect 8582 26922 8610 26927
rect 8582 26865 8610 26894
rect 8582 26839 8583 26865
rect 8609 26839 8610 26865
rect 8582 26081 8610 26839
rect 8582 26055 8583 26081
rect 8609 26055 8610 26081
rect 8022 25271 8023 25297
rect 8049 25271 8050 25297
rect 8022 25241 8050 25271
rect 8414 25690 8442 25695
rect 8414 25297 8442 25662
rect 8414 25271 8415 25297
rect 8441 25271 8442 25297
rect 8414 25265 8442 25271
rect 8022 25215 8023 25241
rect 8049 25215 8050 25241
rect 8022 24513 8050 25215
rect 8582 25186 8610 26055
rect 8582 25153 8610 25158
rect 8862 26866 8890 26871
rect 8974 26866 9002 27622
rect 11046 27649 11074 27655
rect 11046 27623 11047 27649
rect 11073 27623 11074 27649
rect 9918 27454 10050 27459
rect 9946 27426 9970 27454
rect 9998 27426 10022 27454
rect 9918 27421 10050 27426
rect 8862 26865 9002 26866
rect 8862 26839 8863 26865
rect 8889 26839 8975 26865
rect 9001 26839 9002 26865
rect 8862 26838 9002 26839
rect 8862 26081 8890 26838
rect 8974 26833 9002 26838
rect 10038 27313 10066 27319
rect 10038 27287 10039 27313
rect 10065 27287 10066 27313
rect 10038 27257 10066 27287
rect 10038 27231 10039 27257
rect 10065 27231 10066 27257
rect 10038 26754 10066 27231
rect 10038 26721 10066 26726
rect 10598 27257 10626 27263
rect 10598 27231 10599 27257
rect 10625 27231 10626 27257
rect 10598 27202 10626 27231
rect 10598 26922 10626 27174
rect 9918 26670 10050 26675
rect 9946 26642 9970 26670
rect 9998 26642 10022 26670
rect 9918 26637 10050 26642
rect 10038 26529 10066 26535
rect 10038 26503 10039 26529
rect 10065 26503 10066 26529
rect 8862 26055 8863 26081
rect 8889 26055 8890 26081
rect 8862 26026 8890 26055
rect 8862 25298 8890 25998
rect 8022 24487 8023 24513
rect 8049 24487 8050 24513
rect 8022 24457 8050 24487
rect 8022 24431 8023 24457
rect 8049 24431 8050 24457
rect 8022 24234 8050 24431
rect 7126 23683 7154 23702
rect 8022 23729 8050 24206
rect 8022 23703 8023 23729
rect 8049 23703 8050 23729
rect 8022 23674 8050 23703
rect 8582 24513 8610 24519
rect 8582 24487 8583 24513
rect 8609 24487 8610 24513
rect 8582 23730 8610 24487
rect 8862 24234 8890 25270
rect 8918 26473 8946 26479
rect 8918 26447 8919 26473
rect 8945 26447 8946 26473
rect 8918 25690 8946 26447
rect 10038 26473 10066 26503
rect 10038 26447 10039 26473
rect 10065 26447 10066 26473
rect 8974 26081 9002 26087
rect 8974 26055 8975 26081
rect 9001 26055 9002 26081
rect 8974 26026 9002 26055
rect 8974 25993 9002 25998
rect 10038 25970 10066 26447
rect 10598 26473 10626 26894
rect 11046 26922 11074 27623
rect 11382 27650 11410 27655
rect 11494 27650 11522 27655
rect 11382 27649 11522 27650
rect 11382 27623 11383 27649
rect 11409 27623 11495 27649
rect 11521 27623 11522 27649
rect 11382 27622 11522 27623
rect 11382 27617 11410 27622
rect 11494 27313 11522 27622
rect 11494 27287 11495 27313
rect 11521 27287 11522 27313
rect 11494 27258 11522 27287
rect 11494 27257 11746 27258
rect 11494 27231 11495 27257
rect 11521 27231 11746 27257
rect 11494 27230 11746 27231
rect 11494 27225 11522 27230
rect 11046 26865 11074 26894
rect 11046 26839 11047 26865
rect 11073 26839 11074 26865
rect 10990 26754 11018 26759
rect 10598 26447 10599 26473
rect 10625 26447 10626 26473
rect 10598 26441 10626 26447
rect 10878 26474 10906 26479
rect 10990 26474 11018 26726
rect 10878 26473 10990 26474
rect 10878 26447 10879 26473
rect 10905 26447 10990 26473
rect 10878 26446 10990 26447
rect 10878 26441 10906 26446
rect 10990 26408 11018 26446
rect 11046 26026 11074 26839
rect 11718 26865 11746 27230
rect 11718 26839 11719 26865
rect 11745 26839 11746 26865
rect 11718 26810 11746 26839
rect 11774 26810 11802 26815
rect 11718 26809 11802 26810
rect 11718 26783 11775 26809
rect 11801 26783 11802 26809
rect 11718 26782 11802 26783
rect 11046 25993 11074 25998
rect 11102 26081 11130 26087
rect 11102 26055 11103 26081
rect 11129 26055 11130 26081
rect 10038 25942 10122 25970
rect 9918 25886 10050 25891
rect 9946 25858 9970 25886
rect 9998 25858 10022 25886
rect 9918 25853 10050 25858
rect 10094 25802 10122 25942
rect 10038 25774 10122 25802
rect 10038 25745 10066 25774
rect 10038 25719 10039 25745
rect 10065 25719 10066 25745
rect 8918 24905 8946 25662
rect 9142 25689 9170 25695
rect 9142 25663 9143 25689
rect 9169 25663 9170 25689
rect 8974 25298 9002 25303
rect 8974 25251 9002 25270
rect 9142 25186 9170 25663
rect 10038 25689 10066 25719
rect 10038 25663 10039 25689
rect 10065 25663 10066 25689
rect 10038 25186 10066 25663
rect 10598 25690 10626 25695
rect 10598 25643 10626 25662
rect 11102 25690 11130 26055
rect 11718 26081 11746 26782
rect 11774 26777 11802 26782
rect 12726 26474 12754 26479
rect 11718 26055 11719 26081
rect 11745 26055 11746 26081
rect 11718 26026 11746 26055
rect 12558 26081 12586 26087
rect 12558 26055 12559 26081
rect 12585 26055 12586 26081
rect 11774 26026 11802 26031
rect 11718 26025 11802 26026
rect 11718 25999 11775 26025
rect 11801 25999 11802 26025
rect 11718 25998 11802 25999
rect 11102 25297 11130 25662
rect 11494 25745 11522 25751
rect 11494 25719 11495 25745
rect 11521 25719 11522 25745
rect 11494 25690 11522 25719
rect 11718 25690 11746 25998
rect 11774 25993 11802 25998
rect 12558 26026 12586 26055
rect 11494 25689 11746 25690
rect 11494 25663 11495 25689
rect 11521 25663 11746 25689
rect 11494 25662 11746 25663
rect 11494 25657 11522 25662
rect 11102 25271 11103 25297
rect 11129 25271 11130 25297
rect 10318 25186 10346 25191
rect 10038 25158 10122 25186
rect 9142 25153 9170 25158
rect 9918 25102 10050 25107
rect 9946 25074 9970 25102
rect 9998 25074 10022 25102
rect 9918 25069 10050 25074
rect 10094 25018 10122 25158
rect 8918 24879 8919 24905
rect 8945 24879 8946 24905
rect 8918 24873 8946 24879
rect 10038 24990 10122 25018
rect 10038 24961 10066 24990
rect 10038 24935 10039 24961
rect 10065 24935 10066 24961
rect 10038 24905 10066 24935
rect 10038 24879 10039 24905
rect 10065 24879 10066 24905
rect 8862 24201 8890 24206
rect 9478 24513 9506 24519
rect 9478 24487 9479 24513
rect 9505 24487 9506 24513
rect 9478 24457 9506 24487
rect 9478 24431 9479 24457
rect 9505 24431 9506 24457
rect 9478 24234 9506 24431
rect 10038 24402 10066 24879
rect 10318 24905 10346 25158
rect 10318 24879 10319 24905
rect 10345 24879 10346 24905
rect 10318 24514 10346 24879
rect 10318 24481 10346 24486
rect 10822 24514 10850 24519
rect 10822 24467 10850 24486
rect 11102 24402 11130 25271
rect 11718 25297 11746 25662
rect 11718 25271 11719 25297
rect 11745 25271 11746 25297
rect 11718 25242 11746 25271
rect 12558 25297 12586 25998
rect 12558 25271 12559 25297
rect 12585 25271 12586 25297
rect 11774 25242 11802 25247
rect 11718 25241 11802 25242
rect 11718 25215 11775 25241
rect 11801 25215 11802 25241
rect 11718 25214 11802 25215
rect 11494 24962 11522 24967
rect 11718 24962 11746 25214
rect 11774 25209 11802 25214
rect 12558 25242 12586 25271
rect 12726 25298 12754 26446
rect 13342 26081 13370 26087
rect 13342 26055 13343 26081
rect 13369 26055 13370 26081
rect 13342 26025 13370 26055
rect 13342 25999 13343 26025
rect 13369 25999 13370 26025
rect 13118 25689 13146 25695
rect 13118 25663 13119 25689
rect 13145 25663 13146 25689
rect 12950 25298 12978 25303
rect 12726 25297 12950 25298
rect 12726 25271 12727 25297
rect 12753 25271 12950 25297
rect 12726 25270 12950 25271
rect 12726 25265 12754 25270
rect 12950 25232 12978 25270
rect 13118 25242 13146 25663
rect 12558 25209 12586 25214
rect 11494 24961 11746 24962
rect 11494 24935 11495 24961
rect 11521 24935 11746 24961
rect 11494 24934 11746 24935
rect 11494 24905 11522 24934
rect 11494 24879 11495 24905
rect 11521 24879 11522 24905
rect 11382 24514 11410 24519
rect 11494 24514 11522 24879
rect 13118 24905 13146 25214
rect 13118 24879 13119 24905
rect 13145 24879 13146 24905
rect 13118 24873 13146 24879
rect 13342 25690 13370 25999
rect 13510 25690 13538 25695
rect 13342 25689 13538 25690
rect 13342 25663 13343 25689
rect 13369 25663 13511 25689
rect 13537 25663 13538 25689
rect 13342 25662 13538 25663
rect 11382 24513 11522 24514
rect 11382 24487 11383 24513
rect 11409 24487 11495 24513
rect 11521 24487 11522 24513
rect 11382 24486 11522 24487
rect 11382 24481 11410 24486
rect 10038 24374 10122 24402
rect 9918 24318 10050 24323
rect 9946 24290 9970 24318
rect 9998 24290 10022 24318
rect 9918 24285 10050 24290
rect 9086 24121 9114 24127
rect 9086 24095 9087 24121
rect 9113 24095 9114 24121
rect 9086 23730 9114 24095
rect 8610 23702 9114 23730
rect 8582 23664 8610 23702
rect 8022 23608 8050 23646
rect 6678 23311 6679 23337
rect 6705 23311 6706 23337
rect 6678 23305 6706 23311
rect 7014 23562 7042 23567
rect 6174 22945 6258 22946
rect 6174 22919 6175 22945
rect 6201 22919 6258 22945
rect 6174 22918 6258 22919
rect 6174 22913 6202 22918
rect 4998 22863 4999 22889
rect 5025 22863 5026 22889
rect 4998 22554 5026 22863
rect 6230 22889 6258 22918
rect 6230 22863 6231 22889
rect 6257 22863 6258 22889
rect 4998 22161 5026 22526
rect 5838 22553 5866 22559
rect 5838 22527 5839 22553
rect 5865 22527 5866 22553
rect 4998 22135 4999 22161
rect 5025 22135 5026 22161
rect 4998 22105 5026 22135
rect 4998 22079 4999 22105
rect 5025 22079 5026 22105
rect 4998 22073 5026 22079
rect 5278 22161 5306 22167
rect 5278 22135 5279 22161
rect 5305 22135 5306 22161
rect 4382 19809 4578 19810
rect 4382 19783 4383 19809
rect 4409 19783 4551 19809
rect 4577 19783 4578 19809
rect 4382 19782 4578 19783
rect 4382 19777 4410 19782
rect 4438 19473 4466 19782
rect 4550 19777 4578 19782
rect 5278 21377 5306 22135
rect 5278 21351 5279 21377
rect 5305 21351 5306 21377
rect 5278 20593 5306 21351
rect 5278 20567 5279 20593
rect 5305 20567 5306 20593
rect 5278 19809 5306 20567
rect 5278 19783 5279 19809
rect 5305 19783 5306 19809
rect 4438 19447 4439 19473
rect 4465 19447 4466 19473
rect 4438 19417 4466 19447
rect 4438 19391 4439 19417
rect 4465 19391 4466 19417
rect 3822 18999 3823 19025
rect 3849 18999 3850 19025
rect 3822 18242 3850 18999
rect 4382 19026 4410 19031
rect 4438 19026 4466 19391
rect 4494 19026 4522 19031
rect 4382 19025 4522 19026
rect 4382 18999 4383 19025
rect 4409 18999 4495 19025
rect 4521 18999 4522 19025
rect 4382 18998 4522 18999
rect 4382 18993 4410 18998
rect 4438 18689 4466 18998
rect 4494 18993 4522 18998
rect 5278 19025 5306 19783
rect 5278 18999 5279 19025
rect 5305 18999 5306 19025
rect 4438 18663 4439 18689
rect 4465 18663 4466 18689
rect 4438 18633 4466 18663
rect 4438 18607 4439 18633
rect 4465 18607 4466 18633
rect 4382 18242 4410 18247
rect 4438 18242 4466 18607
rect 4494 18242 4522 18247
rect 3598 18241 3850 18242
rect 3598 18215 3823 18241
rect 3849 18215 3850 18241
rect 3598 18214 3850 18215
rect 2478 17401 2506 17430
rect 2478 17375 2479 17401
rect 2505 17375 2506 17401
rect 2478 17369 2506 17375
rect 3038 17905 3066 17911
rect 3038 17879 3039 17905
rect 3065 17879 3066 17905
rect 3038 17849 3066 17879
rect 3038 17823 3039 17849
rect 3065 17823 3066 17849
rect 3038 17458 3066 17823
rect 3038 17121 3066 17430
rect 3038 17095 3039 17121
rect 3065 17095 3066 17121
rect 3038 17065 3066 17095
rect 3038 17039 3039 17065
rect 3065 17039 3066 17065
rect 3038 17033 3066 17039
rect 3598 17850 3626 18214
rect 3822 18209 3850 18214
rect 4326 18241 4522 18242
rect 4326 18215 4383 18241
rect 4409 18215 4495 18241
rect 4521 18215 4522 18241
rect 4326 18214 4522 18215
rect 3598 17066 3626 17822
rect 3878 17850 3906 17855
rect 4158 17850 4186 17855
rect 3878 17849 4186 17850
rect 3878 17823 3879 17849
rect 3905 17823 4159 17849
rect 4185 17823 4186 17849
rect 3878 17822 4186 17823
rect 3878 17817 3906 17822
rect 4158 17738 4186 17822
rect 4158 17705 4186 17710
rect 4102 17457 4130 17463
rect 4102 17431 4103 17457
rect 4129 17431 4130 17457
rect 4102 17066 4130 17431
rect 3598 17065 4130 17066
rect 3598 17039 3599 17065
rect 3625 17039 4130 17065
rect 3598 17038 4130 17039
rect 3598 17033 3626 17038
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2478 16673 2506 16679
rect 2478 16647 2479 16673
rect 2505 16647 2506 16673
rect 2478 16617 2506 16647
rect 4102 16674 4130 17038
rect 4102 16627 4130 16646
rect 2478 16591 2479 16617
rect 2505 16591 2506 16617
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2478 15946 2506 16591
rect 2982 16337 3010 16343
rect 2982 16311 2983 16337
rect 3009 16311 3010 16337
rect 2982 16281 3010 16311
rect 4326 16337 4354 18214
rect 4382 18209 4410 18214
rect 4494 18209 4522 18214
rect 5278 18241 5306 18999
rect 5278 18215 5279 18241
rect 5305 18215 5306 18241
rect 5278 17850 5306 18215
rect 5838 21769 5866 22527
rect 6230 22161 6258 22863
rect 6230 22135 6231 22161
rect 6257 22135 6258 22161
rect 6230 22105 6258 22135
rect 6230 22079 6231 22105
rect 6257 22079 6258 22105
rect 6230 21854 6258 22079
rect 7014 22609 7042 23534
rect 7518 23562 7546 23567
rect 7518 23393 7546 23534
rect 7518 23367 7519 23393
rect 7545 23367 7546 23393
rect 7518 23337 7546 23367
rect 7518 23311 7519 23337
rect 7545 23311 7546 23337
rect 7518 23305 7546 23311
rect 9086 23337 9114 23702
rect 9478 23729 9506 24206
rect 10038 24234 10066 24239
rect 10094 24234 10122 24374
rect 10066 24206 10122 24234
rect 10038 24177 10066 24206
rect 10038 24151 10039 24177
rect 10065 24151 10066 24177
rect 10038 24121 10066 24151
rect 10038 24095 10039 24121
rect 10065 24095 10066 24121
rect 10038 24089 10066 24095
rect 10598 24122 10626 24127
rect 10598 24075 10626 24094
rect 11102 24122 11130 24374
rect 9478 23703 9479 23729
rect 9505 23703 9506 23729
rect 9478 23673 9506 23703
rect 11102 23729 11130 24094
rect 11102 23703 11103 23729
rect 11129 23703 11130 23729
rect 11102 23697 11130 23703
rect 11494 24177 11522 24486
rect 11494 24151 11495 24177
rect 11521 24151 11522 24177
rect 11494 24121 11522 24151
rect 11494 24095 11495 24121
rect 11521 24095 11522 24121
rect 11494 23730 11522 24095
rect 12278 24514 12306 24519
rect 11494 23697 11522 23702
rect 11718 23730 11746 23735
rect 9478 23647 9479 23673
rect 9505 23647 9506 23673
rect 9478 23641 9506 23647
rect 11718 23674 11746 23702
rect 12278 23729 12306 24486
rect 12558 24513 12586 24519
rect 12558 24487 12559 24513
rect 12585 24487 12586 24513
rect 12558 24402 12586 24487
rect 13342 24513 13370 25662
rect 13510 25657 13538 25662
rect 13510 25298 13538 25303
rect 13398 24906 13426 24911
rect 13510 24906 13538 25270
rect 13398 24905 13538 24906
rect 13398 24879 13399 24905
rect 13425 24879 13511 24905
rect 13537 24879 13538 24905
rect 13398 24878 13538 24879
rect 13398 24873 13426 24878
rect 13342 24487 13343 24513
rect 13369 24487 13370 24513
rect 13342 24457 13370 24487
rect 13342 24431 13343 24457
rect 13369 24431 13370 24457
rect 12558 24369 12586 24374
rect 13118 24402 13146 24407
rect 13118 24121 13146 24374
rect 13118 24095 13119 24121
rect 13145 24095 13146 24121
rect 13118 24089 13146 24095
rect 13342 24346 13370 24431
rect 13342 24122 13370 24318
rect 13510 24234 13538 24878
rect 13510 24201 13538 24206
rect 13510 24122 13538 24127
rect 13342 24121 13538 24122
rect 13342 24095 13343 24121
rect 13369 24095 13511 24121
rect 13537 24095 13538 24121
rect 13342 24094 13538 24095
rect 13342 24089 13370 24094
rect 12278 23703 12279 23729
rect 12305 23703 12306 23729
rect 11774 23674 11802 23679
rect 11718 23673 11802 23674
rect 11718 23647 11775 23673
rect 11801 23647 11802 23673
rect 11718 23646 11802 23647
rect 11774 23641 11802 23646
rect 10990 23618 11018 23623
rect 9086 23311 9087 23337
rect 9113 23311 9114 23337
rect 7014 22583 7015 22609
rect 7041 22583 7042 22609
rect 7014 22553 7042 22583
rect 8134 22945 8162 22951
rect 8134 22919 8135 22945
rect 8161 22919 8162 22945
rect 7014 22527 7015 22553
rect 7041 22527 7042 22553
rect 7014 21854 7042 22527
rect 7574 22554 7602 22559
rect 7574 22507 7602 22526
rect 8134 22554 8162 22919
rect 9030 22945 9058 22951
rect 9030 22919 9031 22945
rect 9057 22919 9058 22945
rect 9030 22889 9058 22919
rect 9030 22863 9031 22889
rect 9057 22863 9058 22889
rect 8134 22161 8162 22526
rect 8134 22135 8135 22161
rect 8161 22135 8162 22161
rect 6230 21826 6426 21854
rect 5838 21743 5839 21769
rect 5865 21743 5866 21769
rect 5838 20985 5866 21743
rect 6398 21770 6426 21826
rect 6510 21826 7042 21854
rect 7294 21882 7322 21887
rect 6510 21770 6538 21826
rect 6398 21769 6538 21770
rect 6398 21743 6399 21769
rect 6425 21743 6511 21769
rect 6537 21743 6538 21769
rect 6398 21742 6538 21743
rect 6398 21377 6426 21742
rect 6510 21737 6538 21742
rect 7294 21769 7322 21854
rect 7294 21743 7295 21769
rect 7321 21743 7322 21769
rect 6398 21351 6399 21377
rect 6425 21351 6426 21377
rect 6398 21321 6426 21351
rect 6398 21295 6399 21321
rect 6425 21295 6426 21321
rect 6398 21289 6426 21295
rect 5838 20959 5839 20985
rect 5865 20959 5866 20985
rect 5838 20201 5866 20959
rect 7014 21041 7042 21047
rect 7014 21015 7015 21041
rect 7041 21015 7042 21041
rect 7014 20985 7042 21015
rect 7014 20959 7015 20985
rect 7041 20959 7042 20985
rect 5838 20175 5839 20201
rect 5865 20175 5866 20201
rect 5838 19417 5866 20175
rect 5838 19391 5839 19417
rect 5865 19391 5866 19417
rect 5838 18633 5866 19391
rect 5838 18607 5839 18633
rect 5865 18607 5866 18633
rect 5838 18522 5866 18607
rect 5838 17850 5866 18494
rect 5278 17849 5866 17850
rect 5278 17823 5839 17849
rect 5865 17823 5866 17849
rect 5278 17822 5866 17823
rect 4382 17458 4410 17463
rect 4494 17458 4522 17463
rect 4410 17457 4522 17458
rect 4410 17431 4495 17457
rect 4521 17431 4522 17457
rect 4410 17430 4522 17431
rect 4382 17392 4410 17430
rect 4438 17121 4466 17430
rect 4494 17425 4522 17430
rect 5278 17457 5306 17822
rect 5838 17817 5866 17822
rect 6454 20593 6482 20599
rect 6454 20567 6455 20593
rect 6481 20567 6482 20593
rect 6454 20537 6482 20567
rect 6454 20511 6455 20537
rect 6481 20511 6482 20537
rect 6454 19809 6482 20511
rect 6454 19783 6455 19809
rect 6481 19783 6482 19809
rect 6454 19753 6482 19783
rect 6454 19727 6455 19753
rect 6481 19727 6482 19753
rect 6454 19025 6482 19727
rect 6454 18999 6455 19025
rect 6481 18999 6482 19025
rect 6454 18969 6482 18999
rect 6454 18943 6455 18969
rect 6481 18943 6482 18969
rect 6454 18241 6482 18943
rect 6454 18215 6455 18241
rect 6481 18215 6482 18241
rect 6454 18185 6482 18215
rect 6454 18159 6455 18185
rect 6481 18159 6482 18185
rect 5278 17431 5279 17457
rect 5305 17431 5306 17457
rect 4438 17095 4439 17121
rect 4465 17095 4466 17121
rect 4438 17065 4466 17095
rect 4438 17039 4439 17065
rect 4465 17039 4466 17065
rect 4382 16674 4410 16679
rect 4438 16674 4466 17039
rect 4550 16674 4578 16679
rect 4382 16673 4578 16674
rect 4382 16647 4383 16673
rect 4409 16647 4551 16673
rect 4577 16647 4578 16673
rect 4382 16646 4578 16647
rect 4382 16641 4410 16646
rect 4326 16311 4327 16337
rect 4353 16311 4354 16337
rect 2982 16255 2983 16281
rect 3009 16255 3010 16281
rect 2982 15974 3010 16255
rect 3598 16281 3626 16287
rect 3598 16255 3599 16281
rect 3625 16255 3626 16281
rect 2982 15946 3066 15974
rect 2422 15890 2450 15895
rect 2478 15890 2506 15918
rect 3038 15913 3066 15918
rect 2422 15889 2506 15890
rect 2422 15863 2423 15889
rect 2449 15863 2506 15889
rect 2422 15862 2506 15863
rect 2422 15833 2450 15862
rect 2422 15807 2423 15833
rect 2449 15807 2450 15833
rect 2422 15498 2450 15807
rect 2534 15498 2562 15503
rect 2422 15497 2562 15498
rect 2422 15471 2423 15497
rect 2449 15471 2535 15497
rect 2561 15471 2562 15497
rect 2422 15470 2562 15471
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2422 15162 2450 15470
rect 2534 15465 2562 15470
rect 3598 15498 3626 16255
rect 4326 16281 4354 16311
rect 4326 16255 4327 16281
rect 4353 16255 4354 16281
rect 4326 15974 4354 16255
rect 4326 15946 4410 15974
rect 3822 15889 3850 15895
rect 3822 15863 3823 15889
rect 3849 15863 3850 15889
rect 3822 15498 3850 15863
rect 4382 15554 4410 15946
rect 4550 15946 4578 16646
rect 5278 16674 5306 17431
rect 6454 17682 6482 18159
rect 6454 17457 6482 17654
rect 6454 17431 6455 17457
rect 6481 17431 6482 17457
rect 6454 17401 6482 17431
rect 6454 17375 6455 17401
rect 6481 17375 6482 17401
rect 6454 17369 6482 17375
rect 7014 20257 7042 20959
rect 7014 20231 7015 20257
rect 7041 20231 7042 20257
rect 7014 20201 7042 20231
rect 7014 20175 7015 20201
rect 7041 20175 7042 20201
rect 7014 19473 7042 20175
rect 7014 19447 7015 19473
rect 7041 19447 7042 19473
rect 7014 19417 7042 19447
rect 7014 19391 7015 19417
rect 7041 19391 7042 19417
rect 7014 18689 7042 19391
rect 7014 18663 7015 18689
rect 7041 18663 7042 18689
rect 7014 18633 7042 18663
rect 7014 18607 7015 18633
rect 7041 18607 7042 18633
rect 7014 17905 7042 18607
rect 7014 17879 7015 17905
rect 7041 17879 7042 17905
rect 7014 17849 7042 17879
rect 7014 17823 7015 17849
rect 7041 17823 7042 17849
rect 7014 17682 7042 17823
rect 7294 20985 7322 21743
rect 7294 20959 7295 20985
rect 7321 20959 7322 20985
rect 7294 20201 7322 20959
rect 7294 20175 7295 20201
rect 7321 20175 7322 20201
rect 7294 19417 7322 20175
rect 7294 19391 7295 19417
rect 7321 19391 7322 19417
rect 7294 18633 7322 19391
rect 7294 18607 7295 18633
rect 7321 18607 7322 18633
rect 7294 18522 7322 18607
rect 7294 17849 7322 18494
rect 7294 17823 7295 17849
rect 7321 17823 7322 17849
rect 7294 17817 7322 17823
rect 8134 21882 8162 22135
rect 8134 21377 8162 21854
rect 8134 21351 8135 21377
rect 8161 21351 8162 21377
rect 8134 20593 8162 21351
rect 8134 20567 8135 20593
rect 8161 20567 8162 20593
rect 8134 19809 8162 20567
rect 8134 19783 8135 19809
rect 8161 19783 8162 19809
rect 8134 19025 8162 19783
rect 8246 22609 8274 22615
rect 8246 22583 8247 22609
rect 8273 22583 8274 22609
rect 8246 22553 8274 22583
rect 8246 22527 8247 22553
rect 8273 22527 8274 22553
rect 8246 21825 8274 22527
rect 8246 21799 8247 21825
rect 8273 21799 8274 21825
rect 8246 21769 8274 21799
rect 8246 21743 8247 21769
rect 8273 21743 8274 21769
rect 8246 21041 8274 21743
rect 8246 21015 8247 21041
rect 8273 21015 8274 21041
rect 8246 20985 8274 21015
rect 8246 20959 8247 20985
rect 8273 20959 8274 20985
rect 8246 20257 8274 20959
rect 8246 20231 8247 20257
rect 8273 20231 8274 20257
rect 8246 20201 8274 20231
rect 8246 20175 8247 20201
rect 8273 20175 8274 20201
rect 8246 19473 8274 20175
rect 8246 19447 8247 19473
rect 8273 19447 8274 19473
rect 8246 19417 8274 19447
rect 8246 19391 8247 19417
rect 8273 19391 8274 19417
rect 8246 19334 8274 19391
rect 9030 22161 9058 22863
rect 9030 22135 9031 22161
rect 9057 22135 9058 22161
rect 9030 22105 9058 22135
rect 9030 22079 9031 22105
rect 9057 22079 9058 22105
rect 9030 21770 9058 22079
rect 9030 21377 9058 21742
rect 9030 21351 9031 21377
rect 9057 21351 9058 21377
rect 9030 21321 9058 21351
rect 9030 21295 9031 21321
rect 9057 21295 9058 21321
rect 9030 20593 9058 21295
rect 9086 22553 9114 23311
rect 9310 23562 9338 23567
rect 9310 23338 9338 23534
rect 9918 23534 10050 23539
rect 9946 23506 9970 23534
rect 9998 23506 10022 23534
rect 9918 23501 10050 23506
rect 9534 23338 9562 23343
rect 9310 23337 9562 23338
rect 9310 23311 9311 23337
rect 9337 23311 9535 23337
rect 9561 23311 9562 23337
rect 9310 23310 9562 23311
rect 9310 23305 9338 23310
rect 9534 23305 9562 23310
rect 10318 23337 10346 23343
rect 10318 23311 10319 23337
rect 10345 23311 10346 23337
rect 9918 22750 10050 22755
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 9918 22717 10050 22722
rect 9086 22527 9087 22553
rect 9113 22527 9114 22553
rect 9086 21769 9114 22527
rect 9086 21743 9087 21769
rect 9113 21743 9114 21769
rect 9086 20986 9114 21743
rect 9310 22554 9338 22559
rect 9534 22554 9562 22559
rect 9310 22553 9562 22554
rect 9310 22527 9311 22553
rect 9337 22527 9535 22553
rect 9561 22527 9562 22553
rect 9310 22526 9562 22527
rect 9310 21770 9338 22526
rect 9534 22521 9562 22526
rect 10318 22553 10346 23311
rect 10878 23338 10906 23343
rect 10990 23338 11018 23590
rect 10878 23337 11018 23338
rect 10878 23311 10879 23337
rect 10905 23311 10991 23337
rect 11017 23311 11018 23337
rect 10878 23310 11018 23311
rect 10878 23305 10906 23310
rect 10990 23305 11018 23310
rect 11270 23618 11298 23623
rect 10318 22527 10319 22553
rect 10345 22527 10346 22553
rect 9918 21966 10050 21971
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 9918 21933 10050 21938
rect 9310 21723 9338 21742
rect 9534 21770 9562 21775
rect 9534 21723 9562 21742
rect 10318 21769 10346 22527
rect 10318 21743 10319 21769
rect 10345 21743 10346 21769
rect 9918 21182 10050 21187
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 9918 21149 10050 21154
rect 9814 21041 9842 21047
rect 9814 21015 9815 21041
rect 9841 21015 9842 21041
rect 9142 20986 9170 20991
rect 9086 20985 9170 20986
rect 9086 20959 9143 20985
rect 9169 20959 9170 20985
rect 9086 20958 9170 20959
rect 9030 20567 9031 20593
rect 9057 20567 9058 20593
rect 9030 20537 9058 20567
rect 9030 20511 9031 20537
rect 9057 20511 9058 20537
rect 9030 19809 9058 20511
rect 9030 19783 9031 19809
rect 9057 19783 9058 19809
rect 9030 19753 9058 19783
rect 9030 19727 9031 19753
rect 9057 19727 9058 19753
rect 8246 19306 8442 19334
rect 8134 18999 8135 19025
rect 8161 18999 8162 19025
rect 8134 18241 8162 18999
rect 8134 18215 8135 18241
rect 8161 18215 8162 18241
rect 7014 17121 7042 17654
rect 7014 17095 7015 17121
rect 7041 17095 7042 17121
rect 5838 17065 5866 17071
rect 5838 17039 5839 17065
rect 5865 17039 5866 17065
rect 5278 16627 5306 16646
rect 5558 16674 5586 16679
rect 4550 15913 4578 15918
rect 4942 15889 4970 15895
rect 4942 15863 4943 15889
rect 4969 15863 4970 15889
rect 4942 15833 4970 15863
rect 5558 15890 5586 16646
rect 5558 15843 5586 15862
rect 5838 16281 5866 17039
rect 7014 17065 7042 17095
rect 8134 17457 8162 18215
rect 8134 17431 8135 17457
rect 8161 17431 8162 17457
rect 7014 17039 7015 17065
rect 7041 17039 7042 17065
rect 5838 16255 5839 16281
rect 5865 16255 5866 16281
rect 5838 15890 5866 16255
rect 6454 16673 6482 16679
rect 6454 16647 6455 16673
rect 6481 16647 6482 16673
rect 6454 16617 6482 16647
rect 6454 16591 6455 16617
rect 6481 16591 6482 16617
rect 4942 15807 4943 15833
rect 4969 15807 4970 15833
rect 4494 15554 4522 15559
rect 4382 15553 4522 15554
rect 4382 15527 4495 15553
rect 4521 15527 4522 15553
rect 4382 15526 4522 15527
rect 3598 15497 3850 15498
rect 3598 15471 3599 15497
rect 3625 15471 3850 15497
rect 3598 15470 3850 15471
rect 2366 15106 2394 15111
rect 2422 15106 2450 15134
rect 2366 15105 2450 15106
rect 2366 15079 2367 15105
rect 2393 15079 2450 15105
rect 2366 15078 2450 15079
rect 2366 15049 2394 15078
rect 2366 15023 2367 15049
rect 2393 15023 2394 15049
rect 2366 14713 2394 15023
rect 2366 14687 2367 14713
rect 2393 14687 2394 14713
rect 2366 14602 2394 14687
rect 2590 14713 2618 14719
rect 2590 14687 2591 14713
rect 2617 14687 2618 14713
rect 2590 14602 2618 14687
rect 2366 14574 2618 14602
rect 3374 14714 3402 14719
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2142 14321 2282 14322
rect 2142 14295 2143 14321
rect 2169 14295 2282 14321
rect 2142 14294 2282 14295
rect 2142 14289 2170 14294
rect 2254 14266 2282 14294
rect 2254 14265 2338 14266
rect 2254 14239 2255 14265
rect 2281 14239 2338 14265
rect 2254 14238 2338 14239
rect 2254 14233 2282 14238
rect 1582 10375 1583 10401
rect 1609 10375 1610 10401
rect 1582 10122 1610 10375
rect 1358 10066 1610 10094
rect 1694 10962 1722 10967
rect 1358 9617 1386 10066
rect 1358 9591 1359 9617
rect 1385 9591 1386 9617
rect 1358 8833 1386 9591
rect 1358 8807 1359 8833
rect 1385 8807 1386 8833
rect 1358 8049 1386 8807
rect 1358 8023 1359 8049
rect 1385 8023 1386 8049
rect 1358 7265 1386 8023
rect 1358 7239 1359 7265
rect 1385 7239 1386 7265
rect 1358 7233 1386 7239
rect 1022 6594 1050 6599
rect 1022 4522 1050 6566
rect 1582 6482 1610 6487
rect 1582 6435 1610 6454
rect 1022 4129 1050 4494
rect 1190 6090 1218 6095
rect 1190 5697 1218 6062
rect 1694 6090 1722 10934
rect 1862 10122 1890 10127
rect 1862 10010 1890 10094
rect 1862 9977 1890 9982
rect 1918 6873 1946 11830
rect 2142 13929 2170 13935
rect 2142 13903 2143 13929
rect 2169 13903 2170 13929
rect 2142 13145 2170 13903
rect 2310 13930 2338 14238
rect 2310 13864 2338 13902
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2422 13650 2450 14574
rect 2142 13119 2143 13145
rect 2169 13119 2170 13145
rect 2142 12361 2170 13119
rect 2366 13622 2450 13650
rect 2534 13930 2562 13935
rect 2366 13034 2394 13622
rect 2478 13538 2506 13543
rect 2534 13538 2562 13902
rect 2478 13537 2562 13538
rect 2478 13511 2479 13537
rect 2505 13511 2562 13537
rect 2478 13510 2562 13511
rect 2478 13481 2506 13510
rect 2478 13455 2479 13481
rect 2505 13455 2506 13481
rect 2478 13449 2506 13455
rect 2422 13146 2450 13151
rect 2534 13146 2562 13510
rect 2422 13145 2562 13146
rect 2422 13119 2423 13145
rect 2449 13119 2535 13145
rect 2561 13119 2562 13145
rect 2422 13118 2562 13119
rect 2422 13113 2450 13118
rect 2366 13006 2450 13034
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12335 2143 12361
rect 2169 12335 2170 12361
rect 2142 11970 2170 12335
rect 2366 12754 2394 12759
rect 2422 12754 2450 13006
rect 2366 12753 2450 12754
rect 2366 12727 2367 12753
rect 2393 12727 2450 12753
rect 2366 12726 2450 12727
rect 2366 12697 2394 12726
rect 2366 12671 2367 12697
rect 2393 12671 2394 12697
rect 2366 12250 2394 12671
rect 2422 12362 2450 12367
rect 2534 12362 2562 13118
rect 3374 13929 3402 14686
rect 3598 14713 3626 15470
rect 3598 14687 3599 14713
rect 3625 14687 3626 14713
rect 3598 14681 3626 14687
rect 3822 15105 3850 15470
rect 3822 15079 3823 15105
rect 3849 15079 3850 15105
rect 3374 13903 3375 13929
rect 3401 13903 3402 13929
rect 3374 13145 3402 13903
rect 3822 14321 3850 15079
rect 3822 14295 3823 14321
rect 3849 14295 3850 14321
rect 3822 14266 3850 14295
rect 3822 13538 3850 14238
rect 3374 13119 3375 13145
rect 3401 13119 3402 13145
rect 3374 12586 3402 13119
rect 3374 12553 3402 12558
rect 3598 13537 3850 13538
rect 3598 13511 3823 13537
rect 3849 13511 3850 13537
rect 3598 13510 3850 13511
rect 2422 12361 2534 12362
rect 2422 12335 2423 12361
rect 2449 12335 2534 12361
rect 2422 12334 2534 12335
rect 2422 12329 2450 12334
rect 2534 12296 2562 12334
rect 3598 12361 3626 13510
rect 3822 13505 3850 13510
rect 4494 15497 4522 15526
rect 4494 15471 4495 15497
rect 4521 15471 4522 15497
rect 4494 15162 4522 15471
rect 4494 14769 4522 15134
rect 4494 14743 4495 14769
rect 4521 14743 4522 14769
rect 4494 14713 4522 14743
rect 4494 14687 4495 14713
rect 4521 14687 4522 14713
rect 4494 13985 4522 14687
rect 4942 15105 4970 15807
rect 5838 15498 5866 15862
rect 5950 15946 5978 15951
rect 5950 15889 5978 15918
rect 5950 15863 5951 15889
rect 5977 15863 5978 15889
rect 5950 15857 5978 15863
rect 6230 15946 6258 15951
rect 6230 15834 6258 15918
rect 6454 15946 6482 16591
rect 7014 16337 7042 17039
rect 7014 16311 7015 16337
rect 7041 16311 7042 16337
rect 6734 16282 6762 16287
rect 6734 15974 6762 16254
rect 7014 16282 7042 16311
rect 7014 16235 7042 16254
rect 7294 17065 7322 17071
rect 7294 17039 7295 17065
rect 7321 17039 7322 17065
rect 7294 16281 7322 17039
rect 8134 17066 8162 17431
rect 8134 16674 8162 17038
rect 7294 16255 7295 16281
rect 7321 16255 7322 16281
rect 6230 15833 6314 15834
rect 6230 15807 6231 15833
rect 6257 15807 6314 15833
rect 6230 15806 6314 15807
rect 6230 15801 6258 15806
rect 5838 15465 5866 15470
rect 6118 15498 6146 15503
rect 6118 15451 6146 15470
rect 6286 15497 6314 15806
rect 6286 15471 6287 15497
rect 6313 15471 6314 15497
rect 6286 15465 6314 15471
rect 6454 15498 6482 15918
rect 6622 15946 6762 15974
rect 6510 15498 6538 15503
rect 6454 15497 6538 15498
rect 6454 15471 6511 15497
rect 6537 15471 6538 15497
rect 6454 15470 6538 15471
rect 6510 15162 6538 15470
rect 6510 15129 6538 15134
rect 4942 15079 4943 15105
rect 4969 15079 4970 15105
rect 4942 15049 4970 15079
rect 4942 15023 4943 15049
rect 4969 15023 4970 15049
rect 4942 14322 4970 15023
rect 5278 15105 5306 15111
rect 5278 15079 5279 15105
rect 5305 15079 5306 15105
rect 5278 14713 5306 15079
rect 6454 15105 6482 15111
rect 6454 15079 6455 15105
rect 6481 15079 6482 15105
rect 6454 15050 6482 15079
rect 6622 15050 6650 15946
rect 5278 14687 5279 14713
rect 5305 14687 5306 14713
rect 4998 14322 5026 14327
rect 4942 14321 5026 14322
rect 4942 14295 4999 14321
rect 5025 14295 5026 14321
rect 4942 14294 5026 14295
rect 4494 13959 4495 13985
rect 4521 13959 4522 13985
rect 4494 13929 4522 13959
rect 4494 13903 4495 13929
rect 4521 13903 4522 13929
rect 4494 13201 4522 13903
rect 4494 13175 4495 13201
rect 4521 13175 4522 13201
rect 4494 13146 4522 13175
rect 4494 13099 4522 13118
rect 4998 14265 5026 14294
rect 4998 14239 4999 14265
rect 5025 14239 5026 14265
rect 4998 13537 5026 14239
rect 5278 14266 5306 14687
rect 6174 15049 6650 15050
rect 6174 15023 6455 15049
rect 6481 15023 6650 15049
rect 6174 15022 6650 15023
rect 6846 15498 6874 15503
rect 7294 15498 7322 16255
rect 6874 15497 7322 15498
rect 6874 15471 7295 15497
rect 7321 15471 7322 15497
rect 6874 15470 7322 15471
rect 6174 14769 6202 15022
rect 6454 15017 6482 15022
rect 6174 14743 6175 14769
rect 6201 14743 6202 14769
rect 6174 14713 6202 14743
rect 6174 14687 6175 14713
rect 6201 14687 6202 14713
rect 5278 14233 5306 14238
rect 5558 14321 5586 14327
rect 5558 14295 5559 14321
rect 5585 14295 5586 14321
rect 5558 14266 5586 14295
rect 6174 14322 6202 14687
rect 6734 14714 6762 14719
rect 6846 14714 6874 15470
rect 7294 15465 7322 15470
rect 7910 16673 8162 16674
rect 7910 16647 8135 16673
rect 8161 16647 8162 16673
rect 7910 16646 8162 16647
rect 7910 15889 7938 16646
rect 8134 16641 8162 16646
rect 8414 18689 8442 19306
rect 8414 18663 8415 18689
rect 8441 18663 8442 18689
rect 8414 18633 8442 18663
rect 8414 18607 8415 18633
rect 8441 18607 8442 18633
rect 8414 17905 8442 18607
rect 9030 19025 9058 19727
rect 9030 18999 9031 19025
rect 9057 18999 9058 19025
rect 9030 18969 9058 18999
rect 9030 18943 9031 18969
rect 9057 18943 9058 18969
rect 9030 18241 9058 18943
rect 9030 18215 9031 18241
rect 9057 18215 9058 18241
rect 9030 18186 9058 18215
rect 9030 18139 9058 18158
rect 9142 20201 9170 20958
rect 9142 20175 9143 20201
rect 9169 20175 9170 20201
rect 9142 19417 9170 20175
rect 9142 19391 9143 19417
rect 9169 19391 9170 19417
rect 9142 18633 9170 19391
rect 9814 20985 9842 21015
rect 9814 20959 9815 20985
rect 9841 20959 9842 20985
rect 9814 20257 9842 20959
rect 10318 20985 10346 21743
rect 10318 20959 10319 20985
rect 10345 20959 10346 20985
rect 9918 20398 10050 20403
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 9918 20365 10050 20370
rect 9814 20231 9815 20257
rect 9841 20231 9842 20257
rect 9814 20201 9842 20231
rect 9814 20175 9815 20201
rect 9841 20175 9842 20201
rect 9814 19473 9842 20175
rect 10318 20201 10346 20959
rect 10318 20175 10319 20201
rect 10345 20175 10346 20201
rect 9918 19614 10050 19619
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 9918 19581 10050 19586
rect 9814 19447 9815 19473
rect 9841 19447 9842 19473
rect 9814 19417 9842 19447
rect 9814 19391 9815 19417
rect 9841 19391 9842 19417
rect 9814 19334 9842 19391
rect 10318 19417 10346 20175
rect 10318 19391 10319 19417
rect 10345 19391 10346 19417
rect 9814 19306 10066 19334
rect 10038 18914 10066 19306
rect 10038 18886 10122 18914
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10094 18746 10122 18886
rect 9142 18607 9143 18633
rect 9169 18607 9170 18633
rect 8414 17879 8415 17905
rect 8441 17879 8442 17905
rect 8414 17849 8442 17879
rect 8414 17823 8415 17849
rect 8441 17823 8442 17849
rect 8414 17458 8442 17823
rect 9142 17849 9170 18607
rect 10038 18718 10122 18746
rect 10038 18689 10066 18718
rect 10038 18663 10039 18689
rect 10065 18663 10066 18689
rect 10038 18633 10066 18663
rect 10038 18607 10039 18633
rect 10065 18607 10066 18633
rect 9142 17823 9143 17849
rect 9169 17823 9170 17849
rect 8526 17458 8554 17463
rect 8414 17457 8554 17458
rect 8414 17431 8415 17457
rect 8441 17431 8527 17457
rect 8553 17431 8554 17457
rect 8414 17430 8554 17431
rect 8414 17121 8442 17430
rect 8526 17425 8554 17430
rect 8414 17095 8415 17121
rect 8441 17095 8442 17121
rect 8414 17065 8442 17095
rect 8414 17039 8415 17065
rect 8441 17039 8442 17065
rect 8414 16674 8442 17039
rect 9142 17066 9170 17823
rect 8526 16674 8554 16679
rect 8414 16673 8554 16674
rect 8414 16647 8415 16673
rect 8441 16647 8527 16673
rect 8553 16647 8554 16673
rect 8414 16646 8554 16647
rect 8414 16337 8442 16646
rect 8526 16641 8554 16646
rect 8414 16311 8415 16337
rect 8441 16311 8442 16337
rect 7910 15863 7911 15889
rect 7937 15863 7938 15889
rect 6734 14713 6874 14714
rect 6734 14687 6735 14713
rect 6761 14687 6874 14713
rect 6734 14686 6874 14687
rect 6734 14681 6762 14686
rect 6174 14321 6258 14322
rect 6174 14295 6175 14321
rect 6201 14295 6258 14321
rect 6174 14294 6258 14295
rect 6174 14289 6202 14294
rect 5558 13930 5586 14238
rect 6230 14265 6258 14294
rect 6846 14321 6874 14686
rect 6902 15162 6930 15167
rect 6902 14714 6930 15134
rect 7910 15105 7938 15863
rect 8302 16282 8330 16287
rect 8414 16282 8442 16311
rect 8330 16281 8442 16282
rect 8330 16255 8415 16281
rect 8441 16255 8442 16281
rect 8330 16254 8442 16255
rect 8302 15554 8330 16254
rect 8414 16249 8442 16254
rect 9142 16281 9170 17038
rect 9142 16255 9143 16281
rect 9169 16255 9170 16281
rect 9142 15974 9170 16255
rect 9814 18186 9842 18191
rect 9814 17962 9842 18158
rect 10038 18130 10066 18607
rect 10318 18633 10346 19391
rect 10318 18607 10319 18633
rect 10345 18607 10346 18633
rect 10038 18102 10122 18130
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 10094 17962 10122 18102
rect 9814 17934 10122 17962
rect 9814 17905 9842 17934
rect 9814 17879 9815 17905
rect 9841 17879 9842 17905
rect 9814 17849 9842 17879
rect 9814 17823 9815 17849
rect 9841 17823 9842 17849
rect 9814 17121 9842 17823
rect 10038 17850 10066 17934
rect 10038 17817 10066 17822
rect 10318 17849 10346 18607
rect 10318 17823 10319 17849
rect 10345 17823 10346 17849
rect 10318 17458 10346 17823
rect 10822 22945 10850 22951
rect 10822 22919 10823 22945
rect 10849 22919 10850 22945
rect 10822 22161 10850 22919
rect 10822 22135 10823 22161
rect 10849 22135 10850 22161
rect 10822 21377 10850 22135
rect 10822 21351 10823 21377
rect 10849 21351 10850 21377
rect 10822 20593 10850 21351
rect 11270 22946 11298 23590
rect 12278 23338 12306 23703
rect 13454 23730 13482 24094
rect 13510 24089 13538 24094
rect 13454 23673 13482 23702
rect 13454 23647 13455 23673
rect 13481 23647 13482 23673
rect 11494 22946 11522 22951
rect 11270 22945 11522 22946
rect 11270 22919 11271 22945
rect 11297 22919 11495 22945
rect 11521 22919 11522 22945
rect 11270 22918 11522 22919
rect 11270 22609 11298 22918
rect 11494 22913 11522 22918
rect 12278 22945 12306 23310
rect 12278 22919 12279 22945
rect 12305 22919 12306 22945
rect 11270 22583 11271 22609
rect 11297 22583 11298 22609
rect 11270 22553 11298 22583
rect 11270 22527 11271 22553
rect 11297 22527 11298 22553
rect 11270 22162 11298 22527
rect 11494 22162 11522 22167
rect 11270 22161 11522 22162
rect 11270 22135 11271 22161
rect 11297 22135 11495 22161
rect 11521 22135 11522 22161
rect 11270 22134 11522 22135
rect 11270 21825 11298 22134
rect 11494 22129 11522 22134
rect 12278 22161 12306 22919
rect 12278 22135 12279 22161
rect 12305 22135 12306 22161
rect 12278 22129 12306 22135
rect 12838 23338 12866 23343
rect 12838 22553 12866 23310
rect 13454 22946 13482 23647
rect 13958 23393 13986 23399
rect 13958 23367 13959 23393
rect 13985 23367 13986 23393
rect 13958 23337 13986 23367
rect 13958 23311 13959 23337
rect 13985 23311 13986 23337
rect 13958 22946 13986 23311
rect 13454 22945 13986 22946
rect 13454 22919 13455 22945
rect 13481 22919 13986 22945
rect 13454 22918 13986 22919
rect 13454 22889 13482 22918
rect 13454 22863 13455 22889
rect 13481 22863 13482 22889
rect 13454 22857 13482 22863
rect 12838 22527 12839 22553
rect 12865 22527 12866 22553
rect 11270 21799 11271 21825
rect 11297 21799 11298 21825
rect 11270 21769 11298 21799
rect 11270 21743 11271 21769
rect 11297 21743 11298 21769
rect 11270 21378 11298 21743
rect 12838 21770 12866 22527
rect 13958 22609 13986 22918
rect 13958 22583 13959 22609
rect 13985 22583 13986 22609
rect 13958 22553 13986 22583
rect 13958 22527 13959 22553
rect 13985 22527 13986 22553
rect 13230 22161 13258 22167
rect 13230 22135 13231 22161
rect 13257 22135 13258 22161
rect 13230 22106 13258 22135
rect 13230 22040 13258 22078
rect 12838 21704 12866 21742
rect 13118 21770 13146 21775
rect 11494 21378 11522 21383
rect 11270 21377 11522 21378
rect 11270 21351 11271 21377
rect 11297 21351 11495 21377
rect 11521 21351 11522 21377
rect 11270 21350 11522 21351
rect 11270 21345 11298 21350
rect 11494 21345 11522 21350
rect 12278 21377 12306 21383
rect 12278 21351 12279 21377
rect 12305 21351 12306 21377
rect 10822 20567 10823 20593
rect 10849 20567 10850 20593
rect 10822 19809 10850 20567
rect 10822 19783 10823 19809
rect 10849 19783 10850 19809
rect 10822 19025 10850 19783
rect 10822 18999 10823 19025
rect 10849 18999 10850 19025
rect 10822 18242 10850 18999
rect 11270 21041 11298 21047
rect 11270 21015 11271 21041
rect 11297 21015 11298 21041
rect 11270 20985 11298 21015
rect 11270 20959 11271 20985
rect 11297 20959 11298 20985
rect 11270 20594 11298 20959
rect 11494 20594 11522 20599
rect 11270 20593 11522 20594
rect 11270 20567 11271 20593
rect 11297 20567 11495 20593
rect 11521 20567 11522 20593
rect 11270 20566 11522 20567
rect 11270 20257 11298 20566
rect 11494 20561 11522 20566
rect 12278 20593 12306 21351
rect 12278 20567 12279 20593
rect 12305 20567 12306 20593
rect 11270 20231 11271 20257
rect 11297 20231 11298 20257
rect 11270 20201 11298 20231
rect 11270 20175 11271 20201
rect 11297 20175 11298 20201
rect 11270 19810 11298 20175
rect 11494 19810 11522 19815
rect 11270 19809 11522 19810
rect 11270 19783 11271 19809
rect 11297 19783 11495 19809
rect 11521 19783 11522 19809
rect 11270 19782 11522 19783
rect 11270 19473 11298 19782
rect 11494 19777 11522 19782
rect 12278 19809 12306 20567
rect 12278 19783 12279 19809
rect 12305 19783 12306 19809
rect 11270 19447 11271 19473
rect 11297 19447 11298 19473
rect 11270 19417 11298 19447
rect 11270 19391 11271 19417
rect 11297 19391 11298 19417
rect 11270 19026 11298 19391
rect 11494 19026 11522 19031
rect 11270 19025 11522 19026
rect 11270 18999 11271 19025
rect 11297 18999 11495 19025
rect 11521 18999 11522 19025
rect 11270 18998 11522 18999
rect 11270 18689 11298 18998
rect 11494 18993 11522 18998
rect 12278 19025 12306 19783
rect 12950 20985 12978 20991
rect 12950 20959 12951 20985
rect 12977 20959 12978 20985
rect 12950 20258 12978 20959
rect 12950 20201 12978 20230
rect 12950 20175 12951 20201
rect 12977 20175 12978 20201
rect 12950 19417 12978 20175
rect 12950 19391 12951 19417
rect 12977 19391 12978 19417
rect 12950 19334 12978 19391
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11270 18663 11271 18689
rect 11297 18663 11298 18689
rect 11270 18633 11298 18663
rect 11270 18607 11271 18633
rect 11297 18607 11298 18633
rect 10934 18242 10962 18247
rect 10822 18241 10934 18242
rect 10822 18215 10823 18241
rect 10849 18215 10934 18241
rect 10822 18214 10934 18215
rect 10822 17458 10850 18214
rect 10934 18209 10962 18214
rect 11270 18242 11298 18607
rect 12278 18466 12306 18999
rect 12838 19306 12978 19334
rect 13118 19418 13146 21742
rect 13398 21770 13426 21775
rect 13510 21770 13538 21775
rect 13398 21769 13510 21770
rect 13398 21743 13399 21769
rect 13425 21743 13510 21769
rect 13398 21742 13510 21743
rect 13398 21737 13426 21742
rect 13454 21377 13482 21383
rect 13454 21351 13455 21377
rect 13481 21351 13482 21377
rect 13454 21321 13482 21351
rect 13454 21295 13455 21321
rect 13481 21295 13482 21321
rect 13454 20593 13482 21295
rect 13454 20567 13455 20593
rect 13481 20567 13482 20593
rect 13454 20538 13482 20567
rect 13454 20491 13482 20510
rect 12838 18633 12866 19306
rect 12838 18607 12839 18633
rect 12865 18607 12866 18633
rect 12838 18522 12866 18607
rect 12838 18489 12866 18494
rect 11494 18242 11522 18247
rect 11270 18241 11522 18242
rect 11270 18215 11271 18241
rect 11297 18215 11495 18241
rect 11521 18215 11522 18241
rect 11270 18214 11522 18215
rect 10318 17457 10850 17458
rect 10318 17431 10823 17457
rect 10849 17431 10850 17457
rect 10318 17430 10850 17431
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9814 17095 9815 17121
rect 9841 17095 9842 17121
rect 9814 17065 9842 17095
rect 9814 17039 9815 17065
rect 9841 17039 9842 17065
rect 9814 16337 9842 17039
rect 10318 17066 10346 17430
rect 10822 17425 10850 17430
rect 11270 17905 11298 18214
rect 11494 18209 11522 18214
rect 12278 18242 12306 18438
rect 12278 18195 12306 18214
rect 11270 17879 11271 17905
rect 11297 17879 11298 17905
rect 11270 17850 11298 17879
rect 11270 17458 11298 17822
rect 13118 17849 13146 19390
rect 13454 19810 13482 19815
rect 13510 19810 13538 21742
rect 13958 21042 13986 22527
rect 14014 22106 14042 22111
rect 14014 21770 14042 22078
rect 14014 21737 14042 21742
rect 14014 21042 14042 21047
rect 13958 21041 14042 21042
rect 13958 21015 14015 21041
rect 14041 21015 14042 21041
rect 13958 21014 14042 21015
rect 14014 20985 14042 21014
rect 14014 20959 14015 20985
rect 14041 20959 14042 20985
rect 14014 20538 14042 20959
rect 14014 20257 14042 20510
rect 14014 20231 14015 20257
rect 14041 20231 14042 20257
rect 14014 20202 14042 20231
rect 14014 20155 14042 20174
rect 13454 19809 13538 19810
rect 13454 19783 13455 19809
rect 13481 19783 13538 19809
rect 13454 19782 13538 19783
rect 13454 19753 13482 19782
rect 13454 19727 13455 19753
rect 13481 19727 13482 19753
rect 13454 19474 13482 19727
rect 13454 19025 13482 19446
rect 14014 19474 14042 19479
rect 14014 19417 14042 19446
rect 14014 19391 14015 19417
rect 14041 19391 14042 19417
rect 14014 19385 14042 19391
rect 13454 18999 13455 19025
rect 13481 18999 13482 19025
rect 13454 18969 13482 18999
rect 13454 18943 13455 18969
rect 13481 18943 13482 18969
rect 13398 18634 13426 18639
rect 13454 18634 13482 18943
rect 13510 18634 13538 18639
rect 13398 18633 13538 18634
rect 13398 18607 13399 18633
rect 13425 18607 13511 18633
rect 13537 18607 13538 18633
rect 13398 18606 13538 18607
rect 13398 18601 13426 18606
rect 13454 18241 13482 18606
rect 13510 18601 13538 18606
rect 13454 18215 13455 18241
rect 13481 18215 13482 18241
rect 13454 18186 13482 18215
rect 13454 18185 13538 18186
rect 13454 18159 13455 18185
rect 13481 18159 13538 18185
rect 13454 18158 13538 18159
rect 13454 18153 13482 18158
rect 13118 17823 13119 17849
rect 13145 17823 13146 17849
rect 13118 17817 13146 17823
rect 13398 17850 13426 17855
rect 13510 17850 13538 18158
rect 13398 17849 13538 17850
rect 13398 17823 13399 17849
rect 13425 17823 13511 17849
rect 13537 17823 13538 17849
rect 13398 17822 13538 17823
rect 13398 17817 13426 17822
rect 11494 17458 11522 17463
rect 11270 17457 11522 17458
rect 11270 17431 11271 17457
rect 11297 17431 11495 17457
rect 11521 17431 11522 17457
rect 11270 17430 11522 17431
rect 10318 17019 10346 17038
rect 11270 17121 11298 17430
rect 11494 17425 11522 17430
rect 12558 17457 12586 17463
rect 12558 17431 12559 17457
rect 12585 17431 12586 17457
rect 11270 17095 11271 17121
rect 11297 17095 11298 17121
rect 11270 17065 11298 17095
rect 11270 17039 11271 17065
rect 11297 17039 11298 17065
rect 10822 16673 10850 16679
rect 10822 16647 10823 16673
rect 10849 16647 10850 16673
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9814 16311 9815 16337
rect 9841 16311 9842 16337
rect 9814 16281 9842 16311
rect 9814 16255 9815 16281
rect 9841 16255 9842 16281
rect 9814 15974 9842 16255
rect 8862 15946 9170 15974
rect 9310 15946 9842 15974
rect 10598 16282 10626 16287
rect 10822 16282 10850 16647
rect 10598 16281 10850 16282
rect 10598 16255 10599 16281
rect 10625 16255 10850 16281
rect 10598 16254 10850 16255
rect 8470 15554 8498 15559
rect 8302 15553 8498 15554
rect 8302 15527 8471 15553
rect 8497 15527 8498 15553
rect 8302 15526 8498 15527
rect 8470 15498 8498 15526
rect 8470 15451 8498 15470
rect 8862 15497 8890 15946
rect 8862 15471 8863 15497
rect 8889 15471 8890 15497
rect 8862 15465 8890 15471
rect 9030 15889 9058 15895
rect 9030 15863 9031 15889
rect 9057 15863 9058 15889
rect 9030 15833 9058 15863
rect 9030 15807 9031 15833
rect 9057 15807 9058 15833
rect 9030 15498 9058 15807
rect 7910 15079 7911 15105
rect 7937 15079 7938 15105
rect 7910 15073 7938 15079
rect 9030 15105 9058 15470
rect 9030 15079 9031 15105
rect 9057 15079 9058 15105
rect 9030 15049 9058 15079
rect 9030 15023 9031 15049
rect 9057 15023 9058 15049
rect 7126 14714 7154 14719
rect 6902 14713 7154 14714
rect 6902 14687 6903 14713
rect 6929 14687 7127 14713
rect 7153 14687 7154 14713
rect 6902 14686 7154 14687
rect 6902 14681 6930 14686
rect 6846 14295 6847 14321
rect 6873 14295 6874 14321
rect 6846 14289 6874 14295
rect 7126 14322 7154 14686
rect 8862 14713 8890 14719
rect 8862 14687 8863 14713
rect 8889 14687 8890 14713
rect 7294 14322 7322 14327
rect 7518 14322 7546 14327
rect 7126 14321 7546 14322
rect 7126 14295 7295 14321
rect 7321 14295 7519 14321
rect 7545 14295 7546 14321
rect 7126 14294 7546 14295
rect 7294 14289 7322 14294
rect 7518 14289 7546 14294
rect 8414 14321 8442 14327
rect 8414 14295 8415 14321
rect 8441 14295 8442 14321
rect 6230 14239 6231 14265
rect 6257 14239 6258 14265
rect 4998 13511 4999 13537
rect 5025 13511 5026 13537
rect 4998 13481 5026 13511
rect 4998 13455 4999 13481
rect 5025 13455 5026 13481
rect 4998 13146 5026 13455
rect 3822 12753 3850 12759
rect 3822 12727 3823 12753
rect 3849 12727 3850 12753
rect 3822 12586 3850 12727
rect 4998 12753 5026 13118
rect 4998 12727 4999 12753
rect 5025 12727 5026 12753
rect 4998 12697 5026 12727
rect 4998 12671 4999 12697
rect 5025 12671 5026 12697
rect 4998 12642 5026 12671
rect 4998 12609 5026 12614
rect 5502 13929 5586 13930
rect 5502 13903 5559 13929
rect 5585 13903 5586 13929
rect 5502 13902 5586 13903
rect 5502 13537 5530 13902
rect 5558 13897 5586 13902
rect 6118 13930 6146 13935
rect 6230 13930 6258 14239
rect 8190 13985 8218 13991
rect 8190 13959 8191 13985
rect 8217 13959 8218 13985
rect 6118 13929 6258 13930
rect 6118 13903 6119 13929
rect 6145 13903 6231 13929
rect 6257 13903 6258 13929
rect 6118 13902 6258 13903
rect 5502 13511 5503 13537
rect 5529 13511 5530 13537
rect 5502 13482 5530 13511
rect 6118 13538 6146 13902
rect 6230 13897 6258 13902
rect 7014 13930 7042 13935
rect 7014 13538 7042 13902
rect 6118 13537 6258 13538
rect 6118 13511 6119 13537
rect 6145 13511 6258 13537
rect 6118 13510 6258 13511
rect 6118 13505 6146 13510
rect 5502 13145 5530 13454
rect 6230 13481 6258 13510
rect 6230 13455 6231 13481
rect 6257 13455 6258 13481
rect 5502 13119 5503 13145
rect 5529 13119 5530 13145
rect 5502 12753 5530 13119
rect 5502 12727 5503 12753
rect 5529 12727 5530 12753
rect 3822 12553 3850 12558
rect 4494 12586 4522 12591
rect 3598 12335 3599 12361
rect 3625 12335 3626 12361
rect 2366 12222 2506 12250
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11577 2170 11942
rect 2142 11551 2143 11577
rect 2169 11551 2170 11577
rect 2142 10793 2170 11551
rect 2478 11969 2506 12222
rect 2478 11943 2479 11969
rect 2505 11943 2506 11969
rect 2478 11913 2506 11943
rect 3318 11970 3346 11975
rect 3318 11923 3346 11942
rect 3598 11970 3626 12335
rect 3598 11937 3626 11942
rect 3766 12362 3794 12367
rect 3766 11969 3794 12334
rect 3766 11943 3767 11969
rect 3793 11943 3794 11969
rect 3766 11937 3794 11943
rect 3990 12362 4018 12367
rect 2478 11887 2479 11913
rect 2505 11887 2506 11913
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 2478 11185 2506 11887
rect 3990 11914 4018 12334
rect 4494 11969 4522 12558
rect 5502 12362 5530 12727
rect 6062 13146 6090 13151
rect 6230 13146 6258 13455
rect 6062 13145 6258 13146
rect 6062 13119 6063 13145
rect 6089 13119 6231 13145
rect 6257 13119 6258 13145
rect 6062 13118 6258 13119
rect 6062 12753 6090 13118
rect 6062 12727 6063 12753
rect 6089 12727 6090 12753
rect 4494 11943 4495 11969
rect 4521 11943 4522 11969
rect 4494 11937 4522 11943
rect 5054 12361 5530 12362
rect 5054 12335 5503 12361
rect 5529 12335 5530 12361
rect 5054 12334 5530 12335
rect 3990 11913 4130 11914
rect 3990 11887 3991 11913
rect 4017 11887 4130 11913
rect 3990 11886 4130 11887
rect 3990 11881 4018 11886
rect 4102 11774 4130 11886
rect 4102 11746 4242 11774
rect 2478 11159 2479 11185
rect 2505 11159 2506 11185
rect 2478 11130 2506 11159
rect 2478 11083 2506 11102
rect 2870 11633 2898 11639
rect 2870 11607 2871 11633
rect 2897 11607 2898 11633
rect 2870 11577 2898 11607
rect 4214 11634 4242 11746
rect 4494 11634 4522 11639
rect 4214 11633 4522 11634
rect 4214 11607 4495 11633
rect 4521 11607 4522 11633
rect 4214 11606 4522 11607
rect 2870 11551 2871 11577
rect 2897 11551 2898 11577
rect 2870 11130 2898 11551
rect 2142 10767 2143 10793
rect 2169 10767 2170 10793
rect 2142 10761 2170 10767
rect 2814 10849 2842 10855
rect 2814 10823 2815 10849
rect 2841 10823 2842 10849
rect 2814 10793 2842 10823
rect 2814 10767 2815 10793
rect 2841 10767 2842 10793
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2478 10402 2506 10407
rect 2814 10402 2842 10767
rect 2478 10401 2842 10402
rect 2478 10375 2479 10401
rect 2505 10375 2842 10401
rect 2478 10374 2842 10375
rect 2478 10345 2506 10374
rect 2478 10319 2479 10345
rect 2505 10319 2506 10345
rect 2142 10010 2170 10015
rect 2142 9225 2170 9982
rect 2422 10010 2450 10015
rect 2478 10010 2506 10319
rect 2534 10010 2562 10015
rect 2422 10009 2562 10010
rect 2422 9983 2423 10009
rect 2449 9983 2535 10009
rect 2561 9983 2562 10009
rect 2422 9982 2562 9983
rect 2422 9977 2450 9982
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 2478 9617 2506 9982
rect 2534 9977 2562 9982
rect 2478 9591 2479 9617
rect 2505 9591 2506 9617
rect 2478 9561 2506 9591
rect 2478 9535 2479 9561
rect 2505 9535 2506 9561
rect 2142 9199 2143 9225
rect 2169 9199 2170 9225
rect 2142 8441 2170 9199
rect 2422 9226 2450 9231
rect 2478 9226 2506 9535
rect 2534 9226 2562 9231
rect 2422 9225 2562 9226
rect 2422 9199 2423 9225
rect 2449 9199 2535 9225
rect 2561 9199 2562 9225
rect 2422 9198 2562 9199
rect 2422 9193 2450 9198
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 2478 8833 2506 9198
rect 2534 9193 2562 9198
rect 2478 8807 2479 8833
rect 2505 8807 2506 8833
rect 2478 8777 2506 8807
rect 2478 8751 2479 8777
rect 2505 8751 2506 8777
rect 2142 8415 2143 8441
rect 2169 8415 2170 8441
rect 2142 7657 2170 8415
rect 2422 8442 2450 8447
rect 2478 8442 2506 8751
rect 2534 8442 2562 8447
rect 2422 8441 2534 8442
rect 2422 8415 2423 8441
rect 2449 8415 2534 8441
rect 2422 8414 2534 8415
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 2422 8050 2450 8414
rect 2534 8376 2562 8414
rect 2478 8050 2506 8055
rect 2422 8049 2506 8050
rect 2422 8023 2479 8049
rect 2505 8023 2506 8049
rect 2422 8022 2506 8023
rect 2478 7993 2506 8022
rect 2478 7967 2479 7993
rect 2505 7967 2506 7993
rect 2142 7631 2143 7657
rect 2169 7631 2170 7657
rect 2142 7602 2170 7631
rect 2142 7569 2170 7574
rect 2422 7658 2450 7663
rect 2478 7658 2506 7967
rect 2534 7658 2562 7663
rect 2422 7657 2562 7658
rect 2422 7631 2423 7657
rect 2449 7631 2535 7657
rect 2561 7631 2562 7657
rect 2422 7630 2562 7631
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 1918 6847 1919 6873
rect 1945 6847 1946 6873
rect 1918 6482 1946 6847
rect 1918 6449 1946 6454
rect 2030 7265 2058 7271
rect 2030 7239 2031 7265
rect 2057 7239 2058 7265
rect 2030 7210 2058 7239
rect 2254 7210 2282 7215
rect 2422 7210 2450 7630
rect 2534 7625 2562 7630
rect 2030 7209 2450 7210
rect 2030 7183 2255 7209
rect 2281 7183 2450 7209
rect 2030 7182 2450 7183
rect 1694 6057 1722 6062
rect 1190 5671 1191 5697
rect 1217 5671 1218 5697
rect 1190 5305 1218 5671
rect 1190 5279 1191 5305
rect 1217 5279 1218 5305
rect 1190 4913 1218 5279
rect 1190 4887 1191 4913
rect 1217 4887 1218 4913
rect 1190 4521 1218 4887
rect 1190 4495 1191 4521
rect 1217 4495 1218 4521
rect 1190 4489 1218 4495
rect 2030 5306 2058 7182
rect 2254 7177 2282 7182
rect 2870 6929 2898 11102
rect 3430 11577 3458 11583
rect 3430 11551 3431 11577
rect 3457 11551 3458 11577
rect 3430 11185 3458 11551
rect 3430 11159 3431 11185
rect 3457 11159 3458 11185
rect 3430 10793 3458 11159
rect 3430 10767 3431 10793
rect 3457 10767 3458 10793
rect 3430 10401 3458 10767
rect 4494 11577 4522 11606
rect 4494 11551 4495 11577
rect 4521 11551 4522 11577
rect 4494 10849 4522 11551
rect 5054 11577 5082 12334
rect 5502 12329 5530 12334
rect 5670 12642 5698 12647
rect 5670 11969 5698 12614
rect 6062 12642 6090 12727
rect 6062 12361 6090 12614
rect 6062 12335 6063 12361
rect 6089 12335 6090 12361
rect 6062 12329 6090 12335
rect 6230 12697 6258 13118
rect 6230 12671 6231 12697
rect 6257 12671 6258 12697
rect 6230 12361 6258 12671
rect 6230 12335 6231 12361
rect 6257 12335 6258 12361
rect 6230 12329 6258 12335
rect 6958 13537 7042 13538
rect 6958 13511 7015 13537
rect 7041 13511 7042 13537
rect 6958 13510 7042 13511
rect 6958 13482 6986 13510
rect 7014 13505 7042 13510
rect 8190 13929 8218 13959
rect 8190 13903 8191 13929
rect 8217 13903 8218 13929
rect 8190 13537 8218 13903
rect 8190 13511 8191 13537
rect 8217 13511 8218 13537
rect 6958 13145 6986 13454
rect 8190 13481 8218 13511
rect 8190 13455 8191 13481
rect 8217 13455 8218 13481
rect 6958 13119 6959 13145
rect 6985 13119 6986 13145
rect 6958 12754 6986 13119
rect 8134 13201 8162 13207
rect 8134 13175 8135 13201
rect 8161 13175 8162 13201
rect 8134 13146 8162 13175
rect 8190 13146 8218 13455
rect 8134 13145 8218 13146
rect 8134 13119 8135 13145
rect 8161 13119 8218 13145
rect 8134 13118 8218 13119
rect 8134 13113 8162 13118
rect 7014 12754 7042 12759
rect 6958 12753 7042 12754
rect 6958 12727 7015 12753
rect 7041 12727 7042 12753
rect 6958 12726 7042 12727
rect 6958 12361 6986 12726
rect 7014 12721 7042 12726
rect 8190 12753 8218 13118
rect 8190 12727 8191 12753
rect 8217 12727 8218 12753
rect 8190 12697 8218 12727
rect 8190 12671 8191 12697
rect 8217 12671 8218 12697
rect 6958 12335 6959 12361
rect 6985 12335 6986 12361
rect 5670 11943 5671 11969
rect 5697 11943 5698 11969
rect 5670 11913 5698 11943
rect 6958 11970 6986 12335
rect 8134 12417 8162 12423
rect 8134 12391 8135 12417
rect 8161 12391 8162 12417
rect 8134 12362 8162 12391
rect 8190 12362 8218 12671
rect 8134 12361 8218 12362
rect 8134 12335 8135 12361
rect 8161 12335 8218 12361
rect 8134 12334 8218 12335
rect 8134 12329 8162 12334
rect 7014 11970 7042 11975
rect 6958 11969 7042 11970
rect 6958 11943 7015 11969
rect 7041 11943 7042 11969
rect 6958 11942 7042 11943
rect 7014 11937 7042 11942
rect 8190 11969 8218 12334
rect 8190 11943 8191 11969
rect 8217 11943 8218 11969
rect 5670 11887 5671 11913
rect 5697 11887 5698 11913
rect 5670 11881 5698 11887
rect 8190 11913 8218 11943
rect 8414 13930 8442 14295
rect 8414 13538 8442 13902
rect 8862 13930 8890 14687
rect 9030 14714 9058 15023
rect 9310 15498 9338 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9534 15498 9562 15503
rect 9310 15497 9562 15498
rect 9310 15471 9311 15497
rect 9337 15471 9535 15497
rect 9561 15471 9562 15497
rect 9310 15470 9562 15471
rect 9310 14714 9338 15470
rect 9534 15465 9562 15470
rect 10598 15497 10626 16254
rect 10822 15890 10850 16254
rect 11270 16674 11298 17039
rect 11494 16674 11522 16679
rect 11270 16673 11522 16674
rect 11270 16647 11271 16673
rect 11297 16647 11495 16673
rect 11521 16647 11522 16673
rect 11270 16646 11522 16647
rect 11270 16337 11298 16646
rect 11494 16641 11522 16646
rect 12558 16673 12586 17431
rect 13454 17457 13482 17822
rect 13510 17817 13538 17822
rect 13454 17431 13455 17457
rect 13481 17431 13482 17457
rect 13454 17402 13482 17431
rect 13454 17401 13538 17402
rect 13454 17375 13455 17401
rect 13481 17375 13538 17401
rect 13454 17374 13538 17375
rect 13454 17369 13482 17374
rect 12558 16647 12559 16673
rect 12585 16647 12586 16673
rect 11270 16311 11271 16337
rect 11297 16311 11298 16337
rect 11270 16281 11298 16311
rect 11270 16255 11271 16281
rect 11297 16255 11298 16281
rect 11102 15890 11130 15895
rect 10822 15889 11130 15890
rect 10822 15863 11103 15889
rect 11129 15863 11130 15889
rect 10822 15862 11130 15863
rect 11270 15890 11298 16255
rect 11382 15890 11410 15895
rect 11494 15890 11522 15895
rect 11270 15889 11522 15890
rect 11270 15863 11383 15889
rect 11409 15863 11495 15889
rect 11521 15863 11522 15889
rect 11270 15862 11522 15863
rect 10598 15471 10599 15497
rect 10625 15471 10626 15497
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9422 14714 9450 14719
rect 9534 14714 9562 14719
rect 9030 14713 9562 14714
rect 9030 14687 9423 14713
rect 9449 14687 9535 14713
rect 9561 14687 9562 14713
rect 9030 14686 9562 14687
rect 8862 13883 8890 13902
rect 9422 14321 9450 14686
rect 9534 14681 9562 14686
rect 10598 14713 10626 15471
rect 10598 14687 10599 14713
rect 10625 14687 10626 14713
rect 9422 14295 9423 14321
rect 9449 14295 9450 14321
rect 9422 14265 9450 14295
rect 9422 14239 9423 14265
rect 9449 14239 9450 14265
rect 9422 13930 9450 14239
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9534 13930 9562 13935
rect 9422 13929 9562 13930
rect 9422 13903 9423 13929
rect 9449 13903 9535 13929
rect 9561 13903 9562 13929
rect 9422 13902 9562 13903
rect 8470 13538 8498 13543
rect 8414 13537 8498 13538
rect 8414 13511 8471 13537
rect 8497 13511 8498 13537
rect 8414 13510 8498 13511
rect 8414 12754 8442 13510
rect 8470 13505 8498 13510
rect 9422 13537 9450 13902
rect 9534 13897 9562 13902
rect 10598 13929 10626 14687
rect 10598 13903 10599 13929
rect 10625 13903 10626 13929
rect 9422 13511 9423 13537
rect 9449 13511 9450 13537
rect 9422 13481 9450 13511
rect 9422 13455 9423 13481
rect 9449 13455 9450 13481
rect 8862 13145 8890 13151
rect 8862 13119 8863 13145
rect 8889 13119 8890 13145
rect 8470 12754 8498 12759
rect 8414 12753 8498 12754
rect 8414 12727 8471 12753
rect 8497 12727 8498 12753
rect 8414 12726 8498 12727
rect 8414 12362 8442 12726
rect 8470 12721 8498 12726
rect 8862 12362 8890 13119
rect 8414 12334 8862 12362
rect 8414 11970 8442 12334
rect 8862 12296 8890 12334
rect 9422 13146 9450 13455
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9534 13146 9562 13151
rect 9422 13145 9562 13146
rect 9422 13119 9423 13145
rect 9449 13119 9535 13145
rect 9561 13119 9562 13145
rect 9422 13118 9562 13119
rect 9422 12753 9450 13118
rect 9534 13113 9562 13118
rect 10598 13145 10626 13903
rect 10598 13119 10599 13145
rect 10625 13119 10626 13145
rect 9422 12727 9423 12753
rect 9449 12727 9450 12753
rect 9422 12697 9450 12727
rect 9422 12671 9423 12697
rect 9449 12671 9450 12697
rect 9422 12362 9450 12671
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9534 12362 9562 12367
rect 9422 12361 9562 12362
rect 9422 12335 9423 12361
rect 9449 12335 9535 12361
rect 9561 12335 9562 12361
rect 9422 12334 9562 12335
rect 8470 11970 8498 11975
rect 8414 11969 8498 11970
rect 8414 11943 8471 11969
rect 8497 11943 8498 11969
rect 8414 11942 8498 11943
rect 8470 11937 8498 11942
rect 9422 11969 9450 12334
rect 9534 12329 9562 12334
rect 10598 12362 10626 13119
rect 9422 11943 9423 11969
rect 9449 11943 9450 11969
rect 8190 11887 8191 11913
rect 8217 11887 8218 11913
rect 8190 11802 8218 11887
rect 5054 11551 5055 11577
rect 5081 11551 5082 11577
rect 4494 10823 4495 10849
rect 4521 10823 4522 10849
rect 4494 10794 4522 10823
rect 4606 11185 4634 11191
rect 4606 11159 4607 11185
rect 4633 11159 4634 11185
rect 4606 11129 4634 11159
rect 4606 11103 4607 11129
rect 4633 11103 4634 11129
rect 4606 10794 4634 11103
rect 4494 10793 4634 10794
rect 4494 10767 4495 10793
rect 4521 10767 4634 10793
rect 4494 10766 4634 10767
rect 4494 10761 4522 10766
rect 3430 10375 3431 10401
rect 3457 10375 3458 10401
rect 3430 10010 3458 10375
rect 4606 10401 4634 10766
rect 4606 10375 4607 10401
rect 4633 10375 4634 10401
rect 4270 10346 4298 10351
rect 4270 10094 4298 10318
rect 4606 10346 4634 10375
rect 4606 10299 4634 10318
rect 5054 11185 5082 11551
rect 5054 11159 5055 11185
rect 5081 11159 5082 11185
rect 5054 10793 5082 11159
rect 5054 10767 5055 10793
rect 5081 10767 5082 10793
rect 5054 10401 5082 10767
rect 5054 10375 5055 10401
rect 5081 10375 5082 10401
rect 5054 10094 5082 10375
rect 5838 11633 5866 11639
rect 5838 11607 5839 11633
rect 5865 11607 5866 11633
rect 5838 11577 5866 11607
rect 8190 11633 8218 11774
rect 8190 11607 8191 11633
rect 8217 11607 8218 11633
rect 5838 11551 5839 11577
rect 5865 11551 5866 11577
rect 5838 11185 5866 11551
rect 7294 11577 7322 11583
rect 7294 11551 7295 11577
rect 7321 11551 7322 11577
rect 5838 11159 5839 11185
rect 5865 11159 5866 11185
rect 5838 11129 5866 11159
rect 5838 11103 5839 11129
rect 5865 11103 5866 11129
rect 5838 10849 5866 11103
rect 5838 10823 5839 10849
rect 5865 10823 5866 10849
rect 5838 10793 5866 10823
rect 5838 10767 5839 10793
rect 5865 10767 5866 10793
rect 5838 10401 5866 10767
rect 5838 10375 5839 10401
rect 5865 10375 5866 10401
rect 5838 10346 5866 10375
rect 5838 10280 5866 10318
rect 7238 11185 7266 11191
rect 7238 11159 7239 11185
rect 7265 11159 7266 11185
rect 7238 10793 7266 11159
rect 7294 11186 7322 11551
rect 8190 11577 8218 11607
rect 9422 11913 9450 11943
rect 9422 11887 9423 11913
rect 9449 11887 9450 11913
rect 9422 11802 9450 11887
rect 8190 11551 8191 11577
rect 8217 11551 8218 11577
rect 8190 11545 8218 11551
rect 8862 11577 8890 11583
rect 8862 11551 8863 11577
rect 8889 11551 8890 11577
rect 7294 11153 7322 11158
rect 8078 11185 8106 11191
rect 8078 11159 8079 11185
rect 8105 11159 8106 11185
rect 7238 10767 7239 10793
rect 7265 10767 7266 10793
rect 7238 10401 7266 10767
rect 7238 10375 7239 10401
rect 7265 10375 7266 10401
rect 4270 10066 4522 10094
rect 5054 10066 5530 10094
rect 4494 10065 4522 10066
rect 4494 10039 4495 10065
rect 4521 10039 4522 10065
rect 3598 10010 3626 10015
rect 3430 10009 3626 10010
rect 3430 9983 3599 10009
rect 3625 9983 3626 10009
rect 3430 9982 3626 9983
rect 2870 6903 2871 6929
rect 2897 6903 2898 6929
rect 2870 6873 2898 6903
rect 2870 6847 2871 6873
rect 2897 6847 2898 6873
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2478 6482 2506 6487
rect 2870 6482 2898 6847
rect 3598 9225 3626 9982
rect 4494 10009 4522 10039
rect 4494 9983 4495 10009
rect 4521 9983 4522 10009
rect 3598 9199 3599 9225
rect 3625 9199 3626 9225
rect 3598 8441 3626 9199
rect 3822 9617 3850 9623
rect 3822 9591 3823 9617
rect 3849 9591 3850 9617
rect 3822 8833 3850 9591
rect 4382 9618 4410 9623
rect 4494 9618 4522 9983
rect 5502 10009 5530 10066
rect 5502 9983 5503 10009
rect 5529 9983 5530 10009
rect 4382 9617 4522 9618
rect 4382 9591 4383 9617
rect 4409 9591 4495 9617
rect 4521 9591 4522 9617
rect 4382 9590 4522 9591
rect 4382 9585 4410 9590
rect 4494 9281 4522 9590
rect 4494 9255 4495 9281
rect 4521 9255 4522 9281
rect 4494 9225 4522 9255
rect 4494 9199 4495 9225
rect 4521 9199 4522 9225
rect 3822 8807 3823 8833
rect 3849 8807 3850 8833
rect 3598 8415 3599 8441
rect 3625 8415 3626 8441
rect 3598 7657 3626 8415
rect 3766 8442 3794 8447
rect 3766 8395 3794 8414
rect 3598 7631 3599 7657
rect 3625 7631 3626 7657
rect 3598 7546 3626 7631
rect 3598 7266 3626 7518
rect 3598 6873 3626 7238
rect 3822 8049 3850 8807
rect 4382 8834 4410 8839
rect 4494 8834 4522 9199
rect 5446 9618 5474 9623
rect 5502 9618 5530 9983
rect 6678 10065 6706 10071
rect 6678 10039 6679 10065
rect 6705 10039 6706 10065
rect 6678 10009 6706 10039
rect 6678 9983 6679 10009
rect 6705 9983 6706 10009
rect 5446 9617 5530 9618
rect 5446 9591 5447 9617
rect 5473 9591 5530 9617
rect 5446 9590 5530 9591
rect 6454 9617 6482 9623
rect 6454 9591 6455 9617
rect 6481 9591 6482 9617
rect 5446 9226 5474 9590
rect 6454 9562 6482 9591
rect 6678 9562 6706 9983
rect 7238 10009 7266 10375
rect 8078 11129 8106 11159
rect 8078 11103 8079 11129
rect 8105 11103 8106 11129
rect 8078 10849 8106 11103
rect 8078 10823 8079 10849
rect 8105 10823 8106 10849
rect 8078 10793 8106 10823
rect 8078 10767 8079 10793
rect 8105 10767 8106 10793
rect 8078 10401 8106 10767
rect 8078 10375 8079 10401
rect 8105 10375 8106 10401
rect 8078 10345 8106 10375
rect 8414 11186 8442 11191
rect 8414 10401 8442 11158
rect 8862 11186 8890 11551
rect 8862 10794 8890 11158
rect 9422 11185 9450 11774
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9422 11159 9423 11185
rect 9449 11159 9450 11185
rect 9422 11129 9450 11159
rect 9422 11103 9423 11129
rect 9449 11103 9450 11129
rect 9422 10794 9450 11103
rect 10038 11633 10066 11639
rect 10038 11607 10039 11633
rect 10065 11607 10066 11633
rect 10038 11577 10066 11607
rect 10038 11551 10039 11577
rect 10065 11551 10066 11577
rect 10038 11074 10066 11551
rect 10598 11577 10626 12334
rect 10598 11551 10599 11577
rect 10625 11551 10626 11577
rect 10038 11046 10122 11074
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10094 10906 10122 11046
rect 9590 10878 10122 10906
rect 9590 10794 9618 10878
rect 8862 10793 9170 10794
rect 8862 10767 8863 10793
rect 8889 10767 9170 10793
rect 8862 10766 9170 10767
rect 8862 10761 8890 10766
rect 8414 10375 8415 10401
rect 8441 10375 8442 10401
rect 8414 10369 8442 10375
rect 8078 10319 8079 10345
rect 8105 10319 8106 10345
rect 8078 10094 8106 10319
rect 8078 10066 8162 10094
rect 7238 9983 7239 10009
rect 7265 9983 7266 10009
rect 7182 9618 7210 9623
rect 7238 9618 7266 9983
rect 8134 10065 8162 10066
rect 8134 10039 8135 10065
rect 8161 10039 8162 10065
rect 8134 10009 8162 10039
rect 8134 9983 8135 10009
rect 8161 9983 8162 10009
rect 7182 9617 7266 9618
rect 7182 9591 7183 9617
rect 7209 9591 7266 9617
rect 7182 9590 7266 9591
rect 7182 9585 7210 9590
rect 6454 9561 6706 9562
rect 6454 9535 6455 9561
rect 6481 9535 6706 9561
rect 6454 9534 6706 9535
rect 6454 9529 6482 9534
rect 6678 9281 6706 9534
rect 6678 9255 6679 9281
rect 6705 9255 6706 9281
rect 5502 9226 5530 9231
rect 5446 9225 5530 9226
rect 5446 9199 5503 9225
rect 5529 9199 5530 9225
rect 5446 9198 5530 9199
rect 4382 8833 4522 8834
rect 4382 8807 4383 8833
rect 4409 8807 4495 8833
rect 4521 8807 4522 8833
rect 4382 8806 4522 8807
rect 4382 8801 4410 8806
rect 3822 8023 3823 8049
rect 3849 8023 3850 8049
rect 3822 7266 3850 8023
rect 3822 7233 3850 7238
rect 4494 8442 4522 8806
rect 4494 7713 4522 8414
rect 5278 8833 5306 8839
rect 5278 8807 5279 8833
rect 5305 8807 5306 8833
rect 5278 8442 5306 8807
rect 5446 8442 5474 9198
rect 5502 9193 5530 9198
rect 6678 9225 6706 9255
rect 6678 9199 6679 9225
rect 6705 9199 6706 9225
rect 5278 8441 5474 8442
rect 5278 8415 5447 8441
rect 5473 8415 5474 8441
rect 5278 8414 5474 8415
rect 4494 7687 4495 7713
rect 4521 7687 4522 7713
rect 4494 7657 4522 7687
rect 4494 7631 4495 7657
rect 4521 7631 4522 7657
rect 4494 7602 4522 7631
rect 4494 7265 4522 7574
rect 4998 8049 5026 8055
rect 5278 8050 5306 8414
rect 5446 8409 5474 8414
rect 6454 8833 6482 8839
rect 6454 8807 6455 8833
rect 6481 8807 6482 8833
rect 6454 8777 6482 8807
rect 6454 8751 6455 8777
rect 6481 8751 6482 8777
rect 4998 8023 4999 8049
rect 5025 8023 5026 8049
rect 4998 7993 5026 8023
rect 4998 7967 4999 7993
rect 5025 7967 5026 7993
rect 4998 7602 5026 7967
rect 5166 8049 5306 8050
rect 5166 8023 5279 8049
rect 5305 8023 5306 8049
rect 5166 8022 5306 8023
rect 5166 7657 5194 8022
rect 5278 8017 5306 8022
rect 6454 8386 6482 8751
rect 6622 8497 6650 8503
rect 6622 8471 6623 8497
rect 6649 8471 6650 8497
rect 6622 8442 6650 8471
rect 6678 8442 6706 9199
rect 7238 9225 7266 9590
rect 8078 9617 8106 9623
rect 8078 9591 8079 9617
rect 8105 9591 8106 9617
rect 8078 9562 8106 9591
rect 8134 9562 8162 9983
rect 9142 10009 9170 10766
rect 9422 10793 9618 10794
rect 9422 10767 9423 10793
rect 9449 10767 9591 10793
rect 9617 10767 9618 10793
rect 9422 10766 9618 10767
rect 9422 10761 9450 10766
rect 9142 9983 9143 10009
rect 9169 9983 9170 10009
rect 8078 9561 8162 9562
rect 8078 9535 8079 9561
rect 8105 9535 8162 9561
rect 8078 9534 8162 9535
rect 8078 9529 8106 9534
rect 7238 9199 7239 9225
rect 7265 9199 7266 9225
rect 7182 8834 7210 8839
rect 7238 8834 7266 9199
rect 8134 9281 8162 9534
rect 8134 9255 8135 9281
rect 8161 9255 8162 9281
rect 8134 9225 8162 9255
rect 8134 9199 8135 9225
rect 8161 9199 8162 9225
rect 7182 8833 7266 8834
rect 7182 8807 7183 8833
rect 7209 8807 7266 8833
rect 7182 8806 7266 8807
rect 7182 8801 7210 8806
rect 6622 8441 6706 8442
rect 6622 8415 6623 8441
rect 6649 8415 6706 8441
rect 6622 8414 6706 8415
rect 6622 8409 6650 8414
rect 6454 8049 6482 8358
rect 6678 8386 6706 8414
rect 7182 8442 7210 8447
rect 7238 8442 7266 8806
rect 8078 8833 8106 8839
rect 8078 8807 8079 8833
rect 8105 8807 8106 8833
rect 8078 8778 8106 8807
rect 8134 8778 8162 9199
rect 8638 9617 8666 9623
rect 8638 9591 8639 9617
rect 8665 9591 8666 9617
rect 8638 8834 8666 9591
rect 9142 9225 9170 9983
rect 9590 10401 9618 10766
rect 9590 10375 9591 10401
rect 9617 10375 9618 10401
rect 9590 10345 9618 10375
rect 9590 10319 9591 10345
rect 9617 10319 9618 10345
rect 9142 9199 9143 9225
rect 9169 9199 9170 9225
rect 8638 8833 8722 8834
rect 8638 8807 8639 8833
rect 8665 8807 8722 8833
rect 8638 8806 8722 8807
rect 8638 8801 8666 8806
rect 8078 8777 8162 8778
rect 8078 8751 8079 8777
rect 8105 8751 8162 8777
rect 8078 8750 8162 8751
rect 8078 8745 8106 8750
rect 7182 8441 7266 8442
rect 7182 8415 7183 8441
rect 7209 8415 7266 8441
rect 7182 8414 7266 8415
rect 7182 8409 7210 8414
rect 6678 8353 6706 8358
rect 6454 8023 6455 8049
rect 6481 8023 6482 8049
rect 6454 7993 6482 8023
rect 6454 7967 6455 7993
rect 6481 7967 6482 7993
rect 6454 7961 6482 7967
rect 7238 8049 7266 8414
rect 8078 8497 8106 8503
rect 8078 8471 8079 8497
rect 8105 8471 8106 8497
rect 8078 8442 8106 8471
rect 8134 8442 8162 8750
rect 8078 8441 8162 8442
rect 8078 8415 8079 8441
rect 8105 8415 8162 8441
rect 8078 8414 8162 8415
rect 8078 8409 8106 8414
rect 7238 8023 7239 8049
rect 7265 8023 7266 8049
rect 5166 7631 5167 7657
rect 5193 7631 5194 7657
rect 5166 7625 5194 7631
rect 5838 7713 5866 7719
rect 5838 7687 5839 7713
rect 5865 7687 5866 7713
rect 5838 7657 5866 7687
rect 5838 7631 5839 7657
rect 5865 7631 5866 7657
rect 4998 7569 5026 7574
rect 5838 7602 5866 7631
rect 4494 7239 4495 7265
rect 4521 7239 4522 7265
rect 3598 6847 3599 6873
rect 3625 6847 3626 6873
rect 3598 6841 3626 6847
rect 4494 7209 4522 7239
rect 4494 7183 4495 7209
rect 4521 7183 4522 7209
rect 4494 6929 4522 7183
rect 4494 6903 4495 6929
rect 4521 6903 4522 6929
rect 4494 6873 4522 6903
rect 4494 6847 4495 6873
rect 4521 6847 4522 6873
rect 4494 6841 4522 6847
rect 4886 7266 4914 7271
rect 4886 6873 4914 7238
rect 4886 6847 4887 6873
rect 4913 6847 4914 6873
rect 4886 6841 4914 6847
rect 5838 7265 5866 7574
rect 5838 7239 5839 7265
rect 5865 7239 5866 7265
rect 5838 7209 5866 7239
rect 5838 7183 5839 7209
rect 5865 7183 5866 7209
rect 5838 6929 5866 7183
rect 5838 6903 5839 6929
rect 5865 6903 5866 6929
rect 5838 6873 5866 6903
rect 7238 7657 7266 8023
rect 7238 7631 7239 7657
rect 7265 7631 7266 7657
rect 7238 7266 7266 7631
rect 5838 6847 5839 6873
rect 5865 6847 5866 6873
rect 5838 6841 5866 6847
rect 7182 6874 7210 6879
rect 7238 6874 7266 7238
rect 8134 8386 8162 8414
rect 8134 8050 8162 8358
rect 8134 7993 8162 8022
rect 8134 7967 8135 7993
rect 8161 7967 8162 7993
rect 8134 7713 8162 7967
rect 8134 7687 8135 7713
rect 8161 7687 8162 7713
rect 8134 7657 8162 7687
rect 8134 7631 8135 7657
rect 8161 7631 8162 7657
rect 8134 7265 8162 7631
rect 8134 7239 8135 7265
rect 8161 7239 8162 7265
rect 8134 7210 8162 7239
rect 7182 6873 7266 6874
rect 7182 6847 7183 6873
rect 7209 6847 7266 6873
rect 7182 6846 7266 6847
rect 8078 7209 8162 7210
rect 8078 7183 8135 7209
rect 8161 7183 8162 7209
rect 8694 8162 8722 8806
rect 9142 8441 9170 9199
rect 9534 9618 9562 9623
rect 9590 9618 9618 10319
rect 10598 10793 10626 11551
rect 10598 10767 10599 10793
rect 10625 10767 10626 10793
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10598 10094 10626 10767
rect 9814 10065 9842 10071
rect 9814 10039 9815 10065
rect 9841 10039 9842 10065
rect 9814 10010 9842 10039
rect 10318 10066 10626 10094
rect 11102 15105 11130 15862
rect 11382 15857 11410 15862
rect 11494 15553 11522 15862
rect 11494 15527 11495 15553
rect 11521 15527 11522 15553
rect 11494 15497 11522 15527
rect 11494 15471 11495 15497
rect 11521 15471 11522 15497
rect 11102 15079 11103 15105
rect 11129 15079 11130 15105
rect 11102 14321 11130 15079
rect 11382 15106 11410 15111
rect 11494 15106 11522 15471
rect 11382 15105 11522 15106
rect 11382 15079 11383 15105
rect 11409 15079 11495 15105
rect 11521 15079 11522 15105
rect 11382 15078 11522 15079
rect 11382 15073 11410 15078
rect 11494 14769 11522 15078
rect 11494 14743 11495 14769
rect 11521 14743 11522 14769
rect 11494 14713 11522 14743
rect 11494 14687 11495 14713
rect 11521 14687 11522 14713
rect 11102 14295 11103 14321
rect 11129 14295 11130 14321
rect 11102 13537 11130 14295
rect 11382 14322 11410 14327
rect 11494 14322 11522 14687
rect 11382 14321 11522 14322
rect 11382 14295 11383 14321
rect 11409 14295 11495 14321
rect 11521 14295 11522 14321
rect 11382 14294 11522 14295
rect 11382 14289 11410 14294
rect 11494 13985 11522 14294
rect 11494 13959 11495 13985
rect 11521 13959 11522 13985
rect 11494 13929 11522 13959
rect 11494 13903 11495 13929
rect 11521 13903 11522 13929
rect 11102 13511 11103 13537
rect 11129 13511 11130 13537
rect 11102 12753 11130 13511
rect 11382 13538 11410 13543
rect 11494 13538 11522 13903
rect 11382 13537 11522 13538
rect 11382 13511 11383 13537
rect 11409 13511 11495 13537
rect 11521 13511 11522 13537
rect 11382 13510 11522 13511
rect 11382 13505 11410 13510
rect 11494 13201 11522 13510
rect 11494 13175 11495 13201
rect 11521 13175 11522 13201
rect 11494 13145 11522 13175
rect 11494 13119 11495 13145
rect 11521 13119 11522 13145
rect 11102 12727 11103 12753
rect 11129 12727 11130 12753
rect 11102 11969 11130 12727
rect 11382 12754 11410 12759
rect 11494 12754 11522 13119
rect 11382 12753 11522 12754
rect 11382 12727 11383 12753
rect 11409 12727 11495 12753
rect 11521 12727 11522 12753
rect 11382 12726 11522 12727
rect 11382 12721 11410 12726
rect 11494 12417 11522 12726
rect 11494 12391 11495 12417
rect 11521 12391 11522 12417
rect 11494 12361 11522 12391
rect 11494 12335 11495 12361
rect 11521 12335 11522 12361
rect 11102 11943 11103 11969
rect 11129 11943 11130 11969
rect 11102 11185 11130 11943
rect 11382 11970 11410 11975
rect 11494 11970 11522 12335
rect 11382 11969 11522 11970
rect 11382 11943 11383 11969
rect 11409 11943 11495 11969
rect 11521 11943 11522 11969
rect 11382 11942 11522 11943
rect 11382 11937 11410 11942
rect 11494 11802 11522 11942
rect 11494 11633 11522 11774
rect 11494 11607 11495 11633
rect 11521 11607 11522 11633
rect 11494 11577 11522 11607
rect 11494 11551 11495 11577
rect 11521 11551 11522 11577
rect 11102 11159 11103 11185
rect 11129 11159 11130 11185
rect 11102 10401 11130 11159
rect 11382 11186 11410 11191
rect 11494 11186 11522 11551
rect 11382 11185 11522 11186
rect 11382 11159 11383 11185
rect 11409 11159 11495 11185
rect 11521 11159 11522 11185
rect 11382 11158 11522 11159
rect 11382 11153 11410 11158
rect 11494 10849 11522 11158
rect 12558 15889 12586 16647
rect 12894 17065 12922 17071
rect 12894 17039 12895 17065
rect 12921 17039 12922 17065
rect 12894 16281 12922 17039
rect 13398 17066 13426 17071
rect 13510 17066 13538 17374
rect 13398 17065 13538 17066
rect 13398 17039 13399 17065
rect 13425 17039 13511 17065
rect 13537 17039 13538 17065
rect 13398 17038 13538 17039
rect 13398 17033 13426 17038
rect 13454 16673 13482 17038
rect 13510 17033 13538 17038
rect 13454 16647 13455 16673
rect 13481 16647 13482 16673
rect 13454 16618 13482 16647
rect 13454 16617 13538 16618
rect 13454 16591 13455 16617
rect 13481 16591 13538 16617
rect 13454 16590 13538 16591
rect 13454 16585 13482 16590
rect 12894 16255 12895 16281
rect 12921 16255 12922 16281
rect 12894 15974 12922 16255
rect 13398 16282 13426 16287
rect 13510 16282 13538 16590
rect 13398 16281 13538 16282
rect 13398 16255 13399 16281
rect 13425 16255 13511 16281
rect 13537 16255 13538 16281
rect 13398 16254 13538 16255
rect 13398 16249 13426 16254
rect 12894 15946 13146 15974
rect 12558 15863 12559 15889
rect 12585 15863 12586 15889
rect 12558 15105 12586 15863
rect 12558 15079 12559 15105
rect 12585 15079 12586 15105
rect 12558 14321 12586 15079
rect 12558 14295 12559 14321
rect 12585 14295 12586 14321
rect 12558 13537 12586 14295
rect 12558 13511 12559 13537
rect 12585 13511 12586 13537
rect 12558 12753 12586 13511
rect 12558 12727 12559 12753
rect 12585 12727 12586 12753
rect 12558 11969 12586 12727
rect 12558 11943 12559 11969
rect 12585 11943 12586 11969
rect 12558 11186 12586 11943
rect 12558 11139 12586 11158
rect 12726 15890 12754 15895
rect 12950 15890 12978 15895
rect 12726 15889 12978 15890
rect 12726 15863 12727 15889
rect 12753 15863 12951 15889
rect 12977 15863 12978 15889
rect 12726 15862 12978 15863
rect 12726 15106 12754 15862
rect 12950 15857 12978 15862
rect 13118 15497 13146 15946
rect 13118 15471 13119 15497
rect 13145 15471 13146 15497
rect 12950 15106 12978 15111
rect 12726 15105 12978 15106
rect 12726 15079 12727 15105
rect 12753 15079 12951 15105
rect 12977 15079 12978 15105
rect 12726 15078 12978 15079
rect 12726 14322 12754 15078
rect 12950 15073 12978 15078
rect 13118 14713 13146 15471
rect 13118 14687 13119 14713
rect 13145 14687 13146 14713
rect 12950 14322 12978 14327
rect 12726 14321 12978 14322
rect 12726 14295 12727 14321
rect 12753 14295 12951 14321
rect 12977 14295 12978 14321
rect 12726 14294 12978 14295
rect 12726 13538 12754 14294
rect 12950 14289 12978 14294
rect 13118 13929 13146 14687
rect 13118 13903 13119 13929
rect 13145 13903 13146 13929
rect 12950 13538 12978 13543
rect 12726 13537 12978 13538
rect 12726 13511 12727 13537
rect 12753 13511 12951 13537
rect 12977 13511 12978 13537
rect 12726 13510 12978 13511
rect 12726 12754 12754 13510
rect 12950 13505 12978 13510
rect 13118 13145 13146 13903
rect 13118 13119 13119 13145
rect 13145 13119 13146 13145
rect 12950 12754 12978 12759
rect 12726 12753 12978 12754
rect 12726 12727 12727 12753
rect 12753 12727 12951 12753
rect 12977 12727 12978 12753
rect 12726 12726 12978 12727
rect 12726 11969 12754 12726
rect 12950 12721 12978 12726
rect 13118 12362 13146 13119
rect 13118 12315 13146 12334
rect 13286 15498 13314 15503
rect 13510 15498 13538 16254
rect 13286 15497 13538 15498
rect 13286 15471 13287 15497
rect 13313 15471 13511 15497
rect 13537 15471 13538 15497
rect 13286 15470 13538 15471
rect 13286 14714 13314 15470
rect 13510 15465 13538 15470
rect 13510 14714 13538 14719
rect 13286 14713 13538 14714
rect 13286 14687 13287 14713
rect 13313 14687 13511 14713
rect 13537 14687 13538 14713
rect 13286 14686 13538 14687
rect 13286 13930 13314 14686
rect 13510 14681 13538 14686
rect 13510 13930 13538 13935
rect 13286 13929 13538 13930
rect 13286 13903 13287 13929
rect 13313 13903 13511 13929
rect 13537 13903 13538 13929
rect 13286 13902 13538 13903
rect 13286 13146 13314 13902
rect 13510 13897 13538 13902
rect 13510 13146 13538 13151
rect 13286 13145 13538 13146
rect 13286 13119 13287 13145
rect 13313 13119 13511 13145
rect 13537 13119 13538 13145
rect 13286 13118 13538 13119
rect 13286 12362 13314 13118
rect 13510 13113 13538 13118
rect 13510 12362 13538 12367
rect 13286 12361 13538 12362
rect 13286 12335 13287 12361
rect 13313 12335 13511 12361
rect 13537 12335 13538 12361
rect 13286 12334 13538 12335
rect 12726 11943 12727 11969
rect 12753 11943 12754 11969
rect 12726 11802 12754 11943
rect 12726 11186 12754 11774
rect 12950 11969 12978 11975
rect 12950 11943 12951 11969
rect 12977 11943 12978 11969
rect 12950 11802 12978 11943
rect 12950 11769 12978 11774
rect 13286 11802 13314 12334
rect 13510 12306 13538 12334
rect 13510 12273 13538 12278
rect 13118 11577 13146 11583
rect 13118 11551 13119 11577
rect 13145 11551 13146 11577
rect 12950 11186 12978 11191
rect 12726 11185 12978 11186
rect 12726 11159 12727 11185
rect 12753 11159 12951 11185
rect 12977 11159 12978 11185
rect 12726 11158 12978 11159
rect 12726 11153 12754 11158
rect 12950 11153 12978 11158
rect 13118 11186 13146 11551
rect 13286 11578 13314 11774
rect 13510 11578 13538 11583
rect 13286 11577 13538 11578
rect 13286 11551 13287 11577
rect 13313 11551 13511 11577
rect 13537 11551 13538 11577
rect 13286 11550 13538 11551
rect 13286 11545 13314 11550
rect 13510 11545 13538 11550
rect 11494 10823 11495 10849
rect 11521 10823 11522 10849
rect 11494 10793 11522 10823
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11102 10375 11103 10401
rect 11129 10375 11130 10401
rect 9814 9944 9842 9982
rect 10038 10010 10066 10015
rect 9534 9617 9618 9618
rect 9534 9591 9535 9617
rect 9561 9591 9618 9617
rect 9534 9590 9618 9591
rect 9534 9561 9562 9590
rect 9534 9535 9535 9561
rect 9561 9535 9562 9561
rect 9534 8833 9562 9535
rect 10038 9506 10066 9982
rect 10318 10009 10346 10066
rect 10318 9983 10319 10009
rect 10345 9983 10346 10009
rect 10038 9478 10122 9506
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 10094 9338 10122 9478
rect 10038 9310 10122 9338
rect 10038 9281 10066 9310
rect 10038 9255 10039 9281
rect 10065 9255 10066 9281
rect 10038 9225 10066 9255
rect 10038 9199 10039 9225
rect 10065 9199 10066 9225
rect 10038 9193 10066 9199
rect 10318 9225 10346 9983
rect 10878 10010 10906 10015
rect 10990 10010 11018 10015
rect 10878 10009 10990 10010
rect 10878 9983 10879 10009
rect 10905 9983 10990 10009
rect 10878 9982 10990 9983
rect 10878 9977 10906 9982
rect 10990 9963 11018 9982
rect 10318 9199 10319 9225
rect 10345 9199 10346 9225
rect 9534 8807 9535 8833
rect 9561 8807 9562 8833
rect 9534 8777 9562 8807
rect 9534 8751 9535 8777
rect 9561 8751 9562 8777
rect 9142 8415 9143 8441
rect 9169 8415 9170 8441
rect 9142 8162 9170 8415
rect 8694 8134 9170 8162
rect 8694 8049 8722 8134
rect 8694 8023 8695 8049
rect 8721 8023 8722 8049
rect 8694 7266 8722 8023
rect 9142 7658 9170 8134
rect 9422 8442 9450 8447
rect 9534 8442 9562 8751
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9422 8441 9562 8442
rect 9422 8415 9423 8441
rect 9449 8415 9535 8441
rect 9561 8415 9562 8441
rect 9422 8414 9562 8415
rect 9422 8050 9450 8414
rect 9534 8409 9562 8414
rect 10318 8441 10346 9199
rect 10318 8415 10319 8441
rect 10345 8415 10346 8441
rect 9422 7993 9450 8022
rect 9422 7967 9423 7993
rect 9449 7967 9450 7993
rect 9422 7961 9450 7967
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9142 7611 9170 7630
rect 10038 7713 10066 7719
rect 10038 7687 10039 7713
rect 10065 7687 10066 7713
rect 10038 7657 10066 7687
rect 10038 7631 10039 7657
rect 10065 7631 10066 7657
rect 8694 7200 8722 7238
rect 9590 7602 9618 7607
rect 9590 7265 9618 7574
rect 10038 7602 10066 7631
rect 10318 7658 10346 8415
rect 10318 7611 10346 7630
rect 11102 9617 11130 10375
rect 11102 9591 11103 9617
rect 11129 9591 11130 9617
rect 11102 9282 11130 9591
rect 11382 10402 11410 10407
rect 11494 10402 11522 10767
rect 13118 10793 13146 11158
rect 14182 11186 14210 33586
rect 14518 25242 14546 25247
rect 14518 24905 14546 25214
rect 15246 24961 15274 24967
rect 15246 24935 15247 24961
rect 15273 24935 15274 24961
rect 14518 24879 14519 24905
rect 14545 24879 14546 24905
rect 14518 24121 14546 24879
rect 15134 24906 15162 24911
rect 15246 24906 15274 24935
rect 15134 24905 15274 24906
rect 15134 24879 15135 24905
rect 15161 24879 15274 24905
rect 15134 24878 15274 24879
rect 15078 24513 15106 24519
rect 15078 24487 15079 24513
rect 15105 24487 15106 24513
rect 14518 24095 14519 24121
rect 14545 24095 14546 24121
rect 14518 23506 14546 24095
rect 14518 23473 14546 23478
rect 14574 24402 14602 24407
rect 14574 23337 14602 24374
rect 14574 23311 14575 23337
rect 14601 23311 14602 23337
rect 14574 22554 14602 23311
rect 15078 23729 15106 24487
rect 15134 24514 15162 24878
rect 15246 24514 15274 24519
rect 15470 24514 15498 24519
rect 15134 24513 15498 24514
rect 15134 24487 15247 24513
rect 15273 24487 15471 24513
rect 15497 24487 15498 24513
rect 15134 24486 15498 24487
rect 15134 24346 15162 24486
rect 15246 24481 15274 24486
rect 15470 24481 15498 24486
rect 15134 24313 15162 24318
rect 15134 24234 15162 24239
rect 15134 24178 15162 24206
rect 15246 24178 15274 24183
rect 15134 24177 15274 24178
rect 15134 24151 15247 24177
rect 15273 24151 15274 24177
rect 15134 24150 15274 24151
rect 15134 24121 15162 24150
rect 15134 24095 15135 24121
rect 15161 24095 15162 24121
rect 15134 24089 15162 24095
rect 15078 23703 15079 23729
rect 15105 23703 15106 23729
rect 15078 23506 15106 23703
rect 15246 23730 15274 24150
rect 15470 23730 15498 23735
rect 15246 23729 15470 23730
rect 15246 23703 15247 23729
rect 15273 23703 15470 23729
rect 15246 23702 15470 23703
rect 15246 23697 15274 23702
rect 15470 23664 15498 23702
rect 16814 23730 16842 23735
rect 14798 22945 14826 22951
rect 14798 22919 14799 22945
rect 14825 22919 14826 22945
rect 14798 22554 14826 22919
rect 15078 22946 15106 23478
rect 15078 22913 15106 22918
rect 15302 23393 15330 23399
rect 15302 23367 15303 23393
rect 15329 23367 15330 23393
rect 15302 23337 15330 23367
rect 15302 23311 15303 23337
rect 15329 23311 15330 23337
rect 15302 22946 15330 23311
rect 15470 22946 15498 22951
rect 15302 22945 15498 22946
rect 15302 22919 15303 22945
rect 15329 22919 15471 22945
rect 15497 22919 15498 22945
rect 15302 22918 15498 22919
rect 14350 22553 14826 22554
rect 14350 22527 14575 22553
rect 14601 22527 14826 22553
rect 14350 22526 14826 22527
rect 14350 21042 14378 22526
rect 14574 22521 14602 22526
rect 14798 22161 14826 22526
rect 14798 22135 14799 22161
rect 14825 22135 14826 22161
rect 14798 22129 14826 22135
rect 15302 22609 15330 22918
rect 15470 22913 15498 22918
rect 16254 22946 16282 22951
rect 15302 22583 15303 22609
rect 15329 22583 15330 22609
rect 15302 22553 15330 22583
rect 15302 22527 15303 22553
rect 15329 22527 15330 22553
rect 15302 22162 15330 22527
rect 16254 22554 16282 22918
rect 16814 22946 16842 23702
rect 16926 22946 16954 22951
rect 16814 22945 16954 22946
rect 16814 22919 16815 22945
rect 16841 22919 16927 22945
rect 16953 22919 16954 22945
rect 16814 22918 16954 22919
rect 16814 22913 16842 22918
rect 15470 22162 15498 22167
rect 15302 22161 15498 22162
rect 15302 22135 15303 22161
rect 15329 22135 15471 22161
rect 15497 22135 15498 22161
rect 15302 22134 15498 22135
rect 15302 22129 15330 22134
rect 15414 21854 15442 22134
rect 15470 22129 15498 22134
rect 16254 22161 16282 22526
rect 16254 22135 16255 22161
rect 16281 22135 16282 22161
rect 16254 22129 16282 22135
rect 16702 22554 16730 22559
rect 15358 21826 15442 21854
rect 16702 21854 16730 22526
rect 16814 22554 16842 22559
rect 16814 22507 16842 22526
rect 16926 22554 16954 22918
rect 16758 22162 16786 22167
rect 16926 22162 16954 22526
rect 16758 22161 16954 22162
rect 16758 22135 16759 22161
rect 16785 22135 16927 22161
rect 16953 22135 16954 22161
rect 16758 22134 16954 22135
rect 16758 22129 16786 22134
rect 16926 22129 16954 22134
rect 16702 21826 16842 21854
rect 15358 21825 15386 21826
rect 15358 21799 15359 21825
rect 15385 21799 15386 21825
rect 14574 21769 14602 21775
rect 14574 21743 14575 21769
rect 14601 21743 14602 21769
rect 14574 21378 14602 21743
rect 15358 21769 15386 21799
rect 15358 21743 15359 21769
rect 15385 21743 15386 21769
rect 14798 21378 14826 21383
rect 14574 21377 14826 21378
rect 14574 21351 14799 21377
rect 14825 21351 14826 21377
rect 14574 21350 14826 21351
rect 14798 21098 14826 21350
rect 14350 21009 14378 21014
rect 14574 21042 14602 21047
rect 14574 20985 14602 21014
rect 14574 20959 14575 20985
rect 14601 20959 14602 20985
rect 14574 20953 14602 20959
rect 14294 20258 14322 20263
rect 14294 20201 14322 20230
rect 14294 20175 14295 20201
rect 14321 20175 14322 20201
rect 14294 20169 14322 20175
rect 14798 19809 14826 21070
rect 15358 21378 15386 21743
rect 16814 21770 16842 21826
rect 16814 21737 16842 21742
rect 17094 21770 17122 21775
rect 17094 21723 17122 21742
rect 15470 21378 15498 21383
rect 15358 21377 15498 21378
rect 15358 21351 15359 21377
rect 15385 21351 15471 21377
rect 15497 21351 15498 21377
rect 15358 21350 15498 21351
rect 15358 21041 15386 21350
rect 15470 21345 15498 21350
rect 16254 21377 16282 21383
rect 16254 21351 16255 21377
rect 16281 21351 16282 21377
rect 15358 21015 15359 21041
rect 15385 21015 15386 21041
rect 15358 20985 15386 21015
rect 16254 21042 16282 21351
rect 15358 20959 15359 20985
rect 15385 20959 15386 20985
rect 14798 19783 14799 19809
rect 14825 19783 14826 19809
rect 14294 19418 14322 19423
rect 14294 19371 14322 19390
rect 14798 19418 14826 19783
rect 14798 19385 14826 19390
rect 14910 20593 14938 20599
rect 14910 20567 14911 20593
rect 14937 20567 14938 20593
rect 14910 19026 14938 20567
rect 14574 19025 14938 19026
rect 14574 18999 14911 19025
rect 14937 18999 14938 19025
rect 14574 18998 14938 18999
rect 14574 18633 14602 18998
rect 14574 18607 14575 18633
rect 14601 18607 14602 18633
rect 14574 17849 14602 18607
rect 14574 17823 14575 17849
rect 14601 17823 14602 17849
rect 14574 17817 14602 17823
rect 14798 18241 14826 18998
rect 14910 18993 14938 18998
rect 15358 20594 15386 20959
rect 15918 20986 15946 20991
rect 15470 20594 15498 20599
rect 15358 20593 15498 20594
rect 15358 20567 15359 20593
rect 15385 20567 15471 20593
rect 15497 20567 15498 20593
rect 15358 20566 15498 20567
rect 15358 20257 15386 20566
rect 15470 20561 15498 20566
rect 15358 20231 15359 20257
rect 15385 20231 15386 20257
rect 15358 20202 15386 20231
rect 15358 19026 15386 20174
rect 15918 19809 15946 20958
rect 15918 19783 15919 19809
rect 15945 19783 15946 19809
rect 15918 19754 15946 19783
rect 15470 19753 15946 19754
rect 15470 19727 15919 19753
rect 15945 19727 15946 19753
rect 15470 19726 15946 19727
rect 15470 19474 15498 19726
rect 15918 19721 15946 19726
rect 16254 19809 16282 21014
rect 16534 21098 16562 21103
rect 16534 20594 16562 21070
rect 16758 21042 16786 21047
rect 16758 20986 16786 21014
rect 16814 20986 16842 20991
rect 16758 20985 16898 20986
rect 16758 20959 16815 20985
rect 16841 20959 16898 20985
rect 16758 20958 16898 20959
rect 16814 20953 16842 20958
rect 16534 20593 16842 20594
rect 16534 20567 16535 20593
rect 16561 20567 16842 20593
rect 16534 20566 16842 20567
rect 16534 20561 16562 20566
rect 16814 20201 16842 20566
rect 16814 20175 16815 20201
rect 16841 20175 16842 20201
rect 16814 20169 16842 20175
rect 16254 19783 16255 19809
rect 16281 19783 16282 19809
rect 15470 19417 15498 19446
rect 15470 19391 15471 19417
rect 15497 19391 15498 19417
rect 15470 19385 15498 19391
rect 15470 19026 15498 19031
rect 15358 19025 15498 19026
rect 15358 18999 15359 19025
rect 15385 18999 15471 19025
rect 15497 18999 15498 19025
rect 15358 18998 15498 18999
rect 15358 18993 15386 18998
rect 14798 18215 14799 18241
rect 14825 18215 14826 18241
rect 14798 17457 14826 18215
rect 15470 18689 15498 18998
rect 15470 18663 15471 18689
rect 15497 18663 15498 18689
rect 15470 18633 15498 18663
rect 15470 18607 15471 18633
rect 15497 18607 15498 18633
rect 15470 17905 15498 18607
rect 16254 19025 16282 19783
rect 16254 18999 16255 19025
rect 16281 18999 16282 19025
rect 15470 17879 15471 17905
rect 15497 17879 15498 17905
rect 15470 17850 15498 17879
rect 15918 18241 15946 18247
rect 15918 18215 15919 18241
rect 15945 18215 15946 18241
rect 15918 18186 15946 18215
rect 15918 17850 15946 18158
rect 15470 17849 15946 17850
rect 15470 17823 15471 17849
rect 15497 17823 15946 17849
rect 15470 17822 15946 17823
rect 15470 17817 15498 17822
rect 14798 17431 14799 17457
rect 14825 17431 14826 17457
rect 14406 17065 14434 17071
rect 14406 17039 14407 17065
rect 14433 17039 14434 17065
rect 14406 16281 14434 17039
rect 14406 16255 14407 16281
rect 14433 16255 14434 16281
rect 14406 15974 14434 16255
rect 14798 16673 14826 17431
rect 15918 17458 15946 17822
rect 15918 17401 15946 17430
rect 15918 17375 15919 17401
rect 15945 17375 15946 17401
rect 15918 17369 15946 17375
rect 16254 18241 16282 18999
rect 16254 18215 16255 18241
rect 16281 18215 16282 18241
rect 16254 17457 16282 18215
rect 16870 19417 16898 20958
rect 16870 19391 16871 19417
rect 16897 19391 16898 19417
rect 16870 18633 16898 19391
rect 16870 18607 16871 18633
rect 16897 18607 16898 18633
rect 16870 17850 16898 18607
rect 16870 17849 17010 17850
rect 16870 17823 16871 17849
rect 16897 17823 17010 17849
rect 16870 17822 17010 17823
rect 16870 17817 16898 17822
rect 16254 17431 16255 17457
rect 16281 17431 16282 17457
rect 14798 16647 14799 16673
rect 14825 16647 14826 16673
rect 14406 15946 14602 15974
rect 14182 11153 14210 11158
rect 14574 15497 14602 15946
rect 14574 15471 14575 15497
rect 14601 15471 14602 15497
rect 14574 14713 14602 15471
rect 14574 14687 14575 14713
rect 14601 14687 14602 14713
rect 14574 13929 14602 14687
rect 14574 13903 14575 13929
rect 14601 13903 14602 13929
rect 14574 13145 14602 13903
rect 14574 13119 14575 13145
rect 14601 13119 14602 13145
rect 14574 12362 14602 13119
rect 14574 11577 14602 12334
rect 14574 11551 14575 11577
rect 14601 11551 14602 11577
rect 13118 10767 13119 10793
rect 13145 10767 13146 10793
rect 11382 10401 11522 10402
rect 11382 10375 11383 10401
rect 11409 10375 11495 10401
rect 11521 10375 11522 10401
rect 11382 10374 11522 10375
rect 11382 10010 11410 10374
rect 11494 10369 11522 10374
rect 12558 10401 12586 10407
rect 12558 10375 12559 10401
rect 12585 10375 12586 10401
rect 11382 9618 11410 9982
rect 11494 9618 11522 9623
rect 11382 9617 11522 9618
rect 11382 9591 11383 9617
rect 11409 9591 11495 9617
rect 11521 9591 11522 9617
rect 11382 9590 11522 9591
rect 11382 9585 11410 9590
rect 11494 9585 11522 9590
rect 12278 9618 12306 9623
rect 11102 8833 11130 9254
rect 11102 8807 11103 8833
rect 11129 8807 11130 8833
rect 11102 8049 11130 8807
rect 11494 9338 11522 9343
rect 11494 9281 11522 9310
rect 11494 9255 11495 9281
rect 11521 9255 11522 9281
rect 11494 9225 11522 9255
rect 11494 9199 11495 9225
rect 11521 9199 11522 9225
rect 11494 8497 11522 9199
rect 11718 9338 11746 9343
rect 11718 8833 11746 9310
rect 11718 8807 11719 8833
rect 11745 8807 11746 8833
rect 11718 8778 11746 8807
rect 12278 9282 12306 9590
rect 12558 9618 12586 10375
rect 12558 9585 12586 9590
rect 12838 10010 12866 10015
rect 12278 8833 12306 9254
rect 12838 9282 12866 9982
rect 13118 10010 13146 10767
rect 13790 10849 13818 10855
rect 13790 10823 13791 10849
rect 13817 10823 13818 10849
rect 13790 10793 13818 10823
rect 13790 10767 13791 10793
rect 13817 10767 13818 10793
rect 13118 9977 13146 9982
rect 13454 10402 13482 10407
rect 13790 10402 13818 10767
rect 13454 10401 13818 10402
rect 13454 10375 13455 10401
rect 13481 10375 13818 10401
rect 13454 10374 13818 10375
rect 14574 10794 14602 11551
rect 14798 15889 14826 16647
rect 14798 15863 14799 15889
rect 14825 15863 14826 15889
rect 14798 15105 14826 15863
rect 14798 15079 14799 15105
rect 14825 15079 14826 15105
rect 14798 14321 14826 15079
rect 14798 14295 14799 14321
rect 14825 14295 14826 14321
rect 14798 13537 14826 14295
rect 14798 13511 14799 13537
rect 14825 13511 14826 13537
rect 14798 12753 14826 13511
rect 14798 12727 14799 12753
rect 14825 12727 14826 12753
rect 14798 12026 14826 12727
rect 15246 17121 15274 17127
rect 15246 17095 15247 17121
rect 15273 17095 15274 17121
rect 15246 17065 15274 17095
rect 15246 17039 15247 17065
rect 15273 17039 15274 17065
rect 15246 16674 15274 17039
rect 15470 16674 15498 16679
rect 15246 16673 15498 16674
rect 15246 16647 15247 16673
rect 15273 16647 15471 16673
rect 15497 16647 15498 16673
rect 15246 16646 15498 16647
rect 15246 16337 15274 16646
rect 15470 16641 15498 16646
rect 16254 16673 16282 17431
rect 16814 17458 16842 17463
rect 16926 17458 16954 17463
rect 16842 17457 16954 17458
rect 16842 17431 16927 17457
rect 16953 17431 16954 17457
rect 16842 17430 16954 17431
rect 16814 17411 16842 17430
rect 16254 16647 16255 16673
rect 16281 16647 16282 16673
rect 15246 16311 15247 16337
rect 15273 16311 15274 16337
rect 15246 16281 15274 16311
rect 15246 16255 15247 16281
rect 15273 16255 15274 16281
rect 15246 15890 15274 16255
rect 15470 15890 15498 15895
rect 15246 15889 15498 15890
rect 15246 15863 15247 15889
rect 15273 15863 15471 15889
rect 15497 15863 15498 15889
rect 15246 15862 15498 15863
rect 15246 15553 15274 15862
rect 15470 15857 15498 15862
rect 16254 15889 16282 16647
rect 16254 15863 16255 15889
rect 16281 15863 16282 15889
rect 15246 15527 15247 15553
rect 15273 15527 15274 15553
rect 15246 15497 15274 15527
rect 15246 15471 15247 15497
rect 15273 15471 15274 15497
rect 15246 15106 15274 15471
rect 15470 15106 15498 15111
rect 15246 15105 15498 15106
rect 15246 15079 15247 15105
rect 15273 15079 15471 15105
rect 15497 15079 15498 15105
rect 15246 15078 15498 15079
rect 15246 14769 15274 15078
rect 15470 15073 15498 15078
rect 16254 15105 16282 15863
rect 16814 16282 16842 16287
rect 16814 15498 16842 16254
rect 16870 15666 16898 17430
rect 16926 17425 16954 17430
rect 16982 17065 17010 17822
rect 16982 17039 16983 17065
rect 17009 17039 17010 17065
rect 16926 16673 16954 16679
rect 16926 16647 16927 16673
rect 16953 16647 16954 16673
rect 16926 15834 16954 16647
rect 16982 16282 17010 17039
rect 16982 16216 17010 16254
rect 16926 15801 16954 15806
rect 16870 15638 17010 15666
rect 16814 15465 16842 15470
rect 16254 15079 16255 15105
rect 16281 15079 16282 15105
rect 15246 14743 15247 14769
rect 15273 14743 15274 14769
rect 15246 14713 15274 14743
rect 15246 14687 15247 14713
rect 15273 14687 15274 14713
rect 15246 14322 15274 14687
rect 15470 14322 15498 14327
rect 15246 14321 15498 14322
rect 15246 14295 15247 14321
rect 15273 14295 15471 14321
rect 15497 14295 15498 14321
rect 15246 14294 15498 14295
rect 15246 13985 15274 14294
rect 15470 14289 15498 14294
rect 16254 14321 16282 15079
rect 16254 14295 16255 14321
rect 16281 14295 16282 14321
rect 15246 13959 15247 13985
rect 15273 13959 15274 13985
rect 15246 13929 15274 13959
rect 15246 13903 15247 13929
rect 15273 13903 15274 13929
rect 15246 13538 15274 13903
rect 15470 13538 15498 13543
rect 15246 13537 15470 13538
rect 15246 13511 15247 13537
rect 15273 13511 15470 13537
rect 15246 13510 15470 13511
rect 15246 13201 15274 13510
rect 15470 13472 15498 13510
rect 16254 13537 16282 14295
rect 16254 13511 16255 13537
rect 16281 13511 16282 13537
rect 15246 13175 15247 13201
rect 15273 13175 15274 13201
rect 15246 13145 15274 13175
rect 15246 13119 15247 13145
rect 15273 13119 15274 13145
rect 15246 12754 15274 13119
rect 15470 12754 15498 12759
rect 15246 12753 15498 12754
rect 15246 12727 15247 12753
rect 15273 12727 15471 12753
rect 15497 12727 15498 12753
rect 15246 12726 15498 12727
rect 15246 12417 15274 12726
rect 15470 12721 15498 12726
rect 16254 12753 16282 13511
rect 16982 13146 17010 15638
rect 16982 13113 17010 13118
rect 17094 15498 17122 15503
rect 17094 14713 17122 15470
rect 17094 14687 17095 14713
rect 17121 14687 17122 14713
rect 17094 13929 17122 14687
rect 17094 13903 17095 13929
rect 17121 13903 17122 13929
rect 17094 13482 17122 13903
rect 17094 13145 17122 13454
rect 17094 13119 17095 13145
rect 17121 13119 17122 13145
rect 16254 12727 16255 12753
rect 16281 12727 16282 12753
rect 15246 12391 15247 12417
rect 15273 12391 15274 12417
rect 15134 12362 15162 12367
rect 15246 12362 15274 12391
rect 15134 12361 15274 12362
rect 15134 12335 15135 12361
rect 15161 12335 15274 12361
rect 15134 12334 15274 12335
rect 15134 12306 15162 12334
rect 15134 12273 15162 12278
rect 14798 11969 14826 11998
rect 16254 12026 16282 12727
rect 17094 12361 17122 13119
rect 17094 12335 17095 12361
rect 17121 12335 17122 12361
rect 17094 12329 17122 12335
rect 14798 11943 14799 11969
rect 14825 11943 14826 11969
rect 14798 11185 14826 11943
rect 15470 11970 15498 11975
rect 15470 11633 15498 11942
rect 15918 11970 15946 11975
rect 15918 11913 15946 11942
rect 16254 11969 16282 11998
rect 16254 11943 16255 11969
rect 16281 11943 16282 11969
rect 16254 11937 16282 11943
rect 15918 11887 15919 11913
rect 15945 11887 15946 11913
rect 15918 11881 15946 11887
rect 15470 11607 15471 11633
rect 15497 11607 15498 11633
rect 15470 11577 15498 11607
rect 15470 11551 15471 11577
rect 15497 11551 15498 11577
rect 14798 11159 14799 11185
rect 14825 11159 14826 11185
rect 14798 10794 14826 11159
rect 14574 10793 14826 10794
rect 14574 10767 14575 10793
rect 14601 10767 14826 10793
rect 14574 10766 14826 10767
rect 13454 10345 13482 10374
rect 13454 10319 13455 10345
rect 13481 10319 13482 10345
rect 13454 10066 13482 10319
rect 13454 9617 13482 10038
rect 14014 10066 14042 10071
rect 14014 10009 14042 10038
rect 14014 9983 14015 10009
rect 14041 9983 14042 10009
rect 14014 9977 14042 9983
rect 14294 10010 14322 10015
rect 14294 9963 14322 9982
rect 14574 10010 14602 10766
rect 14798 10401 14826 10766
rect 14798 10375 14799 10401
rect 14825 10375 14826 10401
rect 14798 10369 14826 10375
rect 15358 11186 15386 11191
rect 15470 11186 15498 11551
rect 17094 11858 17122 11863
rect 17094 11578 17122 11830
rect 15358 11185 15498 11186
rect 15358 11159 15359 11185
rect 15385 11159 15471 11185
rect 15497 11159 15498 11185
rect 15358 11158 15498 11159
rect 15358 10849 15386 11158
rect 15470 11153 15498 11158
rect 16534 11185 16562 11191
rect 16534 11159 16535 11185
rect 16561 11159 16562 11185
rect 15358 10823 15359 10849
rect 15385 10823 15386 10849
rect 15358 10793 15386 10823
rect 15358 10767 15359 10793
rect 15385 10767 15386 10793
rect 15358 10402 15386 10767
rect 15470 10402 15498 10407
rect 15358 10401 15498 10402
rect 15358 10375 15359 10401
rect 15385 10375 15471 10401
rect 15497 10375 15498 10401
rect 15358 10374 15498 10375
rect 14574 9977 14602 9982
rect 15358 10066 15386 10374
rect 15470 10369 15498 10374
rect 16478 10401 16506 10407
rect 16478 10375 16479 10401
rect 16505 10375 16506 10401
rect 15358 10009 15386 10038
rect 15358 9983 15359 10009
rect 15385 9983 15386 10009
rect 15358 9977 15386 9983
rect 13454 9591 13455 9617
rect 13481 9591 13482 9617
rect 13454 9562 13482 9591
rect 12838 9225 12866 9254
rect 12838 9199 12839 9225
rect 12865 9199 12866 9225
rect 12838 9193 12866 9199
rect 13398 9561 13482 9562
rect 13398 9535 13455 9561
rect 13481 9535 13482 9561
rect 13398 9534 13482 9535
rect 13398 9338 13426 9534
rect 13454 9529 13482 9534
rect 14798 9617 14826 9623
rect 14798 9591 14799 9617
rect 14825 9591 14826 9617
rect 13398 9226 13426 9310
rect 13510 9226 13538 9231
rect 13398 9225 13538 9226
rect 13398 9199 13399 9225
rect 13425 9199 13511 9225
rect 13537 9199 13538 9225
rect 13398 9198 13538 9199
rect 12278 8807 12279 8833
rect 12305 8807 12306 8833
rect 12278 8801 12306 8807
rect 13398 8833 13426 9198
rect 13510 9193 13538 9198
rect 14574 9226 14602 9231
rect 14798 9226 14826 9591
rect 15750 9617 15778 9623
rect 15750 9591 15751 9617
rect 15777 9591 15778 9617
rect 15750 9562 15778 9591
rect 16478 9618 16506 10375
rect 16534 10094 16562 11159
rect 16814 11186 16842 11191
rect 16926 11186 16954 11191
rect 16842 11185 16954 11186
rect 16842 11159 16927 11185
rect 16953 11159 16954 11185
rect 16842 11158 16954 11159
rect 16814 11139 16842 11158
rect 16814 10402 16842 10407
rect 16926 10402 16954 11158
rect 17094 10793 17122 11550
rect 17094 10767 17095 10793
rect 17121 10767 17122 10793
rect 17094 10761 17122 10767
rect 16814 10401 16954 10402
rect 16814 10375 16815 10401
rect 16841 10375 16927 10401
rect 16953 10375 16954 10401
rect 16814 10374 16954 10375
rect 16814 10369 16842 10374
rect 16534 10066 16786 10094
rect 16534 9618 16562 9623
rect 16478 9617 16562 9618
rect 16478 9591 16535 9617
rect 16561 9591 16562 9617
rect 16478 9590 16562 9591
rect 14574 9225 14826 9226
rect 14574 9199 14575 9225
rect 14601 9199 14826 9225
rect 14574 9198 14826 9199
rect 13398 8807 13399 8833
rect 13425 8807 13426 8833
rect 11774 8778 11802 8783
rect 11718 8777 11802 8778
rect 11718 8751 11775 8777
rect 11801 8751 11802 8777
rect 11718 8750 11802 8751
rect 11774 8745 11802 8750
rect 13398 8777 13426 8807
rect 13398 8751 13399 8777
rect 13425 8751 13426 8777
rect 13398 8745 13426 8751
rect 11494 8471 11495 8497
rect 11521 8471 11522 8497
rect 11494 8441 11522 8471
rect 14014 8497 14042 8503
rect 14014 8471 14015 8497
rect 14041 8471 14042 8497
rect 11494 8415 11495 8441
rect 11521 8415 11522 8441
rect 11102 8023 11103 8049
rect 11129 8023 11130 8049
rect 10038 7569 10066 7574
rect 9590 7239 9591 7265
rect 9617 7239 9618 7265
rect 9590 7209 9618 7239
rect 11102 7265 11130 8023
rect 11382 8050 11410 8055
rect 11494 8050 11522 8415
rect 13118 8441 13146 8447
rect 13118 8415 13119 8441
rect 13145 8415 13146 8441
rect 11382 8049 11522 8050
rect 11382 8023 11383 8049
rect 11409 8023 11495 8049
rect 11521 8023 11522 8049
rect 11382 8022 11522 8023
rect 11382 8017 11410 8022
rect 11494 7713 11522 8022
rect 11494 7687 11495 7713
rect 11521 7687 11522 7713
rect 11494 7657 11522 7687
rect 11494 7631 11495 7657
rect 11521 7631 11522 7657
rect 11494 7602 11522 7631
rect 11102 7239 11103 7265
rect 11129 7239 11130 7265
rect 11102 7233 11130 7239
rect 11382 7266 11410 7271
rect 11494 7266 11522 7574
rect 11382 7265 11522 7266
rect 11382 7239 11383 7265
rect 11409 7239 11495 7265
rect 11521 7239 11522 7265
rect 11382 7238 11522 7239
rect 11382 7233 11410 7238
rect 11494 7233 11522 7238
rect 12558 8049 12586 8055
rect 12558 8023 12559 8049
rect 12585 8023 12586 8049
rect 12558 7602 12586 8023
rect 12558 7265 12586 7574
rect 12558 7239 12559 7265
rect 12585 7239 12586 7265
rect 12558 7233 12586 7239
rect 13118 7657 13146 8415
rect 14014 8441 14042 8471
rect 14014 8415 14015 8441
rect 14041 8415 14042 8441
rect 13118 7631 13119 7657
rect 13145 7631 13146 7657
rect 13118 7602 13146 7631
rect 8078 7182 8162 7183
rect 8078 6929 8106 7182
rect 8134 7177 8162 7182
rect 9590 7183 9591 7209
rect 9617 7183 9618 7209
rect 9590 7177 9618 7183
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 8078 6903 8079 6929
rect 8105 6903 8106 6929
rect 8078 6873 8106 6903
rect 10878 6929 10906 6935
rect 10878 6903 10879 6929
rect 10905 6903 10906 6929
rect 8078 6847 8079 6873
rect 8105 6847 8106 6873
rect 7182 6841 7210 6846
rect 8078 6841 8106 6847
rect 9814 6873 9842 6879
rect 9814 6847 9815 6873
rect 9841 6847 9842 6873
rect 2478 6425 2506 6454
rect 2478 6399 2479 6425
rect 2505 6399 2506 6425
rect 2478 6393 2506 6399
rect 2814 6454 2870 6482
rect 2030 4913 2058 5278
rect 2030 4887 2031 4913
rect 2057 4887 2058 4913
rect 2030 4857 2058 4887
rect 2030 4831 2031 4857
rect 2057 4831 2058 4857
rect 2030 4577 2058 4831
rect 2030 4551 2031 4577
rect 2057 4551 2058 4577
rect 2030 4521 2058 4551
rect 2030 4495 2031 4521
rect 2057 4495 2058 4521
rect 2030 4214 2058 4495
rect 1022 4103 1023 4129
rect 1049 4103 1050 4129
rect 1022 3737 1050 4103
rect 1022 3711 1023 3737
rect 1049 3711 1050 3737
rect 1022 3705 1050 3711
rect 1862 4186 2058 4214
rect 2086 6146 2114 6151
rect 2086 6089 2114 6118
rect 2814 6146 2842 6454
rect 2870 6449 2898 6454
rect 4158 6481 4186 6487
rect 4158 6455 4159 6481
rect 4185 6455 4186 6481
rect 4046 6426 4074 6431
rect 4158 6426 4186 6455
rect 4046 6425 4158 6426
rect 4046 6399 4047 6425
rect 4073 6399 4158 6425
rect 4046 6398 4158 6399
rect 4046 6393 4074 6398
rect 4158 6393 4186 6398
rect 4998 6481 5026 6487
rect 4998 6455 4999 6481
rect 5025 6455 5026 6481
rect 2086 6063 2087 6089
rect 2113 6063 2114 6089
rect 2086 5697 2114 6063
rect 2534 6090 2562 6095
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2086 5671 2087 5697
rect 2113 5671 2114 5697
rect 2086 5641 2114 5671
rect 2086 5615 2087 5641
rect 2113 5615 2114 5641
rect 2086 5361 2114 5615
rect 2086 5335 2087 5361
rect 2113 5335 2114 5361
rect 2086 5305 2114 5335
rect 2086 5279 2087 5305
rect 2113 5279 2114 5305
rect 2086 4914 2114 5279
rect 2534 5305 2562 6062
rect 2814 6089 2842 6118
rect 3038 6146 3066 6151
rect 2814 6063 2815 6089
rect 2841 6063 2842 6089
rect 2814 6057 2842 6063
rect 2870 6090 2898 6095
rect 2870 5697 2898 6062
rect 3038 6089 3066 6118
rect 3038 6063 3039 6089
rect 3065 6063 3066 6089
rect 3038 6057 3066 6063
rect 2870 5671 2871 5697
rect 2897 5671 2898 5697
rect 2870 5665 2898 5671
rect 3318 5698 3346 5703
rect 3542 5698 3570 5703
rect 3318 5697 3570 5698
rect 3318 5671 3319 5697
rect 3345 5671 3543 5697
rect 3569 5671 3570 5697
rect 3318 5670 3570 5671
rect 2534 5279 2535 5305
rect 2561 5279 2562 5305
rect 2534 5273 2562 5279
rect 2814 5306 2842 5311
rect 2814 5259 2842 5278
rect 3038 5306 3066 5311
rect 3038 5259 3066 5278
rect 3318 5306 3346 5670
rect 3542 5665 3570 5670
rect 4998 5698 5026 6455
rect 5278 6481 5306 6487
rect 5278 6455 5279 6481
rect 5305 6455 5306 6481
rect 5278 6426 5306 6455
rect 6454 6482 6482 6487
rect 6454 6435 6482 6454
rect 7014 6482 7042 6487
rect 5278 6379 5306 6398
rect 5838 6426 5866 6431
rect 5838 6145 5866 6398
rect 5838 6119 5839 6145
rect 5865 6119 5866 6145
rect 5838 6090 5866 6119
rect 4998 5665 5026 5670
rect 5558 5698 5586 5703
rect 5558 5651 5586 5670
rect 3318 5273 3346 5278
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2086 4214 2114 4886
rect 2870 4913 2898 4919
rect 2870 4887 2871 4913
rect 2897 4887 2898 4913
rect 2534 4522 2562 4527
rect 2534 4475 2562 4494
rect 2870 4522 2898 4887
rect 2870 4489 2898 4494
rect 3318 4914 3346 4919
rect 3318 4577 3346 4886
rect 3542 4914 3570 4919
rect 3542 4867 3570 4886
rect 3318 4551 3319 4577
rect 3345 4551 3346 4577
rect 3318 4521 3346 4551
rect 3318 4495 3319 4521
rect 3345 4495 3346 4521
rect 3318 4489 3346 4495
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 5838 4214 5866 6062
rect 7014 6089 7042 6454
rect 7798 6481 7826 6487
rect 7798 6455 7799 6481
rect 7825 6455 7826 6481
rect 7798 6425 7826 6455
rect 7798 6399 7799 6425
rect 7825 6399 7826 6425
rect 7518 6146 7546 6151
rect 7518 6145 7602 6146
rect 7518 6119 7519 6145
rect 7545 6119 7602 6145
rect 7518 6118 7602 6119
rect 7518 6113 7546 6118
rect 7014 6063 7015 6089
rect 7041 6063 7042 6089
rect 6118 5698 6146 5703
rect 6118 5305 6146 5670
rect 6454 5697 6482 5703
rect 6454 5671 6455 5697
rect 6481 5671 6482 5697
rect 6454 5641 6482 5671
rect 6454 5615 6455 5641
rect 6481 5615 6482 5641
rect 6118 5279 6119 5305
rect 6145 5279 6146 5305
rect 6118 4410 6146 5279
rect 6398 5306 6426 5311
rect 6454 5306 6482 5615
rect 6510 5306 6538 5311
rect 6398 5305 6538 5306
rect 6398 5279 6399 5305
rect 6425 5279 6511 5305
rect 6537 5279 6538 5305
rect 6398 5278 6538 5279
rect 6398 5273 6426 5278
rect 6510 5082 6538 5278
rect 7014 5138 7042 6063
rect 7574 6090 7602 6118
rect 7574 6043 7602 6062
rect 7798 6090 7826 6399
rect 8974 6481 9002 6487
rect 8974 6455 8975 6481
rect 9001 6455 9002 6481
rect 7798 5697 7826 6062
rect 8470 6089 8498 6095
rect 8470 6063 8471 6089
rect 8497 6063 8498 6089
rect 8470 5922 8498 6063
rect 8470 5889 8498 5894
rect 8974 5922 9002 6455
rect 7798 5671 7799 5697
rect 7825 5671 7826 5697
rect 7798 5641 7826 5671
rect 8974 5697 9002 5894
rect 8974 5671 8975 5697
rect 9001 5671 9002 5697
rect 8974 5665 9002 5671
rect 9534 6482 9562 6487
rect 9534 5922 9562 6454
rect 9534 5697 9562 5894
rect 9534 5671 9535 5697
rect 9561 5671 9562 5697
rect 7798 5615 7799 5641
rect 7825 5615 7826 5641
rect 7014 5105 7042 5110
rect 7518 5305 7546 5311
rect 7798 5306 7826 5615
rect 7966 5306 7994 5311
rect 7518 5279 7519 5305
rect 7545 5279 7546 5305
rect 7518 5138 7546 5279
rect 7518 5105 7546 5110
rect 7686 5305 7994 5306
rect 7686 5279 7799 5305
rect 7825 5279 7967 5305
rect 7993 5279 7994 5305
rect 7686 5278 7994 5279
rect 6342 4522 6370 4527
rect 6510 4522 6538 5054
rect 6342 4521 6538 4522
rect 6342 4495 6343 4521
rect 6369 4495 6511 4521
rect 6537 4495 6538 4521
rect 6342 4494 6538 4495
rect 6342 4489 6370 4494
rect 6510 4489 6538 4494
rect 7014 4521 7042 4527
rect 7014 4495 7015 4521
rect 7041 4495 7042 4521
rect 6118 4377 6146 4382
rect 2086 4186 2170 4214
rect 1862 4129 1890 4186
rect 1862 4103 1863 4129
rect 1889 4103 1890 4129
rect 1862 4073 1890 4103
rect 1862 4047 1863 4073
rect 1889 4047 1890 4073
rect 1862 3793 1890 4047
rect 1862 3767 1863 3793
rect 1889 3767 1890 3793
rect 1862 3737 1890 3767
rect 1862 3711 1863 3737
rect 1889 3711 1890 3737
rect 1862 3009 1890 3711
rect 1862 2983 1863 3009
rect 1889 2983 1890 3009
rect 910 2953 938 2959
rect 910 2927 911 2953
rect 937 2927 938 2953
rect 910 2561 938 2927
rect 1862 2953 1890 2983
rect 1862 2927 1863 2953
rect 1889 2927 1890 2953
rect 1862 2921 1890 2927
rect 910 2535 911 2561
rect 937 2535 938 2561
rect 910 2226 938 2535
rect 2086 2562 2114 2567
rect 2142 2562 2170 4186
rect 5782 4186 5866 4214
rect 5782 4130 5810 4186
rect 5894 4130 5922 4135
rect 5782 4129 5922 4130
rect 5782 4103 5783 4129
rect 5809 4103 5895 4129
rect 5921 4103 5922 4129
rect 5782 4102 5922 4103
rect 5782 3794 5810 4102
rect 5894 4097 5922 4102
rect 6454 4130 6482 4135
rect 6454 4083 6482 4102
rect 7014 4130 7042 4495
rect 7518 4521 7546 4527
rect 7518 4495 7519 4521
rect 7545 4495 7546 4521
rect 7518 4410 7546 4495
rect 7518 4377 7546 4382
rect 7686 4214 7714 5278
rect 7798 5273 7826 5278
rect 7966 5273 7994 5278
rect 8078 5138 8106 5143
rect 7742 5082 7770 5087
rect 7742 4522 7770 5054
rect 8078 4913 8106 5110
rect 9478 5138 9506 5143
rect 8078 4887 8079 4913
rect 8105 4887 8106 4913
rect 8078 4881 8106 4887
rect 8246 5082 8274 5087
rect 8246 4914 8274 5054
rect 8470 4914 8498 4919
rect 8246 4913 8498 4914
rect 8246 4887 8247 4913
rect 8273 4887 8471 4913
rect 8497 4887 8498 4913
rect 8246 4886 8498 4887
rect 8246 4881 8274 4886
rect 7966 4522 7994 4527
rect 7742 4521 7994 4522
rect 7742 4495 7743 4521
rect 7769 4495 7967 4521
rect 7993 4495 7994 4521
rect 7742 4494 7994 4495
rect 7742 4489 7770 4494
rect 7966 4489 7994 4494
rect 7798 4410 7826 4415
rect 7686 4186 7770 4214
rect 5838 3794 5866 3799
rect 5782 3793 5866 3794
rect 5782 3767 5839 3793
rect 5865 3767 5866 3793
rect 5782 3766 5866 3767
rect 5838 3737 5866 3766
rect 5838 3711 5839 3737
rect 5865 3711 5866 3737
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 5838 3009 5866 3711
rect 7014 3738 7042 4102
rect 7014 3691 7042 3710
rect 7518 3738 7546 3743
rect 5838 2983 5839 3009
rect 5865 2983 5866 3009
rect 5838 2953 5866 2983
rect 5838 2927 5839 2953
rect 5865 2927 5866 2953
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 2086 2561 2170 2562
rect 2086 2535 2087 2561
rect 2113 2535 2170 2561
rect 2086 2534 2170 2535
rect 3766 2562 3794 2567
rect 2086 2505 2114 2534
rect 2086 2479 2087 2505
rect 2113 2479 2114 2505
rect 2086 2473 2114 2479
rect 910 2193 938 2198
rect 3766 2225 3794 2534
rect 5278 2562 5306 2567
rect 5278 2505 5306 2534
rect 5838 2562 5866 2927
rect 7014 2953 7042 2959
rect 7014 2927 7015 2953
rect 7041 2927 7042 2953
rect 5838 2529 5866 2534
rect 6230 2562 6258 2567
rect 5278 2479 5279 2505
rect 5305 2479 5306 2505
rect 5278 2473 5306 2479
rect 3766 2199 3767 2225
rect 3793 2199 3794 2225
rect 2870 2169 2898 2175
rect 2870 2143 2871 2169
rect 2897 2143 2898 2169
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 2086 1778 2114 1783
rect 2086 400 2114 1750
rect 2870 1778 2898 2143
rect 3766 2169 3794 2199
rect 3766 2143 3767 2169
rect 3793 2143 3794 2169
rect 3766 2137 3794 2143
rect 2870 1731 2898 1750
rect 3822 1777 3850 1783
rect 3822 1751 3823 1777
rect 3849 1751 3850 1777
rect 3822 1722 3850 1751
rect 3822 1656 3850 1694
rect 6230 400 6258 2534
rect 7014 2562 7042 2927
rect 7518 2954 7546 3710
rect 7742 3010 7770 4186
rect 7798 4130 7826 4382
rect 7798 4064 7826 4102
rect 8246 4130 8274 4135
rect 8358 4130 8386 4886
rect 8470 4881 8498 4886
rect 9478 4214 9506 5110
rect 9534 4913 9562 5671
rect 9814 6482 9842 6847
rect 10878 6873 10906 6903
rect 12446 6929 12474 6935
rect 12446 6903 12447 6929
rect 12473 6903 12474 6929
rect 10878 6847 10879 6873
rect 10905 6847 10906 6873
rect 9814 6146 9842 6454
rect 10430 6481 10458 6487
rect 10430 6455 10431 6481
rect 10457 6455 10458 6481
rect 10430 6426 10458 6455
rect 10430 6379 10458 6398
rect 10878 6426 10906 6847
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9814 6089 9842 6118
rect 9814 6063 9815 6089
rect 9841 6063 9842 6089
rect 9814 5305 9842 6063
rect 10878 6145 10906 6398
rect 10878 6119 10879 6145
rect 10905 6119 10906 6145
rect 10878 6090 10906 6119
rect 10878 6043 10906 6062
rect 11550 6873 11578 6879
rect 11550 6847 11551 6873
rect 11577 6847 11578 6873
rect 11550 6146 11578 6847
rect 12446 6873 12474 6903
rect 12446 6847 12447 6873
rect 12473 6847 12474 6873
rect 11550 6089 11578 6118
rect 11550 6063 11551 6089
rect 11577 6063 11578 6089
rect 10430 5697 10458 5703
rect 10430 5671 10431 5697
rect 10457 5671 10458 5697
rect 10430 5641 10458 5671
rect 10430 5615 10431 5641
rect 10457 5615 10458 5641
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9814 5279 9815 5305
rect 9841 5279 9842 5305
rect 9814 5273 9842 5279
rect 10374 5306 10402 5311
rect 10430 5306 10458 5615
rect 10486 5306 10514 5311
rect 10374 5305 10514 5306
rect 10374 5279 10375 5305
rect 10401 5279 10487 5305
rect 10513 5279 10514 5305
rect 10374 5278 10514 5279
rect 10374 5273 10402 5278
rect 9534 4887 9535 4913
rect 9561 4887 9562 4913
rect 9534 4881 9562 4887
rect 10430 4914 10458 4919
rect 10486 4914 10514 5278
rect 10430 4913 10514 4914
rect 10430 4887 10431 4913
rect 10457 4887 10514 4913
rect 10430 4886 10514 4887
rect 11550 5305 11578 6063
rect 11550 5279 11551 5305
rect 11577 5279 11578 5305
rect 10430 4857 10458 4886
rect 10430 4831 10431 4857
rect 10457 4831 10458 4857
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10038 4521 10066 4527
rect 10038 4495 10039 4521
rect 10065 4495 10066 4521
rect 10038 4466 10066 4495
rect 10038 4433 10066 4438
rect 10430 4522 10458 4831
rect 8470 4186 8498 4191
rect 9478 4186 9562 4214
rect 8470 4130 8498 4158
rect 8246 4129 8498 4130
rect 8246 4103 8247 4129
rect 8273 4103 8471 4129
rect 8497 4103 8498 4129
rect 8246 4102 8498 4103
rect 7742 2977 7770 2982
rect 7798 3738 7826 3743
rect 7966 3738 7994 3743
rect 7798 3737 7994 3738
rect 7798 3711 7799 3737
rect 7825 3711 7967 3737
rect 7993 3711 7994 3737
rect 7798 3710 7994 3711
rect 7798 3402 7826 3710
rect 7966 3705 7994 3710
rect 7574 2954 7602 2959
rect 7518 2926 7574 2954
rect 7574 2907 7602 2926
rect 7014 2169 7042 2534
rect 7014 2143 7015 2169
rect 7041 2143 7042 2169
rect 7014 1777 7042 2143
rect 7574 2170 7602 2175
rect 7686 2170 7714 2175
rect 7798 2170 7826 3374
rect 8246 3402 8274 4102
rect 8470 4097 8498 4102
rect 9254 4130 9282 4135
rect 8078 3345 8106 3351
rect 8078 3319 8079 3345
rect 8105 3319 8106 3345
rect 8078 2954 8106 3319
rect 8246 3345 8274 3374
rect 8246 3319 8247 3345
rect 8273 3319 8274 3345
rect 8246 3313 8274 3319
rect 8470 3402 8498 3407
rect 8470 3345 8498 3374
rect 8470 3319 8471 3345
rect 8497 3319 8498 3345
rect 8470 3313 8498 3319
rect 8078 2618 8106 2926
rect 8078 2561 8106 2590
rect 8078 2535 8079 2561
rect 8105 2535 8106 2561
rect 8078 2529 8106 2535
rect 8470 3010 8498 3015
rect 8470 2953 8498 2982
rect 8470 2927 8471 2953
rect 8497 2927 8498 2953
rect 8470 2562 8498 2927
rect 8470 2529 8498 2534
rect 8974 2562 9002 2567
rect 8974 2505 9002 2534
rect 8974 2479 8975 2505
rect 9001 2479 9002 2505
rect 8974 2473 9002 2479
rect 9254 2561 9282 4102
rect 9534 4129 9562 4186
rect 9534 4103 9535 4129
rect 9561 4103 9562 4129
rect 9534 3346 9562 4103
rect 10374 4130 10402 4135
rect 10374 4073 10402 4102
rect 10374 4047 10375 4073
rect 10401 4047 10402 4073
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9534 3299 9562 3318
rect 9814 3737 9842 3743
rect 9814 3711 9815 3737
rect 9841 3711 9842 3737
rect 9814 3346 9842 3711
rect 10374 3738 10402 4047
rect 10374 3705 10402 3710
rect 9814 2954 9842 3318
rect 10430 3345 10458 4494
rect 10878 4577 10906 4583
rect 10878 4551 10879 4577
rect 10905 4551 10906 4577
rect 10878 4522 10906 4551
rect 11550 4522 11578 5279
rect 12054 6481 12082 6487
rect 12054 6455 12055 6481
rect 12081 6455 12082 6481
rect 12054 5697 12082 6455
rect 12054 5671 12055 5697
rect 12081 5671 12082 5697
rect 11774 4914 11802 4919
rect 11774 4522 11802 4886
rect 12054 4914 12082 5671
rect 12446 6482 12474 6847
rect 13118 6873 13146 7574
rect 13118 6847 13119 6873
rect 13145 6847 13146 6873
rect 12446 6145 12474 6454
rect 12950 6482 12978 6487
rect 12950 6425 12978 6454
rect 12950 6399 12951 6425
rect 12977 6399 12978 6425
rect 12950 6393 12978 6399
rect 12446 6119 12447 6145
rect 12473 6119 12474 6145
rect 12446 6090 12474 6119
rect 12446 5361 12474 6062
rect 13118 6089 13146 6847
rect 13454 8049 13482 8055
rect 13454 8023 13455 8049
rect 13481 8023 13482 8049
rect 13454 7993 13482 8023
rect 13454 7967 13455 7993
rect 13481 7967 13482 7993
rect 13454 7265 13482 7967
rect 13454 7239 13455 7265
rect 13481 7239 13482 7265
rect 13454 7209 13482 7239
rect 13454 7183 13455 7209
rect 13481 7183 13482 7209
rect 13118 6063 13119 6089
rect 13145 6063 13146 6089
rect 12446 5335 12447 5361
rect 12473 5335 12474 5361
rect 12446 5305 12474 5335
rect 12446 5279 12447 5305
rect 12473 5279 12474 5305
rect 12446 5273 12474 5279
rect 12894 5697 12922 5703
rect 12894 5671 12895 5697
rect 12921 5671 12922 5697
rect 12894 5641 12922 5671
rect 12894 5615 12895 5641
rect 12921 5615 12922 5641
rect 12054 4867 12082 4886
rect 12838 4914 12866 4919
rect 10878 4475 10906 4494
rect 11270 4521 11802 4522
rect 11270 4495 11551 4521
rect 11577 4495 11802 4521
rect 11270 4494 11802 4495
rect 11270 4466 11298 4494
rect 11550 4489 11578 4494
rect 10878 3793 10906 3799
rect 10878 3767 10879 3793
rect 10905 3767 10906 3793
rect 10878 3738 10906 3767
rect 10878 3691 10906 3710
rect 11270 3737 11298 4438
rect 11270 3711 11271 3737
rect 11297 3711 11298 3737
rect 11270 3705 11298 3711
rect 11774 4129 11802 4494
rect 12390 4577 12418 4583
rect 12390 4551 12391 4577
rect 12417 4551 12418 4577
rect 12390 4522 12418 4551
rect 11774 4103 11775 4129
rect 11801 4103 11802 4129
rect 10430 3319 10431 3345
rect 10457 3319 10458 3345
rect 10430 3289 10458 3319
rect 10430 3263 10431 3289
rect 10457 3263 10458 3289
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9814 2921 9842 2926
rect 10038 2954 10066 2959
rect 10038 2907 10066 2926
rect 9254 2535 9255 2561
rect 9281 2535 9282 2561
rect 7574 2169 7826 2170
rect 7574 2143 7575 2169
rect 7601 2143 7687 2169
rect 7713 2143 7826 2169
rect 7574 2142 7826 2143
rect 9254 2170 9282 2535
rect 7574 2137 7602 2142
rect 7014 1751 7015 1777
rect 7041 1751 7042 1777
rect 7014 1745 7042 1751
rect 7574 1778 7602 1783
rect 7686 1778 7714 2142
rect 9254 2137 9282 2142
rect 9422 2618 9450 2623
rect 7574 1777 7714 1778
rect 7574 1751 7575 1777
rect 7601 1751 7687 1777
rect 7713 1751 7714 1777
rect 7574 1750 7714 1751
rect 7574 1722 7602 1750
rect 7686 1745 7714 1750
rect 9422 1778 9450 2590
rect 10430 2562 10458 3263
rect 11774 3345 11802 4103
rect 11774 3319 11775 3345
rect 11801 3319 11802 3345
rect 10430 2505 10458 2534
rect 10430 2479 10431 2505
rect 10457 2479 10458 2505
rect 10430 2473 10458 2479
rect 10766 3009 10794 3015
rect 10766 2983 10767 3009
rect 10793 2983 10794 3009
rect 10766 2953 10794 2983
rect 10766 2927 10767 2953
rect 10793 2927 10794 2953
rect 10766 2562 10794 2927
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10766 2225 10794 2534
rect 10766 2199 10767 2225
rect 10793 2199 10794 2225
rect 9814 2170 9842 2175
rect 9814 2123 9842 2142
rect 10766 2169 10794 2199
rect 10766 2143 10767 2169
rect 10793 2143 10794 2169
rect 10766 2137 10794 2143
rect 11550 2954 11578 2959
rect 11550 2562 11578 2926
rect 11550 2169 11578 2534
rect 11774 2561 11802 3319
rect 11774 2535 11775 2561
rect 11801 2535 11802 2561
rect 11774 2529 11802 2535
rect 12334 4186 12362 4191
rect 12334 3738 12362 4158
rect 12390 3794 12418 4494
rect 12446 3794 12474 3799
rect 12390 3793 12474 3794
rect 12390 3767 12447 3793
rect 12473 3767 12474 3793
rect 12390 3766 12474 3767
rect 12334 3009 12362 3710
rect 12334 2983 12335 3009
rect 12361 2983 12362 3009
rect 12334 2953 12362 2983
rect 12334 2927 12335 2953
rect 12361 2927 12362 2953
rect 11550 2143 11551 2169
rect 11577 2143 11578 2169
rect 11550 2137 11578 2143
rect 11102 2058 11130 2063
rect 9422 1731 9450 1750
rect 9590 1777 9618 1783
rect 9590 1751 9591 1777
rect 9617 1751 9618 1777
rect 7574 1689 7602 1694
rect 9590 1722 9618 1751
rect 9590 1689 9618 1694
rect 9814 1777 9842 1783
rect 9814 1751 9815 1777
rect 9841 1751 9842 1777
rect 9814 1722 9842 1751
rect 9814 1689 9842 1694
rect 10374 1778 10402 1783
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10374 400 10402 1750
rect 11102 1777 11130 2030
rect 11102 1751 11103 1777
rect 11129 1751 11130 1777
rect 11102 1745 11130 1751
rect 12278 1778 12306 1783
rect 12334 1778 12362 2927
rect 12446 3737 12474 3766
rect 12446 3711 12447 3737
rect 12473 3711 12474 3737
rect 12446 2225 12474 3711
rect 12838 3737 12866 4886
rect 12894 4913 12922 5615
rect 12894 4887 12895 4913
rect 12921 4887 12922 4913
rect 12894 4857 12922 4887
rect 12894 4831 12895 4857
rect 12921 4831 12922 4857
rect 12894 4214 12922 4831
rect 13118 5305 13146 6063
rect 13118 5279 13119 5305
rect 13145 5279 13146 5305
rect 13118 4914 13146 5279
rect 13118 4522 13146 4886
rect 13398 6481 13426 6487
rect 13398 6455 13399 6481
rect 13425 6455 13426 6481
rect 13398 5697 13426 6455
rect 13454 6482 13482 7183
rect 13454 6449 13482 6454
rect 14014 7713 14042 8415
rect 14014 7687 14015 7713
rect 14041 7687 14042 7713
rect 14014 7657 14042 7687
rect 14014 7631 14015 7657
rect 14041 7631 14042 7657
rect 14014 6929 14042 7631
rect 14014 6903 14015 6929
rect 14041 6903 14042 6929
rect 14014 6873 14042 6903
rect 14014 6847 14015 6873
rect 14041 6847 14042 6873
rect 14014 6482 14042 6847
rect 14574 8441 14602 9198
rect 14574 8415 14575 8441
rect 14601 8415 14602 8441
rect 14574 7657 14602 8415
rect 14574 7631 14575 7657
rect 14601 7631 14602 7657
rect 14574 6873 14602 7631
rect 14574 6847 14575 6873
rect 14601 6847 14602 6873
rect 14014 6145 14042 6454
rect 14238 6482 14266 6487
rect 14238 6425 14266 6454
rect 14238 6399 14239 6425
rect 14265 6399 14266 6425
rect 14238 6393 14266 6399
rect 14014 6119 14015 6145
rect 14041 6119 14042 6145
rect 14014 6089 14042 6119
rect 14014 6063 14015 6089
rect 14041 6063 14042 6089
rect 14014 6057 14042 6063
rect 14574 6089 14602 6847
rect 14574 6063 14575 6089
rect 14601 6063 14602 6089
rect 13398 5671 13399 5697
rect 13425 5671 13426 5697
rect 13398 4914 13426 5671
rect 13398 4867 13426 4886
rect 14014 5697 14042 5703
rect 14014 5671 14015 5697
rect 14041 5671 14042 5697
rect 14014 5642 14042 5671
rect 14182 5642 14210 5647
rect 14014 5641 14210 5642
rect 14014 5615 14183 5641
rect 14209 5615 14210 5641
rect 14014 5614 14210 5615
rect 14014 5361 14042 5614
rect 14182 5609 14210 5614
rect 14014 5335 14015 5361
rect 14041 5335 14042 5361
rect 14014 5305 14042 5335
rect 14014 5279 14015 5305
rect 14041 5279 14042 5305
rect 13958 4577 13986 4583
rect 13958 4551 13959 4577
rect 13985 4551 13986 4577
rect 13958 4522 13986 4551
rect 13118 4521 13258 4522
rect 13118 4495 13119 4521
rect 13145 4495 13258 4521
rect 13118 4494 13258 4495
rect 13118 4489 13146 4494
rect 12894 4186 12978 4214
rect 12950 4129 12978 4158
rect 12950 4103 12951 4129
rect 12977 4103 12978 4129
rect 12950 4073 12978 4103
rect 13230 4129 13258 4494
rect 13230 4103 13231 4129
rect 13257 4103 13258 4129
rect 13230 4097 13258 4103
rect 12950 4047 12951 4073
rect 12977 4047 12978 4073
rect 12950 4041 12978 4047
rect 12838 3711 12839 3737
rect 12865 3711 12866 3737
rect 12838 3705 12866 3711
rect 13958 3793 13986 4494
rect 14014 4214 14042 5279
rect 14574 5305 14602 6063
rect 14574 5279 14575 5305
rect 14601 5279 14602 5305
rect 14238 5026 14266 5031
rect 14238 4913 14266 4998
rect 14238 4887 14239 4913
rect 14265 4887 14266 4913
rect 14238 4857 14266 4887
rect 14238 4831 14239 4857
rect 14265 4831 14266 4857
rect 14238 4522 14266 4831
rect 14014 4186 14154 4214
rect 13958 3767 13959 3793
rect 13985 3767 13986 3793
rect 13958 3737 13986 3767
rect 13958 3711 13959 3737
rect 13985 3711 13986 3737
rect 13958 3705 13986 3711
rect 12446 2199 12447 2225
rect 12473 2199 12474 2225
rect 12446 2170 12474 2199
rect 12446 2123 12474 2142
rect 12894 3345 12922 3351
rect 12894 3319 12895 3345
rect 12921 3319 12922 3345
rect 12894 3289 12922 3319
rect 12894 3263 12895 3289
rect 12921 3263 12922 3289
rect 12894 2561 12922 3263
rect 12894 2535 12895 2561
rect 12921 2535 12922 2561
rect 12894 2505 12922 2535
rect 12894 2479 12895 2505
rect 12921 2479 12922 2505
rect 12894 2170 12922 2479
rect 12278 1777 12362 1778
rect 12278 1751 12279 1777
rect 12305 1751 12362 1777
rect 12278 1750 12362 1751
rect 12894 1778 12922 2142
rect 13118 3346 13146 3351
rect 13118 2953 13146 3318
rect 13398 3346 13426 3351
rect 13398 3299 13426 3318
rect 14126 3345 14154 4158
rect 14182 4130 14210 4135
rect 14238 4130 14266 4494
rect 14574 4914 14602 5279
rect 14574 4521 14602 4886
rect 14798 8833 14826 9198
rect 15470 9561 15778 9562
rect 15470 9535 15751 9561
rect 15777 9535 15778 9561
rect 15470 9534 15778 9535
rect 15470 9281 15498 9534
rect 15750 9529 15778 9534
rect 15470 9255 15471 9281
rect 15497 9255 15498 9281
rect 15470 9225 15498 9255
rect 15470 9199 15471 9225
rect 15497 9199 15498 9225
rect 14798 8807 14799 8833
rect 14825 8807 14826 8833
rect 14798 8049 14826 8807
rect 14798 8023 14799 8049
rect 14825 8023 14826 8049
rect 14798 7602 14826 8023
rect 15358 8834 15386 8839
rect 15470 8834 15498 9199
rect 15358 8833 15498 8834
rect 15358 8807 15359 8833
rect 15385 8807 15471 8833
rect 15497 8807 15498 8833
rect 15358 8806 15498 8807
rect 15358 8497 15386 8806
rect 15470 8801 15498 8806
rect 16534 8833 16562 9590
rect 16534 8807 16535 8833
rect 16561 8807 16562 8833
rect 15358 8471 15359 8497
rect 15385 8471 15386 8497
rect 15358 8441 15386 8471
rect 15358 8415 15359 8441
rect 15385 8415 15386 8441
rect 15358 8050 15386 8415
rect 15470 8050 15498 8055
rect 15358 8049 15498 8050
rect 15358 8023 15359 8049
rect 15385 8023 15471 8049
rect 15497 8023 15498 8049
rect 15358 8022 15498 8023
rect 15358 8017 15386 8022
rect 14798 7265 14826 7574
rect 15470 7994 15498 8022
rect 15470 7713 15498 7966
rect 15470 7687 15471 7713
rect 15497 7687 15498 7713
rect 15470 7657 15498 7687
rect 15470 7631 15471 7657
rect 15497 7631 15498 7657
rect 14798 7239 14799 7265
rect 14825 7239 14826 7265
rect 14798 6481 14826 7239
rect 14798 6455 14799 6481
rect 14825 6455 14826 6481
rect 14798 5697 14826 6455
rect 15358 7266 15386 7271
rect 15470 7266 15498 7631
rect 15358 7265 15498 7266
rect 15358 7239 15359 7265
rect 15385 7239 15471 7265
rect 15497 7239 15498 7265
rect 15358 7238 15498 7239
rect 15358 6929 15386 7238
rect 15470 7233 15498 7238
rect 16534 8050 16562 8807
rect 16534 7602 16562 8022
rect 16534 7265 16562 7574
rect 16534 7239 16535 7265
rect 16561 7239 16562 7265
rect 15358 6903 15359 6929
rect 15385 6903 15386 6929
rect 15358 6873 15386 6903
rect 15358 6847 15359 6873
rect 15385 6847 15386 6873
rect 15358 6482 15386 6847
rect 15470 6482 15498 6487
rect 15386 6481 15498 6482
rect 15386 6455 15471 6481
rect 15497 6455 15498 6481
rect 15386 6454 15498 6455
rect 15358 6145 15386 6454
rect 15470 6449 15498 6454
rect 16534 6481 16562 7239
rect 16534 6455 16535 6481
rect 16561 6455 16562 6481
rect 16534 6449 16562 6455
rect 15358 6119 15359 6145
rect 15385 6119 15386 6145
rect 15358 6089 15386 6119
rect 15358 6063 15359 6089
rect 15385 6063 15386 6089
rect 15358 6057 15386 6063
rect 16758 6090 16786 10066
rect 16926 9562 16954 10374
rect 16926 9529 16954 9534
rect 17094 10009 17122 10015
rect 17094 9983 17095 10009
rect 17121 9983 17122 10009
rect 17094 9225 17122 9983
rect 17094 9199 17095 9225
rect 17121 9199 17122 9225
rect 17094 8441 17122 9199
rect 17150 8834 17178 33586
rect 17598 33334 17730 33339
rect 17626 33306 17650 33334
rect 17678 33306 17702 33334
rect 17598 33301 17730 33306
rect 17598 32550 17730 32555
rect 17626 32522 17650 32550
rect 17678 32522 17702 32550
rect 17598 32517 17730 32522
rect 17598 31766 17730 31771
rect 17626 31738 17650 31766
rect 17678 31738 17702 31766
rect 17598 31733 17730 31738
rect 17598 30982 17730 30987
rect 17626 30954 17650 30982
rect 17678 30954 17702 30982
rect 17598 30949 17730 30954
rect 17598 30198 17730 30203
rect 17626 30170 17650 30198
rect 17678 30170 17702 30198
rect 17598 30165 17730 30170
rect 17598 29414 17730 29419
rect 17626 29386 17650 29414
rect 17678 29386 17702 29414
rect 17598 29381 17730 29386
rect 17598 28630 17730 28635
rect 17626 28602 17650 28630
rect 17678 28602 17702 28630
rect 17598 28597 17730 28602
rect 19782 27986 19810 27991
rect 17598 27846 17730 27851
rect 17626 27818 17650 27846
rect 17678 27818 17702 27846
rect 17598 27813 17730 27818
rect 17598 27062 17730 27067
rect 17626 27034 17650 27062
rect 17678 27034 17702 27062
rect 17598 27029 17730 27034
rect 19782 26866 19810 27958
rect 19950 26866 19978 26871
rect 19782 26865 19950 26866
rect 19782 26839 19783 26865
rect 19809 26839 19950 26865
rect 19782 26838 19950 26839
rect 19782 26833 19810 26838
rect 19950 26800 19978 26838
rect 20118 26809 20146 26815
rect 20118 26783 20119 26809
rect 20145 26783 20146 26809
rect 17598 26278 17730 26283
rect 17626 26250 17650 26278
rect 17678 26250 17702 26278
rect 17598 26245 17730 26250
rect 20118 26026 20146 26783
rect 20118 25993 20146 25998
rect 17598 25494 17730 25499
rect 17626 25466 17650 25494
rect 17678 25466 17702 25494
rect 17598 25461 17730 25466
rect 17598 24710 17730 24715
rect 17626 24682 17650 24710
rect 17678 24682 17702 24710
rect 17598 24677 17730 24682
rect 17598 23926 17730 23931
rect 17626 23898 17650 23926
rect 17678 23898 17702 23926
rect 17598 23893 17730 23898
rect 17598 23142 17730 23147
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17598 23109 17730 23114
rect 17262 22554 17290 22559
rect 17262 22507 17290 22526
rect 17486 22554 17514 22559
rect 17486 21826 17514 22526
rect 17598 22358 17730 22363
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17598 22325 17730 22330
rect 17990 21826 18018 21831
rect 17486 21825 18018 21826
rect 17486 21799 17991 21825
rect 18017 21799 18018 21825
rect 17486 21798 18018 21799
rect 17990 21769 18018 21798
rect 19278 21825 19306 21831
rect 19278 21799 19279 21825
rect 19305 21799 19306 21825
rect 17990 21743 17991 21769
rect 18017 21743 18018 21769
rect 17598 21574 17730 21579
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17598 21541 17730 21546
rect 17430 21377 17458 21383
rect 17430 21351 17431 21377
rect 17457 21351 17458 21377
rect 17430 21321 17458 21351
rect 17430 21295 17431 21321
rect 17457 21295 17458 21321
rect 17430 20593 17458 21295
rect 17934 21041 17962 21047
rect 17934 21015 17935 21041
rect 17961 21015 17962 21041
rect 17934 20985 17962 21015
rect 17934 20959 17935 20985
rect 17961 20959 17962 20985
rect 17598 20790 17730 20795
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17598 20757 17730 20762
rect 17430 20567 17431 20593
rect 17457 20567 17458 20593
rect 17430 20537 17458 20567
rect 17430 20511 17431 20537
rect 17457 20511 17458 20537
rect 17430 19809 17458 20511
rect 17934 20258 17962 20959
rect 17990 20986 18018 21743
rect 18438 21770 18466 21775
rect 18550 21770 18578 21775
rect 18466 21769 18578 21770
rect 18466 21743 18551 21769
rect 18577 21743 18578 21769
rect 18466 21742 18578 21743
rect 18438 21737 18466 21742
rect 17990 20953 18018 20958
rect 18550 20985 18578 21742
rect 19278 21769 19306 21799
rect 19278 21743 19279 21769
rect 19305 21743 19306 21769
rect 18550 20959 18551 20985
rect 18577 20959 18578 20985
rect 18550 20930 18578 20959
rect 18550 20897 18578 20902
rect 19054 21377 19082 21383
rect 19054 21351 19055 21377
rect 19081 21351 19082 21377
rect 19054 20930 19082 21351
rect 19054 20594 19082 20902
rect 19054 20547 19082 20566
rect 19278 21378 19306 21743
rect 19446 21378 19474 21383
rect 19278 21377 19474 21378
rect 19278 21351 19279 21377
rect 19305 21351 19447 21377
rect 19473 21351 19474 21377
rect 19278 21350 19474 21351
rect 17990 20258 18018 20263
rect 17934 20257 18018 20258
rect 17934 20231 17991 20257
rect 18017 20231 18018 20257
rect 17934 20230 18018 20231
rect 17990 20201 18018 20230
rect 19278 20257 19306 21350
rect 19446 21345 19474 21350
rect 19446 21041 19474 21047
rect 19446 21015 19447 21041
rect 19473 21015 19474 21041
rect 19446 20986 19474 21015
rect 19446 20538 19474 20958
rect 19446 20505 19474 20510
rect 19950 20593 19978 20599
rect 19950 20567 19951 20593
rect 19977 20567 19978 20593
rect 19950 20538 19978 20567
rect 19950 20491 19978 20510
rect 19278 20231 19279 20257
rect 19305 20231 19306 20257
rect 17990 20175 17991 20201
rect 18017 20175 18018 20201
rect 17598 20006 17730 20011
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17598 19973 17730 19978
rect 17430 19783 17431 19809
rect 17457 19783 17458 19809
rect 17430 19753 17458 19783
rect 17430 19727 17431 19753
rect 17457 19727 17458 19753
rect 17430 19025 17458 19727
rect 17990 19473 18018 20175
rect 17990 19447 17991 19473
rect 18017 19447 18018 19473
rect 17990 19417 18018 19447
rect 17990 19391 17991 19417
rect 18017 19391 18018 19417
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 17430 18999 17431 19025
rect 17457 18999 17458 19025
rect 17430 18969 17458 18999
rect 17430 18943 17431 18969
rect 17457 18943 17458 18969
rect 17430 18242 17458 18943
rect 17990 18689 18018 19391
rect 17990 18663 17991 18689
rect 18017 18663 18018 18689
rect 17990 18633 18018 18663
rect 17990 18607 17991 18633
rect 18017 18607 18018 18633
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17430 18185 17458 18214
rect 17430 18159 17431 18185
rect 17457 18159 17458 18185
rect 17430 18153 17458 18159
rect 17990 18242 18018 18607
rect 17990 17905 18018 18214
rect 17990 17879 17991 17905
rect 18017 17879 18018 17905
rect 17990 17850 18018 17879
rect 17990 17803 18018 17822
rect 18550 20201 18578 20207
rect 18550 20175 18551 20201
rect 18577 20175 18578 20201
rect 18550 19417 18578 20175
rect 19278 20201 19306 20231
rect 19278 20175 19279 20201
rect 19305 20175 19306 20201
rect 18550 19391 18551 19417
rect 18577 19391 18578 19417
rect 18550 18633 18578 19391
rect 18550 18607 18551 18633
rect 18577 18607 18578 18633
rect 18550 18522 18578 18607
rect 19054 19809 19082 19815
rect 19054 19783 19055 19809
rect 19081 19783 19082 19809
rect 19054 19025 19082 19783
rect 19278 19810 19306 20175
rect 19334 19810 19362 19815
rect 19446 19810 19474 19815
rect 19278 19809 19474 19810
rect 19278 19783 19335 19809
rect 19361 19783 19447 19809
rect 19473 19783 19474 19809
rect 19278 19782 19474 19783
rect 19054 18999 19055 19025
rect 19081 18999 19082 19025
rect 19054 18522 19082 18999
rect 18550 18494 19082 18522
rect 18550 17849 18578 18494
rect 18550 17823 18551 17849
rect 18577 17823 18578 17849
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17990 17121 18018 17127
rect 17990 17095 17991 17121
rect 18017 17095 18018 17121
rect 17990 17065 18018 17095
rect 17990 17039 17991 17065
rect 18017 17039 18018 17065
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17318 16617 17346 16623
rect 17318 16591 17319 16617
rect 17345 16591 17346 16617
rect 17318 16282 17346 16591
rect 17486 16282 17514 16287
rect 17318 16281 17514 16282
rect 17318 16255 17319 16281
rect 17345 16255 17487 16281
rect 17513 16255 17514 16281
rect 17318 16254 17514 16255
rect 17318 15974 17346 16254
rect 17486 16249 17514 16254
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17206 15946 17346 15974
rect 17206 15834 17234 15946
rect 17206 15801 17234 15806
rect 17430 15889 17458 15895
rect 17430 15863 17431 15889
rect 17457 15863 17458 15889
rect 17430 15834 17458 15863
rect 17430 15105 17458 15806
rect 17990 15834 18018 17039
rect 18550 17065 18578 17823
rect 18550 17039 18551 17065
rect 18577 17039 18578 17065
rect 18550 16282 18578 17039
rect 19054 18242 19082 18494
rect 19054 17457 19082 18214
rect 19054 17431 19055 17457
rect 19081 17431 19082 17457
rect 19054 16673 19082 17431
rect 19054 16647 19055 16673
rect 19081 16647 19082 16673
rect 19054 16641 19082 16647
rect 19334 19473 19362 19782
rect 19446 19777 19474 19782
rect 19334 19447 19335 19473
rect 19361 19447 19362 19473
rect 19334 19417 19362 19447
rect 19334 19391 19335 19417
rect 19361 19391 19362 19417
rect 19334 19026 19362 19391
rect 19446 19026 19474 19031
rect 19334 19025 19474 19026
rect 19334 18999 19335 19025
rect 19361 18999 19447 19025
rect 19473 18999 19474 19025
rect 19334 18998 19474 18999
rect 19334 18689 19362 18998
rect 19446 18993 19474 18998
rect 19334 18663 19335 18689
rect 19361 18663 19362 18689
rect 19334 18633 19362 18663
rect 19334 18607 19335 18633
rect 19361 18607 19362 18633
rect 19334 18242 19362 18607
rect 19446 18242 19474 18247
rect 19334 18241 19474 18242
rect 19334 18215 19335 18241
rect 19361 18215 19447 18241
rect 19473 18215 19474 18241
rect 19334 18214 19474 18215
rect 19334 17905 19362 18214
rect 19446 18209 19474 18214
rect 19334 17879 19335 17905
rect 19361 17879 19362 17905
rect 19334 17850 19362 17879
rect 19334 17458 19362 17822
rect 19446 17458 19474 17463
rect 19334 17457 19474 17458
rect 19334 17431 19335 17457
rect 19361 17431 19447 17457
rect 19473 17431 19474 17457
rect 19334 17430 19474 17431
rect 19334 17121 19362 17430
rect 19446 17425 19474 17430
rect 19334 17095 19335 17121
rect 19361 17095 19362 17121
rect 19334 17065 19362 17095
rect 19334 17039 19335 17065
rect 19361 17039 19362 17065
rect 19334 16674 19362 17039
rect 19446 16674 19474 16679
rect 19334 16673 19474 16674
rect 19334 16647 19335 16673
rect 19361 16647 19447 16673
rect 19473 16647 19474 16673
rect 19334 16646 19474 16647
rect 19222 16337 19250 16343
rect 19222 16311 19223 16337
rect 19249 16311 19250 16337
rect 17990 15553 18018 15806
rect 17990 15527 17991 15553
rect 18017 15527 18018 15553
rect 17990 15498 18018 15527
rect 17990 15451 18018 15470
rect 18270 16281 18802 16282
rect 18270 16255 18551 16281
rect 18577 16255 18802 16281
rect 18270 16254 18802 16255
rect 18270 15497 18298 16254
rect 18550 16249 18578 16254
rect 18774 15890 18802 16254
rect 19222 16281 19250 16311
rect 19222 16255 19223 16281
rect 19249 16255 19250 16281
rect 19222 15974 19250 16255
rect 19222 15946 19306 15974
rect 19054 15890 19082 15895
rect 18774 15889 19082 15890
rect 18774 15863 19055 15889
rect 19081 15863 19082 15889
rect 18774 15862 19082 15863
rect 18270 15471 18271 15497
rect 18297 15471 18298 15497
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17430 15079 17431 15105
rect 17457 15079 17458 15105
rect 17430 15050 17458 15079
rect 17430 15049 17514 15050
rect 17430 15023 17431 15049
rect 17457 15023 17514 15049
rect 17430 15022 17514 15023
rect 17430 15017 17458 15022
rect 17374 14714 17402 14719
rect 17486 14714 17514 15022
rect 17374 14713 17514 14714
rect 17374 14687 17375 14713
rect 17401 14687 17487 14713
rect 17513 14687 17514 14713
rect 17374 14686 17514 14687
rect 17374 14681 17402 14686
rect 17430 14321 17458 14686
rect 17486 14681 17514 14686
rect 18270 14713 18298 15471
rect 18270 14687 18271 14713
rect 18297 14687 18298 14713
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17430 14295 17431 14321
rect 17457 14295 17458 14321
rect 17430 14266 17458 14295
rect 17430 14265 17514 14266
rect 17430 14239 17431 14265
rect 17457 14239 17514 14265
rect 17430 14238 17514 14239
rect 17430 14233 17458 14238
rect 17374 13930 17402 13935
rect 17486 13930 17514 14238
rect 17374 13929 17514 13930
rect 17374 13903 17375 13929
rect 17401 13903 17487 13929
rect 17513 13903 17514 13929
rect 17374 13902 17514 13903
rect 17374 13897 17402 13902
rect 17430 13538 17458 13902
rect 17486 13897 17514 13902
rect 18270 13929 18298 14687
rect 18270 13903 18271 13929
rect 18297 13903 18298 13929
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 17430 13482 17458 13510
rect 18270 13482 18298 13903
rect 19054 15105 19082 15862
rect 19278 15834 19306 15946
rect 19278 15553 19306 15806
rect 19278 15527 19279 15553
rect 19305 15527 19306 15553
rect 19278 15498 19306 15527
rect 19278 15432 19306 15470
rect 19054 15079 19055 15105
rect 19081 15079 19082 15105
rect 19054 14322 19082 15079
rect 19334 15106 19362 16646
rect 19446 16641 19474 16646
rect 19950 15889 19978 15895
rect 19950 15863 19951 15889
rect 19977 15863 19978 15889
rect 19950 15834 19978 15863
rect 19950 15787 19978 15806
rect 19446 15106 19474 15111
rect 19334 15105 19474 15106
rect 19334 15079 19335 15105
rect 19361 15079 19447 15105
rect 19473 15079 19474 15105
rect 19334 15078 19474 15079
rect 19334 15073 19362 15078
rect 19446 14769 19474 15078
rect 19446 14743 19447 14769
rect 19473 14743 19474 14769
rect 19446 14713 19474 14743
rect 19446 14687 19447 14713
rect 19473 14687 19474 14713
rect 19446 14434 19474 14687
rect 19054 13537 19082 14294
rect 19334 14322 19362 14327
rect 19446 14322 19474 14406
rect 20174 14378 20202 34600
rect 22638 33642 22666 33647
rect 22470 30954 22498 30959
rect 22414 29386 22442 29391
rect 21910 28882 21938 28887
rect 21686 28378 21714 28383
rect 20958 28042 20986 28047
rect 20958 27594 20986 28014
rect 21406 28042 21434 28047
rect 21406 27995 21434 28014
rect 21518 28042 21546 28047
rect 21686 28042 21714 28350
rect 21518 28041 21714 28042
rect 21518 28015 21519 28041
rect 21545 28015 21687 28041
rect 21713 28015 21714 28041
rect 21518 28014 21714 28015
rect 21518 28009 21546 28014
rect 21350 27762 21378 27767
rect 20902 27593 20986 27594
rect 20902 27567 20959 27593
rect 20985 27567 20986 27593
rect 20902 27566 20986 27567
rect 20678 26922 20706 26927
rect 20342 26866 20370 26871
rect 20342 26819 20370 26838
rect 20510 26866 20538 26871
rect 20510 26819 20538 26838
rect 20678 26865 20706 26894
rect 20678 26839 20679 26865
rect 20705 26839 20706 26865
rect 20678 26833 20706 26839
rect 20902 26026 20930 27566
rect 20958 27561 20986 27566
rect 21126 27649 21154 27655
rect 21126 27623 21127 27649
rect 21153 27623 21154 27649
rect 21126 27594 21154 27623
rect 21238 27594 21266 27599
rect 21126 27593 21266 27594
rect 21126 27567 21239 27593
rect 21265 27567 21266 27593
rect 21126 27566 21266 27567
rect 21070 27314 21098 27319
rect 20958 27286 21070 27314
rect 20958 26922 20986 27286
rect 21070 27267 21098 27286
rect 21126 27258 21154 27566
rect 21238 27561 21266 27566
rect 21182 27258 21210 27263
rect 21350 27258 21378 27734
rect 21630 27762 21658 28014
rect 21686 28009 21714 28014
rect 21910 28042 21938 28854
rect 22414 28882 22442 29358
rect 22414 28816 22442 28854
rect 22134 28602 22162 28607
rect 22134 28434 22162 28574
rect 21910 28009 21938 28014
rect 21966 28433 22162 28434
rect 21966 28407 22135 28433
rect 22161 28407 22162 28433
rect 21966 28406 22162 28407
rect 21966 28041 21994 28406
rect 22134 28401 22162 28406
rect 22470 28434 22498 30926
rect 22638 29218 22666 33614
rect 22694 33614 22722 34622
rect 23086 34538 23114 34622
rect 23240 34600 23296 35000
rect 23254 34538 23282 34600
rect 23086 34510 23282 34538
rect 22694 33586 22834 33614
rect 22190 28378 22218 28383
rect 22190 28331 22218 28350
rect 22358 28378 22386 28383
rect 22358 28331 22386 28350
rect 22470 28210 22498 28406
rect 22302 28182 22498 28210
rect 22526 29190 22638 29218
rect 22526 28602 22554 29190
rect 22638 29185 22666 29190
rect 22694 29610 22722 29615
rect 22694 28881 22722 29582
rect 22694 28855 22695 28881
rect 22721 28855 22722 28881
rect 22582 28826 22610 28831
rect 22694 28826 22722 28855
rect 22582 28825 22722 28826
rect 22582 28799 22583 28825
rect 22609 28799 22722 28825
rect 22582 28798 22722 28799
rect 22582 28793 22610 28798
rect 21966 28015 21967 28041
rect 21993 28015 21994 28041
rect 21126 27257 21378 27258
rect 21126 27231 21183 27257
rect 21209 27231 21351 27257
rect 21377 27231 21378 27257
rect 21574 27650 21602 27655
rect 21574 27314 21602 27622
rect 21630 27650 21658 27734
rect 21966 27734 21994 28015
rect 22078 28042 22106 28047
rect 22246 28042 22274 28047
rect 22078 28041 22246 28042
rect 22078 28015 22079 28041
rect 22105 28015 22246 28041
rect 22078 28014 22246 28015
rect 22078 28009 22106 28014
rect 21966 27706 22050 27734
rect 21798 27650 21826 27655
rect 21630 27649 21826 27650
rect 21630 27623 21631 27649
rect 21657 27623 21799 27649
rect 21825 27623 21826 27649
rect 21630 27622 21826 27623
rect 21630 27617 21658 27622
rect 21798 27617 21826 27622
rect 22022 27650 22050 27706
rect 22022 27594 22050 27622
rect 22078 27594 22106 27599
rect 22022 27593 22106 27594
rect 22022 27567 22079 27593
rect 22105 27567 22106 27593
rect 22022 27566 22106 27567
rect 21630 27314 21658 27319
rect 21602 27313 21658 27314
rect 21602 27287 21631 27313
rect 21657 27287 21658 27313
rect 21602 27286 21658 27287
rect 21574 27248 21602 27286
rect 21630 27281 21658 27286
rect 21742 27258 21770 27263
rect 21798 27258 21826 27263
rect 21966 27258 21994 27263
rect 21742 27257 21798 27258
rect 21126 27230 21378 27231
rect 21126 27202 21154 27230
rect 21182 27225 21210 27230
rect 21350 27225 21378 27230
rect 21742 27231 21743 27257
rect 21769 27231 21798 27257
rect 21742 27230 21798 27231
rect 21826 27230 21882 27258
rect 20958 26865 20986 26894
rect 20958 26839 20959 26865
rect 20985 26839 20986 26865
rect 20958 26833 20986 26839
rect 21070 27174 21154 27202
rect 21070 26866 21098 27174
rect 21742 27090 21770 27230
rect 21798 27192 21826 27230
rect 21462 27062 21770 27090
rect 21014 26530 21042 26535
rect 21070 26530 21098 26838
rect 21126 26866 21154 26871
rect 21238 26866 21266 26871
rect 21462 26866 21490 27062
rect 21126 26865 21490 26866
rect 21126 26839 21127 26865
rect 21153 26839 21239 26865
rect 21265 26839 21490 26865
rect 21126 26838 21490 26839
rect 21630 26866 21658 26871
rect 21126 26833 21154 26838
rect 21238 26833 21266 26838
rect 21630 26819 21658 26838
rect 21798 26866 21826 26871
rect 21798 26819 21826 26838
rect 21014 26529 21098 26530
rect 21014 26503 21015 26529
rect 21041 26503 21098 26529
rect 21014 26502 21098 26503
rect 21014 26497 21042 26502
rect 21070 26474 21098 26502
rect 21518 26809 21546 26815
rect 21518 26783 21519 26809
rect 21545 26783 21546 26809
rect 21126 26474 21154 26479
rect 21070 26473 21154 26474
rect 21070 26447 21127 26473
rect 21153 26447 21154 26473
rect 21070 26446 21154 26447
rect 21070 26082 21098 26446
rect 21126 26441 21154 26446
rect 21294 26474 21322 26479
rect 21294 26427 21322 26446
rect 21518 26474 21546 26783
rect 21854 26530 21882 27230
rect 21966 27211 21994 27230
rect 21742 26529 21882 26530
rect 21742 26503 21855 26529
rect 21881 26503 21882 26529
rect 21742 26502 21882 26503
rect 21238 26082 21266 26087
rect 21070 26081 21238 26082
rect 21070 26055 21071 26081
rect 21097 26055 21238 26081
rect 21070 26054 21238 26055
rect 21070 26049 21098 26054
rect 20958 26026 20986 26031
rect 20902 25998 20958 26026
rect 21238 26016 21266 26054
rect 21518 26081 21546 26446
rect 21630 26474 21658 26479
rect 21630 26427 21658 26446
rect 21742 26473 21770 26502
rect 21742 26447 21743 26473
rect 21769 26447 21770 26473
rect 21742 26441 21770 26447
rect 21518 26055 21519 26081
rect 21545 26055 21546 26081
rect 21518 26049 21546 26055
rect 21630 26082 21658 26087
rect 21630 26035 21658 26054
rect 21798 26082 21826 26087
rect 21798 26035 21826 26054
rect 21574 26026 21602 26031
rect 20958 25979 20986 25998
rect 21574 25745 21602 25998
rect 21854 25746 21882 26502
rect 21574 25719 21575 25745
rect 21601 25719 21602 25745
rect 21574 25713 21602 25719
rect 21742 25745 21882 25746
rect 21742 25719 21855 25745
rect 21881 25719 21882 25745
rect 21742 25718 21882 25719
rect 21742 25689 21770 25718
rect 21742 25663 21743 25689
rect 21769 25663 21770 25689
rect 21854 25680 21882 25718
rect 21742 25657 21770 25663
rect 22022 25298 22050 27566
rect 22078 27561 22106 27566
rect 22190 27594 22218 28014
rect 22246 27995 22274 28014
rect 22302 27734 22330 28182
rect 22526 28041 22554 28574
rect 22526 28015 22527 28041
rect 22553 28015 22554 28041
rect 22526 28009 22554 28015
rect 22638 28098 22666 28798
rect 22750 28098 22778 28103
rect 22638 28097 22778 28098
rect 22638 28071 22751 28097
rect 22777 28071 22778 28097
rect 22638 28070 22778 28071
rect 22638 28042 22666 28070
rect 22750 28065 22778 28070
rect 22638 27976 22666 28014
rect 22190 27547 22218 27566
rect 22246 27706 22330 27734
rect 22190 27258 22218 27263
rect 22246 27258 22274 27706
rect 22414 27649 22442 27655
rect 22414 27623 22415 27649
rect 22441 27623 22442 27649
rect 22414 27594 22442 27623
rect 22134 27257 22274 27258
rect 22134 27231 22191 27257
rect 22217 27231 22274 27257
rect 22134 27230 22274 27231
rect 22358 27258 22386 27263
rect 22414 27258 22442 27566
rect 22750 27594 22778 27599
rect 22526 27258 22554 27263
rect 22358 27257 22526 27258
rect 22358 27231 22359 27257
rect 22385 27231 22526 27257
rect 22358 27230 22526 27231
rect 22134 26865 22162 27230
rect 22190 27225 22218 27230
rect 22358 27225 22386 27230
rect 22134 26839 22135 26865
rect 22161 26839 22162 26865
rect 22134 26474 22162 26839
rect 22246 26866 22274 26871
rect 22414 26866 22442 26871
rect 22470 26866 22498 27230
rect 22526 27211 22554 27230
rect 22750 27257 22778 27566
rect 22750 27231 22751 27257
rect 22777 27231 22778 27257
rect 22246 26865 22498 26866
rect 22246 26839 22247 26865
rect 22273 26839 22415 26865
rect 22441 26839 22498 26865
rect 22246 26838 22498 26839
rect 22246 26833 22274 26838
rect 22414 26833 22442 26838
rect 22134 26082 22162 26446
rect 22302 26474 22330 26479
rect 22470 26474 22498 26838
rect 22302 26473 22498 26474
rect 22302 26447 22303 26473
rect 22329 26447 22471 26473
rect 22497 26447 22498 26473
rect 22302 26446 22498 26447
rect 22302 26441 22330 26446
rect 22134 25745 22162 26054
rect 22246 26082 22274 26087
rect 22414 26082 22442 26087
rect 22470 26082 22498 26446
rect 22246 26081 22498 26082
rect 22246 26055 22247 26081
rect 22273 26055 22415 26081
rect 22441 26055 22498 26081
rect 22246 26054 22498 26055
rect 22694 26866 22722 26871
rect 22694 26530 22722 26838
rect 22750 26865 22778 27231
rect 22750 26839 22751 26865
rect 22777 26839 22778 26865
rect 22750 26833 22778 26839
rect 22246 26049 22274 26054
rect 22414 26049 22442 26054
rect 22134 25719 22135 25745
rect 22161 25719 22162 25745
rect 22134 25713 22162 25719
rect 22694 25745 22722 26502
rect 22694 25719 22695 25745
rect 22721 25719 22722 25745
rect 22302 25690 22330 25695
rect 22470 25690 22498 25695
rect 22694 25690 22722 25719
rect 22302 25689 22722 25690
rect 22302 25663 22303 25689
rect 22329 25663 22471 25689
rect 22497 25663 22722 25689
rect 22302 25662 22722 25663
rect 22302 25657 22330 25662
rect 22134 25298 22162 25303
rect 22022 25297 22162 25298
rect 22022 25271 22135 25297
rect 22161 25271 22162 25297
rect 22022 25270 22162 25271
rect 22134 24962 22162 25270
rect 22246 25298 22274 25303
rect 22358 25298 22386 25662
rect 22470 25657 22498 25662
rect 22246 25297 22386 25298
rect 22246 25271 22247 25297
rect 22273 25271 22359 25297
rect 22385 25271 22386 25297
rect 22246 25270 22386 25271
rect 22246 25265 22274 25270
rect 22358 25265 22386 25270
rect 22470 24962 22498 24967
rect 22134 24961 22498 24962
rect 22134 24935 22471 24961
rect 22497 24935 22498 24961
rect 22134 24934 22498 24935
rect 22470 24929 22498 24934
rect 22582 24962 22610 25662
rect 22750 24962 22778 24967
rect 22582 24961 22750 24962
rect 22582 24935 22583 24961
rect 22609 24935 22750 24961
rect 22582 24934 22750 24935
rect 22582 24929 22610 24934
rect 22750 24896 22778 24934
rect 22806 21854 22834 33586
rect 23086 29610 23114 29615
rect 23030 29218 23058 29223
rect 23030 28882 23058 29190
rect 23030 28825 23058 28854
rect 23086 28882 23114 29582
rect 23310 29609 23338 29615
rect 23310 29583 23311 29609
rect 23337 29583 23338 29609
rect 23310 29386 23338 29583
rect 23366 29610 23394 29615
rect 23366 29563 23394 29582
rect 23590 29610 23618 29615
rect 23590 29609 23730 29610
rect 23590 29583 23591 29609
rect 23617 29583 23730 29609
rect 23590 29582 23730 29583
rect 23590 29577 23618 29582
rect 23310 29353 23338 29358
rect 23590 29386 23618 29391
rect 23198 29218 23226 29223
rect 23198 29217 23338 29218
rect 23198 29191 23199 29217
rect 23225 29191 23338 29217
rect 23198 29190 23338 29191
rect 23198 29185 23226 29190
rect 23310 29161 23338 29190
rect 23310 29135 23311 29161
rect 23337 29135 23338 29161
rect 23254 28882 23282 28887
rect 23086 28881 23282 28882
rect 23086 28855 23087 28881
rect 23113 28855 23255 28881
rect 23281 28855 23282 28881
rect 23086 28854 23282 28855
rect 23086 28849 23114 28854
rect 23254 28849 23282 28854
rect 23030 28799 23031 28825
rect 23057 28799 23058 28825
rect 23030 28793 23058 28799
rect 23310 28826 23338 29135
rect 23590 29161 23618 29358
rect 23702 29218 23730 29582
rect 23870 29218 23898 29223
rect 23702 29217 23898 29218
rect 23702 29191 23703 29217
rect 23729 29191 23871 29217
rect 23897 29191 23898 29217
rect 23702 29190 23898 29191
rect 23702 29185 23730 29190
rect 23590 29135 23591 29161
rect 23617 29135 23618 29161
rect 23030 28434 23058 28439
rect 23030 28098 23058 28406
rect 22974 28097 23058 28098
rect 22974 28071 23031 28097
rect 23057 28071 23058 28097
rect 22974 28070 23058 28071
rect 22974 27594 23002 28070
rect 23030 28065 23058 28070
rect 23142 28378 23170 28383
rect 23310 28378 23338 28798
rect 23534 28882 23562 28887
rect 23534 28434 23562 28854
rect 23590 28602 23618 29135
rect 23646 28826 23674 28831
rect 23646 28779 23674 28798
rect 23590 28569 23618 28574
rect 23590 28434 23618 28439
rect 23534 28433 23618 28434
rect 23534 28407 23591 28433
rect 23617 28407 23618 28433
rect 23534 28406 23618 28407
rect 23170 28377 23338 28378
rect 23170 28351 23311 28377
rect 23337 28351 23338 28377
rect 23170 28350 23338 28351
rect 23142 28097 23170 28350
rect 23142 28071 23143 28097
rect 23169 28071 23170 28097
rect 23142 28065 23170 28071
rect 23310 28097 23338 28350
rect 23310 28071 23311 28097
rect 23337 28071 23338 28097
rect 23310 27734 23338 28071
rect 23590 28097 23618 28406
rect 23590 28071 23591 28097
rect 23617 28071 23618 28097
rect 23590 28065 23618 28071
rect 23758 28434 23786 29190
rect 23870 29185 23898 29190
rect 23814 28826 23842 28831
rect 23814 28779 23842 28798
rect 23870 28434 23898 28439
rect 23758 28433 23898 28434
rect 23758 28407 23759 28433
rect 23785 28407 23871 28433
rect 23897 28407 23898 28433
rect 23758 28406 23898 28407
rect 23758 28098 23786 28406
rect 23870 28401 23898 28406
rect 23870 28098 23898 28103
rect 23758 28097 23898 28098
rect 23758 28071 23871 28097
rect 23897 28071 23898 28097
rect 23758 28070 23898 28071
rect 23758 28041 23786 28070
rect 23870 28065 23898 28070
rect 23758 28015 23759 28041
rect 23785 28015 23786 28041
rect 23758 27734 23786 28015
rect 23254 27706 23282 27711
rect 23310 27706 23674 27734
rect 22974 27547 23002 27566
rect 23086 27594 23114 27599
rect 23254 27594 23282 27678
rect 23086 27593 23282 27594
rect 23086 27567 23087 27593
rect 23113 27567 23255 27593
rect 23281 27567 23282 27593
rect 23086 27566 23282 27567
rect 22918 27258 22946 27263
rect 23030 27258 23058 27263
rect 23086 27258 23114 27566
rect 23254 27561 23282 27566
rect 23534 27594 23562 27599
rect 23534 27547 23562 27566
rect 23646 27594 23674 27706
rect 23702 27706 23786 27734
rect 23702 27673 23730 27678
rect 23814 27594 23842 27599
rect 23646 27593 23842 27594
rect 23646 27567 23647 27593
rect 23673 27567 23815 27593
rect 23841 27567 23842 27593
rect 23646 27566 23842 27567
rect 22946 27257 23114 27258
rect 22946 27231 23031 27257
rect 23057 27231 23114 27257
rect 22946 27230 23114 27231
rect 23310 27257 23338 27263
rect 23310 27231 23311 27257
rect 23337 27231 23338 27257
rect 22918 26922 22946 27230
rect 23030 27225 23058 27230
rect 22918 26865 22946 26894
rect 22918 26839 22919 26865
rect 22945 26839 22946 26865
rect 22918 26833 22946 26839
rect 23086 26922 23114 26927
rect 23086 26865 23114 26894
rect 23086 26839 23087 26865
rect 23113 26839 23114 26865
rect 23086 26833 23114 26839
rect 23310 26809 23338 27231
rect 23422 27257 23450 27263
rect 23422 27231 23423 27257
rect 23449 27231 23450 27257
rect 23422 26866 23450 27231
rect 23646 27257 23674 27566
rect 23814 27561 23842 27566
rect 23646 27231 23647 27257
rect 23673 27231 23674 27257
rect 23422 26819 23450 26838
rect 23478 26922 23506 26927
rect 23310 26783 23311 26809
rect 23337 26783 23338 26809
rect 22862 26530 22890 26535
rect 22862 25745 22890 26502
rect 22862 25719 22863 25745
rect 22889 25719 22890 25745
rect 22862 25713 22890 25719
rect 22974 26473 23002 26479
rect 22974 26447 22975 26473
rect 23001 26447 23002 26473
rect 22974 25689 23002 26447
rect 23310 26473 23338 26783
rect 23310 26447 23311 26473
rect 23337 26447 23338 26473
rect 22974 25663 22975 25689
rect 23001 25663 23002 25689
rect 22974 25578 23002 25663
rect 22974 25545 23002 25550
rect 23030 26082 23058 26087
rect 23030 24961 23058 26054
rect 23310 26081 23338 26447
rect 23310 26055 23311 26081
rect 23337 26055 23338 26081
rect 23310 25689 23338 26055
rect 23310 25663 23311 25689
rect 23337 25663 23338 25689
rect 23310 25578 23338 25663
rect 23310 25297 23338 25550
rect 23310 25271 23311 25297
rect 23337 25271 23338 25297
rect 23310 25265 23338 25271
rect 23422 26474 23450 26479
rect 23478 26474 23506 26894
rect 23646 26866 23674 27231
rect 23646 26865 23786 26866
rect 23646 26839 23647 26865
rect 23673 26839 23786 26865
rect 23646 26838 23786 26839
rect 23646 26833 23674 26838
rect 23534 26474 23562 26479
rect 23422 26473 23562 26474
rect 23422 26447 23423 26473
rect 23449 26447 23535 26473
rect 23561 26447 23562 26473
rect 23422 26446 23562 26447
rect 23422 26081 23450 26446
rect 23534 26441 23562 26446
rect 23422 26055 23423 26081
rect 23449 26055 23450 26081
rect 23422 25690 23450 26055
rect 23534 26025 23562 26031
rect 23534 25999 23535 26025
rect 23561 25999 23562 26025
rect 23534 25690 23562 25999
rect 23422 25689 23562 25690
rect 23422 25663 23423 25689
rect 23449 25663 23535 25689
rect 23561 25663 23562 25689
rect 23422 25662 23562 25663
rect 23422 25298 23450 25662
rect 23534 25657 23562 25662
rect 23590 25298 23618 25303
rect 23422 25297 23618 25298
rect 23422 25271 23423 25297
rect 23449 25271 23591 25297
rect 23617 25271 23618 25297
rect 23422 25270 23618 25271
rect 23422 25265 23450 25270
rect 23030 24935 23031 24961
rect 23057 24935 23058 24961
rect 23030 24929 23058 24935
rect 23142 24962 23170 24967
rect 23310 24962 23338 24967
rect 23170 24961 23338 24962
rect 23170 24935 23311 24961
rect 23337 24935 23338 24961
rect 23170 24934 23338 24935
rect 23142 24513 23170 24934
rect 23142 24487 23143 24513
rect 23169 24487 23170 24513
rect 23142 24481 23170 24487
rect 23310 24513 23338 24934
rect 23590 24794 23618 25270
rect 23758 24906 23786 26838
rect 23926 24906 23954 24911
rect 23758 24905 24010 24906
rect 23758 24879 23759 24905
rect 23785 24879 23927 24905
rect 23953 24879 24010 24905
rect 23758 24878 24010 24879
rect 23758 24873 23786 24878
rect 23926 24873 23954 24878
rect 23590 24766 23786 24794
rect 23310 24487 23311 24513
rect 23337 24487 23338 24513
rect 23310 24481 23338 24487
rect 23758 24514 23786 24766
rect 23870 24514 23898 24519
rect 23758 24513 23898 24514
rect 23758 24487 23759 24513
rect 23785 24487 23871 24513
rect 23897 24487 23898 24513
rect 23758 24486 23898 24487
rect 23758 24481 23786 24486
rect 23478 24458 23506 24463
rect 23478 24411 23506 24430
rect 23870 24234 23898 24486
rect 23758 24206 23954 24234
rect 23758 24121 23786 24206
rect 23926 24177 23954 24206
rect 23926 24151 23927 24177
rect 23953 24151 23954 24177
rect 23926 24145 23954 24151
rect 23758 24095 23759 24121
rect 23785 24095 23786 24121
rect 23758 24066 23786 24095
rect 23758 24038 23842 24066
rect 23702 23338 23730 23343
rect 23198 22890 23226 22895
rect 23198 22843 23226 22862
rect 23366 22890 23394 22895
rect 23366 22843 23394 22862
rect 23478 22890 23506 22895
rect 23702 22890 23730 23310
rect 23814 22946 23842 24038
rect 23982 24010 24010 24878
rect 23870 23982 24010 24010
rect 24038 24905 24066 24911
rect 24038 24879 24039 24905
rect 24065 24879 24066 24905
rect 24038 24458 24066 24879
rect 24038 24121 24066 24430
rect 24038 24095 24039 24121
rect 24065 24095 24066 24121
rect 23870 23338 23898 23982
rect 23870 23291 23898 23310
rect 23982 23337 24010 23343
rect 23982 23311 23983 23337
rect 24009 23311 24010 23337
rect 23870 22946 23898 22951
rect 23814 22945 23898 22946
rect 23814 22919 23871 22945
rect 23897 22919 23898 22945
rect 23814 22918 23898 22919
rect 23478 22889 23562 22890
rect 23478 22863 23479 22889
rect 23505 22863 23562 22889
rect 23478 22862 23562 22863
rect 23478 22857 23506 22862
rect 23534 22722 23562 22862
rect 22806 21826 22890 21854
rect 20510 20594 20538 20599
rect 20510 19810 20538 20566
rect 21238 20593 21266 20599
rect 21238 20567 21239 20593
rect 21265 20567 21266 20593
rect 21182 20538 21210 20543
rect 20510 19763 20538 19782
rect 20958 20201 20986 20207
rect 20958 20175 20959 20201
rect 20985 20175 20986 20201
rect 20958 19810 20986 20175
rect 20958 19418 20986 19782
rect 21182 19809 21210 20510
rect 21182 19783 21183 19809
rect 21209 19783 21210 19809
rect 21182 19753 21210 19783
rect 21182 19727 21183 19753
rect 21209 19727 21210 19753
rect 21182 19721 21210 19727
rect 21238 20537 21266 20567
rect 21238 20511 21239 20537
rect 21265 20511 21266 20537
rect 21238 20202 21266 20511
rect 21462 20202 21490 20207
rect 21238 20201 21490 20202
rect 21238 20175 21239 20201
rect 21265 20175 21463 20201
rect 21489 20175 21490 20201
rect 21238 20174 21490 20175
rect 20958 19371 20986 19390
rect 20230 19025 20258 19031
rect 20230 18999 20231 19025
rect 20257 18999 20258 19025
rect 20230 18242 20258 18999
rect 21238 19025 21266 20174
rect 21462 20169 21490 20174
rect 21798 19473 21826 19479
rect 21798 19447 21799 19473
rect 21825 19447 21826 19473
rect 21798 19417 21826 19447
rect 21798 19391 21799 19417
rect 21825 19391 21826 19417
rect 21798 19362 21826 19391
rect 21798 19329 21826 19334
rect 22526 19418 22554 19423
rect 21238 18999 21239 19025
rect 21265 18999 21266 19025
rect 21238 18969 21266 18999
rect 21238 18943 21239 18969
rect 21265 18943 21266 18969
rect 20230 18176 20258 18214
rect 20958 18633 20986 18639
rect 20958 18607 20959 18633
rect 20985 18607 20986 18633
rect 20958 17849 20986 18607
rect 20958 17823 20959 17849
rect 20985 17823 20986 17849
rect 20174 14345 20202 14350
rect 20230 17457 20258 17463
rect 20230 17431 20231 17457
rect 20257 17431 20258 17457
rect 20230 16673 20258 17431
rect 20230 16647 20231 16673
rect 20257 16647 20258 16673
rect 20230 15889 20258 16647
rect 20958 17065 20986 17823
rect 20958 17039 20959 17065
rect 20985 17039 20986 17065
rect 20230 15863 20231 15889
rect 20257 15863 20258 15889
rect 20230 15105 20258 15863
rect 20230 15079 20231 15105
rect 20257 15079 20258 15105
rect 20230 14714 20258 15079
rect 20790 16282 20818 16287
rect 20790 15497 20818 16254
rect 20958 16282 20986 17039
rect 20958 16235 20986 16254
rect 21238 18634 21266 18943
rect 21462 18634 21490 18639
rect 21238 18633 21490 18634
rect 21238 18607 21239 18633
rect 21265 18607 21463 18633
rect 21489 18607 21490 18633
rect 21238 18606 21490 18607
rect 21238 18241 21266 18606
rect 21462 18601 21490 18606
rect 22526 18633 22554 19390
rect 22526 18607 22527 18633
rect 22553 18607 22554 18633
rect 21238 18215 21239 18241
rect 21265 18215 21266 18241
rect 21238 18185 21266 18215
rect 21238 18159 21239 18185
rect 21265 18159 21266 18185
rect 21238 17850 21266 18159
rect 21462 17850 21490 17855
rect 21238 17849 21490 17850
rect 21238 17823 21239 17849
rect 21265 17823 21463 17849
rect 21489 17823 21490 17849
rect 21238 17822 21490 17823
rect 21238 17457 21266 17822
rect 21462 17817 21490 17822
rect 22526 17850 22554 18607
rect 22750 19025 22778 19031
rect 22750 18999 22751 19025
rect 22777 18999 22778 19025
rect 22750 18241 22778 18999
rect 22750 18215 22751 18241
rect 22777 18215 22778 18241
rect 22750 17850 22778 18215
rect 22526 17849 22778 17850
rect 22526 17823 22527 17849
rect 22553 17823 22778 17849
rect 22526 17822 22778 17823
rect 22526 17817 22554 17822
rect 21238 17431 21239 17457
rect 21265 17431 21266 17457
rect 21238 17401 21266 17431
rect 22750 17457 22778 17822
rect 22750 17431 22751 17457
rect 22777 17431 22778 17457
rect 22750 17425 22778 17431
rect 21238 17375 21239 17401
rect 21265 17375 21266 17401
rect 21238 17066 21266 17375
rect 22862 17346 22890 21826
rect 23534 20202 23562 22694
rect 23534 20169 23562 20174
rect 22694 17318 22890 17346
rect 23254 19473 23282 19479
rect 23254 19447 23255 19473
rect 23281 19447 23282 19473
rect 23254 19417 23282 19447
rect 23254 19391 23255 19417
rect 23281 19391 23282 19417
rect 23254 19026 23282 19391
rect 23702 19418 23730 22862
rect 23758 22889 23786 22895
rect 23758 22863 23759 22889
rect 23785 22863 23786 22889
rect 23758 22554 23786 22863
rect 23870 22554 23898 22918
rect 23758 22553 23898 22554
rect 23758 22527 23759 22553
rect 23785 22527 23871 22553
rect 23897 22527 23898 22553
rect 23758 22526 23898 22527
rect 23758 19810 23786 22526
rect 23870 22521 23898 22526
rect 23982 22945 24010 23311
rect 23982 22919 23983 22945
rect 24009 22919 24010 22945
rect 23982 22722 24010 22919
rect 24038 22890 24066 24095
rect 24038 22857 24066 22862
rect 23982 22553 24010 22694
rect 23982 22527 23983 22553
rect 24009 22527 24010 22553
rect 23982 22521 24010 22527
rect 23870 19810 23898 19815
rect 23758 19809 23898 19810
rect 23758 19783 23759 19809
rect 23785 19783 23871 19809
rect 23897 19783 23898 19809
rect 23758 19782 23898 19783
rect 23758 19777 23786 19782
rect 23870 19777 23898 19782
rect 24038 19753 24066 19759
rect 24038 19727 24039 19753
rect 24065 19727 24066 19753
rect 23870 19418 23898 19423
rect 23702 19417 23898 19418
rect 23702 19391 23703 19417
rect 23729 19391 23871 19417
rect 23897 19391 23898 19417
rect 23702 19390 23898 19391
rect 23702 19385 23730 19390
rect 23870 19385 23898 19390
rect 24038 19417 24066 19727
rect 24038 19391 24039 19417
rect 24065 19391 24066 19417
rect 23478 19362 23506 19367
rect 23422 19026 23450 19031
rect 23254 19025 23450 19026
rect 23254 18999 23255 19025
rect 23281 18999 23423 19025
rect 23449 18999 23450 19025
rect 23254 18998 23450 18999
rect 23254 18242 23282 18998
rect 23422 18993 23450 18998
rect 23422 18689 23450 18695
rect 23422 18663 23423 18689
rect 23449 18663 23450 18689
rect 23422 18634 23450 18663
rect 23478 18634 23506 19334
rect 23422 18633 23506 18634
rect 23422 18607 23423 18633
rect 23449 18607 23506 18633
rect 23422 18606 23506 18607
rect 23422 18601 23450 18606
rect 23422 18242 23450 18247
rect 23254 18241 23450 18242
rect 23254 18215 23255 18241
rect 23281 18215 23423 18241
rect 23449 18215 23450 18241
rect 23254 18214 23450 18215
rect 23254 17458 23282 18214
rect 23422 18209 23450 18214
rect 23422 17905 23450 17911
rect 23422 17879 23423 17905
rect 23449 17879 23450 17905
rect 23422 17850 23450 17879
rect 23478 17850 23506 18606
rect 23422 17849 23506 17850
rect 23422 17823 23423 17849
rect 23449 17823 23506 17849
rect 23422 17822 23506 17823
rect 23422 17817 23450 17822
rect 23422 17458 23450 17463
rect 23254 17457 23450 17458
rect 23254 17431 23255 17457
rect 23281 17431 23423 17457
rect 23449 17431 23450 17457
rect 23254 17430 23450 17431
rect 21462 17066 21490 17071
rect 21238 17065 21490 17066
rect 21238 17039 21239 17065
rect 21265 17039 21463 17065
rect 21489 17039 21490 17065
rect 21238 17038 21490 17039
rect 21238 16673 21266 17038
rect 21462 17033 21490 17038
rect 22246 17065 22274 17071
rect 22246 17039 22247 17065
rect 22273 17039 22274 17065
rect 21238 16647 21239 16673
rect 21265 16647 21266 16673
rect 21238 16617 21266 16647
rect 21238 16591 21239 16617
rect 21265 16591 21266 16617
rect 21238 16282 21266 16591
rect 22246 16674 22274 17039
rect 21462 16282 21490 16287
rect 21238 16281 21490 16282
rect 21238 16255 21239 16281
rect 21265 16255 21463 16281
rect 21489 16255 21490 16281
rect 21238 16254 21490 16255
rect 20790 15471 20791 15497
rect 20817 15471 20818 15497
rect 20790 14714 20818 15471
rect 20230 14713 20818 14714
rect 20230 14687 20791 14713
rect 20817 14687 20818 14713
rect 20230 14686 20818 14687
rect 19334 14321 19474 14322
rect 19334 14295 19335 14321
rect 19361 14295 19447 14321
rect 19473 14295 19474 14321
rect 19334 14294 19474 14295
rect 19334 14289 19362 14294
rect 19446 13985 19474 14294
rect 20230 14322 20258 14686
rect 20790 14681 20818 14686
rect 21014 15889 21042 15895
rect 21014 15863 21015 15889
rect 21041 15863 21042 15889
rect 21014 15834 21042 15863
rect 21182 15834 21210 15839
rect 21238 15834 21266 16254
rect 21462 16249 21490 16254
rect 22246 16282 22274 16646
rect 22246 16235 22274 16254
rect 22694 15946 22722 17318
rect 23254 17121 23282 17430
rect 23422 17425 23450 17430
rect 23254 17095 23255 17121
rect 23281 17095 23282 17121
rect 23254 17065 23282 17095
rect 23254 17039 23255 17065
rect 23281 17039 23282 17065
rect 22750 16674 22778 16679
rect 22750 16627 22778 16646
rect 23254 16674 23282 17039
rect 23422 16674 23450 16679
rect 23254 16673 23450 16674
rect 23254 16647 23255 16673
rect 23281 16647 23423 16673
rect 23449 16647 23450 16673
rect 23254 16646 23450 16647
rect 23254 16337 23282 16646
rect 23422 16641 23450 16646
rect 23254 16311 23255 16337
rect 23281 16311 23282 16337
rect 23254 16282 23282 16311
rect 22638 15918 22722 15946
rect 22806 16281 23282 16282
rect 22806 16255 23255 16281
rect 23281 16255 23282 16281
rect 22806 16254 23282 16255
rect 21014 15833 21266 15834
rect 21014 15807 21183 15833
rect 21209 15807 21266 15833
rect 21014 15806 21266 15807
rect 21014 15105 21042 15806
rect 21182 15801 21210 15806
rect 21238 15498 21266 15806
rect 21518 15834 21546 15839
rect 21462 15498 21490 15503
rect 21238 15497 21490 15498
rect 21238 15471 21239 15497
rect 21265 15471 21463 15497
rect 21489 15471 21490 15497
rect 21238 15470 21490 15471
rect 21238 15465 21266 15470
rect 21462 15465 21490 15470
rect 21014 15079 21015 15105
rect 21041 15079 21042 15105
rect 21014 15050 21042 15079
rect 21182 15050 21210 15055
rect 21014 15049 21210 15050
rect 21014 15023 21183 15049
rect 21209 15023 21210 15049
rect 21014 15022 21210 15023
rect 20230 14275 20258 14294
rect 21014 14434 21042 15022
rect 21182 15017 21210 15022
rect 21014 14322 21042 14406
rect 21238 14714 21266 14719
rect 21462 14714 21490 14719
rect 21238 14713 21462 14714
rect 21238 14687 21239 14713
rect 21265 14687 21462 14713
rect 21238 14686 21462 14687
rect 21014 14321 21210 14322
rect 21014 14295 21015 14321
rect 21041 14295 21210 14321
rect 21014 14294 21210 14295
rect 21014 14289 21042 14294
rect 21182 14266 21210 14294
rect 21238 14266 21266 14686
rect 21462 14648 21490 14686
rect 21182 14265 21266 14266
rect 21182 14239 21183 14265
rect 21209 14239 21266 14265
rect 21182 14238 21266 14239
rect 21182 14233 21210 14238
rect 19446 13959 19447 13985
rect 19473 13959 19474 13985
rect 19446 13929 19474 13959
rect 19446 13903 19447 13929
rect 19473 13903 19474 13929
rect 19054 13511 19055 13537
rect 19081 13511 19082 13537
rect 19054 13505 19082 13511
rect 19334 13538 19362 13543
rect 19446 13538 19474 13903
rect 20958 13930 20986 13935
rect 19334 13537 19474 13538
rect 19334 13511 19335 13537
rect 19361 13511 19447 13537
rect 19473 13511 19474 13537
rect 19334 13510 19474 13511
rect 19334 13505 19362 13510
rect 19446 13505 19474 13510
rect 20510 13538 20538 13543
rect 17430 13481 17794 13482
rect 17430 13455 17431 13481
rect 17457 13455 17794 13481
rect 17430 13454 17794 13455
rect 17430 13449 17458 13454
rect 17262 13146 17290 13151
rect 17262 12753 17290 13118
rect 17486 13146 17514 13151
rect 17486 13099 17514 13118
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 17262 12727 17263 12753
rect 17289 12727 17290 12753
rect 17262 12697 17290 12727
rect 17262 12671 17263 12697
rect 17289 12671 17290 12697
rect 17262 12362 17290 12671
rect 17766 12586 17794 13454
rect 18270 13145 18298 13454
rect 18270 13119 18271 13145
rect 18297 13119 18298 13145
rect 18270 13113 18298 13119
rect 18718 13146 18746 13151
rect 18942 13146 18970 13151
rect 18718 13145 18970 13146
rect 18718 13119 18719 13145
rect 18745 13119 18943 13145
rect 18969 13119 18970 13145
rect 18718 13118 18970 13119
rect 17794 12558 17850 12586
rect 17766 12553 17794 12558
rect 17486 12362 17514 12367
rect 17262 12361 17514 12362
rect 17262 12335 17263 12361
rect 17289 12335 17487 12361
rect 17513 12335 17514 12361
rect 17262 12334 17514 12335
rect 17262 12329 17290 12334
rect 17430 11970 17458 12334
rect 17486 12329 17514 12334
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 17430 11913 17458 11942
rect 17430 11887 17431 11913
rect 17457 11887 17458 11913
rect 17430 11881 17458 11887
rect 17766 11970 17794 11975
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 17766 10849 17794 11942
rect 17822 11633 17850 12558
rect 17822 11607 17823 11633
rect 17849 11607 17850 11633
rect 17822 11577 17850 11607
rect 17822 11551 17823 11577
rect 17849 11551 17850 11577
rect 17822 11545 17850 11551
rect 18438 12362 18466 12367
rect 18438 11578 18466 12334
rect 18550 12362 18578 12367
rect 18550 12315 18578 12334
rect 18438 11512 18466 11550
rect 18718 11970 18746 13118
rect 18942 13113 18970 13118
rect 18718 11578 18746 11942
rect 19054 12754 19082 12759
rect 19054 12362 19082 12726
rect 19334 12754 19362 12759
rect 19446 12754 19474 12759
rect 19334 12753 19474 12754
rect 19334 12727 19335 12753
rect 19361 12727 19447 12753
rect 19473 12727 19474 12753
rect 19334 12726 19474 12727
rect 19334 12586 19362 12726
rect 19446 12721 19474 12726
rect 20510 12754 20538 13510
rect 20958 13538 20986 13902
rect 20958 13145 20986 13510
rect 20958 13119 20959 13145
rect 20985 13119 20986 13145
rect 20958 13113 20986 13119
rect 21238 13930 21266 14238
rect 21462 13930 21490 13935
rect 21238 13929 21490 13930
rect 21238 13903 21239 13929
rect 21265 13903 21463 13929
rect 21489 13903 21490 13929
rect 21238 13902 21490 13903
rect 21238 13146 21266 13902
rect 21462 13897 21490 13902
rect 21518 13818 21546 15806
rect 22246 15497 22274 15503
rect 22246 15471 22247 15497
rect 22273 15471 22274 15497
rect 22246 15106 22274 15471
rect 22638 15386 22666 15918
rect 22750 15889 22778 15895
rect 22750 15863 22751 15889
rect 22777 15863 22778 15889
rect 22694 15834 22722 15839
rect 22694 15498 22722 15806
rect 22694 15432 22722 15470
rect 22638 15358 22722 15386
rect 22246 14713 22274 15078
rect 22246 14687 22247 14713
rect 22273 14687 22274 14713
rect 22246 13930 22274 14687
rect 22246 13897 22274 13902
rect 21406 13790 21546 13818
rect 21406 13537 21434 13790
rect 21406 13511 21407 13537
rect 21433 13511 21434 13537
rect 21406 13481 21434 13511
rect 21406 13455 21407 13481
rect 21433 13455 21434 13481
rect 21406 13449 21434 13455
rect 21462 13146 21490 13151
rect 21238 13145 21490 13146
rect 21238 13119 21239 13145
rect 21265 13119 21463 13145
rect 21489 13119 21490 13145
rect 21238 13118 21490 13119
rect 20510 12688 20538 12726
rect 21238 12753 21266 13118
rect 21462 13113 21490 13118
rect 21238 12727 21239 12753
rect 21265 12727 21266 12753
rect 21238 12697 21266 12727
rect 21238 12671 21239 12697
rect 21265 12671 21266 12697
rect 21238 12665 21266 12671
rect 19054 11969 19082 12334
rect 19278 12558 19334 12586
rect 19278 12417 19306 12558
rect 19334 12553 19362 12558
rect 19278 12391 19279 12417
rect 19305 12391 19306 12417
rect 19278 12361 19306 12391
rect 19278 12335 19279 12361
rect 19305 12335 19306 12361
rect 19278 12329 19306 12335
rect 21630 12362 21658 12367
rect 19054 11943 19055 11969
rect 19081 11943 19082 11969
rect 19054 11937 19082 11943
rect 19222 11970 19250 11975
rect 19222 11923 19250 11942
rect 19446 11970 19474 11975
rect 19446 11923 19474 11942
rect 21630 11970 21658 12334
rect 22134 12362 22162 12367
rect 22134 12315 22162 12334
rect 22582 12361 22610 12367
rect 22582 12335 22583 12361
rect 22609 12335 22610 12361
rect 21798 11970 21826 11975
rect 21630 11969 21826 11970
rect 21630 11943 21631 11969
rect 21657 11943 21799 11969
rect 21825 11943 21826 11969
rect 21630 11942 21826 11943
rect 21630 11634 21658 11942
rect 21798 11937 21826 11942
rect 22358 11970 22386 11975
rect 22582 11970 22610 12335
rect 22694 12362 22722 15358
rect 22750 15106 22778 15863
rect 22750 15059 22778 15078
rect 22750 14714 22778 14719
rect 22806 14714 22834 16254
rect 23254 16249 23282 16254
rect 23198 15889 23226 15895
rect 23198 15863 23199 15889
rect 23225 15863 23226 15889
rect 23198 15834 23226 15863
rect 23198 15801 23226 15806
rect 23422 15890 23450 15895
rect 23478 15890 23506 17822
rect 24038 17514 24066 19391
rect 24038 17481 24066 17486
rect 23422 15889 23506 15890
rect 23422 15863 23423 15889
rect 23449 15863 23506 15889
rect 23422 15862 23506 15863
rect 23422 15834 23450 15862
rect 23422 15801 23450 15806
rect 22918 15498 22946 15503
rect 22918 15451 22946 15470
rect 23198 15106 23226 15111
rect 23422 15106 23450 15111
rect 23198 15105 23450 15106
rect 23198 15079 23199 15105
rect 23225 15079 23423 15105
rect 23449 15079 23450 15105
rect 23198 15078 23450 15079
rect 22778 14686 22834 14714
rect 22918 14714 22946 14719
rect 22750 14667 22778 14686
rect 22918 14667 22946 14686
rect 23198 14714 23226 15078
rect 23422 15073 23450 15078
rect 23198 14681 23226 14686
rect 24038 14826 24066 14831
rect 22694 12329 22722 12334
rect 22862 14378 22890 14383
rect 22862 14321 22890 14350
rect 22862 14295 22863 14321
rect 22889 14295 22890 14321
rect 22862 14265 22890 14295
rect 22862 14239 22863 14265
rect 22889 14239 22890 14265
rect 22862 13985 22890 14239
rect 22862 13959 22863 13985
rect 22889 13959 22890 13985
rect 22862 13929 22890 13959
rect 22862 13903 22863 13929
rect 22889 13903 22890 13929
rect 22862 13537 22890 13903
rect 22862 13511 22863 13537
rect 22889 13511 22890 13537
rect 22862 13481 22890 13511
rect 22862 13455 22863 13481
rect 22889 13455 22890 13481
rect 22862 13201 22890 13455
rect 22862 13175 22863 13201
rect 22889 13175 22890 13201
rect 22862 13145 22890 13175
rect 22862 13119 22863 13145
rect 22889 13119 22890 13145
rect 22862 12753 22890 13119
rect 22862 12727 22863 12753
rect 22889 12727 22890 12753
rect 22862 12697 22890 12727
rect 22862 12671 22863 12697
rect 22889 12671 22890 12697
rect 22862 12417 22890 12671
rect 22862 12391 22863 12417
rect 22889 12391 22890 12417
rect 22862 12361 22890 12391
rect 22862 12335 22863 12361
rect 22889 12335 22890 12361
rect 22358 11969 22610 11970
rect 22358 11943 22359 11969
rect 22385 11943 22610 11969
rect 22358 11942 22610 11943
rect 22358 11937 22386 11942
rect 21630 11633 21714 11634
rect 21630 11607 21631 11633
rect 21657 11607 21714 11633
rect 21630 11606 21714 11607
rect 21630 11601 21658 11606
rect 18942 11578 18970 11583
rect 18718 11577 18970 11578
rect 18718 11551 18719 11577
rect 18745 11551 18943 11577
rect 18969 11551 18970 11577
rect 18718 11550 18970 11551
rect 18718 11545 18746 11550
rect 18942 11545 18970 11550
rect 21686 11577 21714 11606
rect 22582 11578 22610 11942
rect 21686 11551 21687 11577
rect 21713 11551 21714 11577
rect 20902 11354 20930 11359
rect 20230 11186 20258 11191
rect 20398 11186 20426 11191
rect 20230 11185 20426 11186
rect 20230 11159 20231 11185
rect 20257 11159 20399 11185
rect 20425 11159 20426 11185
rect 20230 11158 20426 11159
rect 20230 11153 20258 11158
rect 17766 10823 17767 10849
rect 17793 10823 17794 10849
rect 17766 10793 17794 10823
rect 20398 10849 20426 11158
rect 20902 11185 20930 11326
rect 20902 11159 20903 11185
rect 20929 11159 20930 11185
rect 20902 11153 20930 11159
rect 21630 11354 21658 11359
rect 20398 10823 20399 10849
rect 20425 10823 20426 10849
rect 17766 10767 17767 10793
rect 17793 10767 17794 10793
rect 17766 10761 17794 10767
rect 19446 10793 19474 10799
rect 19446 10767 19447 10793
rect 19473 10767 19474 10793
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 17990 10065 18018 10071
rect 17990 10039 17991 10065
rect 18017 10039 18018 10065
rect 17990 10009 18018 10039
rect 19446 10066 19474 10767
rect 20398 10793 20426 10823
rect 20398 10767 20399 10793
rect 20425 10767 20426 10793
rect 19446 10033 19474 10038
rect 20006 10401 20034 10407
rect 20006 10375 20007 10401
rect 20033 10375 20034 10401
rect 20006 10066 20034 10375
rect 20398 10346 20426 10767
rect 21630 10793 21658 11326
rect 21686 11186 21714 11551
rect 22470 11550 22582 11578
rect 21798 11186 21826 11191
rect 21686 11185 21826 11186
rect 21686 11159 21687 11185
rect 21713 11159 21799 11185
rect 21825 11159 21826 11185
rect 21686 11158 21826 11159
rect 21686 11153 21714 11158
rect 21798 10962 21826 11158
rect 22358 11186 22386 11191
rect 22470 11186 22498 11550
rect 22582 11531 22610 11550
rect 22862 11969 22890 12335
rect 24038 14321 24066 14798
rect 24038 14295 24039 14321
rect 24065 14295 24066 14321
rect 24038 13929 24066 14295
rect 24038 13903 24039 13929
rect 24065 13903 24066 13929
rect 24038 13537 24066 13903
rect 24038 13511 24039 13537
rect 24065 13511 24066 13537
rect 24038 13145 24066 13511
rect 24038 13119 24039 13145
rect 24065 13119 24066 13145
rect 24038 12753 24066 13119
rect 24038 12727 24039 12753
rect 24065 12727 24066 12753
rect 24038 12361 24066 12727
rect 24038 12335 24039 12361
rect 24065 12335 24066 12361
rect 22862 11943 22863 11969
rect 22889 11943 22890 11969
rect 22862 11913 22890 11943
rect 22862 11887 22863 11913
rect 22889 11887 22890 11913
rect 22862 11633 22890 11887
rect 22862 11607 22863 11633
rect 22889 11607 22890 11633
rect 22862 11577 22890 11607
rect 22862 11551 22863 11577
rect 22889 11551 22890 11577
rect 22358 11185 22498 11186
rect 22358 11159 22359 11185
rect 22385 11159 22498 11185
rect 22358 11158 22498 11159
rect 22358 11153 22386 11158
rect 21798 10929 21826 10934
rect 21630 10767 21631 10793
rect 21657 10767 21658 10793
rect 20398 10313 20426 10318
rect 20902 10401 20930 10407
rect 20902 10375 20903 10401
rect 20929 10375 20930 10401
rect 20902 10346 20930 10375
rect 21462 10402 21490 10407
rect 21630 10402 21658 10767
rect 21854 10906 21882 10911
rect 21854 10793 21882 10878
rect 21854 10767 21855 10793
rect 21881 10767 21882 10793
rect 21854 10761 21882 10767
rect 22078 10906 22106 10911
rect 22078 10793 22106 10878
rect 22078 10767 22079 10793
rect 22105 10767 22106 10793
rect 21462 10401 21714 10402
rect 21462 10375 21463 10401
rect 21489 10375 21714 10401
rect 21462 10374 21714 10375
rect 21462 10369 21490 10374
rect 20902 10299 20930 10318
rect 20006 10033 20034 10038
rect 21182 10066 21210 10071
rect 17990 9983 17991 10009
rect 18017 9983 18018 10009
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 17430 9617 17458 9623
rect 17430 9591 17431 9617
rect 17457 9591 17458 9617
rect 17430 9562 17458 9591
rect 17430 9515 17458 9534
rect 17990 9562 18018 9983
rect 17990 9281 18018 9534
rect 21182 9617 21210 10038
rect 21686 10009 21714 10374
rect 22078 10401 22106 10767
rect 22078 10375 22079 10401
rect 22105 10375 22106 10401
rect 22078 10346 22106 10375
rect 22134 10346 22162 10351
rect 22526 10346 22554 10351
rect 22078 10345 22386 10346
rect 22078 10319 22135 10345
rect 22161 10319 22386 10345
rect 22078 10318 22386 10319
rect 22134 10313 22162 10318
rect 21686 9983 21687 10009
rect 21713 9983 21714 10009
rect 21686 9977 21714 9983
rect 21182 9591 21183 9617
rect 21209 9591 21210 9617
rect 21182 9450 21210 9591
rect 17990 9255 17991 9281
rect 18017 9255 18018 9281
rect 17990 9225 18018 9255
rect 19222 9281 19250 9287
rect 19222 9255 19223 9281
rect 19249 9255 19250 9281
rect 17990 9199 17991 9225
rect 18017 9199 18018 9225
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 17150 8833 17234 8834
rect 17150 8807 17151 8833
rect 17177 8807 17234 8833
rect 17150 8806 17234 8807
rect 17150 8801 17178 8806
rect 17206 8778 17234 8806
rect 17206 8777 17290 8778
rect 17206 8751 17207 8777
rect 17233 8751 17290 8777
rect 17206 8750 17290 8751
rect 17206 8745 17234 8750
rect 17094 8415 17095 8441
rect 17121 8415 17122 8441
rect 17094 8050 17122 8415
rect 17262 8442 17290 8750
rect 17486 8442 17514 8447
rect 17262 8441 17514 8442
rect 17262 8415 17263 8441
rect 17289 8415 17487 8441
rect 17513 8415 17514 8441
rect 17262 8414 17514 8415
rect 17262 8409 17290 8414
rect 17094 7658 17122 8022
rect 17430 8049 17458 8414
rect 17486 8409 17514 8414
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 17430 8023 17431 8049
rect 17457 8023 17458 8049
rect 17430 7994 17458 8023
rect 17430 7928 17458 7966
rect 17766 7994 17794 7999
rect 17094 6873 17122 7630
rect 17374 7658 17402 7663
rect 17486 7658 17514 7663
rect 17374 7657 17514 7658
rect 17374 7631 17375 7657
rect 17401 7631 17487 7657
rect 17513 7631 17514 7657
rect 17374 7630 17514 7631
rect 17374 7625 17402 7630
rect 17486 7602 17514 7630
rect 17430 7266 17458 7271
rect 17486 7266 17514 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 17430 7265 17514 7266
rect 17430 7239 17431 7265
rect 17457 7239 17514 7265
rect 17430 7238 17514 7239
rect 17430 7209 17458 7238
rect 17430 7183 17431 7209
rect 17457 7183 17458 7209
rect 17262 6874 17290 6879
rect 17430 6874 17458 7183
rect 17486 6874 17514 6879
rect 17094 6847 17095 6873
rect 17121 6847 17122 6873
rect 17094 6841 17122 6847
rect 17206 6873 17514 6874
rect 17206 6847 17263 6873
rect 17289 6847 17487 6873
rect 17513 6847 17514 6873
rect 17206 6846 17514 6847
rect 17206 6481 17234 6846
rect 17262 6841 17290 6846
rect 17486 6841 17514 6846
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17206 6455 17207 6481
rect 17233 6455 17234 6481
rect 17206 6425 17234 6455
rect 17206 6399 17207 6425
rect 17233 6399 17234 6425
rect 17206 6146 17234 6399
rect 16814 6090 16842 6095
rect 16758 6062 16814 6090
rect 14798 5671 14799 5697
rect 14825 5671 14826 5697
rect 14798 4913 14826 5671
rect 15918 5810 15946 5815
rect 15918 5697 15946 5782
rect 15918 5671 15919 5697
rect 15945 5671 15946 5697
rect 15918 5641 15946 5671
rect 15918 5615 15919 5641
rect 15945 5615 15946 5641
rect 14798 4887 14799 4913
rect 14825 4887 14826 4913
rect 14798 4881 14826 4887
rect 15470 5361 15498 5367
rect 15470 5335 15471 5361
rect 15497 5335 15498 5361
rect 15470 5305 15498 5335
rect 15470 5279 15471 5305
rect 15497 5279 15498 5305
rect 15470 5026 15498 5279
rect 14574 4495 14575 4521
rect 14601 4495 14602 4521
rect 14574 4489 14602 4495
rect 15470 4577 15498 4998
rect 15918 5026 15946 5615
rect 15918 4913 15946 4998
rect 15918 4887 15919 4913
rect 15945 4887 15946 4913
rect 15918 4857 15946 4887
rect 15918 4831 15919 4857
rect 15945 4831 15946 4857
rect 15918 4825 15946 4831
rect 16534 5698 16562 5703
rect 16758 5698 16786 6062
rect 16814 6024 16842 6062
rect 17206 5922 17234 6118
rect 17766 6145 17794 7966
rect 17990 7602 18018 9199
rect 18550 9225 18578 9231
rect 18550 9199 18551 9225
rect 18577 9199 18578 9225
rect 18550 8441 18578 9199
rect 19222 9225 19250 9255
rect 19222 9199 19223 9225
rect 19249 9199 19250 9225
rect 18550 8415 18551 8441
rect 18577 8415 18578 8441
rect 18550 8386 18578 8415
rect 18550 7658 18578 8358
rect 19054 8833 19082 8839
rect 19054 8807 19055 8833
rect 19081 8807 19082 8833
rect 19054 8386 19082 8807
rect 19054 8050 19082 8358
rect 19054 8003 19082 8022
rect 19222 8834 19250 9199
rect 21182 9226 21210 9422
rect 22358 9617 22386 10318
rect 22526 10094 22554 10318
rect 22526 10066 22610 10094
rect 22582 10009 22610 10038
rect 22582 9983 22583 10009
rect 22609 9983 22610 10009
rect 22582 9977 22610 9983
rect 22862 10066 22890 11551
rect 23814 12138 23842 12143
rect 23814 11354 23842 12110
rect 22974 11185 23002 11191
rect 22974 11159 22975 11185
rect 23001 11159 23002 11185
rect 22974 11129 23002 11159
rect 22974 11103 22975 11129
rect 23001 11103 23002 11129
rect 22974 10849 23002 11103
rect 22974 10823 22975 10849
rect 23001 10823 23002 10849
rect 22974 10793 23002 10823
rect 22974 10767 22975 10793
rect 23001 10767 23002 10793
rect 22974 10401 23002 10767
rect 22974 10375 22975 10401
rect 23001 10375 23002 10401
rect 22974 10345 23002 10375
rect 22974 10319 22975 10345
rect 23001 10319 23002 10345
rect 22974 10094 23002 10319
rect 22358 9591 22359 9617
rect 22385 9591 22386 9617
rect 22358 9561 22386 9591
rect 22358 9535 22359 9561
rect 22385 9535 22386 9561
rect 21406 9226 21434 9231
rect 21182 9225 21434 9226
rect 21182 9199 21407 9225
rect 21433 9199 21434 9225
rect 21182 9198 21434 9199
rect 21406 9193 21434 9198
rect 22358 9226 22386 9535
rect 22358 9193 22386 9198
rect 22582 9281 22610 9287
rect 22582 9255 22583 9281
rect 22609 9255 22610 9281
rect 22582 9226 22610 9255
rect 22582 9179 22610 9198
rect 19446 8834 19474 8839
rect 19222 8833 19474 8834
rect 19222 8807 19223 8833
rect 19249 8807 19447 8833
rect 19473 8807 19474 8833
rect 19222 8806 19474 8807
rect 19222 8497 19250 8806
rect 19446 8801 19474 8806
rect 22862 8833 22890 10038
rect 22862 8807 22863 8833
rect 22889 8807 22890 8833
rect 19222 8471 19223 8497
rect 19249 8471 19250 8497
rect 19222 8441 19250 8471
rect 19222 8415 19223 8441
rect 19249 8415 19250 8441
rect 19222 8050 19250 8415
rect 22862 8777 22890 8807
rect 22862 8751 22863 8777
rect 22889 8751 22890 8777
rect 22862 8497 22890 8751
rect 22862 8471 22863 8497
rect 22889 8471 22890 8497
rect 22862 8441 22890 8471
rect 22862 8415 22863 8441
rect 22889 8415 22890 8441
rect 19446 8050 19474 8055
rect 19222 8049 19474 8050
rect 19222 8023 19223 8049
rect 19249 8023 19447 8049
rect 19473 8023 19474 8049
rect 19222 8022 19474 8023
rect 18550 7592 18578 7630
rect 18718 7657 18746 7663
rect 18718 7631 18719 7657
rect 18745 7631 18746 7657
rect 18718 7602 18746 7631
rect 17990 7569 18018 7574
rect 18718 7569 18746 7574
rect 18942 7657 18970 7663
rect 18942 7631 18943 7657
rect 18969 7631 18970 7657
rect 18942 7602 18970 7631
rect 18942 7569 18970 7574
rect 19222 7602 19250 8022
rect 19446 8017 19474 8022
rect 20230 8049 20258 8055
rect 20230 8023 20231 8049
rect 20257 8023 20258 8049
rect 19222 7569 19250 7574
rect 20230 7546 20258 8023
rect 21014 8049 21042 8055
rect 21014 8023 21015 8049
rect 21041 8023 21042 8049
rect 21014 7994 21042 8023
rect 22806 8050 22834 8055
rect 21182 7994 21210 7999
rect 21014 7993 21266 7994
rect 21014 7967 21183 7993
rect 21209 7967 21266 7993
rect 21014 7966 21266 7967
rect 18774 7266 18802 7271
rect 17766 6119 17767 6145
rect 17793 6119 17794 6145
rect 17766 6089 17794 6119
rect 17766 6063 17767 6089
rect 17793 6063 17794 6089
rect 16534 5697 16842 5698
rect 16534 5671 16535 5697
rect 16561 5671 16842 5697
rect 16534 5670 16842 5671
rect 16534 4913 16562 5670
rect 16814 5305 16842 5670
rect 16814 5279 16815 5305
rect 16841 5279 16842 5305
rect 16814 5273 16842 5279
rect 17094 5306 17122 5311
rect 16534 4887 16535 4913
rect 16561 4887 16562 4913
rect 15470 4551 15471 4577
rect 15497 4551 15498 4577
rect 15470 4522 15498 4551
rect 15470 4521 15610 4522
rect 15470 4495 15471 4521
rect 15497 4495 15610 4521
rect 15470 4494 15610 4495
rect 15470 4489 15498 4494
rect 15470 4186 15498 4191
rect 14182 4129 14266 4130
rect 14182 4103 14183 4129
rect 14209 4103 14266 4129
rect 14182 4102 14266 4103
rect 15078 4130 15106 4135
rect 14182 4073 14210 4102
rect 14182 4047 14183 4073
rect 14209 4047 14210 4073
rect 14182 4041 14210 4047
rect 14126 3319 14127 3345
rect 14153 3319 14154 3345
rect 14126 3290 14154 3319
rect 13118 2927 13119 2953
rect 13145 2927 13146 2953
rect 13118 2562 13146 2927
rect 14014 3289 14154 3290
rect 14014 3263 14127 3289
rect 14153 3263 14154 3289
rect 14014 3262 14154 3263
rect 14014 3009 14042 3262
rect 14126 3257 14154 3262
rect 14574 3738 14602 3743
rect 14574 3346 14602 3710
rect 14014 2983 14015 3009
rect 14041 2983 14042 3009
rect 14014 2953 14042 2983
rect 14014 2927 14015 2953
rect 14041 2927 14042 2953
rect 13174 2562 13202 2567
rect 13146 2561 13202 2562
rect 13146 2535 13175 2561
rect 13201 2535 13202 2561
rect 13146 2534 13202 2535
rect 13118 2169 13146 2534
rect 13174 2529 13202 2534
rect 14014 2562 14042 2927
rect 14574 2953 14602 3318
rect 15078 3738 15106 4102
rect 15078 3345 15106 3710
rect 15470 3793 15498 4158
rect 15470 3767 15471 3793
rect 15497 3767 15498 3793
rect 15470 3737 15498 3767
rect 15470 3711 15471 3737
rect 15497 3711 15498 3737
rect 15470 3705 15498 3711
rect 15582 3346 15610 4494
rect 16534 4214 16562 4887
rect 17094 4522 17122 5278
rect 15918 4186 15946 4191
rect 15918 4129 15946 4158
rect 15918 4103 15919 4129
rect 15945 4103 15946 4129
rect 15918 4073 15946 4103
rect 15918 4047 15919 4073
rect 15945 4047 15946 4073
rect 16254 4186 16562 4214
rect 16814 4521 17122 4522
rect 16814 4495 17095 4521
rect 17121 4495 17122 4521
rect 16814 4494 17122 4495
rect 16254 4130 16282 4186
rect 16254 4064 16282 4102
rect 15918 4041 15946 4047
rect 16814 3737 16842 4494
rect 17094 4489 17122 4494
rect 16814 3711 16815 3737
rect 16841 3711 16842 3737
rect 16254 3346 16282 3351
rect 15078 3319 15079 3345
rect 15105 3319 15106 3345
rect 15078 3313 15106 3319
rect 15470 3345 15778 3346
rect 15470 3319 15583 3345
rect 15609 3319 15778 3345
rect 15470 3318 15778 3319
rect 14574 2927 14575 2953
rect 14601 2927 14602 2953
rect 14574 2921 14602 2927
rect 15470 3009 15498 3318
rect 15582 3313 15610 3318
rect 15750 3289 15778 3318
rect 15750 3263 15751 3289
rect 15777 3263 15778 3289
rect 15750 3257 15778 3263
rect 15470 2983 15471 3009
rect 15497 2983 15498 3009
rect 15470 2953 15498 2983
rect 15470 2927 15471 2953
rect 15497 2927 15498 2953
rect 14798 2562 14826 2567
rect 14014 2561 14154 2562
rect 14014 2535 14015 2561
rect 14041 2535 14154 2561
rect 14014 2534 14154 2535
rect 13118 2143 13119 2169
rect 13145 2143 13146 2169
rect 12278 1721 12306 1750
rect 12894 1745 12922 1750
rect 12950 1778 12978 1783
rect 13118 1778 13146 2143
rect 14014 2225 14042 2534
rect 14126 2505 14154 2534
rect 14126 2479 14127 2505
rect 14153 2479 14154 2505
rect 14126 2473 14154 2479
rect 14014 2199 14015 2225
rect 14041 2199 14042 2225
rect 14014 2169 14042 2199
rect 14014 2143 14015 2169
rect 14041 2143 14042 2169
rect 14014 2137 14042 2143
rect 14294 2169 14322 2175
rect 14294 2143 14295 2169
rect 14321 2143 14322 2169
rect 14294 2058 14322 2143
rect 14294 2025 14322 2030
rect 14518 2058 14546 2063
rect 12950 1777 13146 1778
rect 12950 1751 12951 1777
rect 12977 1751 13146 1777
rect 12950 1750 13146 1751
rect 13846 1778 13874 1783
rect 12950 1745 12978 1750
rect 12278 1695 12279 1721
rect 12305 1695 12306 1721
rect 12278 1689 12306 1695
rect 13846 1721 13874 1750
rect 13846 1695 13847 1721
rect 13873 1695 13874 1721
rect 13846 1689 13874 1695
rect 14518 400 14546 2030
rect 14798 2058 14826 2534
rect 14798 2025 14826 2030
rect 15358 2562 15386 2567
rect 15470 2562 15498 2927
rect 15358 2561 15498 2562
rect 15358 2535 15359 2561
rect 15385 2535 15471 2561
rect 15497 2535 15498 2561
rect 15358 2534 15498 2535
rect 15358 2225 15386 2534
rect 15470 2529 15498 2534
rect 16254 2562 16282 3318
rect 16814 3346 16842 3711
rect 16814 3313 16842 3318
rect 17206 4129 17234 5894
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17430 5698 17458 5703
rect 17430 5641 17458 5670
rect 17430 5615 17431 5641
rect 17457 5615 17458 5641
rect 17430 4913 17458 5615
rect 17766 5698 17794 6063
rect 18270 6873 18298 6879
rect 18270 6847 18271 6873
rect 18297 6847 18298 6873
rect 18270 6090 18298 6847
rect 18718 6874 18746 6879
rect 18270 6043 18298 6062
rect 18662 6090 18690 6095
rect 17766 5362 17794 5670
rect 17766 5305 17794 5334
rect 17766 5279 17767 5305
rect 17793 5279 17794 5305
rect 17766 5273 17794 5279
rect 18550 5698 18578 5703
rect 18550 5306 18578 5670
rect 18550 5240 18578 5278
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17430 4887 17431 4913
rect 17457 4887 17458 4913
rect 17430 4858 17458 4887
rect 17430 4857 17514 4858
rect 17430 4831 17431 4857
rect 17457 4831 17514 4857
rect 17430 4830 17514 4831
rect 17430 4825 17458 4830
rect 17374 4522 17402 4527
rect 17486 4522 17514 4830
rect 17374 4521 17514 4522
rect 17374 4495 17375 4521
rect 17401 4495 17487 4521
rect 17513 4495 17514 4521
rect 17374 4494 17514 4495
rect 17374 4489 17402 4494
rect 17430 4186 17458 4494
rect 17486 4489 17514 4494
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17430 4153 17458 4158
rect 17206 4103 17207 4129
rect 17233 4103 17234 4129
rect 17206 4073 17234 4103
rect 17206 4047 17207 4073
rect 17233 4047 17234 4073
rect 17206 3738 17234 4047
rect 17262 3738 17290 3743
rect 17486 3738 17514 3743
rect 17206 3737 17514 3738
rect 17206 3711 17263 3737
rect 17289 3711 17487 3737
rect 17513 3711 17514 3737
rect 17206 3710 17514 3711
rect 17206 3345 17234 3710
rect 17262 3705 17290 3710
rect 17486 3705 17514 3710
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17206 3319 17207 3345
rect 17233 3319 17234 3345
rect 17206 3289 17234 3319
rect 17206 3263 17207 3289
rect 17233 3263 17234 3289
rect 17206 3257 17234 3263
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 16254 2529 16282 2534
rect 15358 2199 15359 2225
rect 15385 2199 15386 2225
rect 15358 2169 15386 2199
rect 15358 2143 15359 2169
rect 15385 2143 15386 2169
rect 15358 1778 15386 2143
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 15358 1745 15386 1750
rect 18662 400 18690 6062
rect 18718 5362 18746 6846
rect 18774 6481 18802 7238
rect 19222 7266 19250 7271
rect 19446 7266 19474 7271
rect 19222 7265 19474 7266
rect 19222 7239 19223 7265
rect 19249 7239 19447 7265
rect 19473 7239 19474 7265
rect 19222 7238 19474 7239
rect 18942 6874 18970 6879
rect 18942 6827 18970 6846
rect 19222 6874 19250 7238
rect 19446 7233 19474 7238
rect 20230 7266 20258 7518
rect 20790 7657 20818 7663
rect 20790 7631 20791 7657
rect 20817 7631 20818 7657
rect 20790 7546 20818 7631
rect 20790 7513 20818 7518
rect 20230 7219 20258 7238
rect 21014 7265 21042 7966
rect 21182 7961 21210 7966
rect 21238 7658 21266 7966
rect 21462 7658 21490 7663
rect 21238 7657 21490 7658
rect 21238 7631 21239 7657
rect 21265 7631 21463 7657
rect 21489 7631 21490 7657
rect 21238 7630 21490 7631
rect 21238 7625 21266 7630
rect 21462 7625 21490 7630
rect 21014 7239 21015 7265
rect 21041 7239 21042 7265
rect 19222 6841 19250 6846
rect 21014 7210 21042 7239
rect 21182 7210 21210 7215
rect 21014 7209 21210 7210
rect 21014 7183 21183 7209
rect 21209 7183 21210 7209
rect 21014 7182 21210 7183
rect 18774 6455 18775 6481
rect 18801 6455 18802 6481
rect 18774 6090 18802 6455
rect 19222 6482 19250 6487
rect 19446 6482 19474 6487
rect 19222 6481 19446 6482
rect 19222 6455 19223 6481
rect 19249 6455 19446 6481
rect 19222 6454 19446 6455
rect 18774 6057 18802 6062
rect 18830 6146 18858 6151
rect 18830 6090 18858 6118
rect 19222 6146 19250 6454
rect 19446 6416 19474 6454
rect 20230 6481 20258 6487
rect 20230 6455 20231 6481
rect 20257 6455 20258 6481
rect 19222 6113 19250 6118
rect 18942 6090 18970 6095
rect 18830 6089 18970 6090
rect 18830 6063 18831 6089
rect 18857 6063 18943 6089
rect 18969 6063 18970 6089
rect 18830 6062 18970 6063
rect 18830 6057 18858 6062
rect 18942 6057 18970 6062
rect 19054 5698 19082 5703
rect 19054 5651 19082 5670
rect 19222 5698 19250 5703
rect 19446 5698 19474 5703
rect 19222 5697 19474 5698
rect 19222 5671 19223 5697
rect 19249 5671 19447 5697
rect 19473 5671 19474 5697
rect 19222 5670 19474 5671
rect 18718 5305 18746 5334
rect 18718 5279 18719 5305
rect 18745 5279 18746 5305
rect 18718 5273 18746 5279
rect 18942 5362 18970 5367
rect 18942 5305 18970 5334
rect 19222 5362 19250 5670
rect 19446 5665 19474 5670
rect 20230 5698 20258 6455
rect 20678 6482 20706 6487
rect 20678 6435 20706 6454
rect 21014 6482 21042 7182
rect 21182 7177 21210 7182
rect 21014 6435 21042 6454
rect 20230 5665 20258 5670
rect 19222 5329 19250 5334
rect 18942 5279 18943 5305
rect 18969 5279 18970 5305
rect 18942 5273 18970 5279
rect 22806 400 22834 8022
rect 22862 7713 22890 8415
rect 22862 7687 22863 7713
rect 22889 7687 22890 7713
rect 22862 7657 22890 7687
rect 22862 7631 22863 7657
rect 22889 7631 22890 7657
rect 22862 6929 22890 7631
rect 22862 6903 22863 6929
rect 22889 6903 22890 6929
rect 22862 6873 22890 6903
rect 22862 6847 22863 6873
rect 22889 6847 22890 6873
rect 22862 6481 22890 6847
rect 22862 6455 22863 6481
rect 22889 6455 22890 6481
rect 22862 6425 22890 6455
rect 22862 6399 22863 6425
rect 22889 6399 22890 6425
rect 22862 6393 22890 6399
rect 22918 10066 23002 10094
rect 23758 10402 23786 10407
rect 22918 10065 22946 10066
rect 22918 10039 22919 10065
rect 22945 10039 22946 10065
rect 22918 10009 22946 10039
rect 22918 9983 22919 10009
rect 22945 9983 22946 10009
rect 22918 9617 22946 9983
rect 23758 10009 23786 10374
rect 23758 9983 23759 10009
rect 23785 9983 23786 10009
rect 23758 9977 23786 9983
rect 22918 9591 22919 9617
rect 22945 9591 22946 9617
rect 22918 9561 22946 9591
rect 22918 9535 22919 9561
rect 22945 9535 22946 9561
rect 22918 9281 22946 9535
rect 22918 9255 22919 9281
rect 22945 9255 22946 9281
rect 22918 9226 22946 9255
rect 22918 8049 22946 9198
rect 23758 9618 23786 9623
rect 23814 9618 23842 11326
rect 24038 11969 24066 12335
rect 24038 11943 24039 11969
rect 24065 11943 24066 11969
rect 24038 11578 24066 11943
rect 24038 11185 24066 11550
rect 24038 11159 24039 11185
rect 24065 11159 24066 11185
rect 24038 10793 24066 11159
rect 24038 10767 24039 10793
rect 24065 10767 24066 10793
rect 24038 10402 24066 10767
rect 24038 10336 24066 10374
rect 23758 9617 23842 9618
rect 23758 9591 23759 9617
rect 23785 9591 23842 9617
rect 23758 9590 23842 9591
rect 23758 9225 23786 9590
rect 23758 9199 23759 9225
rect 23785 9199 23786 9225
rect 23758 8833 23786 9199
rect 23758 8807 23759 8833
rect 23785 8807 23786 8833
rect 23758 8441 23786 8807
rect 23758 8415 23759 8441
rect 23785 8415 23786 8441
rect 23758 8409 23786 8415
rect 22918 8023 22919 8049
rect 22945 8023 22946 8049
rect 22918 7993 22946 8023
rect 22918 7967 22919 7993
rect 22945 7967 22946 7993
rect 22918 7265 22946 7967
rect 24038 8049 24066 8055
rect 24038 8023 24039 8049
rect 24065 8023 24066 8049
rect 24038 7657 24066 8023
rect 24038 7631 24039 7657
rect 24065 7631 24066 7657
rect 22918 7239 22919 7265
rect 22945 7239 22946 7265
rect 22918 7209 22946 7239
rect 22918 7183 22919 7209
rect 22945 7183 22946 7209
rect 22918 4129 22946 7183
rect 23814 7265 23842 7271
rect 23814 7239 23815 7265
rect 23841 7239 23842 7265
rect 23758 6874 23786 6879
rect 22918 4103 22919 4129
rect 22945 4103 22946 4129
rect 22918 4073 22946 4103
rect 22918 4047 22919 4073
rect 22945 4047 22946 4073
rect 22918 4041 22946 4047
rect 23702 6873 23786 6874
rect 23702 6847 23759 6873
rect 23785 6847 23786 6873
rect 23702 6846 23786 6847
rect 23702 3962 23730 6846
rect 23758 6841 23786 6846
rect 23814 6481 23842 7239
rect 24038 6762 24066 7631
rect 24038 6729 24066 6734
rect 23814 6455 23815 6481
rect 23841 6455 23842 6481
rect 23814 4074 23842 6455
rect 23814 4041 23842 4046
rect 24038 4129 24066 4135
rect 24038 4103 24039 4129
rect 24065 4103 24066 4129
rect 24038 3962 24066 4103
rect 23702 3934 24066 3962
rect 24038 1386 24066 3934
rect 24038 1353 24066 1358
rect 2072 0 2128 400
rect 6216 0 6272 400
rect 10360 0 10416 400
rect 14504 0 14560 400
rect 18648 0 18704 400
rect 22792 0 22848 400
<< via2 >>
rect 1750 32774 1778 32802
rect 1358 26894 1386 26922
rect 1582 25662 1610 25690
rect 1750 25662 1778 25690
rect 1806 28406 1834 28434
rect 1358 24038 1386 24066
rect 1358 23534 1386 23562
rect 2238 33333 2266 33334
rect 2238 33307 2239 33333
rect 2239 33307 2265 33333
rect 2265 33307 2266 33333
rect 2238 33306 2266 33307
rect 2290 33333 2318 33334
rect 2290 33307 2291 33333
rect 2291 33307 2317 33333
rect 2317 33307 2318 33333
rect 2290 33306 2318 33307
rect 2342 33333 2370 33334
rect 2342 33307 2343 33333
rect 2343 33307 2369 33333
rect 2369 33307 2370 33333
rect 2342 33306 2370 33307
rect 2238 32549 2266 32550
rect 2238 32523 2239 32549
rect 2239 32523 2265 32549
rect 2265 32523 2266 32549
rect 2238 32522 2266 32523
rect 2290 32549 2318 32550
rect 2290 32523 2291 32549
rect 2291 32523 2317 32549
rect 2317 32523 2318 32549
rect 2290 32522 2318 32523
rect 2342 32549 2370 32550
rect 2342 32523 2343 32549
rect 2343 32523 2369 32549
rect 2369 32523 2370 32549
rect 2342 32522 2370 32523
rect 2238 31765 2266 31766
rect 2238 31739 2239 31765
rect 2239 31739 2265 31765
rect 2265 31739 2266 31765
rect 2238 31738 2266 31739
rect 2290 31765 2318 31766
rect 2290 31739 2291 31765
rect 2291 31739 2317 31765
rect 2317 31739 2318 31765
rect 2290 31738 2318 31739
rect 2342 31765 2370 31766
rect 2342 31739 2343 31765
rect 2343 31739 2369 31765
rect 2369 31739 2370 31765
rect 2342 31738 2370 31739
rect 2238 30981 2266 30982
rect 2238 30955 2239 30981
rect 2239 30955 2265 30981
rect 2265 30955 2266 30981
rect 2238 30954 2266 30955
rect 2290 30981 2318 30982
rect 2290 30955 2291 30981
rect 2291 30955 2317 30981
rect 2317 30955 2318 30981
rect 2290 30954 2318 30955
rect 2342 30981 2370 30982
rect 2342 30955 2343 30981
rect 2343 30955 2369 30981
rect 2369 30955 2370 30981
rect 2342 30954 2370 30955
rect 2238 30197 2266 30198
rect 2238 30171 2239 30197
rect 2239 30171 2265 30197
rect 2265 30171 2266 30197
rect 2238 30170 2266 30171
rect 2290 30197 2318 30198
rect 2290 30171 2291 30197
rect 2291 30171 2317 30197
rect 2317 30171 2318 30197
rect 2290 30170 2318 30171
rect 2342 30197 2370 30198
rect 2342 30171 2343 30197
rect 2343 30171 2369 30197
rect 2369 30171 2370 30197
rect 2342 30170 2370 30171
rect 2238 29413 2266 29414
rect 2238 29387 2239 29413
rect 2239 29387 2265 29413
rect 2265 29387 2266 29413
rect 2238 29386 2266 29387
rect 2290 29413 2318 29414
rect 2290 29387 2291 29413
rect 2291 29387 2317 29413
rect 2317 29387 2318 29413
rect 2290 29386 2318 29387
rect 2342 29413 2370 29414
rect 2342 29387 2343 29413
rect 2343 29387 2369 29413
rect 2369 29387 2370 29413
rect 2342 29386 2370 29387
rect 2238 28629 2266 28630
rect 2238 28603 2239 28629
rect 2239 28603 2265 28629
rect 2265 28603 2266 28629
rect 2238 28602 2266 28603
rect 2290 28629 2318 28630
rect 2290 28603 2291 28629
rect 2291 28603 2317 28629
rect 2317 28603 2318 28629
rect 2290 28602 2318 28603
rect 2342 28629 2370 28630
rect 2342 28603 2343 28629
rect 2343 28603 2369 28629
rect 2369 28603 2370 28629
rect 2342 28602 2370 28603
rect 2238 27845 2266 27846
rect 2238 27819 2239 27845
rect 2239 27819 2265 27845
rect 2265 27819 2266 27845
rect 2238 27818 2266 27819
rect 2290 27845 2318 27846
rect 2290 27819 2291 27845
rect 2291 27819 2317 27845
rect 2317 27819 2318 27845
rect 2290 27818 2318 27819
rect 2342 27845 2370 27846
rect 2342 27819 2343 27845
rect 2343 27819 2369 27845
rect 2369 27819 2370 27845
rect 2342 27818 2370 27819
rect 9918 32941 9946 32942
rect 9918 32915 9919 32941
rect 9919 32915 9945 32941
rect 9945 32915 9946 32941
rect 9918 32914 9946 32915
rect 9970 32941 9998 32942
rect 9970 32915 9971 32941
rect 9971 32915 9997 32941
rect 9997 32915 9998 32941
rect 9970 32914 9998 32915
rect 10022 32941 10050 32942
rect 10022 32915 10023 32941
rect 10023 32915 10049 32941
rect 10049 32915 10050 32941
rect 10022 32914 10050 32915
rect 9918 32157 9946 32158
rect 9918 32131 9919 32157
rect 9919 32131 9945 32157
rect 9945 32131 9946 32157
rect 9918 32130 9946 32131
rect 9970 32157 9998 32158
rect 9970 32131 9971 32157
rect 9971 32131 9997 32157
rect 9997 32131 9998 32157
rect 9970 32130 9998 32131
rect 10022 32157 10050 32158
rect 10022 32131 10023 32157
rect 10023 32131 10049 32157
rect 10049 32131 10050 32157
rect 10022 32130 10050 32131
rect 9918 31373 9946 31374
rect 9918 31347 9919 31373
rect 9919 31347 9945 31373
rect 9945 31347 9946 31373
rect 9918 31346 9946 31347
rect 9970 31373 9998 31374
rect 9970 31347 9971 31373
rect 9971 31347 9997 31373
rect 9997 31347 9998 31373
rect 9970 31346 9998 31347
rect 10022 31373 10050 31374
rect 10022 31347 10023 31373
rect 10023 31347 10049 31373
rect 10049 31347 10050 31373
rect 10022 31346 10050 31347
rect 9918 30589 9946 30590
rect 9918 30563 9919 30589
rect 9919 30563 9945 30589
rect 9945 30563 9946 30589
rect 9918 30562 9946 30563
rect 9970 30589 9998 30590
rect 9970 30563 9971 30589
rect 9971 30563 9997 30589
rect 9997 30563 9998 30589
rect 9970 30562 9998 30563
rect 10022 30589 10050 30590
rect 10022 30563 10023 30589
rect 10023 30563 10049 30589
rect 10049 30563 10050 30589
rect 10022 30562 10050 30563
rect 9918 29805 9946 29806
rect 9918 29779 9919 29805
rect 9919 29779 9945 29805
rect 9945 29779 9946 29805
rect 9918 29778 9946 29779
rect 9970 29805 9998 29806
rect 9970 29779 9971 29805
rect 9971 29779 9997 29805
rect 9997 29779 9998 29805
rect 9970 29778 9998 29779
rect 10022 29805 10050 29806
rect 10022 29779 10023 29805
rect 10023 29779 10049 29805
rect 10049 29779 10050 29805
rect 10022 29778 10050 29779
rect 7854 29582 7882 29610
rect 9918 29021 9946 29022
rect 9918 28995 9919 29021
rect 9919 28995 9945 29021
rect 9945 28995 9946 29021
rect 9918 28994 9946 28995
rect 9970 29021 9998 29022
rect 9970 28995 9971 29021
rect 9971 28995 9997 29021
rect 9997 28995 9998 29021
rect 9970 28994 9998 28995
rect 10022 29021 10050 29022
rect 10022 28995 10023 29021
rect 10023 28995 10049 29021
rect 10049 28995 10050 29021
rect 10022 28994 10050 28995
rect 1862 26894 1890 26922
rect 2086 27174 2114 27202
rect 1862 24318 1890 24346
rect 1862 23534 1890 23562
rect 1862 21742 1890 21770
rect 2238 27061 2266 27062
rect 2238 27035 2239 27061
rect 2239 27035 2265 27061
rect 2265 27035 2266 27061
rect 2238 27034 2266 27035
rect 2290 27061 2318 27062
rect 2290 27035 2291 27061
rect 2291 27035 2317 27061
rect 2317 27035 2318 27061
rect 2290 27034 2318 27035
rect 2342 27061 2370 27062
rect 2342 27035 2343 27061
rect 2343 27035 2369 27061
rect 2369 27035 2370 27061
rect 2342 27034 2370 27035
rect 2534 26894 2562 26922
rect 3990 27678 4018 27706
rect 2238 26277 2266 26278
rect 2238 26251 2239 26277
rect 2239 26251 2265 26277
rect 2265 26251 2266 26277
rect 2238 26250 2266 26251
rect 2290 26277 2318 26278
rect 2290 26251 2291 26277
rect 2291 26251 2317 26277
rect 2317 26251 2318 26277
rect 2290 26250 2318 26251
rect 2342 26277 2370 26278
rect 2342 26251 2343 26277
rect 2343 26251 2369 26277
rect 2369 26251 2370 26277
rect 2342 26250 2370 26251
rect 3486 26894 3514 26922
rect 3710 26894 3738 26922
rect 2142 25689 2170 25690
rect 2142 25663 2143 25689
rect 2143 25663 2169 25689
rect 2169 25663 2170 25689
rect 2142 25662 2170 25663
rect 2238 25493 2266 25494
rect 2238 25467 2239 25493
rect 2239 25467 2265 25493
rect 2265 25467 2266 25493
rect 2238 25466 2266 25467
rect 2290 25493 2318 25494
rect 2290 25467 2291 25493
rect 2291 25467 2317 25493
rect 2317 25467 2318 25493
rect 2290 25466 2318 25467
rect 2342 25493 2370 25494
rect 2342 25467 2343 25493
rect 2343 25467 2369 25493
rect 2369 25467 2370 25493
rect 2342 25466 2370 25467
rect 2478 25297 2506 25298
rect 2478 25271 2479 25297
rect 2479 25271 2505 25297
rect 2505 25271 2506 25297
rect 2478 25270 2506 25271
rect 3150 25270 3178 25298
rect 2238 24709 2266 24710
rect 2238 24683 2239 24709
rect 2239 24683 2265 24709
rect 2265 24683 2266 24709
rect 2238 24682 2266 24683
rect 2290 24709 2318 24710
rect 2290 24683 2291 24709
rect 2291 24683 2317 24709
rect 2317 24683 2318 24709
rect 2290 24682 2318 24683
rect 2342 24709 2370 24710
rect 2342 24683 2343 24709
rect 2343 24683 2369 24709
rect 2369 24683 2370 24709
rect 2342 24682 2370 24683
rect 2238 23925 2266 23926
rect 2238 23899 2239 23925
rect 2239 23899 2265 23925
rect 2265 23899 2266 23925
rect 2238 23898 2266 23899
rect 2290 23925 2318 23926
rect 2290 23899 2291 23925
rect 2291 23899 2317 23925
rect 2317 23899 2318 23925
rect 2290 23898 2318 23899
rect 2342 23925 2370 23926
rect 2342 23899 2343 23925
rect 2343 23899 2369 23925
rect 2369 23899 2370 23925
rect 2342 23898 2370 23899
rect 2478 23673 2506 23674
rect 2478 23647 2479 23673
rect 2479 23647 2505 23673
rect 2505 23647 2506 23673
rect 2478 23646 2506 23647
rect 2238 23141 2266 23142
rect 2238 23115 2239 23141
rect 2239 23115 2265 23141
rect 2265 23115 2266 23141
rect 2238 23114 2266 23115
rect 2290 23141 2318 23142
rect 2290 23115 2291 23141
rect 2291 23115 2317 23141
rect 2317 23115 2318 23141
rect 2290 23114 2318 23115
rect 2342 23141 2370 23142
rect 2342 23115 2343 23141
rect 2343 23115 2369 23141
rect 2369 23115 2370 23141
rect 2342 23114 2370 23115
rect 3038 24121 3066 24122
rect 3038 24095 3039 24121
rect 3039 24095 3065 24121
rect 3065 24095 3066 24121
rect 3038 24094 3066 24095
rect 3038 23646 3066 23674
rect 9918 28237 9946 28238
rect 9918 28211 9919 28237
rect 9919 28211 9945 28237
rect 9945 28211 9946 28237
rect 9918 28210 9946 28211
rect 9970 28237 9998 28238
rect 9970 28211 9971 28237
rect 9971 28211 9997 28237
rect 9997 28211 9998 28237
rect 9970 28210 9998 28211
rect 10022 28237 10050 28238
rect 10022 28211 10023 28237
rect 10023 28211 10049 28237
rect 10049 28211 10050 28237
rect 10022 28210 10050 28211
rect 5838 27734 5866 27762
rect 4270 27678 4298 27706
rect 4998 27678 5026 27706
rect 5166 27257 5194 27258
rect 5166 27231 5167 27257
rect 5167 27231 5193 27257
rect 5193 27231 5194 27257
rect 5166 27230 5194 27231
rect 6622 27257 6650 27258
rect 6622 27231 6623 27257
rect 6623 27231 6649 27257
rect 6649 27231 6650 27257
rect 6622 27230 6650 27231
rect 7126 27230 7154 27258
rect 7126 26894 7154 26922
rect 10934 27958 10962 27986
rect 3374 24318 3402 24346
rect 3822 25270 3850 25298
rect 4774 25550 4802 25578
rect 4774 25297 4802 25298
rect 4774 25271 4775 25297
rect 4775 25271 4801 25297
rect 4801 25271 4802 25297
rect 4774 25270 4802 25271
rect 4942 26081 4970 26082
rect 4942 26055 4943 26081
rect 4943 26055 4969 26081
rect 4969 26055 4970 26081
rect 4942 26054 4970 26055
rect 5166 26081 5194 26082
rect 5166 26055 5167 26081
rect 5167 26055 5193 26081
rect 5193 26055 5194 26081
rect 5166 26054 5194 26055
rect 5334 26054 5362 26082
rect 6342 25662 6370 25690
rect 5110 25550 5138 25578
rect 3822 24318 3850 24346
rect 4494 24121 4522 24122
rect 4494 24095 4495 24121
rect 4495 24095 4521 24121
rect 4521 24095 4522 24121
rect 4494 24094 4522 24095
rect 3150 23646 3178 23674
rect 4102 23590 4130 23618
rect 4494 23646 4522 23674
rect 2238 22357 2266 22358
rect 2238 22331 2239 22357
rect 2239 22331 2265 22357
rect 2265 22331 2266 22357
rect 2238 22330 2266 22331
rect 2290 22357 2318 22358
rect 2290 22331 2291 22357
rect 2291 22331 2317 22357
rect 2317 22331 2318 22357
rect 2290 22330 2318 22331
rect 2342 22357 2370 22358
rect 2342 22331 2343 22357
rect 2343 22331 2369 22357
rect 2369 22331 2370 22357
rect 2342 22330 2370 22331
rect 2086 19670 2114 19698
rect 2142 21769 2170 21770
rect 2142 21743 2143 21769
rect 2143 21743 2169 21769
rect 2169 21743 2170 21769
rect 2142 21742 2170 21743
rect 4102 22945 4130 22946
rect 4102 22919 4103 22945
rect 4103 22919 4129 22945
rect 4129 22919 4130 22945
rect 4102 22918 4130 22919
rect 4494 22553 4522 22554
rect 4494 22527 4495 22553
rect 4495 22527 4521 22553
rect 4521 22527 4522 22553
rect 4494 22526 4522 22527
rect 2238 21573 2266 21574
rect 2238 21547 2239 21573
rect 2239 21547 2265 21573
rect 2265 21547 2266 21573
rect 2238 21546 2266 21547
rect 2290 21573 2318 21574
rect 2290 21547 2291 21573
rect 2291 21547 2317 21573
rect 2317 21547 2318 21573
rect 2290 21546 2318 21547
rect 2342 21573 2370 21574
rect 2342 21547 2343 21573
rect 2343 21547 2369 21573
rect 2369 21547 2370 21573
rect 2342 21546 2370 21547
rect 2238 20789 2266 20790
rect 2238 20763 2239 20789
rect 2239 20763 2265 20789
rect 2265 20763 2266 20789
rect 2238 20762 2266 20763
rect 2290 20789 2318 20790
rect 2290 20763 2291 20789
rect 2291 20763 2317 20789
rect 2317 20763 2318 20789
rect 2290 20762 2318 20763
rect 2342 20789 2370 20790
rect 2342 20763 2343 20789
rect 2343 20763 2369 20789
rect 2369 20763 2370 20789
rect 2342 20762 2370 20763
rect 2534 20201 2562 20202
rect 2534 20175 2535 20201
rect 2535 20175 2561 20201
rect 2561 20175 2562 20201
rect 2534 20174 2562 20175
rect 2238 20005 2266 20006
rect 2238 19979 2239 20005
rect 2239 19979 2265 20005
rect 2265 19979 2266 20005
rect 2238 19978 2266 19979
rect 2290 20005 2318 20006
rect 2290 19979 2291 20005
rect 2291 19979 2317 20005
rect 2317 19979 2318 20005
rect 2290 19978 2318 19979
rect 2342 20005 2370 20006
rect 2342 19979 2343 20005
rect 2343 19979 2369 20005
rect 2369 19979 2370 20005
rect 2342 19978 2370 19979
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2142 17849 2170 17850
rect 2142 17823 2143 17849
rect 2143 17823 2169 17849
rect 2169 17823 2170 17849
rect 2142 17822 2170 17823
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 1358 14686 1386 14714
rect 2142 17430 2170 17458
rect 1918 15302 1946 15330
rect 1862 14713 1890 14714
rect 1862 14687 1863 14713
rect 1863 14687 1889 14713
rect 1889 14687 1890 14713
rect 1862 14686 1890 14687
rect 1582 11969 1610 11970
rect 1582 11943 1583 11969
rect 1583 11943 1609 11969
rect 1609 11943 1610 11969
rect 1582 11942 1610 11943
rect 4214 20201 4242 20202
rect 4214 20175 4215 20201
rect 4215 20175 4241 20201
rect 4241 20175 4242 20201
rect 4214 20174 4242 20175
rect 4998 23534 5026 23562
rect 6174 24121 6202 24122
rect 6174 24095 6175 24121
rect 6175 24095 6201 24121
rect 6201 24095 6202 24121
rect 6174 24094 6202 24095
rect 5558 23729 5586 23730
rect 5558 23703 5559 23729
rect 5559 23703 5585 23729
rect 5585 23703 5586 23729
rect 5558 23702 5586 23703
rect 5054 23590 5082 23618
rect 6454 24094 6482 24122
rect 6454 23673 6482 23674
rect 6454 23647 6455 23673
rect 6455 23647 6481 23673
rect 6481 23647 6482 23673
rect 6454 23646 6482 23647
rect 6678 23702 6706 23730
rect 6174 23534 6202 23562
rect 8414 27174 8442 27202
rect 8862 27174 8890 27202
rect 7630 24206 7658 24234
rect 8582 26894 8610 26922
rect 8414 25662 8442 25690
rect 8582 25158 8610 25186
rect 9918 27453 9946 27454
rect 9918 27427 9919 27453
rect 9919 27427 9945 27453
rect 9945 27427 9946 27453
rect 9918 27426 9946 27427
rect 9970 27453 9998 27454
rect 9970 27427 9971 27453
rect 9971 27427 9997 27453
rect 9997 27427 9998 27453
rect 9970 27426 9998 27427
rect 10022 27453 10050 27454
rect 10022 27427 10023 27453
rect 10023 27427 10049 27453
rect 10049 27427 10050 27453
rect 10022 27426 10050 27427
rect 10038 26726 10066 26754
rect 10598 27174 10626 27202
rect 10598 26894 10626 26922
rect 9918 26669 9946 26670
rect 9918 26643 9919 26669
rect 9919 26643 9945 26669
rect 9945 26643 9946 26669
rect 9918 26642 9946 26643
rect 9970 26669 9998 26670
rect 9970 26643 9971 26669
rect 9971 26643 9997 26669
rect 9997 26643 9998 26669
rect 9970 26642 9998 26643
rect 10022 26669 10050 26670
rect 10022 26643 10023 26669
rect 10023 26643 10049 26669
rect 10049 26643 10050 26669
rect 10022 26642 10050 26643
rect 8862 25998 8890 26026
rect 8862 25297 8890 25298
rect 8862 25271 8863 25297
rect 8863 25271 8889 25297
rect 8889 25271 8890 25297
rect 8862 25270 8890 25271
rect 8022 24206 8050 24234
rect 7126 23729 7154 23730
rect 7126 23703 7127 23729
rect 7127 23703 7153 23729
rect 7153 23703 7154 23729
rect 7126 23702 7154 23703
rect 8022 23673 8050 23674
rect 8022 23647 8023 23673
rect 8023 23647 8049 23673
rect 8049 23647 8050 23673
rect 8974 25998 9002 26026
rect 11046 26894 11074 26922
rect 10990 26726 11018 26754
rect 10990 26473 11018 26474
rect 10990 26447 10991 26473
rect 10991 26447 11017 26473
rect 11017 26447 11018 26473
rect 10990 26446 11018 26447
rect 11046 25998 11074 26026
rect 9918 25885 9946 25886
rect 9918 25859 9919 25885
rect 9919 25859 9945 25885
rect 9945 25859 9946 25885
rect 9918 25858 9946 25859
rect 9970 25885 9998 25886
rect 9970 25859 9971 25885
rect 9971 25859 9997 25885
rect 9997 25859 9998 25885
rect 9970 25858 9998 25859
rect 10022 25885 10050 25886
rect 10022 25859 10023 25885
rect 10023 25859 10049 25885
rect 10049 25859 10050 25885
rect 10022 25858 10050 25859
rect 8918 25662 8946 25690
rect 8974 25297 9002 25298
rect 8974 25271 8975 25297
rect 8975 25271 9001 25297
rect 9001 25271 9002 25297
rect 8974 25270 9002 25271
rect 9142 25158 9170 25186
rect 10598 25689 10626 25690
rect 10598 25663 10599 25689
rect 10599 25663 10625 25689
rect 10625 25663 10626 25689
rect 10598 25662 10626 25663
rect 12726 26446 12754 26474
rect 11102 25662 11130 25690
rect 12558 25998 12586 26026
rect 9918 25101 9946 25102
rect 9918 25075 9919 25101
rect 9919 25075 9945 25101
rect 9945 25075 9946 25101
rect 9918 25074 9946 25075
rect 9970 25101 9998 25102
rect 9970 25075 9971 25101
rect 9971 25075 9997 25101
rect 9997 25075 9998 25101
rect 9970 25074 9998 25075
rect 10022 25101 10050 25102
rect 10022 25075 10023 25101
rect 10023 25075 10049 25101
rect 10049 25075 10050 25101
rect 10022 25074 10050 25075
rect 10318 25158 10346 25186
rect 8862 24206 8890 24234
rect 10318 24486 10346 24514
rect 10822 24513 10850 24514
rect 10822 24487 10823 24513
rect 10823 24487 10849 24513
rect 10849 24487 10850 24513
rect 10822 24486 10850 24487
rect 12950 25297 12978 25298
rect 12950 25271 12951 25297
rect 12951 25271 12977 25297
rect 12977 25271 12978 25297
rect 12950 25270 12978 25271
rect 12558 25214 12586 25242
rect 13118 25214 13146 25242
rect 9918 24317 9946 24318
rect 9918 24291 9919 24317
rect 9919 24291 9945 24317
rect 9945 24291 9946 24317
rect 9918 24290 9946 24291
rect 9970 24317 9998 24318
rect 9970 24291 9971 24317
rect 9971 24291 9997 24317
rect 9997 24291 9998 24317
rect 9970 24290 9998 24291
rect 10022 24317 10050 24318
rect 10022 24291 10023 24317
rect 10023 24291 10049 24317
rect 10049 24291 10050 24317
rect 10022 24290 10050 24291
rect 9478 24206 9506 24234
rect 8582 23729 8610 23730
rect 8582 23703 8583 23729
rect 8583 23703 8609 23729
rect 8609 23703 8610 23729
rect 8582 23702 8610 23703
rect 8022 23646 8050 23647
rect 7014 23534 7042 23562
rect 4998 22526 5026 22554
rect 2478 17457 2506 17458
rect 2478 17431 2479 17457
rect 2479 17431 2505 17457
rect 2505 17431 2506 17457
rect 2478 17430 2506 17431
rect 3038 17430 3066 17458
rect 3598 17849 3626 17850
rect 3598 17823 3599 17849
rect 3599 17823 3625 17849
rect 3625 17823 3626 17849
rect 3598 17822 3626 17823
rect 4158 17710 4186 17738
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 4102 16673 4130 16674
rect 4102 16647 4103 16673
rect 4103 16647 4129 16673
rect 4129 16647 4130 16673
rect 4102 16646 4130 16647
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 7518 23534 7546 23562
rect 10038 24206 10066 24234
rect 11102 24374 11130 24402
rect 10598 24121 10626 24122
rect 10598 24095 10599 24121
rect 10599 24095 10625 24121
rect 10625 24095 10626 24121
rect 10598 24094 10626 24095
rect 11102 24094 11130 24122
rect 12278 24486 12306 24514
rect 11494 23702 11522 23730
rect 11718 23729 11746 23730
rect 11718 23703 11719 23729
rect 11719 23703 11745 23729
rect 11745 23703 11746 23729
rect 11718 23702 11746 23703
rect 13510 25270 13538 25298
rect 12558 24374 12586 24402
rect 13118 24374 13146 24402
rect 13342 24318 13370 24346
rect 13510 24206 13538 24234
rect 10990 23590 11018 23618
rect 7574 22553 7602 22554
rect 7574 22527 7575 22553
rect 7575 22527 7601 22553
rect 7601 22527 7602 22553
rect 7574 22526 7602 22527
rect 8134 22526 8162 22554
rect 7294 21854 7322 21882
rect 5838 18494 5866 18522
rect 4382 17457 4410 17458
rect 4382 17431 4383 17457
rect 4383 17431 4409 17457
rect 4409 17431 4410 17457
rect 4382 17430 4410 17431
rect 2478 15918 2506 15946
rect 3038 15918 3066 15946
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 6454 17654 6482 17682
rect 7294 18494 7322 18522
rect 8134 21854 8162 21882
rect 9030 21742 9058 21770
rect 9310 23534 9338 23562
rect 9918 23533 9946 23534
rect 9918 23507 9919 23533
rect 9919 23507 9945 23533
rect 9945 23507 9946 23533
rect 9918 23506 9946 23507
rect 9970 23533 9998 23534
rect 9970 23507 9971 23533
rect 9971 23507 9997 23533
rect 9997 23507 9998 23533
rect 9970 23506 9998 23507
rect 10022 23533 10050 23534
rect 10022 23507 10023 23533
rect 10023 23507 10049 23533
rect 10049 23507 10050 23533
rect 10022 23506 10050 23507
rect 9918 22749 9946 22750
rect 9918 22723 9919 22749
rect 9919 22723 9945 22749
rect 9945 22723 9946 22749
rect 9918 22722 9946 22723
rect 9970 22749 9998 22750
rect 9970 22723 9971 22749
rect 9971 22723 9997 22749
rect 9997 22723 9998 22749
rect 9970 22722 9998 22723
rect 10022 22749 10050 22750
rect 10022 22723 10023 22749
rect 10023 22723 10049 22749
rect 10049 22723 10050 22749
rect 10022 22722 10050 22723
rect 11270 23590 11298 23618
rect 9918 21965 9946 21966
rect 9918 21939 9919 21965
rect 9919 21939 9945 21965
rect 9945 21939 9946 21965
rect 9918 21938 9946 21939
rect 9970 21965 9998 21966
rect 9970 21939 9971 21965
rect 9971 21939 9997 21965
rect 9997 21939 9998 21965
rect 9970 21938 9998 21939
rect 10022 21965 10050 21966
rect 10022 21939 10023 21965
rect 10023 21939 10049 21965
rect 10049 21939 10050 21965
rect 10022 21938 10050 21939
rect 9310 21769 9338 21770
rect 9310 21743 9311 21769
rect 9311 21743 9337 21769
rect 9337 21743 9338 21769
rect 9310 21742 9338 21743
rect 9534 21769 9562 21770
rect 9534 21743 9535 21769
rect 9535 21743 9561 21769
rect 9561 21743 9562 21769
rect 9534 21742 9562 21743
rect 9918 21181 9946 21182
rect 9918 21155 9919 21181
rect 9919 21155 9945 21181
rect 9945 21155 9946 21181
rect 9918 21154 9946 21155
rect 9970 21181 9998 21182
rect 9970 21155 9971 21181
rect 9971 21155 9997 21181
rect 9997 21155 9998 21181
rect 9970 21154 9998 21155
rect 10022 21181 10050 21182
rect 10022 21155 10023 21181
rect 10023 21155 10049 21181
rect 10049 21155 10050 21181
rect 10022 21154 10050 21155
rect 7014 17654 7042 17682
rect 5278 16673 5306 16674
rect 5278 16647 5279 16673
rect 5279 16647 5305 16673
rect 5305 16647 5306 16673
rect 5278 16646 5306 16647
rect 5558 16646 5586 16674
rect 4550 15918 4578 15946
rect 5558 15889 5586 15890
rect 5558 15863 5559 15889
rect 5559 15863 5585 15889
rect 5585 15863 5586 15889
rect 5558 15862 5586 15863
rect 5838 15862 5866 15890
rect 2422 15134 2450 15162
rect 3374 14686 3402 14714
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 1918 11830 1946 11858
rect 1582 10094 1610 10122
rect 1694 10934 1722 10962
rect 1022 6566 1050 6594
rect 1582 6481 1610 6482
rect 1582 6455 1583 6481
rect 1583 6455 1609 6481
rect 1609 6455 1610 6481
rect 1582 6454 1610 6455
rect 1022 4494 1050 4522
rect 1190 6089 1218 6090
rect 1190 6063 1191 6089
rect 1191 6063 1217 6089
rect 1217 6063 1218 6089
rect 1190 6062 1218 6063
rect 1862 10094 1890 10122
rect 1862 9982 1890 10010
rect 2310 13929 2338 13930
rect 2310 13903 2311 13929
rect 2311 13903 2337 13929
rect 2337 13903 2338 13929
rect 2310 13902 2338 13903
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2534 13929 2562 13930
rect 2534 13903 2535 13929
rect 2535 13903 2561 13929
rect 2561 13903 2562 13929
rect 2534 13902 2562 13903
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 3822 14238 3850 14266
rect 3374 12558 3402 12586
rect 2534 12361 2562 12362
rect 2534 12335 2535 12361
rect 2535 12335 2561 12361
rect 2561 12335 2562 12361
rect 2534 12334 2562 12335
rect 4494 15134 4522 15162
rect 5950 15918 5978 15946
rect 6230 15918 6258 15946
rect 6734 16254 6762 16282
rect 7014 16281 7042 16282
rect 7014 16255 7015 16281
rect 7015 16255 7041 16281
rect 7041 16255 7042 16281
rect 7014 16254 7042 16255
rect 8134 17038 8162 17066
rect 6454 15918 6482 15946
rect 5838 15470 5866 15498
rect 6118 15497 6146 15498
rect 6118 15471 6119 15497
rect 6119 15471 6145 15497
rect 6145 15471 6146 15497
rect 6118 15470 6146 15471
rect 6510 15134 6538 15162
rect 4494 13145 4522 13146
rect 4494 13119 4495 13145
rect 4495 13119 4521 13145
rect 4521 13119 4522 13145
rect 4494 13118 4522 13119
rect 6846 15470 6874 15498
rect 5278 14238 5306 14266
rect 9030 18185 9058 18186
rect 9030 18159 9031 18185
rect 9031 18159 9057 18185
rect 9057 18159 9058 18185
rect 9030 18158 9058 18159
rect 9918 20397 9946 20398
rect 9918 20371 9919 20397
rect 9919 20371 9945 20397
rect 9945 20371 9946 20397
rect 9918 20370 9946 20371
rect 9970 20397 9998 20398
rect 9970 20371 9971 20397
rect 9971 20371 9997 20397
rect 9997 20371 9998 20397
rect 9970 20370 9998 20371
rect 10022 20397 10050 20398
rect 10022 20371 10023 20397
rect 10023 20371 10049 20397
rect 10049 20371 10050 20397
rect 10022 20370 10050 20371
rect 9918 19613 9946 19614
rect 9918 19587 9919 19613
rect 9919 19587 9945 19613
rect 9945 19587 9946 19613
rect 9918 19586 9946 19587
rect 9970 19613 9998 19614
rect 9970 19587 9971 19613
rect 9971 19587 9997 19613
rect 9997 19587 9998 19613
rect 9970 19586 9998 19587
rect 10022 19613 10050 19614
rect 10022 19587 10023 19613
rect 10023 19587 10049 19613
rect 10049 19587 10050 19613
rect 10022 19586 10050 19587
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9142 17065 9170 17066
rect 9142 17039 9143 17065
rect 9143 17039 9169 17065
rect 9169 17039 9170 17065
rect 9142 17038 9170 17039
rect 5558 14238 5586 14266
rect 6902 15134 6930 15162
rect 8302 16254 8330 16282
rect 9814 18158 9842 18186
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 10038 17822 10066 17850
rect 13454 23729 13482 23730
rect 13454 23703 13455 23729
rect 13455 23703 13481 23729
rect 13481 23703 13482 23729
rect 13454 23702 13482 23703
rect 12278 23310 12306 23338
rect 12838 23337 12866 23338
rect 12838 23311 12839 23337
rect 12839 23311 12865 23337
rect 12865 23311 12866 23337
rect 12838 23310 12866 23311
rect 13230 22105 13258 22106
rect 13230 22079 13231 22105
rect 13231 22079 13257 22105
rect 13257 22079 13258 22105
rect 13230 22078 13258 22079
rect 12838 21769 12866 21770
rect 12838 21743 12839 21769
rect 12839 21743 12865 21769
rect 12865 21743 12866 21769
rect 12838 21742 12866 21743
rect 13118 21742 13146 21770
rect 12950 20230 12978 20258
rect 10934 18214 10962 18242
rect 13510 21769 13538 21770
rect 13510 21743 13511 21769
rect 13511 21743 13537 21769
rect 13537 21743 13538 21769
rect 13510 21742 13538 21743
rect 13454 20537 13482 20538
rect 13454 20511 13455 20537
rect 13455 20511 13481 20537
rect 13481 20511 13482 20537
rect 13454 20510 13482 20511
rect 13118 19390 13146 19418
rect 12838 18494 12866 18522
rect 12278 18438 12306 18466
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 12278 18241 12306 18242
rect 12278 18215 12279 18241
rect 12279 18215 12305 18241
rect 12305 18215 12306 18241
rect 12278 18214 12306 18215
rect 11270 17849 11298 17850
rect 11270 17823 11271 17849
rect 11271 17823 11297 17849
rect 11297 17823 11298 17849
rect 11270 17822 11298 17823
rect 14014 22078 14042 22106
rect 14014 21742 14042 21770
rect 14014 20510 14042 20538
rect 14014 20201 14042 20202
rect 14014 20175 14015 20201
rect 14015 20175 14041 20201
rect 14041 20175 14042 20201
rect 14014 20174 14042 20175
rect 13454 19446 13482 19474
rect 14014 19473 14042 19474
rect 14014 19447 14015 19473
rect 14015 19447 14041 19473
rect 14041 19447 14042 19473
rect 14014 19446 14042 19447
rect 10318 17065 10346 17066
rect 10318 17039 10319 17065
rect 10319 17039 10345 17065
rect 10345 17039 10346 17065
rect 10318 17038 10346 17039
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 8470 15497 8498 15498
rect 8470 15471 8471 15497
rect 8471 15471 8497 15497
rect 8497 15471 8498 15497
rect 8470 15470 8498 15471
rect 9030 15470 9058 15498
rect 4998 13118 5026 13146
rect 4998 12614 5026 12642
rect 7014 13929 7042 13930
rect 7014 13903 7015 13929
rect 7015 13903 7041 13929
rect 7041 13903 7042 13929
rect 7014 13902 7042 13903
rect 5502 13454 5530 13482
rect 3822 12558 3850 12586
rect 4494 12558 4522 12586
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11942 2170 11970
rect 3318 11969 3346 11970
rect 3318 11943 3319 11969
rect 3319 11943 3345 11969
rect 3345 11943 3346 11969
rect 3318 11942 3346 11943
rect 3598 11942 3626 11970
rect 3766 12361 3794 12362
rect 3766 12335 3767 12361
rect 3767 12335 3793 12361
rect 3793 12335 3794 12361
rect 3766 12334 3794 12335
rect 3990 12361 4018 12362
rect 3990 12335 3991 12361
rect 3991 12335 4017 12361
rect 4017 12335 4018 12361
rect 3990 12334 4018 12335
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 2478 11129 2506 11130
rect 2478 11103 2479 11129
rect 2479 11103 2505 11129
rect 2505 11103 2506 11129
rect 2478 11102 2506 11103
rect 2870 11102 2898 11130
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 2534 8441 2562 8442
rect 2534 8415 2535 8441
rect 2535 8415 2561 8441
rect 2561 8415 2562 8441
rect 2534 8414 2562 8415
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 2142 7574 2170 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 1918 6454 1946 6482
rect 1694 6062 1722 6090
rect 5670 12614 5698 12642
rect 6062 12614 6090 12642
rect 6958 13454 6986 13482
rect 8414 13902 8442 13930
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 8862 13929 8890 13930
rect 8862 13903 8863 13929
rect 8863 13903 8889 13929
rect 8889 13903 8890 13929
rect 8862 13902 8890 13903
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 8862 12361 8890 12362
rect 8862 12335 8863 12361
rect 8863 12335 8889 12361
rect 8889 12335 8890 12361
rect 8862 12334 8890 12335
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 10598 12361 10626 12362
rect 10598 12335 10599 12361
rect 10599 12335 10625 12361
rect 10625 12335 10626 12361
rect 10598 12334 10626 12335
rect 8190 11774 8218 11802
rect 4270 10318 4298 10346
rect 4606 10345 4634 10346
rect 4606 10319 4607 10345
rect 4607 10319 4633 10345
rect 4633 10319 4634 10345
rect 4606 10318 4634 10319
rect 5838 10345 5866 10346
rect 5838 10319 5839 10345
rect 5839 10319 5865 10345
rect 5865 10319 5866 10345
rect 5838 10318 5866 10319
rect 9422 11774 9450 11802
rect 7294 11158 7322 11186
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 3766 8441 3794 8442
rect 3766 8415 3767 8441
rect 3767 8415 3793 8441
rect 3793 8415 3794 8441
rect 3766 8414 3794 8415
rect 3598 7518 3626 7546
rect 3598 7265 3626 7266
rect 3598 7239 3599 7265
rect 3599 7239 3625 7265
rect 3625 7239 3626 7265
rect 3598 7238 3626 7239
rect 8414 11185 8442 11186
rect 8414 11159 8415 11185
rect 8415 11159 8441 11185
rect 8441 11159 8442 11185
rect 8414 11158 8442 11159
rect 8862 11158 8890 11186
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 3822 7238 3850 7266
rect 4494 8441 4522 8442
rect 4494 8415 4495 8441
rect 4495 8415 4521 8441
rect 4521 8415 4522 8441
rect 4494 8414 4522 8415
rect 4494 7574 4522 7602
rect 6454 8358 6482 8386
rect 6678 8358 6706 8386
rect 4998 7574 5026 7602
rect 5838 7574 5866 7602
rect 4886 7265 4914 7266
rect 4886 7239 4887 7265
rect 4887 7239 4913 7265
rect 4913 7239 4914 7265
rect 4886 7238 4914 7239
rect 7238 7265 7266 7266
rect 7238 7239 7239 7265
rect 7239 7239 7265 7265
rect 7265 7239 7266 7265
rect 7238 7238 7266 7239
rect 8134 8358 8162 8386
rect 8134 8049 8162 8050
rect 8134 8023 8135 8049
rect 8135 8023 8161 8049
rect 8161 8023 8162 8049
rect 8134 8022 8162 8023
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 11494 11774 11522 11802
rect 12558 11185 12586 11186
rect 12558 11159 12559 11185
rect 12559 11159 12585 11185
rect 12585 11159 12586 11185
rect 12558 11158 12586 11159
rect 13118 12361 13146 12362
rect 13118 12335 13119 12361
rect 13119 12335 13145 12361
rect 13145 12335 13146 12361
rect 13118 12334 13146 12335
rect 12726 11774 12754 11802
rect 12950 11774 12978 11802
rect 13510 12278 13538 12306
rect 13286 11774 13314 11802
rect 13118 11158 13146 11186
rect 9814 10009 9842 10010
rect 9814 9983 9815 10009
rect 9815 9983 9841 10009
rect 9841 9983 9842 10009
rect 9814 9982 9842 9983
rect 10038 9982 10066 10010
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10990 10009 11018 10010
rect 10990 9983 10991 10009
rect 10991 9983 11017 10009
rect 11017 9983 11018 10009
rect 10990 9982 11018 9983
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9422 8049 9450 8050
rect 9422 8023 9423 8049
rect 9423 8023 9449 8049
rect 9449 8023 9450 8049
rect 9422 8022 9450 8023
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9142 7657 9170 7658
rect 9142 7631 9143 7657
rect 9143 7631 9169 7657
rect 9169 7631 9170 7657
rect 9142 7630 9170 7631
rect 8694 7265 8722 7266
rect 8694 7239 8695 7265
rect 8695 7239 8721 7265
rect 8721 7239 8722 7265
rect 8694 7238 8722 7239
rect 9590 7574 9618 7602
rect 10318 7657 10346 7658
rect 10318 7631 10319 7657
rect 10319 7631 10345 7657
rect 10345 7631 10346 7657
rect 10318 7630 10346 7631
rect 14518 25214 14546 25242
rect 14518 23478 14546 23506
rect 14574 24374 14602 24402
rect 15134 24318 15162 24346
rect 15134 24206 15162 24234
rect 15470 23729 15498 23730
rect 15470 23703 15471 23729
rect 15471 23703 15497 23729
rect 15497 23703 15498 23729
rect 15470 23702 15498 23703
rect 16814 23702 16842 23730
rect 15078 23478 15106 23506
rect 15078 22918 15106 22946
rect 16254 22945 16282 22946
rect 16254 22919 16255 22945
rect 16255 22919 16281 22945
rect 16281 22919 16282 22945
rect 16254 22918 16282 22919
rect 16254 22526 16282 22554
rect 16702 22526 16730 22554
rect 16814 22553 16842 22554
rect 16814 22527 16815 22553
rect 16815 22527 16841 22553
rect 16841 22527 16842 22553
rect 16814 22526 16842 22527
rect 16926 22526 16954 22554
rect 14798 21070 14826 21098
rect 14350 21014 14378 21042
rect 14574 21014 14602 21042
rect 14294 20230 14322 20258
rect 16814 21742 16842 21770
rect 17094 21769 17122 21770
rect 17094 21743 17095 21769
rect 17095 21743 17121 21769
rect 17121 21743 17122 21769
rect 17094 21742 17122 21743
rect 16254 21014 16282 21042
rect 14294 19417 14322 19418
rect 14294 19391 14295 19417
rect 14295 19391 14321 19417
rect 14321 19391 14322 19417
rect 14294 19390 14322 19391
rect 14798 19390 14826 19418
rect 15918 20958 15946 20986
rect 15358 20201 15386 20202
rect 15358 20175 15359 20201
rect 15359 20175 15385 20201
rect 15385 20175 15386 20201
rect 15358 20174 15386 20175
rect 16534 21070 16562 21098
rect 16758 21014 16786 21042
rect 15470 19473 15498 19474
rect 15470 19447 15471 19473
rect 15471 19447 15497 19473
rect 15497 19447 15498 19473
rect 15470 19446 15498 19447
rect 15918 18185 15946 18186
rect 15918 18159 15919 18185
rect 15919 18159 15945 18185
rect 15945 18159 15946 18185
rect 15918 18158 15946 18159
rect 15918 17457 15946 17458
rect 15918 17431 15919 17457
rect 15919 17431 15945 17457
rect 15945 17431 15946 17457
rect 15918 17430 15946 17431
rect 14182 11158 14210 11186
rect 14574 12361 14602 12362
rect 14574 12335 14575 12361
rect 14575 12335 14601 12361
rect 14601 12335 14602 12361
rect 14574 12334 14602 12335
rect 11382 9982 11410 10010
rect 12278 9617 12306 9618
rect 12278 9591 12279 9617
rect 12279 9591 12305 9617
rect 12305 9591 12306 9617
rect 12278 9590 12306 9591
rect 11102 9254 11130 9282
rect 11494 9310 11522 9338
rect 11718 9310 11746 9338
rect 12558 9590 12586 9618
rect 12838 10009 12866 10010
rect 12838 9983 12839 10009
rect 12839 9983 12865 10009
rect 12865 9983 12866 10009
rect 12838 9982 12866 9983
rect 12278 9254 12306 9282
rect 13118 9982 13146 10010
rect 16814 17457 16842 17458
rect 16814 17431 16815 17457
rect 16815 17431 16841 17457
rect 16841 17431 16842 17457
rect 16814 17430 16842 17431
rect 16814 16254 16842 16282
rect 16982 16281 17010 16282
rect 16982 16255 16983 16281
rect 16983 16255 17009 16281
rect 17009 16255 17010 16281
rect 16982 16254 17010 16255
rect 16926 15806 16954 15834
rect 16814 15470 16842 15498
rect 15470 13537 15498 13538
rect 15470 13511 15471 13537
rect 15471 13511 15497 13537
rect 15497 13511 15498 13537
rect 15470 13510 15498 13511
rect 16982 13118 17010 13146
rect 17094 15497 17122 15498
rect 17094 15471 17095 15497
rect 17095 15471 17121 15497
rect 17121 15471 17122 15497
rect 17094 15470 17122 15471
rect 17094 13454 17122 13482
rect 15134 12278 15162 12306
rect 14798 11998 14826 12026
rect 16254 11998 16282 12026
rect 15470 11942 15498 11970
rect 15918 11969 15946 11970
rect 15918 11943 15919 11969
rect 15919 11943 15945 11969
rect 15945 11943 15946 11969
rect 15918 11942 15946 11943
rect 13454 10038 13482 10066
rect 14014 10065 14042 10066
rect 14014 10039 14015 10065
rect 14015 10039 14041 10065
rect 14041 10039 14042 10065
rect 14014 10038 14042 10039
rect 14294 10009 14322 10010
rect 14294 9983 14295 10009
rect 14295 9983 14321 10009
rect 14321 9983 14322 10009
rect 14294 9982 14322 9983
rect 17094 11830 17122 11858
rect 17094 11577 17122 11578
rect 17094 11551 17095 11577
rect 17095 11551 17121 11577
rect 17121 11551 17122 11577
rect 17094 11550 17122 11551
rect 14574 9982 14602 10010
rect 15358 10065 15386 10066
rect 15358 10039 15359 10065
rect 15359 10039 15385 10065
rect 15385 10039 15386 10065
rect 15358 10038 15386 10039
rect 12838 9254 12866 9282
rect 13398 9310 13426 9338
rect 16814 11185 16842 11186
rect 16814 11159 16815 11185
rect 16815 11159 16841 11185
rect 16841 11159 16842 11185
rect 16814 11158 16842 11159
rect 10038 7574 10066 7602
rect 11494 7574 11522 7602
rect 12558 7574 12586 7602
rect 13118 7574 13146 7602
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 2478 6481 2506 6482
rect 2478 6455 2479 6481
rect 2479 6455 2505 6481
rect 2505 6455 2506 6481
rect 2478 6454 2506 6455
rect 2870 6454 2898 6482
rect 2030 5278 2058 5306
rect 2086 6145 2114 6146
rect 2086 6119 2087 6145
rect 2087 6119 2113 6145
rect 2113 6119 2114 6145
rect 2086 6118 2114 6119
rect 4158 6398 4186 6426
rect 2814 6118 2842 6146
rect 2534 6089 2562 6090
rect 2534 6063 2535 6089
rect 2535 6063 2561 6089
rect 2561 6063 2562 6089
rect 2534 6062 2562 6063
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 3038 6118 3066 6146
rect 2870 6062 2898 6090
rect 2814 5305 2842 5306
rect 2814 5279 2815 5305
rect 2815 5279 2841 5305
rect 2841 5279 2842 5305
rect 2814 5278 2842 5279
rect 3038 5305 3066 5306
rect 3038 5279 3039 5305
rect 3039 5279 3065 5305
rect 3065 5279 3066 5305
rect 3038 5278 3066 5279
rect 6454 6481 6482 6482
rect 6454 6455 6455 6481
rect 6455 6455 6481 6481
rect 6481 6455 6482 6481
rect 6454 6454 6482 6455
rect 7014 6454 7042 6482
rect 5278 6425 5306 6426
rect 5278 6399 5279 6425
rect 5279 6399 5305 6425
rect 5305 6399 5306 6425
rect 5278 6398 5306 6399
rect 5838 6398 5866 6426
rect 5838 6089 5866 6090
rect 5838 6063 5839 6089
rect 5839 6063 5865 6089
rect 5865 6063 5866 6089
rect 5838 6062 5866 6063
rect 4998 5670 5026 5698
rect 5558 5697 5586 5698
rect 5558 5671 5559 5697
rect 5559 5671 5585 5697
rect 5585 5671 5586 5697
rect 5558 5670 5586 5671
rect 3318 5278 3346 5306
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2086 4886 2114 4914
rect 2534 4521 2562 4522
rect 2534 4495 2535 4521
rect 2535 4495 2561 4521
rect 2561 4495 2562 4521
rect 2534 4494 2562 4495
rect 2870 4494 2898 4522
rect 3318 4913 3346 4914
rect 3318 4887 3319 4913
rect 3319 4887 3345 4913
rect 3345 4887 3346 4913
rect 3318 4886 3346 4887
rect 3542 4913 3570 4914
rect 3542 4887 3543 4913
rect 3543 4887 3569 4913
rect 3569 4887 3570 4913
rect 3542 4886 3570 4887
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 6118 5670 6146 5698
rect 7574 6089 7602 6090
rect 7574 6063 7575 6089
rect 7575 6063 7601 6089
rect 7601 6063 7602 6089
rect 7574 6062 7602 6063
rect 7798 6062 7826 6090
rect 8470 5894 8498 5922
rect 8974 5894 9002 5922
rect 9534 6481 9562 6482
rect 9534 6455 9535 6481
rect 9535 6455 9561 6481
rect 9561 6455 9562 6481
rect 9534 6454 9562 6455
rect 9534 5894 9562 5922
rect 7014 5110 7042 5138
rect 7518 5110 7546 5138
rect 6510 5054 6538 5082
rect 6118 4382 6146 4410
rect 6454 4129 6482 4130
rect 6454 4103 6455 4129
rect 6455 4103 6481 4129
rect 6481 4103 6482 4129
rect 6454 4102 6482 4103
rect 7518 4382 7546 4410
rect 8078 5110 8106 5138
rect 7742 5054 7770 5082
rect 9478 5110 9506 5138
rect 8246 5054 8274 5082
rect 7798 4382 7826 4410
rect 7014 4102 7042 4130
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 7014 3737 7042 3738
rect 7014 3711 7015 3737
rect 7015 3711 7041 3737
rect 7041 3711 7042 3737
rect 7014 3710 7042 3711
rect 7518 3737 7546 3738
rect 7518 3711 7519 3737
rect 7519 3711 7545 3737
rect 7545 3711 7546 3737
rect 7518 3710 7546 3711
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 3766 2534 3794 2562
rect 910 2198 938 2226
rect 5278 2561 5306 2562
rect 5278 2535 5279 2561
rect 5279 2535 5305 2561
rect 5305 2535 5306 2561
rect 5278 2534 5306 2535
rect 5838 2534 5866 2562
rect 6230 2561 6258 2562
rect 6230 2535 6231 2561
rect 6231 2535 6257 2561
rect 6257 2535 6258 2561
rect 6230 2534 6258 2535
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 2086 1750 2114 1778
rect 2870 1777 2898 1778
rect 2870 1751 2871 1777
rect 2871 1751 2897 1777
rect 2897 1751 2898 1777
rect 2870 1750 2898 1751
rect 3822 1721 3850 1722
rect 3822 1695 3823 1721
rect 3823 1695 3849 1721
rect 3849 1695 3850 1721
rect 3822 1694 3850 1695
rect 7798 4129 7826 4130
rect 7798 4103 7799 4129
rect 7799 4103 7825 4129
rect 7825 4103 7826 4129
rect 7798 4102 7826 4103
rect 9814 6454 9842 6482
rect 10430 6425 10458 6426
rect 10430 6399 10431 6425
rect 10431 6399 10457 6425
rect 10457 6399 10458 6425
rect 10430 6398 10458 6399
rect 10878 6398 10906 6426
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9814 6118 9842 6146
rect 10878 6089 10906 6090
rect 10878 6063 10879 6089
rect 10879 6063 10905 6089
rect 10905 6063 10906 6089
rect 10878 6062 10906 6063
rect 11550 6118 11578 6146
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 10038 4438 10066 4466
rect 10430 4494 10458 4522
rect 8470 4158 8498 4186
rect 7742 2982 7770 3010
rect 7798 3374 7826 3402
rect 7574 2953 7602 2954
rect 7574 2927 7575 2953
rect 7575 2927 7601 2953
rect 7601 2927 7602 2953
rect 7574 2926 7602 2927
rect 7014 2534 7042 2562
rect 9254 4102 9282 4130
rect 8246 3374 8274 3402
rect 8470 3374 8498 3402
rect 8078 2926 8106 2954
rect 8078 2590 8106 2618
rect 8470 3009 8498 3010
rect 8470 2983 8471 3009
rect 8471 2983 8497 3009
rect 8497 2983 8498 3009
rect 8470 2982 8498 2983
rect 8470 2534 8498 2562
rect 8974 2561 9002 2562
rect 8974 2535 8975 2561
rect 8975 2535 9001 2561
rect 9001 2535 9002 2561
rect 8974 2534 9002 2535
rect 10374 4129 10402 4130
rect 10374 4103 10375 4129
rect 10375 4103 10401 4129
rect 10401 4103 10402 4129
rect 10374 4102 10402 4103
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9534 3345 9562 3346
rect 9534 3319 9535 3345
rect 9535 3319 9561 3345
rect 9561 3319 9562 3345
rect 9534 3318 9562 3319
rect 10374 3710 10402 3738
rect 9814 3318 9842 3346
rect 11774 4886 11802 4914
rect 12446 6454 12474 6482
rect 12950 6481 12978 6482
rect 12950 6455 12951 6481
rect 12951 6455 12977 6481
rect 12977 6455 12978 6481
rect 12950 6454 12978 6455
rect 12446 6089 12474 6090
rect 12446 6063 12447 6089
rect 12447 6063 12473 6089
rect 12473 6063 12474 6089
rect 12446 6062 12474 6063
rect 12054 4913 12082 4914
rect 12054 4887 12055 4913
rect 12055 4887 12081 4913
rect 12081 4887 12082 4913
rect 12054 4886 12082 4887
rect 12838 4886 12866 4914
rect 10878 4521 10906 4522
rect 10878 4495 10879 4521
rect 10879 4495 10905 4521
rect 10905 4495 10906 4521
rect 10878 4494 10906 4495
rect 11270 4438 11298 4466
rect 10878 3737 10906 3738
rect 10878 3711 10879 3737
rect 10879 3711 10905 3737
rect 10905 3711 10906 3737
rect 10878 3710 10906 3711
rect 12390 4521 12418 4522
rect 12390 4495 12391 4521
rect 12391 4495 12417 4521
rect 12417 4495 12418 4521
rect 12390 4494 12418 4495
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9814 2926 9842 2954
rect 10038 2953 10066 2954
rect 10038 2927 10039 2953
rect 10039 2927 10065 2953
rect 10065 2927 10066 2953
rect 10038 2926 10066 2927
rect 9254 2142 9282 2170
rect 9422 2590 9450 2618
rect 10430 2561 10458 2562
rect 10430 2535 10431 2561
rect 10431 2535 10457 2561
rect 10457 2535 10458 2561
rect 10430 2534 10458 2535
rect 10766 2534 10794 2562
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9814 2169 9842 2170
rect 9814 2143 9815 2169
rect 9815 2143 9841 2169
rect 9841 2143 9842 2169
rect 9814 2142 9842 2143
rect 11550 2953 11578 2954
rect 11550 2927 11551 2953
rect 11551 2927 11577 2953
rect 11577 2927 11578 2953
rect 11550 2926 11578 2927
rect 11550 2534 11578 2562
rect 12334 4158 12362 4186
rect 12334 3710 12362 3738
rect 11102 2030 11130 2058
rect 9422 1777 9450 1778
rect 9422 1751 9423 1777
rect 9423 1751 9449 1777
rect 9449 1751 9450 1777
rect 9422 1750 9450 1751
rect 7574 1694 7602 1722
rect 9590 1694 9618 1722
rect 9814 1694 9842 1722
rect 10374 1750 10402 1778
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 13118 4886 13146 4914
rect 13454 6454 13482 6482
rect 14014 6454 14042 6482
rect 14238 6481 14266 6482
rect 14238 6455 14239 6481
rect 14239 6455 14265 6481
rect 14265 6455 14266 6481
rect 14238 6454 14266 6455
rect 13398 4913 13426 4914
rect 13398 4887 13399 4913
rect 13399 4887 13425 4913
rect 13425 4887 13426 4913
rect 13398 4886 13426 4887
rect 12950 4158 12978 4186
rect 13958 4521 13986 4522
rect 13958 4495 13959 4521
rect 13959 4495 13985 4521
rect 13985 4495 13986 4521
rect 13958 4494 13986 4495
rect 14238 4998 14266 5026
rect 14238 4494 14266 4522
rect 14126 4158 14154 4186
rect 12446 2169 12474 2170
rect 12446 2143 12447 2169
rect 12447 2143 12473 2169
rect 12473 2143 12474 2169
rect 12446 2142 12474 2143
rect 12894 2142 12922 2170
rect 13118 3318 13146 3346
rect 13398 3345 13426 3346
rect 13398 3319 13399 3345
rect 13399 3319 13425 3345
rect 13425 3319 13426 3345
rect 13398 3318 13426 3319
rect 14574 4886 14602 4914
rect 14798 7574 14826 7602
rect 15470 7966 15498 7994
rect 16534 8049 16562 8050
rect 16534 8023 16535 8049
rect 16535 8023 16561 8049
rect 16561 8023 16562 8049
rect 16534 8022 16562 8023
rect 16534 7574 16562 7602
rect 15358 6481 15386 6482
rect 15358 6455 15359 6481
rect 15359 6455 15385 6481
rect 15385 6455 15386 6481
rect 15358 6454 15386 6455
rect 16926 9534 16954 9562
rect 17598 33333 17626 33334
rect 17598 33307 17599 33333
rect 17599 33307 17625 33333
rect 17625 33307 17626 33333
rect 17598 33306 17626 33307
rect 17650 33333 17678 33334
rect 17650 33307 17651 33333
rect 17651 33307 17677 33333
rect 17677 33307 17678 33333
rect 17650 33306 17678 33307
rect 17702 33333 17730 33334
rect 17702 33307 17703 33333
rect 17703 33307 17729 33333
rect 17729 33307 17730 33333
rect 17702 33306 17730 33307
rect 17598 32549 17626 32550
rect 17598 32523 17599 32549
rect 17599 32523 17625 32549
rect 17625 32523 17626 32549
rect 17598 32522 17626 32523
rect 17650 32549 17678 32550
rect 17650 32523 17651 32549
rect 17651 32523 17677 32549
rect 17677 32523 17678 32549
rect 17650 32522 17678 32523
rect 17702 32549 17730 32550
rect 17702 32523 17703 32549
rect 17703 32523 17729 32549
rect 17729 32523 17730 32549
rect 17702 32522 17730 32523
rect 17598 31765 17626 31766
rect 17598 31739 17599 31765
rect 17599 31739 17625 31765
rect 17625 31739 17626 31765
rect 17598 31738 17626 31739
rect 17650 31765 17678 31766
rect 17650 31739 17651 31765
rect 17651 31739 17677 31765
rect 17677 31739 17678 31765
rect 17650 31738 17678 31739
rect 17702 31765 17730 31766
rect 17702 31739 17703 31765
rect 17703 31739 17729 31765
rect 17729 31739 17730 31765
rect 17702 31738 17730 31739
rect 17598 30981 17626 30982
rect 17598 30955 17599 30981
rect 17599 30955 17625 30981
rect 17625 30955 17626 30981
rect 17598 30954 17626 30955
rect 17650 30981 17678 30982
rect 17650 30955 17651 30981
rect 17651 30955 17677 30981
rect 17677 30955 17678 30981
rect 17650 30954 17678 30955
rect 17702 30981 17730 30982
rect 17702 30955 17703 30981
rect 17703 30955 17729 30981
rect 17729 30955 17730 30981
rect 17702 30954 17730 30955
rect 17598 30197 17626 30198
rect 17598 30171 17599 30197
rect 17599 30171 17625 30197
rect 17625 30171 17626 30197
rect 17598 30170 17626 30171
rect 17650 30197 17678 30198
rect 17650 30171 17651 30197
rect 17651 30171 17677 30197
rect 17677 30171 17678 30197
rect 17650 30170 17678 30171
rect 17702 30197 17730 30198
rect 17702 30171 17703 30197
rect 17703 30171 17729 30197
rect 17729 30171 17730 30197
rect 17702 30170 17730 30171
rect 17598 29413 17626 29414
rect 17598 29387 17599 29413
rect 17599 29387 17625 29413
rect 17625 29387 17626 29413
rect 17598 29386 17626 29387
rect 17650 29413 17678 29414
rect 17650 29387 17651 29413
rect 17651 29387 17677 29413
rect 17677 29387 17678 29413
rect 17650 29386 17678 29387
rect 17702 29413 17730 29414
rect 17702 29387 17703 29413
rect 17703 29387 17729 29413
rect 17729 29387 17730 29413
rect 17702 29386 17730 29387
rect 17598 28629 17626 28630
rect 17598 28603 17599 28629
rect 17599 28603 17625 28629
rect 17625 28603 17626 28629
rect 17598 28602 17626 28603
rect 17650 28629 17678 28630
rect 17650 28603 17651 28629
rect 17651 28603 17677 28629
rect 17677 28603 17678 28629
rect 17650 28602 17678 28603
rect 17702 28629 17730 28630
rect 17702 28603 17703 28629
rect 17703 28603 17729 28629
rect 17729 28603 17730 28629
rect 17702 28602 17730 28603
rect 19782 27958 19810 27986
rect 17598 27845 17626 27846
rect 17598 27819 17599 27845
rect 17599 27819 17625 27845
rect 17625 27819 17626 27845
rect 17598 27818 17626 27819
rect 17650 27845 17678 27846
rect 17650 27819 17651 27845
rect 17651 27819 17677 27845
rect 17677 27819 17678 27845
rect 17650 27818 17678 27819
rect 17702 27845 17730 27846
rect 17702 27819 17703 27845
rect 17703 27819 17729 27845
rect 17729 27819 17730 27845
rect 17702 27818 17730 27819
rect 17598 27061 17626 27062
rect 17598 27035 17599 27061
rect 17599 27035 17625 27061
rect 17625 27035 17626 27061
rect 17598 27034 17626 27035
rect 17650 27061 17678 27062
rect 17650 27035 17651 27061
rect 17651 27035 17677 27061
rect 17677 27035 17678 27061
rect 17650 27034 17678 27035
rect 17702 27061 17730 27062
rect 17702 27035 17703 27061
rect 17703 27035 17729 27061
rect 17729 27035 17730 27061
rect 17702 27034 17730 27035
rect 19950 26865 19978 26866
rect 19950 26839 19951 26865
rect 19951 26839 19977 26865
rect 19977 26839 19978 26865
rect 19950 26838 19978 26839
rect 17598 26277 17626 26278
rect 17598 26251 17599 26277
rect 17599 26251 17625 26277
rect 17625 26251 17626 26277
rect 17598 26250 17626 26251
rect 17650 26277 17678 26278
rect 17650 26251 17651 26277
rect 17651 26251 17677 26277
rect 17677 26251 17678 26277
rect 17650 26250 17678 26251
rect 17702 26277 17730 26278
rect 17702 26251 17703 26277
rect 17703 26251 17729 26277
rect 17729 26251 17730 26277
rect 17702 26250 17730 26251
rect 20118 25998 20146 26026
rect 17598 25493 17626 25494
rect 17598 25467 17599 25493
rect 17599 25467 17625 25493
rect 17625 25467 17626 25493
rect 17598 25466 17626 25467
rect 17650 25493 17678 25494
rect 17650 25467 17651 25493
rect 17651 25467 17677 25493
rect 17677 25467 17678 25493
rect 17650 25466 17678 25467
rect 17702 25493 17730 25494
rect 17702 25467 17703 25493
rect 17703 25467 17729 25493
rect 17729 25467 17730 25493
rect 17702 25466 17730 25467
rect 17598 24709 17626 24710
rect 17598 24683 17599 24709
rect 17599 24683 17625 24709
rect 17625 24683 17626 24709
rect 17598 24682 17626 24683
rect 17650 24709 17678 24710
rect 17650 24683 17651 24709
rect 17651 24683 17677 24709
rect 17677 24683 17678 24709
rect 17650 24682 17678 24683
rect 17702 24709 17730 24710
rect 17702 24683 17703 24709
rect 17703 24683 17729 24709
rect 17729 24683 17730 24709
rect 17702 24682 17730 24683
rect 17598 23925 17626 23926
rect 17598 23899 17599 23925
rect 17599 23899 17625 23925
rect 17625 23899 17626 23925
rect 17598 23898 17626 23899
rect 17650 23925 17678 23926
rect 17650 23899 17651 23925
rect 17651 23899 17677 23925
rect 17677 23899 17678 23925
rect 17650 23898 17678 23899
rect 17702 23925 17730 23926
rect 17702 23899 17703 23925
rect 17703 23899 17729 23925
rect 17729 23899 17730 23925
rect 17702 23898 17730 23899
rect 17598 23141 17626 23142
rect 17598 23115 17599 23141
rect 17599 23115 17625 23141
rect 17625 23115 17626 23141
rect 17598 23114 17626 23115
rect 17650 23141 17678 23142
rect 17650 23115 17651 23141
rect 17651 23115 17677 23141
rect 17677 23115 17678 23141
rect 17650 23114 17678 23115
rect 17702 23141 17730 23142
rect 17702 23115 17703 23141
rect 17703 23115 17729 23141
rect 17729 23115 17730 23141
rect 17702 23114 17730 23115
rect 17262 22553 17290 22554
rect 17262 22527 17263 22553
rect 17263 22527 17289 22553
rect 17289 22527 17290 22553
rect 17262 22526 17290 22527
rect 17486 22553 17514 22554
rect 17486 22527 17487 22553
rect 17487 22527 17513 22553
rect 17513 22527 17514 22553
rect 17486 22526 17514 22527
rect 17598 22357 17626 22358
rect 17598 22331 17599 22357
rect 17599 22331 17625 22357
rect 17625 22331 17626 22357
rect 17598 22330 17626 22331
rect 17650 22357 17678 22358
rect 17650 22331 17651 22357
rect 17651 22331 17677 22357
rect 17677 22331 17678 22357
rect 17650 22330 17678 22331
rect 17702 22357 17730 22358
rect 17702 22331 17703 22357
rect 17703 22331 17729 22357
rect 17729 22331 17730 22357
rect 17702 22330 17730 22331
rect 17598 21573 17626 21574
rect 17598 21547 17599 21573
rect 17599 21547 17625 21573
rect 17625 21547 17626 21573
rect 17598 21546 17626 21547
rect 17650 21573 17678 21574
rect 17650 21547 17651 21573
rect 17651 21547 17677 21573
rect 17677 21547 17678 21573
rect 17650 21546 17678 21547
rect 17702 21573 17730 21574
rect 17702 21547 17703 21573
rect 17703 21547 17729 21573
rect 17729 21547 17730 21573
rect 17702 21546 17730 21547
rect 17598 20789 17626 20790
rect 17598 20763 17599 20789
rect 17599 20763 17625 20789
rect 17625 20763 17626 20789
rect 17598 20762 17626 20763
rect 17650 20789 17678 20790
rect 17650 20763 17651 20789
rect 17651 20763 17677 20789
rect 17677 20763 17678 20789
rect 17650 20762 17678 20763
rect 17702 20789 17730 20790
rect 17702 20763 17703 20789
rect 17703 20763 17729 20789
rect 17729 20763 17730 20789
rect 17702 20762 17730 20763
rect 18438 21742 18466 21770
rect 17990 20958 18018 20986
rect 18550 20902 18578 20930
rect 19054 20902 19082 20930
rect 19054 20593 19082 20594
rect 19054 20567 19055 20593
rect 19055 20567 19081 20593
rect 19081 20567 19082 20593
rect 19054 20566 19082 20567
rect 19446 20985 19474 20986
rect 19446 20959 19447 20985
rect 19447 20959 19473 20985
rect 19473 20959 19474 20985
rect 19446 20958 19474 20959
rect 19446 20510 19474 20538
rect 19950 20537 19978 20538
rect 19950 20511 19951 20537
rect 19951 20511 19977 20537
rect 19977 20511 19978 20537
rect 19950 20510 19978 20511
rect 17598 20005 17626 20006
rect 17598 19979 17599 20005
rect 17599 19979 17625 20005
rect 17625 19979 17626 20005
rect 17598 19978 17626 19979
rect 17650 20005 17678 20006
rect 17650 19979 17651 20005
rect 17651 19979 17677 20005
rect 17677 19979 17678 20005
rect 17650 19978 17678 19979
rect 17702 20005 17730 20006
rect 17702 19979 17703 20005
rect 17703 19979 17729 20005
rect 17729 19979 17730 20005
rect 17702 19978 17730 19979
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17430 18241 17458 18242
rect 17430 18215 17431 18241
rect 17431 18215 17457 18241
rect 17457 18215 17458 18241
rect 17430 18214 17458 18215
rect 17990 18214 18018 18242
rect 17990 17849 18018 17850
rect 17990 17823 17991 17849
rect 17991 17823 18017 17849
rect 18017 17823 18018 17849
rect 17990 17822 18018 17823
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17206 15806 17234 15834
rect 17430 15833 17458 15834
rect 17430 15807 17431 15833
rect 17431 15807 17457 15833
rect 17457 15807 17458 15833
rect 17430 15806 17458 15807
rect 19054 18241 19082 18242
rect 19054 18215 19055 18241
rect 19055 18215 19081 18241
rect 19081 18215 19082 18241
rect 19054 18214 19082 18215
rect 19334 17849 19362 17850
rect 19334 17823 19335 17849
rect 19335 17823 19361 17849
rect 19361 17823 19362 17849
rect 19334 17822 19362 17823
rect 17990 15806 18018 15834
rect 17990 15497 18018 15498
rect 17990 15471 17991 15497
rect 17991 15471 18017 15497
rect 18017 15471 18018 15497
rect 17990 15470 18018 15471
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 17430 13537 17458 13538
rect 17430 13511 17431 13537
rect 17431 13511 17457 13537
rect 17457 13511 17458 13537
rect 17430 13510 17458 13511
rect 19278 15806 19306 15834
rect 19278 15497 19306 15498
rect 19278 15471 19279 15497
rect 19279 15471 19305 15497
rect 19305 15471 19306 15497
rect 19278 15470 19306 15471
rect 19950 15833 19978 15834
rect 19950 15807 19951 15833
rect 19951 15807 19977 15833
rect 19977 15807 19978 15833
rect 19950 15806 19978 15807
rect 19446 14406 19474 14434
rect 19054 14321 19082 14322
rect 19054 14295 19055 14321
rect 19055 14295 19081 14321
rect 19081 14295 19082 14321
rect 19054 14294 19082 14295
rect 22638 33614 22666 33642
rect 22470 30926 22498 30954
rect 22414 29358 22442 29386
rect 21910 28854 21938 28882
rect 21686 28350 21714 28378
rect 20958 28014 20986 28042
rect 21406 28041 21434 28042
rect 21406 28015 21407 28041
rect 21407 28015 21433 28041
rect 21433 28015 21434 28041
rect 21406 28014 21434 28015
rect 21350 27734 21378 27762
rect 20678 26894 20706 26922
rect 20342 26865 20370 26866
rect 20342 26839 20343 26865
rect 20343 26839 20369 26865
rect 20369 26839 20370 26865
rect 20342 26838 20370 26839
rect 20510 26865 20538 26866
rect 20510 26839 20511 26865
rect 20511 26839 20537 26865
rect 20537 26839 20538 26865
rect 20510 26838 20538 26839
rect 21070 27313 21098 27314
rect 21070 27287 21071 27313
rect 21071 27287 21097 27313
rect 21097 27287 21098 27313
rect 21070 27286 21098 27287
rect 22414 28881 22442 28882
rect 22414 28855 22415 28881
rect 22415 28855 22441 28881
rect 22441 28855 22442 28881
rect 22414 28854 22442 28855
rect 22134 28574 22162 28602
rect 21910 28014 21938 28042
rect 22470 28406 22498 28434
rect 22190 28377 22218 28378
rect 22190 28351 22191 28377
rect 22191 28351 22217 28377
rect 22217 28351 22218 28377
rect 22190 28350 22218 28351
rect 22358 28377 22386 28378
rect 22358 28351 22359 28377
rect 22359 28351 22385 28377
rect 22385 28351 22386 28377
rect 22358 28350 22386 28351
rect 22638 29190 22666 29218
rect 22694 29582 22722 29610
rect 22526 28574 22554 28602
rect 21630 27734 21658 27762
rect 21574 27649 21602 27650
rect 21574 27623 21575 27649
rect 21575 27623 21601 27649
rect 21601 27623 21602 27649
rect 21574 27622 21602 27623
rect 22246 28041 22274 28042
rect 22246 28015 22247 28041
rect 22247 28015 22273 28041
rect 22273 28015 22274 28041
rect 22246 28014 22274 28015
rect 22022 27622 22050 27650
rect 21574 27286 21602 27314
rect 21798 27230 21826 27258
rect 20958 26894 20986 26922
rect 21070 26838 21098 26866
rect 21630 26865 21658 26866
rect 21630 26839 21631 26865
rect 21631 26839 21657 26865
rect 21657 26839 21658 26865
rect 21630 26838 21658 26839
rect 21798 26865 21826 26866
rect 21798 26839 21799 26865
rect 21799 26839 21825 26865
rect 21825 26839 21826 26865
rect 21798 26838 21826 26839
rect 21294 26473 21322 26474
rect 21294 26447 21295 26473
rect 21295 26447 21321 26473
rect 21321 26447 21322 26473
rect 21294 26446 21322 26447
rect 21966 27257 21994 27258
rect 21966 27231 21967 27257
rect 21967 27231 21993 27257
rect 21993 27231 21994 27257
rect 21966 27230 21994 27231
rect 21518 26446 21546 26474
rect 21238 26081 21266 26082
rect 21238 26055 21239 26081
rect 21239 26055 21265 26081
rect 21265 26055 21266 26081
rect 21238 26054 21266 26055
rect 20958 26025 20986 26026
rect 20958 25999 20959 26025
rect 20959 25999 20985 26025
rect 20985 25999 20986 26025
rect 21630 26473 21658 26474
rect 21630 26447 21631 26473
rect 21631 26447 21657 26473
rect 21657 26447 21658 26473
rect 21630 26446 21658 26447
rect 21630 26081 21658 26082
rect 21630 26055 21631 26081
rect 21631 26055 21657 26081
rect 21657 26055 21658 26081
rect 21630 26054 21658 26055
rect 21798 26081 21826 26082
rect 21798 26055 21799 26081
rect 21799 26055 21825 26081
rect 21825 26055 21826 26081
rect 21798 26054 21826 26055
rect 20958 25998 20986 25999
rect 21574 25998 21602 26026
rect 22638 28041 22666 28042
rect 22638 28015 22639 28041
rect 22639 28015 22665 28041
rect 22665 28015 22666 28041
rect 22638 28014 22666 28015
rect 22190 27593 22218 27594
rect 22190 27567 22191 27593
rect 22191 27567 22217 27593
rect 22217 27567 22218 27593
rect 22190 27566 22218 27567
rect 22414 27566 22442 27594
rect 22750 27566 22778 27594
rect 22526 27257 22554 27258
rect 22526 27231 22527 27257
rect 22527 27231 22553 27257
rect 22553 27231 22554 27257
rect 22526 27230 22554 27231
rect 22134 26473 22162 26474
rect 22134 26447 22135 26473
rect 22135 26447 22161 26473
rect 22161 26447 22162 26473
rect 22134 26446 22162 26447
rect 22134 26081 22162 26082
rect 22134 26055 22135 26081
rect 22135 26055 22161 26081
rect 22161 26055 22162 26081
rect 22134 26054 22162 26055
rect 22694 26838 22722 26866
rect 22694 26529 22722 26530
rect 22694 26503 22695 26529
rect 22695 26503 22721 26529
rect 22721 26503 22722 26529
rect 22694 26502 22722 26503
rect 22750 24961 22778 24962
rect 22750 24935 22751 24961
rect 22751 24935 22777 24961
rect 22777 24935 22778 24961
rect 22750 24934 22778 24935
rect 23086 29582 23114 29610
rect 23030 29217 23058 29218
rect 23030 29191 23031 29217
rect 23031 29191 23057 29217
rect 23057 29191 23058 29217
rect 23030 29190 23058 29191
rect 23030 28854 23058 28882
rect 23366 29609 23394 29610
rect 23366 29583 23367 29609
rect 23367 29583 23393 29609
rect 23393 29583 23394 29609
rect 23366 29582 23394 29583
rect 23310 29358 23338 29386
rect 23590 29358 23618 29386
rect 23310 28798 23338 28826
rect 23030 28433 23058 28434
rect 23030 28407 23031 28433
rect 23031 28407 23057 28433
rect 23057 28407 23058 28433
rect 23030 28406 23058 28407
rect 23534 28881 23562 28882
rect 23534 28855 23535 28881
rect 23535 28855 23561 28881
rect 23561 28855 23562 28881
rect 23534 28854 23562 28855
rect 23646 28825 23674 28826
rect 23646 28799 23647 28825
rect 23647 28799 23673 28825
rect 23673 28799 23674 28825
rect 23646 28798 23674 28799
rect 23590 28574 23618 28602
rect 23142 28377 23170 28378
rect 23142 28351 23143 28377
rect 23143 28351 23169 28377
rect 23169 28351 23170 28377
rect 23142 28350 23170 28351
rect 23814 28825 23842 28826
rect 23814 28799 23815 28825
rect 23815 28799 23841 28825
rect 23841 28799 23842 28825
rect 23814 28798 23842 28799
rect 23254 27678 23282 27706
rect 22974 27593 23002 27594
rect 22974 27567 22975 27593
rect 22975 27567 23001 27593
rect 23001 27567 23002 27593
rect 22974 27566 23002 27567
rect 23534 27593 23562 27594
rect 23534 27567 23535 27593
rect 23535 27567 23561 27593
rect 23561 27567 23562 27593
rect 23534 27566 23562 27567
rect 23702 27678 23730 27706
rect 22918 27257 22946 27258
rect 22918 27231 22919 27257
rect 22919 27231 22945 27257
rect 22945 27231 22946 27257
rect 22918 27230 22946 27231
rect 22918 26894 22946 26922
rect 23086 26894 23114 26922
rect 23422 26865 23450 26866
rect 23422 26839 23423 26865
rect 23423 26839 23449 26865
rect 23449 26839 23450 26865
rect 23422 26838 23450 26839
rect 23478 26894 23506 26922
rect 22862 26529 22890 26530
rect 22862 26503 22863 26529
rect 22863 26503 22889 26529
rect 22889 26503 22890 26529
rect 22862 26502 22890 26503
rect 22974 25550 23002 25578
rect 23030 26054 23058 26082
rect 23310 25550 23338 25578
rect 23142 24961 23170 24962
rect 23142 24935 23143 24961
rect 23143 24935 23169 24961
rect 23169 24935 23170 24961
rect 23142 24934 23170 24935
rect 23478 24457 23506 24458
rect 23478 24431 23479 24457
rect 23479 24431 23505 24457
rect 23505 24431 23506 24457
rect 23478 24430 23506 24431
rect 23702 23337 23730 23338
rect 23702 23311 23703 23337
rect 23703 23311 23729 23337
rect 23729 23311 23730 23337
rect 23702 23310 23730 23311
rect 23198 22889 23226 22890
rect 23198 22863 23199 22889
rect 23199 22863 23225 22889
rect 23225 22863 23226 22889
rect 23198 22862 23226 22863
rect 23366 22889 23394 22890
rect 23366 22863 23367 22889
rect 23367 22863 23393 22889
rect 23393 22863 23394 22889
rect 23366 22862 23394 22863
rect 24038 24457 24066 24458
rect 24038 24431 24039 24457
rect 24039 24431 24065 24457
rect 24065 24431 24066 24457
rect 24038 24430 24066 24431
rect 23870 23337 23898 23338
rect 23870 23311 23871 23337
rect 23871 23311 23897 23337
rect 23897 23311 23898 23337
rect 23870 23310 23898 23311
rect 23534 22694 23562 22722
rect 20510 20593 20538 20594
rect 20510 20567 20511 20593
rect 20511 20567 20537 20593
rect 20537 20567 20538 20593
rect 20510 20566 20538 20567
rect 21182 20510 21210 20538
rect 20510 19809 20538 19810
rect 20510 19783 20511 19809
rect 20511 19783 20537 19809
rect 20537 19783 20538 19809
rect 20510 19782 20538 19783
rect 20958 19782 20986 19810
rect 20958 19417 20986 19418
rect 20958 19391 20959 19417
rect 20959 19391 20985 19417
rect 20985 19391 20986 19417
rect 20958 19390 20986 19391
rect 21798 19334 21826 19362
rect 22526 19417 22554 19418
rect 22526 19391 22527 19417
rect 22527 19391 22553 19417
rect 22553 19391 22554 19417
rect 22526 19390 22554 19391
rect 20230 18241 20258 18242
rect 20230 18215 20231 18241
rect 20231 18215 20257 18241
rect 20257 18215 20258 18241
rect 20230 18214 20258 18215
rect 20174 14350 20202 14378
rect 20790 16254 20818 16282
rect 20958 16281 20986 16282
rect 20958 16255 20959 16281
rect 20959 16255 20985 16281
rect 20985 16255 20986 16281
rect 20958 16254 20986 16255
rect 23534 20174 23562 20202
rect 23702 22862 23730 22890
rect 24038 22862 24066 22890
rect 23982 22694 24010 22722
rect 23478 19334 23506 19362
rect 22246 16646 22274 16674
rect 22246 16281 22274 16282
rect 22246 16255 22247 16281
rect 22247 16255 22273 16281
rect 22273 16255 22274 16281
rect 22246 16254 22274 16255
rect 22750 16673 22778 16674
rect 22750 16647 22751 16673
rect 22751 16647 22777 16673
rect 22777 16647 22778 16673
rect 22750 16646 22778 16647
rect 21518 15806 21546 15834
rect 20230 14321 20258 14322
rect 20230 14295 20231 14321
rect 20231 14295 20257 14321
rect 20257 14295 20258 14321
rect 20230 14294 20258 14295
rect 21014 14406 21042 14434
rect 21462 14713 21490 14714
rect 21462 14687 21463 14713
rect 21463 14687 21489 14713
rect 21489 14687 21490 14713
rect 21462 14686 21490 14687
rect 20958 13929 20986 13930
rect 20958 13903 20959 13929
rect 20959 13903 20985 13929
rect 20985 13903 20986 13929
rect 20958 13902 20986 13903
rect 20510 13537 20538 13538
rect 20510 13511 20511 13537
rect 20511 13511 20537 13537
rect 20537 13511 20538 13537
rect 20510 13510 20538 13511
rect 17262 13145 17290 13146
rect 17262 13119 17263 13145
rect 17263 13119 17289 13145
rect 17289 13119 17290 13145
rect 17262 13118 17290 13119
rect 17486 13145 17514 13146
rect 17486 13119 17487 13145
rect 17487 13119 17513 13145
rect 17513 13119 17514 13145
rect 17486 13118 17514 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 18270 13454 18298 13482
rect 17766 12558 17794 12586
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 17430 11969 17458 11970
rect 17430 11943 17431 11969
rect 17431 11943 17457 11969
rect 17457 11943 17458 11969
rect 17430 11942 17458 11943
rect 17766 11942 17794 11970
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18438 12334 18466 12362
rect 18550 12361 18578 12362
rect 18550 12335 18551 12361
rect 18551 12335 18577 12361
rect 18577 12335 18578 12361
rect 18550 12334 18578 12335
rect 18438 11577 18466 11578
rect 18438 11551 18439 11577
rect 18439 11551 18465 11577
rect 18465 11551 18466 11577
rect 18438 11550 18466 11551
rect 18718 11942 18746 11970
rect 19054 12753 19082 12754
rect 19054 12727 19055 12753
rect 19055 12727 19081 12753
rect 19081 12727 19082 12753
rect 19054 12726 19082 12727
rect 20958 13510 20986 13538
rect 22694 15806 22722 15834
rect 22694 15497 22722 15498
rect 22694 15471 22695 15497
rect 22695 15471 22721 15497
rect 22721 15471 22722 15497
rect 22694 15470 22722 15471
rect 22246 15078 22274 15106
rect 22246 13902 22274 13930
rect 20510 12753 20538 12754
rect 20510 12727 20511 12753
rect 20511 12727 20537 12753
rect 20537 12727 20538 12753
rect 20510 12726 20538 12727
rect 19054 12334 19082 12362
rect 19334 12558 19362 12586
rect 21630 12361 21658 12362
rect 21630 12335 21631 12361
rect 21631 12335 21657 12361
rect 21657 12335 21658 12361
rect 21630 12334 21658 12335
rect 19222 11969 19250 11970
rect 19222 11943 19223 11969
rect 19223 11943 19249 11969
rect 19249 11943 19250 11969
rect 19222 11942 19250 11943
rect 19446 11969 19474 11970
rect 19446 11943 19447 11969
rect 19447 11943 19473 11969
rect 19473 11943 19474 11969
rect 19446 11942 19474 11943
rect 22134 12361 22162 12362
rect 22134 12335 22135 12361
rect 22135 12335 22161 12361
rect 22161 12335 22162 12361
rect 22134 12334 22162 12335
rect 22750 15105 22778 15106
rect 22750 15079 22751 15105
rect 22751 15079 22777 15105
rect 22777 15079 22778 15105
rect 22750 15078 22778 15079
rect 23198 15806 23226 15834
rect 24038 17486 24066 17514
rect 23422 15806 23450 15834
rect 22918 15497 22946 15498
rect 22918 15471 22919 15497
rect 22919 15471 22945 15497
rect 22945 15471 22946 15497
rect 22918 15470 22946 15471
rect 22750 14713 22778 14714
rect 22750 14687 22751 14713
rect 22751 14687 22777 14713
rect 22777 14687 22778 14713
rect 22750 14686 22778 14687
rect 22918 14713 22946 14714
rect 22918 14687 22919 14713
rect 22919 14687 22945 14713
rect 22945 14687 22946 14713
rect 22918 14686 22946 14687
rect 23198 14686 23226 14714
rect 24038 14798 24066 14826
rect 22694 12334 22722 12362
rect 22862 14350 22890 14378
rect 20902 11326 20930 11354
rect 21630 11326 21658 11354
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 19446 10038 19474 10066
rect 22582 11577 22610 11578
rect 22582 11551 22583 11577
rect 22583 11551 22609 11577
rect 22609 11551 22610 11577
rect 22582 11550 22610 11551
rect 21798 10934 21826 10962
rect 20398 10318 20426 10346
rect 21854 10878 21882 10906
rect 22078 10878 22106 10906
rect 20902 10345 20930 10346
rect 20902 10319 20903 10345
rect 20903 10319 20929 10345
rect 20929 10319 20930 10345
rect 20902 10318 20930 10319
rect 20006 10038 20034 10066
rect 21182 10038 21210 10066
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 17430 9561 17458 9562
rect 17430 9535 17431 9561
rect 17431 9535 17457 9561
rect 17457 9535 17458 9561
rect 17430 9534 17458 9535
rect 17990 9534 18018 9562
rect 21182 9422 21210 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 17094 8022 17122 8050
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 17430 7993 17458 7994
rect 17430 7967 17431 7993
rect 17431 7967 17457 7993
rect 17457 7967 17458 7993
rect 17430 7966 17458 7967
rect 17766 7966 17794 7994
rect 17094 7657 17122 7658
rect 17094 7631 17095 7657
rect 17095 7631 17121 7657
rect 17121 7631 17122 7657
rect 17094 7630 17122 7631
rect 17486 7574 17514 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17206 6118 17234 6146
rect 16814 6089 16842 6090
rect 16814 6063 16815 6089
rect 16815 6063 16841 6089
rect 16841 6063 16842 6089
rect 16814 6062 16842 6063
rect 15918 5782 15946 5810
rect 15470 4998 15498 5026
rect 15918 4998 15946 5026
rect 17206 5894 17234 5922
rect 17990 7574 18018 7602
rect 18550 8358 18578 8386
rect 19054 8358 19082 8386
rect 19054 8049 19082 8050
rect 19054 8023 19055 8049
rect 19055 8023 19081 8049
rect 19081 8023 19082 8049
rect 19054 8022 19082 8023
rect 22526 10318 22554 10346
rect 22582 10065 22610 10066
rect 22582 10039 22583 10065
rect 22583 10039 22609 10065
rect 22609 10039 22610 10065
rect 22582 10038 22610 10039
rect 23814 12110 23842 12138
rect 23814 11326 23842 11354
rect 22862 10038 22890 10066
rect 22358 9198 22386 9226
rect 22582 9225 22610 9226
rect 22582 9199 22583 9225
rect 22583 9199 22609 9225
rect 22609 9199 22610 9225
rect 22582 9198 22610 9199
rect 18550 7657 18578 7658
rect 18550 7631 18551 7657
rect 18551 7631 18577 7657
rect 18577 7631 18578 7657
rect 18550 7630 18578 7631
rect 18718 7574 18746 7602
rect 18942 7574 18970 7602
rect 19222 7574 19250 7602
rect 22806 8022 22834 8050
rect 20230 7518 20258 7546
rect 18774 7265 18802 7266
rect 18774 7239 18775 7265
rect 18775 7239 18801 7265
rect 18801 7239 18802 7265
rect 18774 7238 18802 7239
rect 17094 5278 17122 5306
rect 15470 4158 15498 4186
rect 15078 4129 15106 4130
rect 15078 4103 15079 4129
rect 15079 4103 15105 4129
rect 15105 4103 15106 4129
rect 15078 4102 15106 4103
rect 14574 3737 14602 3738
rect 14574 3711 14575 3737
rect 14575 3711 14601 3737
rect 14601 3711 14602 3737
rect 14574 3710 14602 3711
rect 14574 3318 14602 3346
rect 13118 2534 13146 2562
rect 15078 3710 15106 3738
rect 15918 4158 15946 4186
rect 16254 4129 16282 4130
rect 16254 4103 16255 4129
rect 16255 4103 16281 4129
rect 16281 4103 16282 4129
rect 16254 4102 16282 4103
rect 16254 3345 16282 3346
rect 16254 3319 16255 3345
rect 16255 3319 16281 3345
rect 16281 3319 16282 3345
rect 16254 3318 16282 3319
rect 12894 1750 12922 1778
rect 14798 2561 14826 2562
rect 14798 2535 14799 2561
rect 14799 2535 14825 2561
rect 14825 2535 14826 2561
rect 14798 2534 14826 2535
rect 14294 2030 14322 2058
rect 14518 2030 14546 2058
rect 13846 1777 13874 1778
rect 13846 1751 13847 1777
rect 13847 1751 13873 1777
rect 13873 1751 13874 1777
rect 13846 1750 13874 1751
rect 14798 2030 14826 2058
rect 16814 3318 16842 3346
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17430 5697 17458 5698
rect 17430 5671 17431 5697
rect 17431 5671 17457 5697
rect 17457 5671 17458 5697
rect 17430 5670 17458 5671
rect 18718 6873 18746 6874
rect 18718 6847 18719 6873
rect 18719 6847 18745 6873
rect 18745 6847 18746 6873
rect 18718 6846 18746 6847
rect 18270 6089 18298 6090
rect 18270 6063 18271 6089
rect 18271 6063 18297 6089
rect 18297 6063 18298 6089
rect 18270 6062 18298 6063
rect 18662 6062 18690 6090
rect 17766 5670 17794 5698
rect 17766 5361 17794 5362
rect 17766 5335 17767 5361
rect 17767 5335 17793 5361
rect 17793 5335 17794 5361
rect 17766 5334 17794 5335
rect 18550 5670 18578 5698
rect 18550 5305 18578 5306
rect 18550 5279 18551 5305
rect 18551 5279 18577 5305
rect 18577 5279 18578 5305
rect 18550 5278 18578 5279
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17430 4158 17458 4186
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 16254 2534 16282 2562
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 15358 1750 15386 1778
rect 18942 6873 18970 6874
rect 18942 6847 18943 6873
rect 18943 6847 18969 6873
rect 18969 6847 18970 6873
rect 18942 6846 18970 6847
rect 20790 7518 20818 7546
rect 20230 7265 20258 7266
rect 20230 7239 20231 7265
rect 20231 7239 20257 7265
rect 20257 7239 20258 7265
rect 20230 7238 20258 7239
rect 19222 6846 19250 6874
rect 19446 6481 19474 6482
rect 19446 6455 19447 6481
rect 19447 6455 19473 6481
rect 19473 6455 19474 6481
rect 19446 6454 19474 6455
rect 18774 6062 18802 6090
rect 18830 6118 18858 6146
rect 19222 6118 19250 6146
rect 19054 5697 19082 5698
rect 19054 5671 19055 5697
rect 19055 5671 19081 5697
rect 19081 5671 19082 5697
rect 19054 5670 19082 5671
rect 18718 5334 18746 5362
rect 18942 5334 18970 5362
rect 20678 6481 20706 6482
rect 20678 6455 20679 6481
rect 20679 6455 20705 6481
rect 20705 6455 20706 6481
rect 20678 6454 20706 6455
rect 21014 6481 21042 6482
rect 21014 6455 21015 6481
rect 21015 6455 21041 6481
rect 21041 6455 21042 6481
rect 21014 6454 21042 6455
rect 20230 5670 20258 5698
rect 19222 5334 19250 5362
rect 23758 10374 23786 10402
rect 22918 9225 22946 9226
rect 22918 9199 22919 9225
rect 22919 9199 22945 9225
rect 22945 9199 22946 9225
rect 22918 9198 22946 9199
rect 24038 11577 24066 11578
rect 24038 11551 24039 11577
rect 24039 11551 24065 11577
rect 24065 11551 24066 11577
rect 24038 11550 24066 11551
rect 24038 10401 24066 10402
rect 24038 10375 24039 10401
rect 24039 10375 24065 10401
rect 24065 10375 24066 10401
rect 24038 10374 24066 10375
rect 24038 6734 24066 6762
rect 23814 4046 23842 4074
rect 24038 1358 24066 1386
<< metal3 >>
rect 24600 33642 25000 33656
rect 22633 33614 22638 33642
rect 22666 33614 25000 33642
rect 24600 33600 25000 33614
rect 2233 33306 2238 33334
rect 2266 33306 2290 33334
rect 2318 33306 2342 33334
rect 2370 33306 2375 33334
rect 17593 33306 17598 33334
rect 17626 33306 17650 33334
rect 17678 33306 17702 33334
rect 17730 33306 17735 33334
rect 9913 32914 9918 32942
rect 9946 32914 9970 32942
rect 9998 32914 10022 32942
rect 10050 32914 10055 32942
rect 0 32802 400 32816
rect 0 32774 1750 32802
rect 1778 32774 1783 32802
rect 0 32760 400 32774
rect 2233 32522 2238 32550
rect 2266 32522 2290 32550
rect 2318 32522 2342 32550
rect 2370 32522 2375 32550
rect 17593 32522 17598 32550
rect 17626 32522 17650 32550
rect 17678 32522 17702 32550
rect 17730 32522 17735 32550
rect 9913 32130 9918 32158
rect 9946 32130 9970 32158
rect 9998 32130 10022 32158
rect 10050 32130 10055 32158
rect 2233 31738 2238 31766
rect 2266 31738 2290 31766
rect 2318 31738 2342 31766
rect 2370 31738 2375 31766
rect 17593 31738 17598 31766
rect 17626 31738 17650 31766
rect 17678 31738 17702 31766
rect 17730 31738 17735 31766
rect 9913 31346 9918 31374
rect 9946 31346 9970 31374
rect 9998 31346 10022 31374
rect 10050 31346 10055 31374
rect 2233 30954 2238 30982
rect 2266 30954 2290 30982
rect 2318 30954 2342 30982
rect 2370 30954 2375 30982
rect 17593 30954 17598 30982
rect 17626 30954 17650 30982
rect 17678 30954 17702 30982
rect 17730 30954 17735 30982
rect 24600 30954 25000 30968
rect 22465 30926 22470 30954
rect 22498 30926 25000 30954
rect 24600 30912 25000 30926
rect 9913 30562 9918 30590
rect 9946 30562 9970 30590
rect 9998 30562 10022 30590
rect 10050 30562 10055 30590
rect 2233 30170 2238 30198
rect 2266 30170 2290 30198
rect 2318 30170 2342 30198
rect 2370 30170 2375 30198
rect 17593 30170 17598 30198
rect 17626 30170 17650 30198
rect 17678 30170 17702 30198
rect 17730 30170 17735 30198
rect 9913 29778 9918 29806
rect 9946 29778 9970 29806
rect 9998 29778 10022 29806
rect 10050 29778 10055 29806
rect 7849 29582 7854 29610
rect 7882 29582 22694 29610
rect 22722 29582 23086 29610
rect 23114 29582 23366 29610
rect 23394 29582 23399 29610
rect 2233 29386 2238 29414
rect 2266 29386 2290 29414
rect 2318 29386 2342 29414
rect 2370 29386 2375 29414
rect 17593 29386 17598 29414
rect 17626 29386 17650 29414
rect 17678 29386 17702 29414
rect 17730 29386 17735 29414
rect 22409 29358 22414 29386
rect 22442 29358 23310 29386
rect 23338 29358 23590 29386
rect 23618 29358 23623 29386
rect 22633 29190 22638 29218
rect 22666 29190 23030 29218
rect 23058 29190 23063 29218
rect 9913 28994 9918 29022
rect 9946 28994 9970 29022
rect 9998 28994 10022 29022
rect 10050 28994 10055 29022
rect 21905 28854 21910 28882
rect 21938 28854 22414 28882
rect 22442 28854 22447 28882
rect 23025 28854 23030 28882
rect 23058 28854 23534 28882
rect 23562 28854 23567 28882
rect 23305 28798 23310 28826
rect 23338 28798 23646 28826
rect 23674 28798 23814 28826
rect 23842 28798 23847 28826
rect 2233 28602 2238 28630
rect 2266 28602 2290 28630
rect 2318 28602 2342 28630
rect 2370 28602 2375 28630
rect 17593 28602 17598 28630
rect 17626 28602 17650 28630
rect 17678 28602 17702 28630
rect 17730 28602 17735 28630
rect 22129 28574 22134 28602
rect 22162 28574 22526 28602
rect 22554 28574 22559 28602
rect 23585 28574 23590 28602
rect 23618 28574 24682 28602
rect 0 28434 400 28448
rect 24654 28434 24682 28574
rect 0 28406 1806 28434
rect 1834 28406 1839 28434
rect 22465 28406 22470 28434
rect 22498 28406 23030 28434
rect 23058 28406 23063 28434
rect 24542 28406 24682 28434
rect 0 28392 400 28406
rect 21681 28350 21686 28378
rect 21714 28350 22190 28378
rect 22218 28350 22358 28378
rect 22386 28350 23142 28378
rect 23170 28350 23175 28378
rect 24542 28266 24570 28406
rect 24600 28266 25000 28280
rect 24542 28238 25000 28266
rect 9913 28210 9918 28238
rect 9946 28210 9970 28238
rect 9998 28210 10022 28238
rect 10050 28210 10055 28238
rect 24600 28224 25000 28238
rect 20953 28014 20958 28042
rect 20986 28014 21406 28042
rect 21434 28014 21910 28042
rect 21938 28014 21943 28042
rect 22241 28014 22246 28042
rect 22274 28014 22638 28042
rect 22666 28014 22671 28042
rect 10929 27958 10934 27986
rect 10962 27958 19782 27986
rect 19810 27958 19815 27986
rect 2233 27818 2238 27846
rect 2266 27818 2290 27846
rect 2318 27818 2342 27846
rect 2370 27818 2375 27846
rect 17593 27818 17598 27846
rect 17626 27818 17650 27846
rect 17678 27818 17702 27846
rect 17730 27818 17735 27846
rect 5334 27734 5838 27762
rect 5866 27734 5871 27762
rect 21345 27734 21350 27762
rect 21378 27734 21630 27762
rect 21658 27734 21663 27762
rect 5334 27706 5362 27734
rect 3985 27678 3990 27706
rect 4018 27678 4270 27706
rect 4298 27678 4998 27706
rect 5026 27678 5362 27706
rect 23249 27678 23254 27706
rect 23282 27678 23702 27706
rect 23730 27678 23735 27706
rect 21569 27622 21574 27650
rect 21602 27622 22022 27650
rect 22050 27622 22055 27650
rect 22185 27566 22190 27594
rect 22218 27566 22414 27594
rect 22442 27566 22447 27594
rect 22745 27566 22750 27594
rect 22778 27566 22974 27594
rect 23002 27566 23534 27594
rect 23562 27566 23567 27594
rect 9913 27426 9918 27454
rect 9946 27426 9970 27454
rect 9998 27426 10022 27454
rect 10050 27426 10055 27454
rect 21065 27286 21070 27314
rect 21098 27286 21574 27314
rect 21602 27286 21607 27314
rect 5161 27230 5166 27258
rect 5194 27230 6622 27258
rect 6650 27230 7126 27258
rect 7154 27230 7159 27258
rect 21793 27230 21798 27258
rect 21826 27230 21966 27258
rect 21994 27230 22526 27258
rect 22554 27230 22918 27258
rect 22946 27230 22951 27258
rect 2081 27174 2086 27202
rect 2114 27174 8414 27202
rect 8442 27174 8862 27202
rect 8890 27174 10598 27202
rect 10626 27174 10631 27202
rect 2233 27034 2238 27062
rect 2266 27034 2290 27062
rect 2318 27034 2342 27062
rect 2370 27034 2375 27062
rect 17593 27034 17598 27062
rect 17626 27034 17650 27062
rect 17678 27034 17702 27062
rect 17730 27034 17735 27062
rect 1353 26894 1358 26922
rect 1386 26894 1862 26922
rect 1890 26894 1895 26922
rect 2529 26894 2534 26922
rect 2562 26894 3486 26922
rect 3514 26894 3710 26922
rect 3738 26894 3743 26922
rect 7121 26894 7126 26922
rect 7154 26894 8582 26922
rect 8610 26894 8615 26922
rect 10593 26894 10598 26922
rect 10626 26894 11046 26922
rect 11074 26894 11079 26922
rect 20673 26894 20678 26922
rect 20706 26894 20958 26922
rect 20986 26894 20991 26922
rect 22913 26894 22918 26922
rect 22946 26894 23086 26922
rect 23114 26894 23478 26922
rect 23506 26894 23511 26922
rect 19945 26838 19950 26866
rect 19978 26838 20342 26866
rect 20370 26838 20510 26866
rect 20538 26838 21070 26866
rect 21098 26838 21630 26866
rect 21658 26838 21798 26866
rect 21826 26838 22694 26866
rect 22722 26838 23422 26866
rect 23450 26838 23455 26866
rect 10033 26726 10038 26754
rect 10066 26726 10990 26754
rect 11018 26726 11023 26754
rect 9913 26642 9918 26670
rect 9946 26642 9970 26670
rect 9998 26642 10022 26670
rect 10050 26642 10055 26670
rect 22689 26502 22694 26530
rect 22722 26502 22862 26530
rect 22890 26502 22895 26530
rect 10985 26446 10990 26474
rect 11018 26446 12726 26474
rect 12754 26446 12759 26474
rect 21289 26446 21294 26474
rect 21322 26446 21518 26474
rect 21546 26446 21630 26474
rect 21658 26446 22134 26474
rect 22162 26446 22167 26474
rect 2233 26250 2238 26278
rect 2266 26250 2290 26278
rect 2318 26250 2342 26278
rect 2370 26250 2375 26278
rect 17593 26250 17598 26278
rect 17626 26250 17650 26278
rect 17678 26250 17702 26278
rect 17730 26250 17735 26278
rect 4937 26054 4942 26082
rect 4970 26054 5166 26082
rect 5194 26054 5334 26082
rect 5362 26054 5367 26082
rect 21233 26054 21238 26082
rect 21266 26054 21630 26082
rect 21658 26054 21798 26082
rect 21826 26054 21831 26082
rect 22129 26054 22134 26082
rect 22162 26054 23030 26082
rect 23058 26054 23063 26082
rect 8857 25998 8862 26026
rect 8890 25998 8974 26026
rect 9002 25998 9007 26026
rect 11041 25998 11046 26026
rect 11074 25998 12558 26026
rect 12586 25998 12591 26026
rect 20113 25998 20118 26026
rect 20146 25998 20958 26026
rect 20986 25998 21574 26026
rect 21602 25998 21607 26026
rect 9913 25858 9918 25886
rect 9946 25858 9970 25886
rect 9998 25858 10022 25886
rect 10050 25858 10055 25886
rect 1577 25662 1582 25690
rect 1610 25662 1750 25690
rect 1778 25662 2142 25690
rect 2170 25662 6342 25690
rect 6370 25662 8414 25690
rect 8442 25662 8918 25690
rect 8946 25662 10598 25690
rect 10626 25662 11102 25690
rect 11130 25662 11135 25690
rect 24600 25578 25000 25592
rect 4769 25550 4774 25578
rect 4802 25550 5110 25578
rect 5138 25550 5143 25578
rect 22969 25550 22974 25578
rect 23002 25550 23310 25578
rect 23338 25550 25000 25578
rect 24600 25536 25000 25550
rect 2233 25466 2238 25494
rect 2266 25466 2290 25494
rect 2318 25466 2342 25494
rect 2370 25466 2375 25494
rect 17593 25466 17598 25494
rect 17626 25466 17650 25494
rect 17678 25466 17702 25494
rect 17730 25466 17735 25494
rect 2473 25270 2478 25298
rect 2506 25270 3150 25298
rect 3178 25270 3183 25298
rect 3817 25270 3822 25298
rect 3850 25270 4774 25298
rect 4802 25270 4807 25298
rect 8857 25270 8862 25298
rect 8890 25270 8974 25298
rect 9002 25270 9007 25298
rect 12945 25270 12950 25298
rect 12978 25270 13510 25298
rect 13538 25270 13543 25298
rect 12553 25214 12558 25242
rect 12586 25214 13118 25242
rect 13146 25214 14518 25242
rect 14546 25214 14551 25242
rect 8577 25158 8582 25186
rect 8610 25158 9142 25186
rect 9170 25158 10318 25186
rect 10346 25158 10351 25186
rect 9913 25074 9918 25102
rect 9946 25074 9970 25102
rect 9998 25074 10022 25102
rect 10050 25074 10055 25102
rect 22745 24934 22750 24962
rect 22778 24934 23142 24962
rect 23170 24934 23175 24962
rect 2233 24682 2238 24710
rect 2266 24682 2290 24710
rect 2318 24682 2342 24710
rect 2370 24682 2375 24710
rect 17593 24682 17598 24710
rect 17626 24682 17650 24710
rect 17678 24682 17702 24710
rect 17730 24682 17735 24710
rect 10313 24486 10318 24514
rect 10346 24486 10822 24514
rect 10850 24486 12278 24514
rect 12306 24486 12311 24514
rect 23473 24430 23478 24458
rect 23506 24430 24038 24458
rect 24066 24430 24071 24458
rect 11097 24374 11102 24402
rect 11130 24374 12558 24402
rect 12586 24374 13118 24402
rect 13146 24374 14574 24402
rect 14602 24374 14607 24402
rect 1857 24318 1862 24346
rect 1890 24318 3374 24346
rect 3402 24318 3822 24346
rect 3850 24318 3855 24346
rect 13337 24318 13342 24346
rect 13370 24318 15134 24346
rect 15162 24318 15167 24346
rect 9913 24290 9918 24318
rect 9946 24290 9970 24318
rect 9998 24290 10022 24318
rect 10050 24290 10055 24318
rect 7625 24206 7630 24234
rect 7658 24206 8022 24234
rect 8050 24206 8862 24234
rect 8890 24206 9478 24234
rect 9506 24206 10038 24234
rect 10066 24206 10071 24234
rect 13505 24206 13510 24234
rect 13538 24206 15134 24234
rect 15162 24206 15167 24234
rect 3033 24094 3038 24122
rect 3066 24094 4494 24122
rect 4522 24094 4527 24122
rect 6169 24094 6174 24122
rect 6202 24094 6454 24122
rect 6482 24094 6487 24122
rect 10593 24094 10598 24122
rect 10626 24094 11102 24122
rect 11130 24094 11135 24122
rect 0 24066 400 24080
rect 0 24038 1358 24066
rect 1386 24038 1391 24066
rect 0 24024 400 24038
rect 2233 23898 2238 23926
rect 2266 23898 2290 23926
rect 2318 23898 2342 23926
rect 2370 23898 2375 23926
rect 17593 23898 17598 23926
rect 17626 23898 17650 23926
rect 17678 23898 17702 23926
rect 17730 23898 17735 23926
rect 5553 23702 5558 23730
rect 5586 23702 6678 23730
rect 6706 23702 7126 23730
rect 7154 23702 8582 23730
rect 8610 23702 8615 23730
rect 11489 23702 11494 23730
rect 11522 23702 11718 23730
rect 11746 23702 13454 23730
rect 13482 23702 13487 23730
rect 15465 23702 15470 23730
rect 15498 23702 16814 23730
rect 16842 23702 16847 23730
rect 2473 23646 2478 23674
rect 2506 23646 3038 23674
rect 3066 23646 3071 23674
rect 3145 23646 3150 23674
rect 3178 23646 4494 23674
rect 4522 23646 4527 23674
rect 6449 23646 6454 23674
rect 6482 23646 8022 23674
rect 8050 23646 8055 23674
rect 4097 23590 4102 23618
rect 4130 23590 4214 23618
rect 4242 23590 5054 23618
rect 5082 23590 5087 23618
rect 9310 23590 10990 23618
rect 11018 23590 11270 23618
rect 11298 23590 11303 23618
rect 9310 23562 9338 23590
rect 1353 23534 1358 23562
rect 1386 23534 1862 23562
rect 1890 23534 1895 23562
rect 4993 23534 4998 23562
rect 5026 23534 6174 23562
rect 6202 23534 6207 23562
rect 7009 23534 7014 23562
rect 7042 23534 7518 23562
rect 7546 23534 9310 23562
rect 9338 23534 9343 23562
rect 9913 23506 9918 23534
rect 9946 23506 9970 23534
rect 9998 23506 10022 23534
rect 10050 23506 10055 23534
rect 14513 23478 14518 23506
rect 14546 23478 15078 23506
rect 15106 23478 15111 23506
rect 12273 23310 12278 23338
rect 12306 23310 12838 23338
rect 12866 23310 12871 23338
rect 23697 23310 23702 23338
rect 23730 23310 23870 23338
rect 23898 23310 23903 23338
rect 2233 23114 2238 23142
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2370 23114 2375 23142
rect 17593 23114 17598 23142
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17730 23114 17735 23142
rect 4097 22918 4102 22946
rect 4130 22918 4214 22946
rect 4242 22918 4247 22946
rect 15073 22918 15078 22946
rect 15106 22918 16254 22946
rect 16282 22918 16287 22946
rect 24600 22890 25000 22904
rect 23193 22862 23198 22890
rect 23226 22862 23366 22890
rect 23394 22862 23702 22890
rect 23730 22862 23735 22890
rect 24033 22862 24038 22890
rect 24066 22862 25000 22890
rect 24600 22848 25000 22862
rect 9913 22722 9918 22750
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 10050 22722 10055 22750
rect 23529 22694 23534 22722
rect 23562 22694 23982 22722
rect 24010 22694 24015 22722
rect 4489 22526 4494 22554
rect 4522 22526 4998 22554
rect 5026 22526 5031 22554
rect 7569 22526 7574 22554
rect 7602 22526 8134 22554
rect 8162 22526 8167 22554
rect 16249 22526 16254 22554
rect 16282 22526 16702 22554
rect 16730 22526 16814 22554
rect 16842 22526 16847 22554
rect 16921 22526 16926 22554
rect 16954 22526 17262 22554
rect 17290 22526 17486 22554
rect 17514 22526 17519 22554
rect 2233 22330 2238 22358
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2370 22330 2375 22358
rect 17593 22330 17598 22358
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17730 22330 17735 22358
rect 13225 22078 13230 22106
rect 13258 22078 14014 22106
rect 14042 22078 14047 22106
rect 9913 21938 9918 21966
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 10050 21938 10055 21966
rect 7289 21854 7294 21882
rect 7322 21854 8134 21882
rect 8162 21854 8167 21882
rect 1857 21742 1862 21770
rect 1890 21742 2142 21770
rect 2170 21742 2175 21770
rect 9025 21742 9030 21770
rect 9058 21742 9310 21770
rect 9338 21742 9534 21770
rect 9562 21742 9567 21770
rect 12833 21742 12838 21770
rect 12866 21742 13118 21770
rect 13146 21742 13151 21770
rect 13505 21742 13510 21770
rect 13538 21742 14014 21770
rect 14042 21742 14047 21770
rect 16809 21742 16814 21770
rect 16842 21742 17094 21770
rect 17122 21742 18438 21770
rect 18466 21742 18471 21770
rect 2233 21546 2238 21574
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2370 21546 2375 21574
rect 17593 21546 17598 21574
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17730 21546 17735 21574
rect 9913 21154 9918 21182
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 10050 21154 10055 21182
rect 14793 21070 14798 21098
rect 14826 21070 16534 21098
rect 16562 21070 16567 21098
rect 14345 21014 14350 21042
rect 14378 21014 14574 21042
rect 14602 21014 16254 21042
rect 16282 21014 16758 21042
rect 16786 21014 16791 21042
rect 15913 20958 15918 20986
rect 15946 20958 17990 20986
rect 18018 20958 19446 20986
rect 19474 20958 19479 20986
rect 18545 20902 18550 20930
rect 18578 20902 19054 20930
rect 19082 20902 19087 20930
rect 2233 20762 2238 20790
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2370 20762 2375 20790
rect 17593 20762 17598 20790
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17730 20762 17735 20790
rect 19049 20566 19054 20594
rect 19082 20566 20510 20594
rect 20538 20566 20543 20594
rect 13449 20510 13454 20538
rect 13482 20510 14014 20538
rect 14042 20510 14047 20538
rect 19441 20510 19446 20538
rect 19474 20510 19950 20538
rect 19978 20510 21182 20538
rect 21210 20510 21215 20538
rect 9913 20370 9918 20398
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 10050 20370 10055 20398
rect 12945 20230 12950 20258
rect 12978 20230 14294 20258
rect 14322 20230 14327 20258
rect 24600 20202 25000 20216
rect 2529 20174 2534 20202
rect 2562 20174 4214 20202
rect 4242 20174 4247 20202
rect 14009 20174 14014 20202
rect 14042 20174 15358 20202
rect 15386 20174 15391 20202
rect 23529 20174 23534 20202
rect 23562 20174 25000 20202
rect 24600 20160 25000 20174
rect 2233 19978 2238 20006
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2370 19978 2375 20006
rect 17593 19978 17598 20006
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17730 19978 17735 20006
rect 20505 19782 20510 19810
rect 20538 19782 20958 19810
rect 20986 19782 20991 19810
rect 0 19698 400 19712
rect 0 19670 2086 19698
rect 2114 19670 2119 19698
rect 0 19656 400 19670
rect 9913 19586 9918 19614
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 10050 19586 10055 19614
rect 13449 19446 13454 19474
rect 13482 19446 14014 19474
rect 14042 19446 15470 19474
rect 15498 19446 15503 19474
rect 13113 19390 13118 19418
rect 13146 19390 14294 19418
rect 14322 19390 14798 19418
rect 14826 19390 14831 19418
rect 20953 19390 20958 19418
rect 20986 19390 22526 19418
rect 22554 19390 22559 19418
rect 21793 19334 21798 19362
rect 21826 19334 23478 19362
rect 23506 19334 23511 19362
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 5833 18494 5838 18522
rect 5866 18494 7294 18522
rect 7322 18494 7327 18522
rect 12833 18494 12838 18522
rect 12866 18494 12871 18522
rect 12838 18466 12866 18494
rect 12273 18438 12278 18466
rect 12306 18438 12866 18466
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 10929 18214 10934 18242
rect 10962 18214 12278 18242
rect 12306 18214 12311 18242
rect 17425 18214 17430 18242
rect 17458 18214 17990 18242
rect 18018 18214 18023 18242
rect 19049 18214 19054 18242
rect 19082 18214 20230 18242
rect 20258 18214 20263 18242
rect 17430 18186 17458 18214
rect 9025 18158 9030 18186
rect 9058 18158 9814 18186
rect 9842 18158 9847 18186
rect 15913 18158 15918 18186
rect 15946 18158 17458 18186
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2137 17822 2142 17850
rect 2170 17822 3598 17850
rect 3626 17822 3631 17850
rect 10033 17822 10038 17850
rect 10066 17822 11270 17850
rect 11298 17822 11303 17850
rect 17985 17822 17990 17850
rect 18018 17822 19334 17850
rect 19362 17822 19367 17850
rect 4153 17710 4158 17738
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 4186 17458 4214 17738
rect 6449 17654 6454 17682
rect 6482 17654 7014 17682
rect 7042 17654 7047 17682
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 24600 17514 25000 17528
rect 24033 17486 24038 17514
rect 24066 17486 25000 17514
rect 24600 17472 25000 17486
rect 2137 17430 2142 17458
rect 2170 17430 2478 17458
rect 2506 17430 3038 17458
rect 3066 17430 4382 17458
rect 4410 17430 4415 17458
rect 15913 17430 15918 17458
rect 15946 17430 16814 17458
rect 16842 17430 16847 17458
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 8129 17038 8134 17066
rect 8162 17038 9142 17066
rect 9170 17038 10318 17066
rect 10346 17038 10351 17066
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 4097 16646 4102 16674
rect 4130 16646 5278 16674
rect 5306 16646 5558 16674
rect 5586 16646 5591 16674
rect 22241 16646 22246 16674
rect 22274 16646 22750 16674
rect 22778 16646 22783 16674
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 6729 16254 6734 16282
rect 6762 16254 7014 16282
rect 7042 16254 8302 16282
rect 8330 16254 8335 16282
rect 16809 16254 16814 16282
rect 16842 16254 16982 16282
rect 17010 16254 17015 16282
rect 20785 16254 20790 16282
rect 20818 16254 20958 16282
rect 20986 16254 22246 16282
rect 22274 16254 22279 16282
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 2473 15918 2478 15946
rect 2506 15918 3038 15946
rect 3066 15918 3071 15946
rect 4545 15918 4550 15946
rect 4578 15918 5950 15946
rect 5978 15918 6230 15946
rect 6258 15918 6454 15946
rect 6482 15918 6487 15946
rect 5553 15862 5558 15890
rect 5586 15862 5838 15890
rect 5866 15862 5871 15890
rect 16921 15806 16926 15834
rect 16954 15806 17206 15834
rect 17234 15806 17430 15834
rect 17458 15806 17990 15834
rect 18018 15806 18023 15834
rect 19273 15806 19278 15834
rect 19306 15806 19950 15834
rect 19978 15806 21518 15834
rect 21546 15806 22694 15834
rect 22722 15806 23198 15834
rect 23226 15806 23422 15834
rect 23450 15806 23455 15834
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 5833 15470 5838 15498
rect 5866 15470 6118 15498
rect 6146 15470 6846 15498
rect 6874 15470 6879 15498
rect 8465 15470 8470 15498
rect 8498 15470 9030 15498
rect 9058 15470 9063 15498
rect 16809 15470 16814 15498
rect 16842 15470 17094 15498
rect 17122 15470 17127 15498
rect 17985 15470 17990 15498
rect 18018 15470 19278 15498
rect 19306 15470 19311 15498
rect 22689 15470 22694 15498
rect 22722 15470 22918 15498
rect 22946 15470 22951 15498
rect 0 15330 400 15344
rect 0 15302 1918 15330
rect 1946 15302 1951 15330
rect 0 15288 400 15302
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 2417 15134 2422 15162
rect 2450 15134 4494 15162
rect 4522 15134 4527 15162
rect 6505 15134 6510 15162
rect 6538 15134 6902 15162
rect 6930 15134 6935 15162
rect 22241 15078 22246 15106
rect 22274 15078 22750 15106
rect 22778 15078 22783 15106
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 24600 14826 25000 14840
rect 24033 14798 24038 14826
rect 24066 14798 25000 14826
rect 24600 14784 25000 14798
rect 1353 14686 1358 14714
rect 1386 14686 1862 14714
rect 1890 14686 3374 14714
rect 3402 14686 3407 14714
rect 21457 14686 21462 14714
rect 21490 14686 22750 14714
rect 22778 14686 22918 14714
rect 22946 14686 23198 14714
rect 23226 14686 23231 14714
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 19441 14406 19446 14434
rect 19474 14406 21014 14434
rect 21042 14406 21047 14434
rect 20169 14350 20174 14378
rect 20202 14350 22862 14378
rect 22890 14350 22895 14378
rect 19049 14294 19054 14322
rect 19082 14294 20230 14322
rect 20258 14294 20263 14322
rect 3817 14238 3822 14266
rect 3850 14238 5278 14266
rect 5306 14238 5558 14266
rect 5586 14238 5591 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2305 13902 2310 13930
rect 2338 13902 2534 13930
rect 2562 13902 2567 13930
rect 7009 13902 7014 13930
rect 7042 13902 8414 13930
rect 8442 13902 8862 13930
rect 8890 13902 8895 13930
rect 20953 13902 20958 13930
rect 20986 13902 22246 13930
rect 22274 13902 22279 13930
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 15465 13510 15470 13538
rect 15498 13510 17430 13538
rect 17458 13510 17463 13538
rect 20505 13510 20510 13538
rect 20538 13510 20958 13538
rect 20986 13510 20991 13538
rect 5497 13454 5502 13482
rect 5530 13454 6958 13482
rect 6986 13454 6991 13482
rect 17089 13454 17094 13482
rect 17122 13454 18270 13482
rect 18298 13454 18303 13482
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 4489 13118 4494 13146
rect 4522 13118 4998 13146
rect 5026 13118 5031 13146
rect 16977 13118 16982 13146
rect 17010 13118 17262 13146
rect 17290 13118 17486 13146
rect 17514 13118 17519 13146
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 19049 12726 19054 12754
rect 19082 12726 20510 12754
rect 20538 12726 20543 12754
rect 4993 12614 4998 12642
rect 5026 12614 5670 12642
rect 5698 12614 6062 12642
rect 6090 12614 6095 12642
rect 3369 12558 3374 12586
rect 3402 12558 3822 12586
rect 3850 12558 4494 12586
rect 4522 12558 4527 12586
rect 17761 12558 17766 12586
rect 17794 12558 19334 12586
rect 19362 12558 19367 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 2529 12334 2534 12362
rect 2562 12334 3766 12362
rect 3794 12334 3990 12362
rect 4018 12334 4023 12362
rect 8857 12334 8862 12362
rect 8890 12334 10598 12362
rect 10626 12334 10631 12362
rect 13113 12334 13118 12362
rect 13146 12334 14574 12362
rect 14602 12334 14607 12362
rect 18433 12334 18438 12362
rect 18466 12334 18550 12362
rect 18578 12334 19054 12362
rect 19082 12334 19087 12362
rect 21625 12334 21630 12362
rect 21658 12334 22134 12362
rect 22162 12334 22694 12362
rect 22722 12334 22727 12362
rect 13505 12278 13510 12306
rect 13538 12278 15134 12306
rect 15162 12278 15167 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 24600 12138 25000 12152
rect 23809 12110 23814 12138
rect 23842 12110 25000 12138
rect 24600 12096 25000 12110
rect 14793 11998 14798 12026
rect 14826 11998 16254 12026
rect 16282 11998 16287 12026
rect 1577 11942 1582 11970
rect 1610 11942 2142 11970
rect 2170 11942 3318 11970
rect 3346 11942 3598 11970
rect 3626 11942 3631 11970
rect 15465 11942 15470 11970
rect 15498 11942 15918 11970
rect 15946 11942 17430 11970
rect 17458 11942 17766 11970
rect 17794 11942 18718 11970
rect 18746 11942 19222 11970
rect 19250 11942 19446 11970
rect 19474 11942 19479 11970
rect 1913 11830 1918 11858
rect 1946 11830 17094 11858
rect 17122 11830 17127 11858
rect 8185 11774 8190 11802
rect 8218 11774 9422 11802
rect 9450 11774 9455 11802
rect 11489 11774 11494 11802
rect 11522 11774 12726 11802
rect 12754 11774 12950 11802
rect 12978 11774 13286 11802
rect 13314 11774 13319 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 17089 11550 17094 11578
rect 17122 11550 18438 11578
rect 18466 11550 18471 11578
rect 22577 11550 22582 11578
rect 22610 11550 24038 11578
rect 24066 11550 24071 11578
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 20897 11326 20902 11354
rect 20930 11326 21630 11354
rect 21658 11326 23814 11354
rect 23842 11326 23847 11354
rect 7289 11158 7294 11186
rect 7322 11158 8414 11186
rect 8442 11158 8862 11186
rect 8890 11158 8895 11186
rect 12553 11158 12558 11186
rect 12586 11158 13118 11186
rect 13146 11158 13151 11186
rect 14177 11158 14182 11186
rect 14210 11158 16814 11186
rect 16842 11158 16847 11186
rect 2473 11102 2478 11130
rect 2506 11102 2870 11130
rect 2898 11102 2903 11130
rect 0 10962 400 10976
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 0 10934 1694 10962
rect 1722 10934 1727 10962
rect 21793 10934 21798 10962
rect 0 10920 400 10934
rect 21826 10878 21854 10962
rect 21882 10878 22078 10906
rect 22106 10878 22111 10906
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 23753 10374 23758 10402
rect 23786 10374 24038 10402
rect 24066 10374 24071 10402
rect 4265 10318 4270 10346
rect 4298 10318 4606 10346
rect 4634 10318 5838 10346
rect 5866 10318 5871 10346
rect 20393 10318 20398 10346
rect 20426 10318 20902 10346
rect 20930 10318 22526 10346
rect 22554 10318 22559 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 1577 10094 1582 10122
rect 1610 10094 1862 10122
rect 1890 10094 1895 10122
rect 13449 10038 13454 10066
rect 13482 10038 14014 10066
rect 14042 10038 15358 10066
rect 15386 10038 15391 10066
rect 19441 10038 19446 10066
rect 19474 10038 20006 10066
rect 20034 10038 21182 10066
rect 21210 10038 21215 10066
rect 22577 10038 22582 10066
rect 22610 10038 22862 10066
rect 22890 10038 22895 10066
rect 1857 9982 1862 10010
rect 1890 9982 2142 10010
rect 2170 9982 2175 10010
rect 9809 9982 9814 10010
rect 9842 9982 10038 10010
rect 10066 9982 10990 10010
rect 11018 9982 11382 10010
rect 11410 9982 11415 10010
rect 12833 9982 12838 10010
rect 12866 9982 13118 10010
rect 13146 9982 14294 10010
rect 14322 9982 14574 10010
rect 14602 9982 14607 10010
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 12273 9590 12278 9618
rect 12306 9590 12558 9618
rect 12586 9590 12591 9618
rect 16921 9534 16926 9562
rect 16954 9534 17430 9562
rect 17458 9534 17990 9562
rect 18018 9534 18023 9562
rect 24600 9450 25000 9464
rect 21177 9422 21182 9450
rect 21210 9422 25000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 24600 9408 25000 9422
rect 11489 9310 11494 9338
rect 11522 9310 11718 9338
rect 11746 9310 13398 9338
rect 13426 9310 13431 9338
rect 11097 9254 11102 9282
rect 11130 9254 12278 9282
rect 12306 9254 12838 9282
rect 12866 9254 12871 9282
rect 22353 9198 22358 9226
rect 22386 9198 22582 9226
rect 22610 9198 22918 9226
rect 22946 9198 22951 9226
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 2529 8414 2534 8442
rect 2562 8414 3766 8442
rect 3794 8414 4494 8442
rect 4522 8414 4527 8442
rect 6449 8358 6454 8386
rect 6482 8358 6678 8386
rect 6706 8358 8134 8386
rect 8162 8358 8167 8386
rect 18545 8358 18550 8386
rect 18578 8358 19054 8386
rect 19082 8358 19087 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 8129 8022 8134 8050
rect 8162 8022 9422 8050
rect 9450 8022 9455 8050
rect 16529 8022 16534 8050
rect 16562 8022 17094 8050
rect 17122 8022 17127 8050
rect 19049 8022 19054 8050
rect 19082 8022 22806 8050
rect 22834 8022 22839 8050
rect 15465 7966 15470 7994
rect 15498 7966 17430 7994
rect 17458 7966 17766 7994
rect 17794 7966 17799 7994
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 9137 7630 9142 7658
rect 9170 7630 10318 7658
rect 10346 7630 10351 7658
rect 17089 7630 17094 7658
rect 17122 7630 18550 7658
rect 18578 7630 18583 7658
rect 2137 7574 2142 7602
rect 2170 7574 2175 7602
rect 4489 7574 4494 7602
rect 4522 7574 4998 7602
rect 5026 7574 5838 7602
rect 5866 7574 9590 7602
rect 9618 7574 10038 7602
rect 10066 7574 11494 7602
rect 11522 7574 11527 7602
rect 12553 7574 12558 7602
rect 12586 7574 13118 7602
rect 13146 7574 13151 7602
rect 14793 7574 14798 7602
rect 14826 7574 16534 7602
rect 16562 7574 16567 7602
rect 17481 7574 17486 7602
rect 17514 7574 17990 7602
rect 18018 7574 18718 7602
rect 18746 7574 18942 7602
rect 18970 7574 19222 7602
rect 19250 7574 19255 7602
rect 2142 7546 2170 7574
rect 2142 7518 3598 7546
rect 3626 7518 3631 7546
rect 20225 7518 20230 7546
rect 20258 7518 20790 7546
rect 20818 7518 20823 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 3593 7238 3598 7266
rect 3626 7238 3822 7266
rect 3850 7238 4886 7266
rect 4914 7238 4919 7266
rect 7233 7238 7238 7266
rect 7266 7238 8694 7266
rect 8722 7238 8727 7266
rect 18769 7238 18774 7266
rect 18802 7238 20230 7266
rect 20258 7238 20263 7266
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 18713 6846 18718 6874
rect 18746 6846 18942 6874
rect 18970 6846 19222 6874
rect 19250 6846 19255 6874
rect 24600 6762 25000 6776
rect 24033 6734 24038 6762
rect 24066 6734 25000 6762
rect 24600 6720 25000 6734
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 0 6594 400 6608
rect 0 6566 1022 6594
rect 1050 6566 1055 6594
rect 0 6552 400 6566
rect 1577 6454 1582 6482
rect 1610 6454 1918 6482
rect 1946 6454 1951 6482
rect 2473 6454 2478 6482
rect 2506 6454 2870 6482
rect 2898 6454 2903 6482
rect 6449 6454 6454 6482
rect 6482 6454 7014 6482
rect 7042 6454 7047 6482
rect 9529 6454 9534 6482
rect 9562 6454 9814 6482
rect 9842 6454 9847 6482
rect 12441 6454 12446 6482
rect 12474 6454 12950 6482
rect 12978 6454 13454 6482
rect 13482 6454 14014 6482
rect 14042 6454 14238 6482
rect 14266 6454 15358 6482
rect 15386 6454 15391 6482
rect 19441 6454 19446 6482
rect 19474 6454 20678 6482
rect 20706 6454 21014 6482
rect 21042 6454 21047 6482
rect 4153 6398 4158 6426
rect 4186 6398 5278 6426
rect 5306 6398 5838 6426
rect 5866 6398 5871 6426
rect 10425 6398 10430 6426
rect 10458 6398 10878 6426
rect 10906 6398 10911 6426
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2081 6118 2086 6146
rect 2114 6118 2814 6146
rect 2842 6118 3038 6146
rect 3066 6118 3071 6146
rect 9809 6118 9814 6146
rect 9842 6118 11550 6146
rect 11578 6118 11583 6146
rect 17201 6118 17206 6146
rect 17234 6118 18830 6146
rect 18858 6118 19222 6146
rect 19250 6118 19255 6146
rect 1185 6062 1190 6090
rect 1218 6062 1694 6090
rect 1722 6062 2534 6090
rect 2562 6062 2870 6090
rect 2898 6062 2903 6090
rect 5833 6062 5838 6090
rect 5866 6062 7574 6090
rect 7602 6062 7798 6090
rect 7826 6062 7831 6090
rect 10873 6062 10878 6090
rect 10906 6062 12446 6090
rect 12474 6062 12479 6090
rect 16809 6062 16814 6090
rect 16842 6062 18270 6090
rect 18298 6062 18662 6090
rect 18690 6062 18774 6090
rect 18802 6062 18807 6090
rect 8465 5894 8470 5922
rect 8498 5894 8974 5922
rect 9002 5894 9534 5922
rect 9562 5894 9567 5922
rect 15946 5894 17206 5922
rect 17234 5894 17239 5922
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 15913 5782 15918 5810
rect 15946 5782 15974 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 4993 5670 4998 5698
rect 5026 5670 5558 5698
rect 5586 5670 6118 5698
rect 6146 5670 6151 5698
rect 17425 5670 17430 5698
rect 17458 5670 17766 5698
rect 17794 5670 17799 5698
rect 18545 5670 18550 5698
rect 18578 5670 19054 5698
rect 19082 5670 20230 5698
rect 20258 5670 20263 5698
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 17761 5334 17766 5362
rect 17794 5334 18718 5362
rect 18746 5334 18942 5362
rect 18970 5334 19222 5362
rect 19250 5334 19255 5362
rect 2025 5278 2030 5306
rect 2058 5278 2814 5306
rect 2842 5278 3038 5306
rect 3066 5278 3318 5306
rect 3346 5278 3351 5306
rect 17089 5278 17094 5306
rect 17122 5278 18550 5306
rect 18578 5278 18583 5306
rect 7009 5110 7014 5138
rect 7042 5110 7518 5138
rect 7546 5110 8078 5138
rect 8106 5110 9478 5138
rect 9506 5110 9511 5138
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 6505 5054 6510 5082
rect 6538 5054 7742 5082
rect 7770 5054 8246 5082
rect 8274 5054 8279 5082
rect 14233 4998 14238 5026
rect 14266 4998 15470 5026
rect 15498 4998 15918 5026
rect 15946 4998 15951 5026
rect 2081 4886 2086 4914
rect 2114 4886 3318 4914
rect 3346 4886 3542 4914
rect 3570 4886 3575 4914
rect 11769 4886 11774 4914
rect 11802 4886 12054 4914
rect 12082 4886 12838 4914
rect 12866 4886 13118 4914
rect 13146 4886 13398 4914
rect 13426 4886 14574 4914
rect 14602 4886 14607 4914
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 1017 4494 1022 4522
rect 1050 4494 2534 4522
rect 2562 4494 2870 4522
rect 2898 4494 2903 4522
rect 10425 4494 10430 4522
rect 10458 4494 10878 4522
rect 10906 4494 12390 4522
rect 12418 4494 12423 4522
rect 13953 4494 13958 4522
rect 13986 4494 14238 4522
rect 14266 4494 14271 4522
rect 10033 4438 10038 4466
rect 10066 4438 11270 4466
rect 11298 4438 11303 4466
rect 6113 4382 6118 4410
rect 6146 4382 7518 4410
rect 7546 4382 7798 4410
rect 7826 4382 7831 4410
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 8465 4158 8470 4186
rect 8498 4158 10094 4186
rect 12329 4158 12334 4186
rect 12362 4158 12950 4186
rect 12978 4158 14126 4186
rect 14154 4158 15470 4186
rect 15498 4158 15918 4186
rect 15946 4158 17430 4186
rect 17458 4158 17463 4186
rect 10066 4130 10094 4158
rect 6449 4102 6454 4130
rect 6482 4102 7014 4130
rect 7042 4102 7047 4130
rect 7793 4102 7798 4130
rect 7826 4102 9254 4130
rect 9282 4102 9287 4130
rect 10066 4102 10374 4130
rect 10402 4102 10407 4130
rect 15073 4102 15078 4130
rect 15106 4102 16254 4130
rect 16282 4102 16287 4130
rect 24600 4074 25000 4088
rect 23809 4046 23814 4074
rect 23842 4046 25000 4074
rect 24600 4032 25000 4046
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 7009 3710 7014 3738
rect 7042 3710 7518 3738
rect 7546 3710 7551 3738
rect 10369 3710 10374 3738
rect 10402 3710 10878 3738
rect 10906 3710 12334 3738
rect 12362 3710 12367 3738
rect 14569 3710 14574 3738
rect 14602 3710 15078 3738
rect 15106 3710 15111 3738
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 7793 3374 7798 3402
rect 7826 3374 8246 3402
rect 8274 3374 8470 3402
rect 8498 3374 8503 3402
rect 9529 3318 9534 3346
rect 9562 3318 9814 3346
rect 9842 3318 9847 3346
rect 13113 3318 13118 3346
rect 13146 3318 13398 3346
rect 13426 3318 14574 3346
rect 14602 3318 14607 3346
rect 16249 3318 16254 3346
rect 16282 3318 16814 3346
rect 16842 3318 16847 3346
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 7737 2982 7742 3010
rect 7770 2982 8470 3010
rect 8498 2982 8503 3010
rect 7569 2926 7574 2954
rect 7602 2926 8078 2954
rect 8106 2926 8111 2954
rect 9809 2926 9814 2954
rect 9842 2926 10038 2954
rect 10066 2926 11550 2954
rect 11578 2926 11583 2954
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 8073 2590 8078 2618
rect 8106 2590 9422 2618
rect 9450 2590 9455 2618
rect 3761 2534 3766 2562
rect 3794 2534 5278 2562
rect 5306 2534 5838 2562
rect 5866 2534 5871 2562
rect 6225 2534 6230 2562
rect 6258 2534 7014 2562
rect 7042 2534 7047 2562
rect 8465 2534 8470 2562
rect 8498 2534 8974 2562
rect 9002 2534 10430 2562
rect 10458 2534 10766 2562
rect 10794 2534 10799 2562
rect 11545 2534 11550 2562
rect 11578 2534 13118 2562
rect 13146 2534 13151 2562
rect 14793 2534 14798 2562
rect 14826 2534 16254 2562
rect 16282 2534 16287 2562
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 0 2226 400 2240
rect 0 2198 910 2226
rect 938 2198 943 2226
rect 0 2184 400 2198
rect 9249 2142 9254 2170
rect 9282 2142 9814 2170
rect 9842 2142 10094 2170
rect 12441 2142 12446 2170
rect 12474 2142 12894 2170
rect 12922 2142 12927 2170
rect 10066 2058 10094 2142
rect 10066 2030 11102 2058
rect 11130 2030 14294 2058
rect 14322 2030 14518 2058
rect 14546 2030 14798 2058
rect 14826 2030 14831 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 2081 1750 2086 1778
rect 2114 1750 2870 1778
rect 2898 1750 2903 1778
rect 9417 1750 9422 1778
rect 9450 1750 10374 1778
rect 10402 1750 10407 1778
rect 12889 1750 12894 1778
rect 12922 1750 13846 1778
rect 13874 1750 15358 1778
rect 15386 1750 15391 1778
rect 3817 1694 3822 1722
rect 3850 1694 7574 1722
rect 7602 1694 9590 1722
rect 9618 1694 9814 1722
rect 9842 1694 9847 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
rect 24600 1386 25000 1400
rect 24033 1358 24038 1386
rect 24066 1358 25000 1386
rect 24600 1344 25000 1358
<< via3 >>
rect 2238 33306 2266 33334
rect 2290 33306 2318 33334
rect 2342 33306 2370 33334
rect 17598 33306 17626 33334
rect 17650 33306 17678 33334
rect 17702 33306 17730 33334
rect 9918 32914 9946 32942
rect 9970 32914 9998 32942
rect 10022 32914 10050 32942
rect 2238 32522 2266 32550
rect 2290 32522 2318 32550
rect 2342 32522 2370 32550
rect 17598 32522 17626 32550
rect 17650 32522 17678 32550
rect 17702 32522 17730 32550
rect 9918 32130 9946 32158
rect 9970 32130 9998 32158
rect 10022 32130 10050 32158
rect 2238 31738 2266 31766
rect 2290 31738 2318 31766
rect 2342 31738 2370 31766
rect 17598 31738 17626 31766
rect 17650 31738 17678 31766
rect 17702 31738 17730 31766
rect 9918 31346 9946 31374
rect 9970 31346 9998 31374
rect 10022 31346 10050 31374
rect 2238 30954 2266 30982
rect 2290 30954 2318 30982
rect 2342 30954 2370 30982
rect 17598 30954 17626 30982
rect 17650 30954 17678 30982
rect 17702 30954 17730 30982
rect 9918 30562 9946 30590
rect 9970 30562 9998 30590
rect 10022 30562 10050 30590
rect 2238 30170 2266 30198
rect 2290 30170 2318 30198
rect 2342 30170 2370 30198
rect 17598 30170 17626 30198
rect 17650 30170 17678 30198
rect 17702 30170 17730 30198
rect 9918 29778 9946 29806
rect 9970 29778 9998 29806
rect 10022 29778 10050 29806
rect 2238 29386 2266 29414
rect 2290 29386 2318 29414
rect 2342 29386 2370 29414
rect 17598 29386 17626 29414
rect 17650 29386 17678 29414
rect 17702 29386 17730 29414
rect 9918 28994 9946 29022
rect 9970 28994 9998 29022
rect 10022 28994 10050 29022
rect 2238 28602 2266 28630
rect 2290 28602 2318 28630
rect 2342 28602 2370 28630
rect 17598 28602 17626 28630
rect 17650 28602 17678 28630
rect 17702 28602 17730 28630
rect 9918 28210 9946 28238
rect 9970 28210 9998 28238
rect 10022 28210 10050 28238
rect 2238 27818 2266 27846
rect 2290 27818 2318 27846
rect 2342 27818 2370 27846
rect 17598 27818 17626 27846
rect 17650 27818 17678 27846
rect 17702 27818 17730 27846
rect 9918 27426 9946 27454
rect 9970 27426 9998 27454
rect 10022 27426 10050 27454
rect 2238 27034 2266 27062
rect 2290 27034 2318 27062
rect 2342 27034 2370 27062
rect 17598 27034 17626 27062
rect 17650 27034 17678 27062
rect 17702 27034 17730 27062
rect 9918 26642 9946 26670
rect 9970 26642 9998 26670
rect 10022 26642 10050 26670
rect 2238 26250 2266 26278
rect 2290 26250 2318 26278
rect 2342 26250 2370 26278
rect 17598 26250 17626 26278
rect 17650 26250 17678 26278
rect 17702 26250 17730 26278
rect 9918 25858 9946 25886
rect 9970 25858 9998 25886
rect 10022 25858 10050 25886
rect 2238 25466 2266 25494
rect 2290 25466 2318 25494
rect 2342 25466 2370 25494
rect 17598 25466 17626 25494
rect 17650 25466 17678 25494
rect 17702 25466 17730 25494
rect 9918 25074 9946 25102
rect 9970 25074 9998 25102
rect 10022 25074 10050 25102
rect 2238 24682 2266 24710
rect 2290 24682 2318 24710
rect 2342 24682 2370 24710
rect 17598 24682 17626 24710
rect 17650 24682 17678 24710
rect 17702 24682 17730 24710
rect 9918 24290 9946 24318
rect 9970 24290 9998 24318
rect 10022 24290 10050 24318
rect 2238 23898 2266 23926
rect 2290 23898 2318 23926
rect 2342 23898 2370 23926
rect 17598 23898 17626 23926
rect 17650 23898 17678 23926
rect 17702 23898 17730 23926
rect 4214 23590 4242 23618
rect 9918 23506 9946 23534
rect 9970 23506 9998 23534
rect 10022 23506 10050 23534
rect 2238 23114 2266 23142
rect 2290 23114 2318 23142
rect 2342 23114 2370 23142
rect 17598 23114 17626 23142
rect 17650 23114 17678 23142
rect 17702 23114 17730 23142
rect 4214 22918 4242 22946
rect 9918 22722 9946 22750
rect 9970 22722 9998 22750
rect 10022 22722 10050 22750
rect 2238 22330 2266 22358
rect 2290 22330 2318 22358
rect 2342 22330 2370 22358
rect 17598 22330 17626 22358
rect 17650 22330 17678 22358
rect 17702 22330 17730 22358
rect 9918 21938 9946 21966
rect 9970 21938 9998 21966
rect 10022 21938 10050 21966
rect 2238 21546 2266 21574
rect 2290 21546 2318 21574
rect 2342 21546 2370 21574
rect 17598 21546 17626 21574
rect 17650 21546 17678 21574
rect 17702 21546 17730 21574
rect 9918 21154 9946 21182
rect 9970 21154 9998 21182
rect 10022 21154 10050 21182
rect 2238 20762 2266 20790
rect 2290 20762 2318 20790
rect 2342 20762 2370 20790
rect 17598 20762 17626 20790
rect 17650 20762 17678 20790
rect 17702 20762 17730 20790
rect 9918 20370 9946 20398
rect 9970 20370 9998 20398
rect 10022 20370 10050 20398
rect 2238 19978 2266 20006
rect 2290 19978 2318 20006
rect 2342 19978 2370 20006
rect 17598 19978 17626 20006
rect 17650 19978 17678 20006
rect 17702 19978 17730 20006
rect 9918 19586 9946 19614
rect 9970 19586 9998 19614
rect 10022 19586 10050 19614
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 33334 2384 33350
rect 2224 33306 2238 33334
rect 2266 33306 2290 33334
rect 2318 33306 2342 33334
rect 2370 33306 2384 33334
rect 2224 32550 2384 33306
rect 2224 32522 2238 32550
rect 2266 32522 2290 32550
rect 2318 32522 2342 32550
rect 2370 32522 2384 32550
rect 2224 31766 2384 32522
rect 2224 31738 2238 31766
rect 2266 31738 2290 31766
rect 2318 31738 2342 31766
rect 2370 31738 2384 31766
rect 2224 30982 2384 31738
rect 2224 30954 2238 30982
rect 2266 30954 2290 30982
rect 2318 30954 2342 30982
rect 2370 30954 2384 30982
rect 2224 30198 2384 30954
rect 2224 30170 2238 30198
rect 2266 30170 2290 30198
rect 2318 30170 2342 30198
rect 2370 30170 2384 30198
rect 2224 29414 2384 30170
rect 2224 29386 2238 29414
rect 2266 29386 2290 29414
rect 2318 29386 2342 29414
rect 2370 29386 2384 29414
rect 2224 28630 2384 29386
rect 2224 28602 2238 28630
rect 2266 28602 2290 28630
rect 2318 28602 2342 28630
rect 2370 28602 2384 28630
rect 2224 27846 2384 28602
rect 2224 27818 2238 27846
rect 2266 27818 2290 27846
rect 2318 27818 2342 27846
rect 2370 27818 2384 27846
rect 2224 27062 2384 27818
rect 2224 27034 2238 27062
rect 2266 27034 2290 27062
rect 2318 27034 2342 27062
rect 2370 27034 2384 27062
rect 2224 26278 2384 27034
rect 2224 26250 2238 26278
rect 2266 26250 2290 26278
rect 2318 26250 2342 26278
rect 2370 26250 2384 26278
rect 2224 25494 2384 26250
rect 2224 25466 2238 25494
rect 2266 25466 2290 25494
rect 2318 25466 2342 25494
rect 2370 25466 2384 25494
rect 2224 24710 2384 25466
rect 2224 24682 2238 24710
rect 2266 24682 2290 24710
rect 2318 24682 2342 24710
rect 2370 24682 2384 24710
rect 2224 23926 2384 24682
rect 2224 23898 2238 23926
rect 2266 23898 2290 23926
rect 2318 23898 2342 23926
rect 2370 23898 2384 23926
rect 2224 23142 2384 23898
rect 9904 32942 10064 33350
rect 9904 32914 9918 32942
rect 9946 32914 9970 32942
rect 9998 32914 10022 32942
rect 10050 32914 10064 32942
rect 9904 32158 10064 32914
rect 9904 32130 9918 32158
rect 9946 32130 9970 32158
rect 9998 32130 10022 32158
rect 10050 32130 10064 32158
rect 9904 31374 10064 32130
rect 9904 31346 9918 31374
rect 9946 31346 9970 31374
rect 9998 31346 10022 31374
rect 10050 31346 10064 31374
rect 9904 30590 10064 31346
rect 9904 30562 9918 30590
rect 9946 30562 9970 30590
rect 9998 30562 10022 30590
rect 10050 30562 10064 30590
rect 9904 29806 10064 30562
rect 9904 29778 9918 29806
rect 9946 29778 9970 29806
rect 9998 29778 10022 29806
rect 10050 29778 10064 29806
rect 9904 29022 10064 29778
rect 9904 28994 9918 29022
rect 9946 28994 9970 29022
rect 9998 28994 10022 29022
rect 10050 28994 10064 29022
rect 9904 28238 10064 28994
rect 9904 28210 9918 28238
rect 9946 28210 9970 28238
rect 9998 28210 10022 28238
rect 10050 28210 10064 28238
rect 9904 27454 10064 28210
rect 9904 27426 9918 27454
rect 9946 27426 9970 27454
rect 9998 27426 10022 27454
rect 10050 27426 10064 27454
rect 9904 26670 10064 27426
rect 9904 26642 9918 26670
rect 9946 26642 9970 26670
rect 9998 26642 10022 26670
rect 10050 26642 10064 26670
rect 9904 25886 10064 26642
rect 9904 25858 9918 25886
rect 9946 25858 9970 25886
rect 9998 25858 10022 25886
rect 10050 25858 10064 25886
rect 9904 25102 10064 25858
rect 9904 25074 9918 25102
rect 9946 25074 9970 25102
rect 9998 25074 10022 25102
rect 10050 25074 10064 25102
rect 9904 24318 10064 25074
rect 9904 24290 9918 24318
rect 9946 24290 9970 24318
rect 9998 24290 10022 24318
rect 10050 24290 10064 24318
rect 2224 23114 2238 23142
rect 2266 23114 2290 23142
rect 2318 23114 2342 23142
rect 2370 23114 2384 23142
rect 2224 22358 2384 23114
rect 4214 23618 4242 23623
rect 4214 22946 4242 23590
rect 4214 22913 4242 22918
rect 9904 23534 10064 24290
rect 9904 23506 9918 23534
rect 9946 23506 9970 23534
rect 9998 23506 10022 23534
rect 10050 23506 10064 23534
rect 2224 22330 2238 22358
rect 2266 22330 2290 22358
rect 2318 22330 2342 22358
rect 2370 22330 2384 22358
rect 2224 21574 2384 22330
rect 2224 21546 2238 21574
rect 2266 21546 2290 21574
rect 2318 21546 2342 21574
rect 2370 21546 2384 21574
rect 2224 20790 2384 21546
rect 2224 20762 2238 20790
rect 2266 20762 2290 20790
rect 2318 20762 2342 20790
rect 2370 20762 2384 20790
rect 2224 20006 2384 20762
rect 2224 19978 2238 20006
rect 2266 19978 2290 20006
rect 2318 19978 2342 20006
rect 2370 19978 2384 20006
rect 2224 19222 2384 19978
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 22750 10064 23506
rect 9904 22722 9918 22750
rect 9946 22722 9970 22750
rect 9998 22722 10022 22750
rect 10050 22722 10064 22750
rect 9904 21966 10064 22722
rect 9904 21938 9918 21966
rect 9946 21938 9970 21966
rect 9998 21938 10022 21966
rect 10050 21938 10064 21966
rect 9904 21182 10064 21938
rect 9904 21154 9918 21182
rect 9946 21154 9970 21182
rect 9998 21154 10022 21182
rect 10050 21154 10064 21182
rect 9904 20398 10064 21154
rect 9904 20370 9918 20398
rect 9946 20370 9970 20398
rect 9998 20370 10022 20398
rect 10050 20370 10064 20398
rect 9904 19614 10064 20370
rect 9904 19586 9918 19614
rect 9946 19586 9970 19614
rect 9998 19586 10022 19614
rect 10050 19586 10064 19614
rect 9904 18830 10064 19586
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 33334 17744 33350
rect 17584 33306 17598 33334
rect 17626 33306 17650 33334
rect 17678 33306 17702 33334
rect 17730 33306 17744 33334
rect 17584 32550 17744 33306
rect 17584 32522 17598 32550
rect 17626 32522 17650 32550
rect 17678 32522 17702 32550
rect 17730 32522 17744 32550
rect 17584 31766 17744 32522
rect 17584 31738 17598 31766
rect 17626 31738 17650 31766
rect 17678 31738 17702 31766
rect 17730 31738 17744 31766
rect 17584 30982 17744 31738
rect 17584 30954 17598 30982
rect 17626 30954 17650 30982
rect 17678 30954 17702 30982
rect 17730 30954 17744 30982
rect 17584 30198 17744 30954
rect 17584 30170 17598 30198
rect 17626 30170 17650 30198
rect 17678 30170 17702 30198
rect 17730 30170 17744 30198
rect 17584 29414 17744 30170
rect 17584 29386 17598 29414
rect 17626 29386 17650 29414
rect 17678 29386 17702 29414
rect 17730 29386 17744 29414
rect 17584 28630 17744 29386
rect 17584 28602 17598 28630
rect 17626 28602 17650 28630
rect 17678 28602 17702 28630
rect 17730 28602 17744 28630
rect 17584 27846 17744 28602
rect 17584 27818 17598 27846
rect 17626 27818 17650 27846
rect 17678 27818 17702 27846
rect 17730 27818 17744 27846
rect 17584 27062 17744 27818
rect 17584 27034 17598 27062
rect 17626 27034 17650 27062
rect 17678 27034 17702 27062
rect 17730 27034 17744 27062
rect 17584 26278 17744 27034
rect 17584 26250 17598 26278
rect 17626 26250 17650 26278
rect 17678 26250 17702 26278
rect 17730 26250 17744 26278
rect 17584 25494 17744 26250
rect 17584 25466 17598 25494
rect 17626 25466 17650 25494
rect 17678 25466 17702 25494
rect 17730 25466 17744 25494
rect 17584 24710 17744 25466
rect 17584 24682 17598 24710
rect 17626 24682 17650 24710
rect 17678 24682 17702 24710
rect 17730 24682 17744 24710
rect 17584 23926 17744 24682
rect 17584 23898 17598 23926
rect 17626 23898 17650 23926
rect 17678 23898 17702 23926
rect 17730 23898 17744 23926
rect 17584 23142 17744 23898
rect 17584 23114 17598 23142
rect 17626 23114 17650 23142
rect 17678 23114 17702 23142
rect 17730 23114 17744 23142
rect 17584 22358 17744 23114
rect 17584 22330 17598 22358
rect 17626 22330 17650 22358
rect 17678 22330 17702 22358
rect 17730 22330 17744 22358
rect 17584 21574 17744 22330
rect 17584 21546 17598 21574
rect 17626 21546 17650 21574
rect 17678 21546 17702 21574
rect 17730 21546 17744 21574
rect 17584 20790 17744 21546
rect 17584 20762 17598 20790
rect 17626 20762 17650 20790
rect 17678 20762 17702 20790
rect 17730 20762 17744 20790
rect 17584 20006 17744 20762
rect 17584 19978 17598 20006
rect 17626 19978 17650 20006
rect 17678 19978 17702 20006
rect 17730 19978 17744 20006
rect 17584 19222 17744 19978
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 4144 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 6664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 6888 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136
timestamp 1667941163
transform 1 0 8288 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142
timestamp 1667941163
transform 1 0 8624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 10416 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_177
timestamp 1667941163
transform 1 0 10584 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1667941163
transform 1 0 12376 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1667941163
transform 1 0 12544 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_237
timestamp 1667941163
transform 1 0 13944 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_247
timestamp 1667941163
transform 1 0 14504 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 16296 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1667941163
transform 1 0 16464 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1667941163
transform 1 0 18256 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317
timestamp 1667941163
transform 1 0 18424 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1667941163
transform 1 0 20216 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_352
timestamp 1667941163
transform 1 0 20384 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1667941163
transform 1 0 22176 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_387
timestamp 1667941163
transform 1 0 22344 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1667941163
transform 1 0 24136 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_18
timestamp 1667941163
transform 1 0 1680 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_26
timestamp 1667941163
transform 1 0 2128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_30 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2352 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_32
timestamp 1667941163
transform 1 0 2464 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_57
timestamp 1667941163
transform 1 0 3864 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_65
timestamp 1667941163
transform 1 0 4312 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_69
timestamp 1667941163
transform 1 0 4536 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_105
timestamp 1667941163
transform 1 0 6552 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_109
timestamp 1667941163
transform 1 0 6776 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 6888 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_136
timestamp 1667941163
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_140
timestamp 1667941163
transform 1 0 8512 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_144
timestamp 1667941163
transform 1 0 8736 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_160
timestamp 1667941163
transform 1 0 9632 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_186
timestamp 1667941163
transform 1 0 11088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 12544 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1667941163
transform 1 0 12712 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_240
timestamp 1667941163
transform 1 0 14112 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_266
timestamp 1667941163
transform 1 0 15568 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_282
timestamp 1667941163
transform 1 0 16464 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 16688 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1667941163
transform 1 0 20272 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1667941163
transform 1 0 20496 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_357
timestamp 1667941163
transform 1 0 20664 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_389
timestamp 1667941163
transform 1 0 22456 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_405
timestamp 1667941163
transform 1 0 23352 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_413
timestamp 1667941163
transform 1 0 23800 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_417
timestamp 1667941163
transform 1 0 24024 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1667941163
transform 1 0 24136 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_27
timestamp 1667941163
transform 1 0 2184 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_69
timestamp 1667941163
transform 1 0 4536 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_77
timestamp 1667941163
transform 1 0 4984 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_108
timestamp 1667941163
transform 1 0 6720 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_124
timestamp 1667941163
transform 1 0 7616 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_150
timestamp 1667941163
transform 1 0 9072 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 10528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_179
timestamp 1667941163
transform 1 0 10696 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 11592 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_220
timestamp 1667941163
transform 1 0 12992 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_246
timestamp 1667941163
transform 1 0 14448 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1667941163
transform 1 0 14672 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_275
timestamp 1667941163
transform 1 0 16072 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_307
timestamp 1667941163
transform 1 0 17864 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_315
timestamp 1667941163
transform 1 0 18312 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1667941163
transform 1 0 18648 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1667941163
transform 1 0 22232 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1667941163
transform 1 0 22456 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1667941163
transform 1 0 22624 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_408
timestamp 1667941163
transform 1 0 23520 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_416
timestamp 1667941163
transform 1 0 23968 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_27
timestamp 1667941163
transform 1 0 2184 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_59
timestamp 1667941163
transform 1 0 3976 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_67
timestamp 1667941163
transform 1 0 4424 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_89
timestamp 1667941163
transform 1 0 5656 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_115
timestamp 1667941163
transform 1 0 7112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 8568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_144
timestamp 1667941163
transform 1 0 8736 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_160
timestamp 1667941163
transform 1 0 9632 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_186
timestamp 1667941163
transform 1 0 11088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1667941163
transform 1 0 12544 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1667941163
transform 1 0 12712 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_240
timestamp 1667941163
transform 1 0 14112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_266
timestamp 1667941163
transform 1 0 15568 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1667941163
transform 1 0 16464 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1667941163
transform 1 0 16688 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1667941163
transform 1 0 20272 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1667941163
transform 1 0 20496 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_357
timestamp 1667941163
transform 1 0 20664 0 -1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_389
timestamp 1667941163
transform 1 0 22456 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_405
timestamp 1667941163
transform 1 0 23352 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1667941163
transform 1 0 23800 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1667941163
transform 1 0 24024 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1667941163
transform 1 0 24136 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1667941163
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_108
timestamp 1667941163
transform 1 0 6720 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_124
timestamp 1667941163
transform 1 0 7616 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_150
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 10528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_179
timestamp 1667941163
transform 1 0 10696 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 11592 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_220
timestamp 1667941163
transform 1 0 12992 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1667941163
transform 1 0 14448 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1667941163
transform 1 0 14672 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_275
timestamp 1667941163
transform 1 0 16072 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_301
timestamp 1667941163
transform 1 0 17528 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_317
timestamp 1667941163
transform 1 0 18424 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1667941163
transform 1 0 18648 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1667941163
transform 1 0 22232 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1667941163
transform 1 0 22456 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_392
timestamp 1667941163
transform 1 0 22624 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_408
timestamp 1667941163
transform 1 0 23520 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_416
timestamp 1667941163
transform 1 0 23968 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_27
timestamp 1667941163
transform 1 0 2184 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_59
timestamp 1667941163
transform 1 0 3976 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_67
timestamp 1667941163
transform 1 0 4424 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_89
timestamp 1667941163
transform 1 0 5656 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_115
timestamp 1667941163
transform 1 0 7112 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 8568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_144
timestamp 1667941163
transform 1 0 8736 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_160
timestamp 1667941163
transform 1 0 9632 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_186
timestamp 1667941163
transform 1 0 11088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1667941163
transform 1 0 12544 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1667941163
transform 1 0 12712 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_240
timestamp 1667941163
transform 1 0 14112 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_266
timestamp 1667941163
transform 1 0 15568 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1667941163
transform 1 0 16464 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_286
timestamp 1667941163
transform 1 0 16688 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_311
timestamp 1667941163
transform 1 0 18088 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_343
timestamp 1667941163
transform 1 0 19880 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_351
timestamp 1667941163
transform 1 0 20328 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_357
timestamp 1667941163
transform 1 0 20664 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_389
timestamp 1667941163
transform 1 0 22456 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_405
timestamp 1667941163
transform 1 0 23352 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1667941163
transform 1 0 23800 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1667941163
transform 1 0 24024 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1667941163
transform 1 0 24136 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_27
timestamp 1667941163
transform 1 0 2184 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_69
timestamp 1667941163
transform 1 0 4536 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_77
timestamp 1667941163
transform 1 0 4984 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 6552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_108
timestamp 1667941163
transform 1 0 6720 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_124
timestamp 1667941163
transform 1 0 7616 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_150
timestamp 1667941163
transform 1 0 9072 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 10528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_179
timestamp 1667941163
transform 1 0 10696 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_195
timestamp 1667941163
transform 1 0 11592 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_221
timestamp 1667941163
transform 1 0 13048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1667941163
transform 1 0 14504 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_250
timestamp 1667941163
transform 1 0 14672 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_275
timestamp 1667941163
transform 1 0 16072 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_301
timestamp 1667941163
transform 1 0 17528 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_317
timestamp 1667941163
transform 1 0 18424 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1667941163
transform 1 0 18648 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1667941163
transform 1 0 22232 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1667941163
transform 1 0 22456 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_392
timestamp 1667941163
transform 1 0 22624 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_394
timestamp 1667941163
transform 1 0 22736 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1667941163
transform 1 0 24136 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1667941163
transform 1 0 784 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_27
timestamp 1667941163
transform 1 0 2184 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_53
timestamp 1667941163
transform 1 0 3640 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1667941163
transform 1 0 4536 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1667941163
transform 1 0 4760 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_89
timestamp 1667941163
transform 1 0 5656 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_115
timestamp 1667941163
transform 1 0 7112 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 8568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_144
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1667941163
transform 1 0 9632 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_186
timestamp 1667941163
transform 1 0 11088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1667941163
transform 1 0 12544 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_215
timestamp 1667941163
transform 1 0 12712 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_240
timestamp 1667941163
transform 1 0 14112 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_266
timestamp 1667941163
transform 1 0 15568 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_282
timestamp 1667941163
transform 1 0 16464 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_311
timestamp 1667941163
transform 1 0 18088 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_343
timestamp 1667941163
transform 1 0 19880 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_351
timestamp 1667941163
transform 1 0 20328 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_357
timestamp 1667941163
transform 1 0 20664 0 -1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_389
timestamp 1667941163
transform 1 0 22456 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_405
timestamp 1667941163
transform 1 0 23352 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_413
timestamp 1667941163
transform 1 0 23800 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1667941163
transform 1 0 24024 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1667941163
transform 1 0 24136 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1667941163
transform 1 0 784 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_27
timestamp 1667941163
transform 1 0 2184 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1667941163
transform 1 0 2744 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_62
timestamp 1667941163
transform 1 0 4144 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_94
timestamp 1667941163
transform 1 0 5936 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_102
timestamp 1667941163
transform 1 0 6384 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_108
timestamp 1667941163
transform 1 0 6720 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_124
timestamp 1667941163
transform 1 0 7616 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_150
timestamp 1667941163
transform 1 0 9072 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 10528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_179
timestamp 1667941163
transform 1 0 10696 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_195
timestamp 1667941163
transform 1 0 11592 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_221
timestamp 1667941163
transform 1 0 13048 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1667941163
transform 1 0 14504 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1667941163
transform 1 0 14672 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_275
timestamp 1667941163
transform 1 0 16072 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_301
timestamp 1667941163
transform 1 0 17528 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_317
timestamp 1667941163
transform 1 0 18424 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1667941163
transform 1 0 18648 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1667941163
transform 1 0 22232 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1667941163
transform 1 0 22456 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_392
timestamp 1667941163
transform 1 0 22624 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_408
timestamp 1667941163
transform 1 0 23520 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_416
timestamp 1667941163
transform 1 0 23968 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1667941163
transform 1 0 784 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_27
timestamp 1667941163
transform 1 0 2184 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_53
timestamp 1667941163
transform 1 0 3640 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_69
timestamp 1667941163
transform 1 0 4536 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_73
timestamp 1667941163
transform 1 0 4760 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_89
timestamp 1667941163
transform 1 0 5656 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_115
timestamp 1667941163
transform 1 0 7112 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 8568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_144
timestamp 1667941163
transform 1 0 8736 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_160
timestamp 1667941163
transform 1 0 9632 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_186
timestamp 1667941163
transform 1 0 11088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1667941163
transform 1 0 12544 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1667941163
transform 1 0 12712 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_240
timestamp 1667941163
transform 1 0 14112 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_266
timestamp 1667941163
transform 1 0 15568 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_282
timestamp 1667941163
transform 1 0 16464 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_286
timestamp 1667941163
transform 1 0 16688 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_311
timestamp 1667941163
transform 1 0 18088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_337
timestamp 1667941163
transform 1 0 19544 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_353
timestamp 1667941163
transform 1 0 20440 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_357
timestamp 1667941163
transform 1 0 20664 0 -1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_389
timestamp 1667941163
transform 1 0 22456 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1667941163
transform 1 0 23352 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1667941163
transform 1 0 23800 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1667941163
transform 1 0 24024 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1667941163
transform 1 0 24136 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1667941163
transform 1 0 784 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_27
timestamp 1667941163
transform 1 0 2184 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1667941163
transform 1 0 2744 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_62
timestamp 1667941163
transform 1 0 4144 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_78
timestamp 1667941163
transform 1 0 5040 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_80
timestamp 1667941163
transform 1 0 5152 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 6552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_108
timestamp 1667941163
transform 1 0 6720 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_124
timestamp 1667941163
transform 1 0 7616 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_150
timestamp 1667941163
transform 1 0 9072 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 10528 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_179
timestamp 1667941163
transform 1 0 10696 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_195
timestamp 1667941163
transform 1 0 11592 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_221
timestamp 1667941163
transform 1 0 13048 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1667941163
transform 1 0 14504 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1667941163
transform 1 0 14672 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_275
timestamp 1667941163
transform 1 0 16072 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_301
timestamp 1667941163
transform 1 0 17528 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_317
timestamp 1667941163
transform 1 0 18424 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1667941163
transform 1 0 18648 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_346
timestamp 1667941163
transform 1 0 20048 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_378
timestamp 1667941163
transform 1 0 21840 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_386
timestamp 1667941163
transform 1 0 22288 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1667941163
transform 1 0 22624 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1667941163
transform 1 0 23520 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1667941163
transform 1 0 23968 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1667941163
transform 1 0 784 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_27
timestamp 1667941163
transform 1 0 2184 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_53
timestamp 1667941163
transform 1 0 3640 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1667941163
transform 1 0 4536 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_73
timestamp 1667941163
transform 1 0 4760 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_89
timestamp 1667941163
transform 1 0 5656 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_115
timestamp 1667941163
transform 1 0 7112 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 8568 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_144
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_160
timestamp 1667941163
transform 1 0 9632 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_186
timestamp 1667941163
transform 1 0 11088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1667941163
transform 1 0 12544 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1667941163
transform 1 0 12712 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_240
timestamp 1667941163
transform 1 0 14112 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_266
timestamp 1667941163
transform 1 0 15568 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1667941163
transform 1 0 16464 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_286
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_311
timestamp 1667941163
transform 1 0 18088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_337
timestamp 1667941163
transform 1 0 19544 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_353
timestamp 1667941163
transform 1 0 20440 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_357
timestamp 1667941163
transform 1 0 20664 0 -1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_389
timestamp 1667941163
transform 1 0 22456 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_405
timestamp 1667941163
transform 1 0 23352 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_413
timestamp 1667941163
transform 1 0 23800 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_417
timestamp 1667941163
transform 1 0 24024 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1667941163
transform 1 0 24136 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_2
timestamp 1667941163
transform 1 0 784 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 2576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_37
timestamp 1667941163
transform 1 0 2744 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_53
timestamp 1667941163
transform 1 0 3640 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_79
timestamp 1667941163
transform 1 0 5096 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 6552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_108
timestamp 1667941163
transform 1 0 6720 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_124
timestamp 1667941163
transform 1 0 7616 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_150
timestamp 1667941163
transform 1 0 9072 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 10528 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_179
timestamp 1667941163
transform 1 0 10696 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_195
timestamp 1667941163
transform 1 0 11592 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_221
timestamp 1667941163
transform 1 0 13048 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1667941163
transform 1 0 14504 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1667941163
transform 1 0 14672 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_275
timestamp 1667941163
transform 1 0 16072 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_301
timestamp 1667941163
transform 1 0 17528 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_317
timestamp 1667941163
transform 1 0 18424 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1667941163
transform 1 0 18648 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_346
timestamp 1667941163
transform 1 0 20048 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_372
timestamp 1667941163
transform 1 0 21504 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_388
timestamp 1667941163
transform 1 0 22400 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_392
timestamp 1667941163
transform 1 0 22624 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_394
timestamp 1667941163
transform 1 0 22736 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_419
timestamp 1667941163
transform 1 0 24136 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1667941163
transform 1 0 784 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_18
timestamp 1667941163
transform 1 0 1680 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_44
timestamp 1667941163
transform 1 0 3136 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 4592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1667941163
transform 1 0 4760 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_98
timestamp 1667941163
transform 1 0 6160 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_106
timestamp 1667941163
transform 1 0 6608 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_134
timestamp 1667941163
transform 1 0 8176 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_144
timestamp 1667941163
transform 1 0 8736 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_160
timestamp 1667941163
transform 1 0 9632 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_186
timestamp 1667941163
transform 1 0 11088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 12544 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1667941163
transform 1 0 12712 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_240
timestamp 1667941163
transform 1 0 14112 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_266
timestamp 1667941163
transform 1 0 15568 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_282
timestamp 1667941163
transform 1 0 16464 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1667941163
transform 1 0 16688 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_311
timestamp 1667941163
transform 1 0 18088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_337
timestamp 1667941163
transform 1 0 19544 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_353
timestamp 1667941163
transform 1 0 20440 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_357
timestamp 1667941163
transform 1 0 20664 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_389
timestamp 1667941163
transform 1 0 22456 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_393
timestamp 1667941163
transform 1 0 22680 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1667941163
transform 1 0 24136 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1667941163
transform 1 0 784 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 2576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_37
timestamp 1667941163
transform 1 0 2744 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_45
timestamp 1667941163
transform 1 0 3192 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_70
timestamp 1667941163
transform 1 0 4592 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_96
timestamp 1667941163
transform 1 0 6048 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_104
timestamp 1667941163
transform 1 0 6496 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_108
timestamp 1667941163
transform 1 0 6720 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_110
timestamp 1667941163
transform 1 0 6832 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_135
timestamp 1667941163
transform 1 0 8232 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_161
timestamp 1667941163
transform 1 0 9688 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1667941163
transform 1 0 10696 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_204
timestamp 1667941163
transform 1 0 12096 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_230
timestamp 1667941163
transform 1 0 13552 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_246
timestamp 1667941163
transform 1 0 14448 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1667941163
transform 1 0 14672 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_275
timestamp 1667941163
transform 1 0 16072 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_301
timestamp 1667941163
transform 1 0 17528 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_317
timestamp 1667941163
transform 1 0 18424 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1667941163
transform 1 0 18648 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_346
timestamp 1667941163
transform 1 0 20048 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_372
timestamp 1667941163
transform 1 0 21504 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_388
timestamp 1667941163
transform 1 0 22400 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_392
timestamp 1667941163
transform 1 0 22624 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_394
timestamp 1667941163
transform 1 0 22736 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_419
timestamp 1667941163
transform 1 0 24136 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_2
timestamp 1667941163
transform 1 0 784 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_18
timestamp 1667941163
transform 1 0 1680 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_44
timestamp 1667941163
transform 1 0 3136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 4592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_73
timestamp 1667941163
transform 1 0 4760 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_98
timestamp 1667941163
transform 1 0 6160 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_106
timestamp 1667941163
transform 1 0 6608 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_110
timestamp 1667941163
transform 1 0 6832 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_135
timestamp 1667941163
transform 1 0 8232 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_139
timestamp 1667941163
transform 1 0 8456 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 8568 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_144
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 10136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_195
timestamp 1667941163
transform 1 0 11592 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_211
timestamp 1667941163
transform 1 0 12488 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_215
timestamp 1667941163
transform 1 0 12712 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_240
timestamp 1667941163
transform 1 0 14112 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_266
timestamp 1667941163
transform 1 0 15568 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_282
timestamp 1667941163
transform 1 0 16464 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_311
timestamp 1667941163
transform 1 0 18088 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_337
timestamp 1667941163
transform 1 0 19544 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_353
timestamp 1667941163
transform 1 0 20440 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_357
timestamp 1667941163
transform 1 0 20664 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_382
timestamp 1667941163
transform 1 0 22064 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_390
timestamp 1667941163
transform 1 0 22512 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_394
timestamp 1667941163
transform 1 0 22736 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1667941163
transform 1 0 24136 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_2
timestamp 1667941163
transform 1 0 784 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1667941163
transform 1 0 2576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_37
timestamp 1667941163
transform 1 0 2744 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_53
timestamp 1667941163
transform 1 0 3640 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_79
timestamp 1667941163
transform 1 0 5096 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1667941163
transform 1 0 6552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_108
timestamp 1667941163
transform 1 0 6720 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_110
timestamp 1667941163
transform 1 0 6832 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_135
timestamp 1667941163
transform 1 0 8232 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_161
timestamp 1667941163
transform 1 0 9688 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_179
timestamp 1667941163
transform 1 0 10696 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_204
timestamp 1667941163
transform 1 0 12096 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_230
timestamp 1667941163
transform 1 0 13552 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_246
timestamp 1667941163
transform 1 0 14448 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1667941163
transform 1 0 14672 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_275
timestamp 1667941163
transform 1 0 16072 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_301
timestamp 1667941163
transform 1 0 17528 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_317
timestamp 1667941163
transform 1 0 18424 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_321
timestamp 1667941163
transform 1 0 18648 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_346
timestamp 1667941163
transform 1 0 20048 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_372
timestamp 1667941163
transform 1 0 21504 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_388
timestamp 1667941163
transform 1 0 22400 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_392
timestamp 1667941163
transform 1 0 22624 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_394
timestamp 1667941163
transform 1 0 22736 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_419
timestamp 1667941163
transform 1 0 24136 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_2
timestamp 1667941163
transform 1 0 784 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_18
timestamp 1667941163
transform 1 0 1680 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_44
timestamp 1667941163
transform 1 0 3136 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1667941163
transform 1 0 4592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_73
timestamp 1667941163
transform 1 0 4760 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_81
timestamp 1667941163
transform 1 0 5208 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_83
timestamp 1667941163
transform 1 0 5320 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_108
timestamp 1667941163
transform 1 0 6720 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_134
timestamp 1667941163
transform 1 0 8176 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1667941163
transform 1 0 8736 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 10136 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_195
timestamp 1667941163
transform 1 0 11592 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_211
timestamp 1667941163
transform 1 0 12488 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1667941163
transform 1 0 12712 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_240
timestamp 1667941163
transform 1 0 14112 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_266
timestamp 1667941163
transform 1 0 15568 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_282
timestamp 1667941163
transform 1 0 16464 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1667941163
transform 1 0 16688 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_311
timestamp 1667941163
transform 1 0 18088 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_337
timestamp 1667941163
transform 1 0 19544 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_353
timestamp 1667941163
transform 1 0 20440 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_357
timestamp 1667941163
transform 1 0 20664 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_389
timestamp 1667941163
transform 1 0 22456 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 22680 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1667941163
transform 1 0 24136 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_2
timestamp 1667941163
transform 1 0 784 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1667941163
transform 1 0 2576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_37
timestamp 1667941163
transform 1 0 2744 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_53
timestamp 1667941163
transform 1 0 3640 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_79
timestamp 1667941163
transform 1 0 5096 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1667941163
transform 1 0 6552 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_108
timestamp 1667941163
transform 1 0 6720 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_134
timestamp 1667941163
transform 1 0 8176 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_160
timestamp 1667941163
transform 1 0 9632 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1667941163
transform 1 0 10528 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1667941163
transform 1 0 10696 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_204
timestamp 1667941163
transform 1 0 12096 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_230
timestamp 1667941163
transform 1 0 13552 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_246
timestamp 1667941163
transform 1 0 14448 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1667941163
transform 1 0 14672 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_275
timestamp 1667941163
transform 1 0 16072 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_301
timestamp 1667941163
transform 1 0 17528 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_317
timestamp 1667941163
transform 1 0 18424 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1667941163
transform 1 0 18648 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_346
timestamp 1667941163
transform 1 0 20048 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_378
timestamp 1667941163
transform 1 0 21840 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_386
timestamp 1667941163
transform 1 0 22288 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_392
timestamp 1667941163
transform 1 0 22624 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_394
timestamp 1667941163
transform 1 0 22736 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_419
timestamp 1667941163
transform 1 0 24136 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_2
timestamp 1667941163
transform 1 0 784 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_18
timestamp 1667941163
transform 1 0 1680 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_44
timestamp 1667941163
transform 1 0 3136 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1667941163
transform 1 0 4592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_73
timestamp 1667941163
transform 1 0 4760 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_81
timestamp 1667941163
transform 1 0 5208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_109
timestamp 1667941163
transform 1 0 6776 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_135
timestamp 1667941163
transform 1 0 8232 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_139
timestamp 1667941163
transform 1 0 8456 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1667941163
transform 1 0 8568 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_144
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 10136 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_195
timestamp 1667941163
transform 1 0 11592 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_211
timestamp 1667941163
transform 1 0 12488 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_215
timestamp 1667941163
transform 1 0 12712 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_240
timestamp 1667941163
transform 1 0 14112 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_266
timestamp 1667941163
transform 1 0 15568 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_282
timestamp 1667941163
transform 1 0 16464 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_286
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_311
timestamp 1667941163
transform 1 0 18088 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_337
timestamp 1667941163
transform 1 0 19544 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_353
timestamp 1667941163
transform 1 0 20440 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_357
timestamp 1667941163
transform 1 0 20664 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_365
timestamp 1667941163
transform 1 0 21112 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_393
timestamp 1667941163
transform 1 0 22680 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_419
timestamp 1667941163
transform 1 0 24136 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_2
timestamp 1667941163
transform 1 0 784 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1667941163
transform 1 0 2576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_37
timestamp 1667941163
transform 1 0 2744 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_53
timestamp 1667941163
transform 1 0 3640 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_79
timestamp 1667941163
transform 1 0 5096 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1667941163
transform 1 0 6552 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_108
timestamp 1667941163
transform 1 0 6720 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_134
timestamp 1667941163
transform 1 0 8176 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_160
timestamp 1667941163
transform 1 0 9632 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1667941163
transform 1 0 10528 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1667941163
transform 1 0 10696 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_204
timestamp 1667941163
transform 1 0 12096 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_230
timestamp 1667941163
transform 1 0 13552 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_246
timestamp 1667941163
transform 1 0 14448 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_250
timestamp 1667941163
transform 1 0 14672 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_275
timestamp 1667941163
transform 1 0 16072 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_301
timestamp 1667941163
transform 1 0 17528 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_317
timestamp 1667941163
transform 1 0 18424 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_321
timestamp 1667941163
transform 1 0 18648 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_353
timestamp 1667941163
transform 1 0 20440 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_361
timestamp 1667941163
transform 1 0 20888 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1667941163
transform 1 0 22456 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_392
timestamp 1667941163
transform 1 0 22624 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_394
timestamp 1667941163
transform 1 0 22736 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_419
timestamp 1667941163
transform 1 0 24136 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_2
timestamp 1667941163
transform 1 0 784 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_18
timestamp 1667941163
transform 1 0 1680 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_44
timestamp 1667941163
transform 1 0 3136 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1667941163
transform 1 0 4592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_73
timestamp 1667941163
transform 1 0 4760 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_81
timestamp 1667941163
transform 1 0 5208 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_109
timestamp 1667941163
transform 1 0 6776 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_135
timestamp 1667941163
transform 1 0 8232 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_139
timestamp 1667941163
transform 1 0 8456 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1667941163
transform 1 0 8568 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_144
timestamp 1667941163
transform 1 0 8736 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 10136 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_195
timestamp 1667941163
transform 1 0 11592 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_211
timestamp 1667941163
transform 1 0 12488 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1667941163
transform 1 0 12712 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_240
timestamp 1667941163
transform 1 0 14112 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_266
timestamp 1667941163
transform 1 0 15568 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_282
timestamp 1667941163
transform 1 0 16464 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1667941163
transform 1 0 16688 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_311
timestamp 1667941163
transform 1 0 18088 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_343
timestamp 1667941163
transform 1 0 19880 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_351
timestamp 1667941163
transform 1 0 20328 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_357
timestamp 1667941163
transform 1 0 20664 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_365
timestamp 1667941163
transform 1 0 21112 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 22680 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_419
timestamp 1667941163
transform 1 0 24136 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_2
timestamp 1667941163
transform 1 0 784 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1667941163
transform 1 0 2576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_37
timestamp 1667941163
transform 1 0 2744 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_45
timestamp 1667941163
transform 1 0 3192 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_47
timestamp 1667941163
transform 1 0 3304 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_72
timestamp 1667941163
transform 1 0 4704 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_98
timestamp 1667941163
transform 1 0 6160 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_108
timestamp 1667941163
transform 1 0 6720 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_110
timestamp 1667941163
transform 1 0 6832 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_135
timestamp 1667941163
transform 1 0 8232 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_161
timestamp 1667941163
transform 1 0 9688 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1667941163
transform 1 0 10696 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_204
timestamp 1667941163
transform 1 0 12096 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_230
timestamp 1667941163
transform 1 0 13552 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_246
timestamp 1667941163
transform 1 0 14448 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1667941163
transform 1 0 14672 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_275
timestamp 1667941163
transform 1 0 16072 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_301
timestamp 1667941163
transform 1 0 17528 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1667941163
transform 1 0 18424 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_321
timestamp 1667941163
transform 1 0 18648 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_337
timestamp 1667941163
transform 1 0 19544 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_363
timestamp 1667941163
transform 1 0 21000 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1667941163
transform 1 0 22456 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_392
timestamp 1667941163
transform 1 0 22624 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_394
timestamp 1667941163
transform 1 0 22736 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_419
timestamp 1667941163
transform 1 0 24136 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_2
timestamp 1667941163
transform 1 0 784 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_18
timestamp 1667941163
transform 1 0 1680 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_44
timestamp 1667941163
transform 1 0 3136 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1667941163
transform 1 0 4592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_73
timestamp 1667941163
transform 1 0 4760 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_98
timestamp 1667941163
transform 1 0 6160 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_106
timestamp 1667941163
transform 1 0 6608 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_110
timestamp 1667941163
transform 1 0 6832 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_135
timestamp 1667941163
transform 1 0 8232 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_139
timestamp 1667941163
transform 1 0 8456 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1667941163
transform 1 0 8568 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_144
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 10136 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_195
timestamp 1667941163
transform 1 0 11592 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_211
timestamp 1667941163
transform 1 0 12488 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_215
timestamp 1667941163
transform 1 0 12712 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_240
timestamp 1667941163
transform 1 0 14112 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_266
timestamp 1667941163
transform 1 0 15568 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_282
timestamp 1667941163
transform 1 0 16464 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_311
timestamp 1667941163
transform 1 0 18088 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_327
timestamp 1667941163
transform 1 0 18984 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_329
timestamp 1667941163
transform 1 0 19096 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1667941163
transform 1 0 20496 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_357
timestamp 1667941163
transform 1 0 20664 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_365
timestamp 1667941163
transform 1 0 21112 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_393
timestamp 1667941163
transform 1 0 22680 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_419
timestamp 1667941163
transform 1 0 24136 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_2
timestamp 1667941163
transform 1 0 784 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1667941163
transform 1 0 2576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_37
timestamp 1667941163
transform 1 0 2744 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_45
timestamp 1667941163
transform 1 0 3192 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_47
timestamp 1667941163
transform 1 0 3304 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_72
timestamp 1667941163
transform 1 0 4704 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_98
timestamp 1667941163
transform 1 0 6160 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_108
timestamp 1667941163
transform 1 0 6720 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_110
timestamp 1667941163
transform 1 0 6832 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_135
timestamp 1667941163
transform 1 0 8232 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_161
timestamp 1667941163
transform 1 0 9688 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_179
timestamp 1667941163
transform 1 0 10696 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_204
timestamp 1667941163
transform 1 0 12096 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_230
timestamp 1667941163
transform 1 0 13552 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_246
timestamp 1667941163
transform 1 0 14448 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_250
timestamp 1667941163
transform 1 0 14672 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_275
timestamp 1667941163
transform 1 0 16072 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_301
timestamp 1667941163
transform 1 0 17528 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_317
timestamp 1667941163
transform 1 0 18424 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_321
timestamp 1667941163
transform 1 0 18648 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_337
timestamp 1667941163
transform 1 0 19544 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_363
timestamp 1667941163
transform 1 0 21000 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1667941163
transform 1 0 22456 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_392
timestamp 1667941163
transform 1 0 22624 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_394
timestamp 1667941163
transform 1 0 22736 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_419
timestamp 1667941163
transform 1 0 24136 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_2
timestamp 1667941163
transform 1 0 784 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_18
timestamp 1667941163
transform 1 0 1680 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_44
timestamp 1667941163
transform 1 0 3136 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1667941163
transform 1 0 4592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1667941163
transform 1 0 4760 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_98
timestamp 1667941163
transform 1 0 6160 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_106
timestamp 1667941163
transform 1 0 6608 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 6832 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_136
timestamp 1667941163
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_140
timestamp 1667941163
transform 1 0 8512 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_144
timestamp 1667941163
transform 1 0 8736 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 10136 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_195
timestamp 1667941163
transform 1 0 11592 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_211
timestamp 1667941163
transform 1 0 12488 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_215
timestamp 1667941163
transform 1 0 12712 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_240
timestamp 1667941163
transform 1 0 14112 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_266
timestamp 1667941163
transform 1 0 15568 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_282
timestamp 1667941163
transform 1 0 16464 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1667941163
transform 1 0 16688 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_311
timestamp 1667941163
transform 1 0 18088 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_337
timestamp 1667941163
transform 1 0 19544 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_353
timestamp 1667941163
transform 1 0 20440 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_357
timestamp 1667941163
transform 1 0 20664 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_365
timestamp 1667941163
transform 1 0 21112 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 22680 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_419
timestamp 1667941163
transform 1 0 24136 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_2
timestamp 1667941163
transform 1 0 784 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1667941163
transform 1 0 2576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_37
timestamp 1667941163
transform 1 0 2744 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_65
timestamp 1667941163
transform 1 0 4312 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_91
timestamp 1667941163
transform 1 0 5768 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_99
timestamp 1667941163
transform 1 0 6216 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_103
timestamp 1667941163
transform 1 0 6440 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1667941163
transform 1 0 6552 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_108
timestamp 1667941163
transform 1 0 6720 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_136
timestamp 1667941163
transform 1 0 8288 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_162
timestamp 1667941163
transform 1 0 9744 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_170
timestamp 1667941163
transform 1 0 10192 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_174
timestamp 1667941163
transform 1 0 10416 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1667941163
transform 1 0 10528 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_179
timestamp 1667941163
transform 1 0 10696 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_204
timestamp 1667941163
transform 1 0 12096 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_230
timestamp 1667941163
transform 1 0 13552 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_246
timestamp 1667941163
transform 1 0 14448 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1667941163
transform 1 0 14672 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_275
timestamp 1667941163
transform 1 0 16072 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_301
timestamp 1667941163
transform 1 0 17528 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_317
timestamp 1667941163
transform 1 0 18424 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1667941163
transform 1 0 18648 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_346
timestamp 1667941163
transform 1 0 20048 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 20944 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_364
timestamp 1667941163
transform 1 0 21056 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1667941163
transform 1 0 22456 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_392
timestamp 1667941163
transform 1 0 22624 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_394
timestamp 1667941163
transform 1 0 22736 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_419
timestamp 1667941163
transform 1 0 24136 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_2
timestamp 1667941163
transform 1 0 784 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_18
timestamp 1667941163
transform 1 0 1680 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_44
timestamp 1667941163
transform 1 0 3136 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1667941163
transform 1 0 4592 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_73
timestamp 1667941163
transform 1 0 4760 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_81
timestamp 1667941163
transform 1 0 5208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_109
timestamp 1667941163
transform 1 0 6776 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_135
timestamp 1667941163
transform 1 0 8232 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_139
timestamp 1667941163
transform 1 0 8456 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1667941163
transform 1 0 8568 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_144
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 10136 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_195
timestamp 1667941163
transform 1 0 11592 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_211
timestamp 1667941163
transform 1 0 12488 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_215
timestamp 1667941163
transform 1 0 12712 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_240
timestamp 1667941163
transform 1 0 14112 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_266
timestamp 1667941163
transform 1 0 15568 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_282
timestamp 1667941163
transform 1 0 16464 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_311
timestamp 1667941163
transform 1 0 18088 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_337
timestamp 1667941163
transform 1 0 19544 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_353
timestamp 1667941163
transform 1 0 20440 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_357
timestamp 1667941163
transform 1 0 20664 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_365
timestamp 1667941163
transform 1 0 21112 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 22680 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1667941163
transform 1 0 24136 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_2
timestamp 1667941163
transform 1 0 784 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1667941163
transform 1 0 2576 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_37
timestamp 1667941163
transform 1 0 2744 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_53
timestamp 1667941163
transform 1 0 3640 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_79
timestamp 1667941163
transform 1 0 5096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1667941163
transform 1 0 6552 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_108
timestamp 1667941163
transform 1 0 6720 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_136
timestamp 1667941163
transform 1 0 8288 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_162
timestamp 1667941163
transform 1 0 9744 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_170
timestamp 1667941163
transform 1 0 10192 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_174
timestamp 1667941163
transform 1 0 10416 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1667941163
transform 1 0 10528 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_179
timestamp 1667941163
transform 1 0 10696 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_204
timestamp 1667941163
transform 1 0 12096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_230
timestamp 1667941163
transform 1 0 13552 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_246
timestamp 1667941163
transform 1 0 14448 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_250
timestamp 1667941163
transform 1 0 14672 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_275
timestamp 1667941163
transform 1 0 16072 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_301
timestamp 1667941163
transform 1 0 17528 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_317
timestamp 1667941163
transform 1 0 18424 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1667941163
transform 1 0 18648 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_346
timestamp 1667941163
transform 1 0 20048 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_372
timestamp 1667941163
transform 1 0 21504 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_388
timestamp 1667941163
transform 1 0 22400 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_392
timestamp 1667941163
transform 1 0 22624 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_394
timestamp 1667941163
transform 1 0 22736 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_419
timestamp 1667941163
transform 1 0 24136 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_2
timestamp 1667941163
transform 1 0 784 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_18
timestamp 1667941163
transform 1 0 1680 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_44
timestamp 1667941163
transform 1 0 3136 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1667941163
transform 1 0 4592 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_73
timestamp 1667941163
transform 1 0 4760 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_81
timestamp 1667941163
transform 1 0 5208 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_109
timestamp 1667941163
transform 1 0 6776 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_135
timestamp 1667941163
transform 1 0 8232 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_139
timestamp 1667941163
transform 1 0 8456 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1667941163
transform 1 0 8568 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_144
timestamp 1667941163
transform 1 0 8736 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 10136 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_195
timestamp 1667941163
transform 1 0 11592 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_211
timestamp 1667941163
transform 1 0 12488 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1667941163
transform 1 0 12712 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_240
timestamp 1667941163
transform 1 0 14112 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_266
timestamp 1667941163
transform 1 0 15568 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_282
timestamp 1667941163
transform 1 0 16464 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1667941163
transform 1 0 16688 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_311
timestamp 1667941163
transform 1 0 18088 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_337
timestamp 1667941163
transform 1 0 19544 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_353
timestamp 1667941163
transform 1 0 20440 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1667941163
transform 1 0 20664 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_382
timestamp 1667941163
transform 1 0 22064 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_390
timestamp 1667941163
transform 1 0 22512 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_394
timestamp 1667941163
transform 1 0 22736 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1667941163
transform 1 0 24136 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_2
timestamp 1667941163
transform 1 0 784 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1667941163
transform 1 0 2576 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_37
timestamp 1667941163
transform 1 0 2744 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_53
timestamp 1667941163
transform 1 0 3640 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_79
timestamp 1667941163
transform 1 0 5096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1667941163
transform 1 0 6552 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_108
timestamp 1667941163
transform 1 0 6720 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_136
timestamp 1667941163
transform 1 0 8288 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_162
timestamp 1667941163
transform 1 0 9744 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_170
timestamp 1667941163
transform 1 0 10192 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_174
timestamp 1667941163
transform 1 0 10416 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1667941163
transform 1 0 10528 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_179
timestamp 1667941163
transform 1 0 10696 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_204
timestamp 1667941163
transform 1 0 12096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_230
timestamp 1667941163
transform 1 0 13552 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_246
timestamp 1667941163
transform 1 0 14448 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_250
timestamp 1667941163
transform 1 0 14672 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_275
timestamp 1667941163
transform 1 0 16072 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_301
timestamp 1667941163
transform 1 0 17528 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_317
timestamp 1667941163
transform 1 0 18424 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1667941163
transform 1 0 18648 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_346
timestamp 1667941163
transform 1 0 20048 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_372
timestamp 1667941163
transform 1 0 21504 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_388
timestamp 1667941163
transform 1 0 22400 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_392
timestamp 1667941163
transform 1 0 22624 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_394
timestamp 1667941163
transform 1 0 22736 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_419
timestamp 1667941163
transform 1 0 24136 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_2
timestamp 1667941163
transform 1 0 784 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_18
timestamp 1667941163
transform 1 0 1680 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_44
timestamp 1667941163
transform 1 0 3136 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1667941163
transform 1 0 4592 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_73
timestamp 1667941163
transform 1 0 4760 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_81
timestamp 1667941163
transform 1 0 5208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_85
timestamp 1667941163
transform 1 0 5432 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 6832 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_136
timestamp 1667941163
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_140
timestamp 1667941163
transform 1 0 8512 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_144
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 10136 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_195
timestamp 1667941163
transform 1 0 11592 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_211
timestamp 1667941163
transform 1 0 12488 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1667941163
transform 1 0 12712 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_240
timestamp 1667941163
transform 1 0 14112 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_266
timestamp 1667941163
transform 1 0 15568 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_282
timestamp 1667941163
transform 1 0 16464 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_286
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_311
timestamp 1667941163
transform 1 0 18088 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_337
timestamp 1667941163
transform 1 0 19544 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_353
timestamp 1667941163
transform 1 0 20440 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1667941163
transform 1 0 20664 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_382
timestamp 1667941163
transform 1 0 22064 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_390
timestamp 1667941163
transform 1 0 22512 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_394
timestamp 1667941163
transform 1 0 22736 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_419
timestamp 1667941163
transform 1 0 24136 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_2
timestamp 1667941163
transform 1 0 784 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1667941163
transform 1 0 2576 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_37
timestamp 1667941163
transform 1 0 2744 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_53
timestamp 1667941163
transform 1 0 3640 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_79
timestamp 1667941163
transform 1 0 5096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1667941163
transform 1 0 6552 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_108
timestamp 1667941163
transform 1 0 6720 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_133
timestamp 1667941163
transform 1 0 8120 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_159
timestamp 1667941163
transform 1 0 9576 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_175
timestamp 1667941163
transform 1 0 10472 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_179
timestamp 1667941163
transform 1 0 10696 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_204
timestamp 1667941163
transform 1 0 12096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_230
timestamp 1667941163
transform 1 0 13552 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_246
timestamp 1667941163
transform 1 0 14448 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1667941163
transform 1 0 14672 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_275
timestamp 1667941163
transform 1 0 16072 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_301
timestamp 1667941163
transform 1 0 17528 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1667941163
transform 1 0 18424 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1667941163
transform 1 0 18648 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_346
timestamp 1667941163
transform 1 0 20048 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_372
timestamp 1667941163
transform 1 0 21504 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_388
timestamp 1667941163
transform 1 0 22400 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_392
timestamp 1667941163
transform 1 0 22624 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_394
timestamp 1667941163
transform 1 0 22736 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_419
timestamp 1667941163
transform 1 0 24136 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_2
timestamp 1667941163
transform 1 0 784 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_18
timestamp 1667941163
transform 1 0 1680 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_44
timestamp 1667941163
transform 1 0 3136 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1667941163
transform 1 0 4592 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_73
timestamp 1667941163
transform 1 0 4760 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_75
timestamp 1667941163
transform 1 0 4872 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_100
timestamp 1667941163
transform 1 0 6272 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_126
timestamp 1667941163
transform 1 0 7728 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_144
timestamp 1667941163
transform 1 0 8736 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_169
timestamp 1667941163
transform 1 0 10136 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_195
timestamp 1667941163
transform 1 0 11592 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_211
timestamp 1667941163
transform 1 0 12488 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1667941163
transform 1 0 12712 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_240
timestamp 1667941163
transform 1 0 14112 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_266
timestamp 1667941163
transform 1 0 15568 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_282
timestamp 1667941163
transform 1 0 16464 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1667941163
transform 1 0 16688 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_311
timestamp 1667941163
transform 1 0 18088 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_337
timestamp 1667941163
transform 1 0 19544 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_353
timestamp 1667941163
transform 1 0 20440 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1667941163
transform 1 0 20664 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_382
timestamp 1667941163
transform 1 0 22064 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_408
timestamp 1667941163
transform 1 0 23520 0 -1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_416
timestamp 1667941163
transform 1 0 23968 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_2
timestamp 1667941163
transform 1 0 784 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1667941163
transform 1 0 2576 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_37
timestamp 1667941163
transform 1 0 2744 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_53
timestamp 1667941163
transform 1 0 3640 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_79
timestamp 1667941163
transform 1 0 5096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1667941163
transform 1 0 6552 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_108
timestamp 1667941163
transform 1 0 6720 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_124
timestamp 1667941163
transform 1 0 7616 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_126
timestamp 1667941163
transform 1 0 7728 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_151
timestamp 1667941163
transform 1 0 9128 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_167
timestamp 1667941163
transform 1 0 10024 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_175
timestamp 1667941163
transform 1 0 10472 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_179
timestamp 1667941163
transform 1 0 10696 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_204
timestamp 1667941163
transform 1 0 12096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_230
timestamp 1667941163
transform 1 0 13552 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_246
timestamp 1667941163
transform 1 0 14448 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1667941163
transform 1 0 14672 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_275
timestamp 1667941163
transform 1 0 16072 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_301
timestamp 1667941163
transform 1 0 17528 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1667941163
transform 1 0 18424 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1667941163
transform 1 0 18648 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_346
timestamp 1667941163
transform 1 0 20048 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_372
timestamp 1667941163
transform 1 0 21504 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_388
timestamp 1667941163
transform 1 0 22400 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_392
timestamp 1667941163
transform 1 0 22624 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_417
timestamp 1667941163
transform 1 0 24024 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_419
timestamp 1667941163
transform 1 0 24136 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_2
timestamp 1667941163
transform 1 0 784 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_18
timestamp 1667941163
transform 1 0 1680 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_44
timestamp 1667941163
transform 1 0 3136 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1667941163
transform 1 0 4592 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_73
timestamp 1667941163
transform 1 0 4760 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_89
timestamp 1667941163
transform 1 0 5656 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_115
timestamp 1667941163
transform 1 0 7112 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1667941163
transform 1 0 8568 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_144
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 10136 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_195
timestamp 1667941163
transform 1 0 11592 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_211
timestamp 1667941163
transform 1 0 12488 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1667941163
transform 1 0 12712 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_240
timestamp 1667941163
transform 1 0 14112 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_266
timestamp 1667941163
transform 1 0 15568 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1667941163
transform 1 0 16464 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_286
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_311
timestamp 1667941163
transform 1 0 18088 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_337
timestamp 1667941163
transform 1 0 19544 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_353
timestamp 1667941163
transform 1 0 20440 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1667941163
transform 1 0 20664 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_382
timestamp 1667941163
transform 1 0 22064 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_408
timestamp 1667941163
transform 1 0 23520 0 -1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_416
timestamp 1667941163
transform 1 0 23968 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_2
timestamp 1667941163
transform 1 0 784 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1667941163
transform 1 0 2576 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_37
timestamp 1667941163
transform 1 0 2744 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_53
timestamp 1667941163
transform 1 0 3640 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_79
timestamp 1667941163
transform 1 0 5096 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1667941163
transform 1 0 6552 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_108
timestamp 1667941163
transform 1 0 6720 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_124
timestamp 1667941163
transform 1 0 7616 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_126
timestamp 1667941163
transform 1 0 7728 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_151
timestamp 1667941163
transform 1 0 9128 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_167
timestamp 1667941163
transform 1 0 10024 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_175
timestamp 1667941163
transform 1 0 10472 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_179
timestamp 1667941163
transform 1 0 10696 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_204
timestamp 1667941163
transform 1 0 12096 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_230
timestamp 1667941163
transform 1 0 13552 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_246
timestamp 1667941163
transform 1 0 14448 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_250
timestamp 1667941163
transform 1 0 14672 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_275
timestamp 1667941163
transform 1 0 16072 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_301
timestamp 1667941163
transform 1 0 17528 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_317
timestamp 1667941163
transform 1 0 18424 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1667941163
transform 1 0 18648 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_346
timestamp 1667941163
transform 1 0 20048 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_372
timestamp 1667941163
transform 1 0 21504 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_388
timestamp 1667941163
transform 1 0 22400 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_392
timestamp 1667941163
transform 1 0 22624 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_417
timestamp 1667941163
transform 1 0 24024 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_419
timestamp 1667941163
transform 1 0 24136 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_2
timestamp 1667941163
transform 1 0 784 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_18
timestamp 1667941163
transform 1 0 1680 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_44
timestamp 1667941163
transform 1 0 3136 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1667941163
transform 1 0 4592 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_73
timestamp 1667941163
transform 1 0 4760 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_89
timestamp 1667941163
transform 1 0 5656 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_115
timestamp 1667941163
transform 1 0 7112 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1667941163
transform 1 0 8568 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1667941163
transform 1 0 8736 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 10136 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_195
timestamp 1667941163
transform 1 0 11592 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_211
timestamp 1667941163
transform 1 0 12488 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_215
timestamp 1667941163
transform 1 0 12712 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_240
timestamp 1667941163
transform 1 0 14112 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_266
timestamp 1667941163
transform 1 0 15568 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1667941163
transform 1 0 16464 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1667941163
transform 1 0 16688 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_311
timestamp 1667941163
transform 1 0 18088 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_337
timestamp 1667941163
transform 1 0 19544 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_353
timestamp 1667941163
transform 1 0 20440 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_357
timestamp 1667941163
transform 1 0 20664 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_382
timestamp 1667941163
transform 1 0 22064 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_408
timestamp 1667941163
transform 1 0 23520 0 -1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_416
timestamp 1667941163
transform 1 0 23968 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_2
timestamp 1667941163
transform 1 0 784 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1667941163
transform 1 0 2576 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_37
timestamp 1667941163
transform 1 0 2744 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_53
timestamp 1667941163
transform 1 0 3640 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_79
timestamp 1667941163
transform 1 0 5096 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1667941163
transform 1 0 6552 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_108
timestamp 1667941163
transform 1 0 6720 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_124
timestamp 1667941163
transform 1 0 7616 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_126
timestamp 1667941163
transform 1 0 7728 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_151
timestamp 1667941163
transform 1 0 9128 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_167
timestamp 1667941163
transform 1 0 10024 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_175
timestamp 1667941163
transform 1 0 10472 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1667941163
transform 1 0 10696 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_204
timestamp 1667941163
transform 1 0 12096 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_230
timestamp 1667941163
transform 1 0 13552 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_246
timestamp 1667941163
transform 1 0 14448 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1667941163
transform 1 0 14672 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_275
timestamp 1667941163
transform 1 0 16072 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_301
timestamp 1667941163
transform 1 0 17528 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_317
timestamp 1667941163
transform 1 0 18424 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1667941163
transform 1 0 18648 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_346
timestamp 1667941163
transform 1 0 20048 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_372
timestamp 1667941163
transform 1 0 21504 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_388
timestamp 1667941163
transform 1 0 22400 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_392
timestamp 1667941163
transform 1 0 22624 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_417
timestamp 1667941163
transform 1 0 24024 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_419
timestamp 1667941163
transform 1 0 24136 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_2
timestamp 1667941163
transform 1 0 784 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_18
timestamp 1667941163
transform 1 0 1680 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_44
timestamp 1667941163
transform 1 0 3136 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1667941163
transform 1 0 4592 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_73
timestamp 1667941163
transform 1 0 4760 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_89
timestamp 1667941163
transform 1 0 5656 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_115
timestamp 1667941163
transform 1 0 7112 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1667941163
transform 1 0 8568 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1667941163
transform 1 0 8736 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 10136 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_195
timestamp 1667941163
transform 1 0 11592 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_211
timestamp 1667941163
transform 1 0 12488 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1667941163
transform 1 0 12712 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_240
timestamp 1667941163
transform 1 0 14112 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_266
timestamp 1667941163
transform 1 0 15568 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_282
timestamp 1667941163
transform 1 0 16464 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1667941163
transform 1 0 16688 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_311
timestamp 1667941163
transform 1 0 18088 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_337
timestamp 1667941163
transform 1 0 19544 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_353
timestamp 1667941163
transform 1 0 20440 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_357
timestamp 1667941163
transform 1 0 20664 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_382
timestamp 1667941163
transform 1 0 22064 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_408
timestamp 1667941163
transform 1 0 23520 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_416
timestamp 1667941163
transform 1 0 23968 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_2
timestamp 1667941163
transform 1 0 784 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1667941163
transform 1 0 2576 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_37
timestamp 1667941163
transform 1 0 2744 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_53
timestamp 1667941163
transform 1 0 3640 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_79
timestamp 1667941163
transform 1 0 5096 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1667941163
transform 1 0 6552 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_108
timestamp 1667941163
transform 1 0 6720 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_124
timestamp 1667941163
transform 1 0 7616 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_126
timestamp 1667941163
transform 1 0 7728 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_151
timestamp 1667941163
transform 1 0 9128 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_167
timestamp 1667941163
transform 1 0 10024 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_175
timestamp 1667941163
transform 1 0 10472 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1667941163
transform 1 0 10696 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_204
timestamp 1667941163
transform 1 0 12096 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_230
timestamp 1667941163
transform 1 0 13552 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_246
timestamp 1667941163
transform 1 0 14448 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1667941163
transform 1 0 14672 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_275
timestamp 1667941163
transform 1 0 16072 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_301
timestamp 1667941163
transform 1 0 17528 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_317
timestamp 1667941163
transform 1 0 18424 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1667941163
transform 1 0 18648 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_346
timestamp 1667941163
transform 1 0 20048 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_372
timestamp 1667941163
transform 1 0 21504 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_388
timestamp 1667941163
transform 1 0 22400 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_392
timestamp 1667941163
transform 1 0 22624 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_417
timestamp 1667941163
transform 1 0 24024 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_419
timestamp 1667941163
transform 1 0 24136 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_2
timestamp 1667941163
transform 1 0 784 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_18
timestamp 1667941163
transform 1 0 1680 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_44
timestamp 1667941163
transform 1 0 3136 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1667941163
transform 1 0 4592 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_73
timestamp 1667941163
transform 1 0 4760 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_89
timestamp 1667941163
transform 1 0 5656 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_115
timestamp 1667941163
transform 1 0 7112 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1667941163
transform 1 0 8568 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1667941163
transform 1 0 8736 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 10136 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_195
timestamp 1667941163
transform 1 0 11592 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_211
timestamp 1667941163
transform 1 0 12488 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1667941163
transform 1 0 12712 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_240
timestamp 1667941163
transform 1 0 14112 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_266
timestamp 1667941163
transform 1 0 15568 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_282
timestamp 1667941163
transform 1 0 16464 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1667941163
transform 1 0 16688 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_311
timestamp 1667941163
transform 1 0 18088 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_337
timestamp 1667941163
transform 1 0 19544 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_353
timestamp 1667941163
transform 1 0 20440 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1667941163
transform 1 0 20664 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_382
timestamp 1667941163
transform 1 0 22064 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_408
timestamp 1667941163
transform 1 0 23520 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_416
timestamp 1667941163
transform 1 0 23968 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_2
timestamp 1667941163
transform 1 0 784 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1667941163
transform 1 0 2576 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_37
timestamp 1667941163
transform 1 0 2744 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_53
timestamp 1667941163
transform 1 0 3640 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_79
timestamp 1667941163
transform 1 0 5096 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1667941163
transform 1 0 6552 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_108
timestamp 1667941163
transform 1 0 6720 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_124
timestamp 1667941163
transform 1 0 7616 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_126
timestamp 1667941163
transform 1 0 7728 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_151
timestamp 1667941163
transform 1 0 9128 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_167
timestamp 1667941163
transform 1 0 10024 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_175
timestamp 1667941163
transform 1 0 10472 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1667941163
transform 1 0 10696 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_204
timestamp 1667941163
transform 1 0 12096 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_230
timestamp 1667941163
transform 1 0 13552 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_246
timestamp 1667941163
transform 1 0 14448 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_250
timestamp 1667941163
transform 1 0 14672 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_275
timestamp 1667941163
transform 1 0 16072 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_301
timestamp 1667941163
transform 1 0 17528 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1667941163
transform 1 0 18424 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1667941163
transform 1 0 18648 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_346
timestamp 1667941163
transform 1 0 20048 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_372
timestamp 1667941163
transform 1 0 21504 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_388
timestamp 1667941163
transform 1 0 22400 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_392
timestamp 1667941163
transform 1 0 22624 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_417
timestamp 1667941163
transform 1 0 24024 0 1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1667941163
transform 1 0 24136 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_2
timestamp 1667941163
transform 1 0 784 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_18
timestamp 1667941163
transform 1 0 1680 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_44
timestamp 1667941163
transform 1 0 3136 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1667941163
transform 1 0 4592 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_73
timestamp 1667941163
transform 1 0 4760 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_89
timestamp 1667941163
transform 1 0 5656 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_115
timestamp 1667941163
transform 1 0 7112 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1667941163
transform 1 0 8568 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1667941163
transform 1 0 8736 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 10136 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_195
timestamp 1667941163
transform 1 0 11592 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_211
timestamp 1667941163
transform 1 0 12488 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_215
timestamp 1667941163
transform 1 0 12712 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_240
timestamp 1667941163
transform 1 0 14112 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_266
timestamp 1667941163
transform 1 0 15568 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_282
timestamp 1667941163
transform 1 0 16464 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_286
timestamp 1667941163
transform 1 0 16688 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_311
timestamp 1667941163
transform 1 0 18088 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_337
timestamp 1667941163
transform 1 0 19544 0 -1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_353
timestamp 1667941163
transform 1 0 20440 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_357
timestamp 1667941163
transform 1 0 20664 0 -1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_382
timestamp 1667941163
transform 1 0 22064 0 -1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_408
timestamp 1667941163
transform 1 0 23520 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_416
timestamp 1667941163
transform 1 0 23968 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_2
timestamp 1667941163
transform 1 0 784 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1667941163
transform 1 0 2576 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_37
timestamp 1667941163
transform 1 0 2744 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_53
timestamp 1667941163
transform 1 0 3640 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_79
timestamp 1667941163
transform 1 0 5096 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1667941163
transform 1 0 6552 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_108
timestamp 1667941163
transform 1 0 6720 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_124
timestamp 1667941163
transform 1 0 7616 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_126
timestamp 1667941163
transform 1 0 7728 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_151
timestamp 1667941163
transform 1 0 9128 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_167
timestamp 1667941163
transform 1 0 10024 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_175
timestamp 1667941163
transform 1 0 10472 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1667941163
transform 1 0 10696 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_204
timestamp 1667941163
transform 1 0 12096 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_230
timestamp 1667941163
transform 1 0 13552 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_246
timestamp 1667941163
transform 1 0 14448 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_250
timestamp 1667941163
transform 1 0 14672 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_275
timestamp 1667941163
transform 1 0 16072 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_301
timestamp 1667941163
transform 1 0 17528 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_317
timestamp 1667941163
transform 1 0 18424 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_321
timestamp 1667941163
transform 1 0 18648 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_346
timestamp 1667941163
transform 1 0 20048 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_372
timestamp 1667941163
transform 1 0 21504 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_388
timestamp 1667941163
transform 1 0 22400 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_392
timestamp 1667941163
transform 1 0 22624 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_417
timestamp 1667941163
transform 1 0 24024 0 1 18816
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_419
timestamp 1667941163
transform 1 0 24136 0 1 18816
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_2
timestamp 1667941163
transform 1 0 784 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_18
timestamp 1667941163
transform 1 0 1680 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_44
timestamp 1667941163
transform 1 0 3136 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1667941163
transform 1 0 4592 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_73
timestamp 1667941163
transform 1 0 4760 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_89
timestamp 1667941163
transform 1 0 5656 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_115
timestamp 1667941163
transform 1 0 7112 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1667941163
transform 1 0 8568 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1667941163
transform 1 0 8736 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 10136 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_195
timestamp 1667941163
transform 1 0 11592 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_211
timestamp 1667941163
transform 1 0 12488 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_215
timestamp 1667941163
transform 1 0 12712 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_240
timestamp 1667941163
transform 1 0 14112 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_266
timestamp 1667941163
transform 1 0 15568 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_282
timestamp 1667941163
transform 1 0 16464 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_286
timestamp 1667941163
transform 1 0 16688 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_311
timestamp 1667941163
transform 1 0 18088 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_337
timestamp 1667941163
transform 1 0 19544 0 -1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_353
timestamp 1667941163
transform 1 0 20440 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_357
timestamp 1667941163
transform 1 0 20664 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_382
timestamp 1667941163
transform 1 0 22064 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_408
timestamp 1667941163
transform 1 0 23520 0 -1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_410
timestamp 1667941163
transform 1 0 23632 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_419
timestamp 1667941163
transform 1 0 24136 0 -1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_2
timestamp 1667941163
transform 1 0 784 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1667941163
transform 1 0 2576 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_37
timestamp 1667941163
transform 1 0 2744 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_53
timestamp 1667941163
transform 1 0 3640 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_79
timestamp 1667941163
transform 1 0 5096 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1667941163
transform 1 0 6552 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_108
timestamp 1667941163
transform 1 0 6720 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_124
timestamp 1667941163
transform 1 0 7616 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_126
timestamp 1667941163
transform 1 0 7728 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_151
timestamp 1667941163
transform 1 0 9128 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_167
timestamp 1667941163
transform 1 0 10024 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_175
timestamp 1667941163
transform 1 0 10472 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1667941163
transform 1 0 10696 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_204
timestamp 1667941163
transform 1 0 12096 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_230
timestamp 1667941163
transform 1 0 13552 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_246
timestamp 1667941163
transform 1 0 14448 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_250
timestamp 1667941163
transform 1 0 14672 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_275
timestamp 1667941163
transform 1 0 16072 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_301
timestamp 1667941163
transform 1 0 17528 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_317
timestamp 1667941163
transform 1 0 18424 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_321
timestamp 1667941163
transform 1 0 18648 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_346
timestamp 1667941163
transform 1 0 20048 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_372
timestamp 1667941163
transform 1 0 21504 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_388
timestamp 1667941163
transform 1 0 22400 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1667941163
transform 1 0 22624 0 1 19600
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_408
timestamp 1667941163
transform 1 0 23520 0 1 19600
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_410
timestamp 1667941163
transform 1 0 23632 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_419
timestamp 1667941163
transform 1 0 24136 0 1 19600
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_2
timestamp 1667941163
transform 1 0 784 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_18
timestamp 1667941163
transform 1 0 1680 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_44
timestamp 1667941163
transform 1 0 3136 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1667941163
transform 1 0 4592 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_73
timestamp 1667941163
transform 1 0 4760 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_89
timestamp 1667941163
transform 1 0 5656 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_115
timestamp 1667941163
transform 1 0 7112 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1667941163
transform 1 0 8568 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_144
timestamp 1667941163
transform 1 0 8736 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 10136 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_195
timestamp 1667941163
transform 1 0 11592 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_211
timestamp 1667941163
transform 1 0 12488 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1667941163
transform 1 0 12712 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_240
timestamp 1667941163
transform 1 0 14112 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_266
timestamp 1667941163
transform 1 0 15568 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_282
timestamp 1667941163
transform 1 0 16464 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_286
timestamp 1667941163
transform 1 0 16688 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_311
timestamp 1667941163
transform 1 0 18088 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_337
timestamp 1667941163
transform 1 0 19544 0 -1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_353
timestamp 1667941163
transform 1 0 20440 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1667941163
transform 1 0 20664 0 -1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_382
timestamp 1667941163
transform 1 0 22064 0 -1 20384
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_414
timestamp 1667941163
transform 1 0 23856 0 -1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_418
timestamp 1667941163
transform 1 0 24080 0 -1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_2
timestamp 1667941163
transform 1 0 784 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1667941163
transform 1 0 2576 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_37
timestamp 1667941163
transform 1 0 2744 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_53
timestamp 1667941163
transform 1 0 3640 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_79
timestamp 1667941163
transform 1 0 5096 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1667941163
transform 1 0 6552 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_108
timestamp 1667941163
transform 1 0 6720 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_124
timestamp 1667941163
transform 1 0 7616 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_126
timestamp 1667941163
transform 1 0 7728 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_151
timestamp 1667941163
transform 1 0 9128 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_167
timestamp 1667941163
transform 1 0 10024 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_175
timestamp 1667941163
transform 1 0 10472 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1667941163
transform 1 0 10696 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_204
timestamp 1667941163
transform 1 0 12096 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_230
timestamp 1667941163
transform 1 0 13552 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_246
timestamp 1667941163
transform 1 0 14448 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_250
timestamp 1667941163
transform 1 0 14672 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_275
timestamp 1667941163
transform 1 0 16072 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_301
timestamp 1667941163
transform 1 0 17528 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_317
timestamp 1667941163
transform 1 0 18424 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_321
timestamp 1667941163
transform 1 0 18648 0 1 20384
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_346
timestamp 1667941163
transform 1 0 20048 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_372
timestamp 1667941163
transform 1 0 21504 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_388
timestamp 1667941163
transform 1 0 22400 0 1 20384
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_392
timestamp 1667941163
transform 1 0 22624 0 1 20384
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_408
timestamp 1667941163
transform 1 0 23520 0 1 20384
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_416
timestamp 1667941163
transform 1 0 23968 0 1 20384
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_2
timestamp 1667941163
transform 1 0 784 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_18
timestamp 1667941163
transform 1 0 1680 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_44
timestamp 1667941163
transform 1 0 3136 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1667941163
transform 1 0 4592 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_73
timestamp 1667941163
transform 1 0 4760 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_89
timestamp 1667941163
transform 1 0 5656 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_115
timestamp 1667941163
transform 1 0 7112 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1667941163
transform 1 0 8568 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1667941163
transform 1 0 8736 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 10136 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_195
timestamp 1667941163
transform 1 0 11592 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_211
timestamp 1667941163
transform 1 0 12488 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1667941163
transform 1 0 12712 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_240
timestamp 1667941163
transform 1 0 14112 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_266
timestamp 1667941163
transform 1 0 15568 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_282
timestamp 1667941163
transform 1 0 16464 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_286
timestamp 1667941163
transform 1 0 16688 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_311
timestamp 1667941163
transform 1 0 18088 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_337
timestamp 1667941163
transform 1 0 19544 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_353
timestamp 1667941163
transform 1 0 20440 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1667941163
transform 1 0 20664 0 -1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1667941163
transform 1 0 22456 0 -1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1667941163
transform 1 0 23352 0 -1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1667941163
transform 1 0 23800 0 -1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1667941163
transform 1 0 24024 0 -1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_419
timestamp 1667941163
transform 1 0 24136 0 -1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_2
timestamp 1667941163
transform 1 0 784 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1667941163
transform 1 0 2576 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_37
timestamp 1667941163
transform 1 0 2744 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_53
timestamp 1667941163
transform 1 0 3640 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_79
timestamp 1667941163
transform 1 0 5096 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1667941163
transform 1 0 6552 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_108
timestamp 1667941163
transform 1 0 6720 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_124
timestamp 1667941163
transform 1 0 7616 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_126
timestamp 1667941163
transform 1 0 7728 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_151
timestamp 1667941163
transform 1 0 9128 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_167
timestamp 1667941163
transform 1 0 10024 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_175
timestamp 1667941163
transform 1 0 10472 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_179
timestamp 1667941163
transform 1 0 10696 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_204
timestamp 1667941163
transform 1 0 12096 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_230
timestamp 1667941163
transform 1 0 13552 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_246
timestamp 1667941163
transform 1 0 14448 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_250
timestamp 1667941163
transform 1 0 14672 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_275
timestamp 1667941163
transform 1 0 16072 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_301
timestamp 1667941163
transform 1 0 17528 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_317
timestamp 1667941163
transform 1 0 18424 0 1 21168
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_321
timestamp 1667941163
transform 1 0 18648 0 1 21168
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_346
timestamp 1667941163
transform 1 0 20048 0 1 21168
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_378
timestamp 1667941163
transform 1 0 21840 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_386
timestamp 1667941163
transform 1 0 22288 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_392
timestamp 1667941163
transform 1 0 22624 0 1 21168
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_408
timestamp 1667941163
transform 1 0 23520 0 1 21168
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_416
timestamp 1667941163
transform 1 0 23968 0 1 21168
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_2
timestamp 1667941163
transform 1 0 784 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_18
timestamp 1667941163
transform 1 0 1680 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_44
timestamp 1667941163
transform 1 0 3136 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1667941163
transform 1 0 4592 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_73
timestamp 1667941163
transform 1 0 4760 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_89
timestamp 1667941163
transform 1 0 5656 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_115
timestamp 1667941163
transform 1 0 7112 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1667941163
transform 1 0 8568 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1667941163
transform 1 0 8736 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 10136 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_195
timestamp 1667941163
transform 1 0 11592 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_211
timestamp 1667941163
transform 1 0 12488 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_215
timestamp 1667941163
transform 1 0 12712 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_240
timestamp 1667941163
transform 1 0 14112 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_266
timestamp 1667941163
transform 1 0 15568 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_282
timestamp 1667941163
transform 1 0 16464 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_286
timestamp 1667941163
transform 1 0 16688 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_311
timestamp 1667941163
transform 1 0 18088 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_337
timestamp 1667941163
transform 1 0 19544 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_353
timestamp 1667941163
transform 1 0 20440 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1667941163
transform 1 0 20664 0 -1 21952
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1667941163
transform 1 0 22456 0 -1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1667941163
transform 1 0 23352 0 -1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1667941163
transform 1 0 23800 0 -1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1667941163
transform 1 0 24024 0 -1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1667941163
transform 1 0 24136 0 -1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_2
timestamp 1667941163
transform 1 0 784 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1667941163
transform 1 0 2576 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_37
timestamp 1667941163
transform 1 0 2744 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_53
timestamp 1667941163
transform 1 0 3640 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_79
timestamp 1667941163
transform 1 0 5096 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1667941163
transform 1 0 6552 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_108
timestamp 1667941163
transform 1 0 6720 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_124
timestamp 1667941163
transform 1 0 7616 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_126
timestamp 1667941163
transform 1 0 7728 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_151
timestamp 1667941163
transform 1 0 9128 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_167
timestamp 1667941163
transform 1 0 10024 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_175
timestamp 1667941163
transform 1 0 10472 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_179
timestamp 1667941163
transform 1 0 10696 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_204
timestamp 1667941163
transform 1 0 12096 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_230
timestamp 1667941163
transform 1 0 13552 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_246
timestamp 1667941163
transform 1 0 14448 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1667941163
transform 1 0 14672 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_275
timestamp 1667941163
transform 1 0 16072 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_301
timestamp 1667941163
transform 1 0 17528 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_317
timestamp 1667941163
transform 1 0 18424 0 1 21952
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1667941163
transform 1 0 18648 0 1 21952
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1667941163
transform 1 0 22232 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1667941163
transform 1 0 22456 0 1 21952
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_392
timestamp 1667941163
transform 1 0 22624 0 1 21952
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_408
timestamp 1667941163
transform 1 0 23520 0 1 21952
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_416
timestamp 1667941163
transform 1 0 23968 0 1 21952
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_2
timestamp 1667941163
transform 1 0 784 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_18
timestamp 1667941163
transform 1 0 1680 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_44
timestamp 1667941163
transform 1 0 3136 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1667941163
transform 1 0 4592 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_73
timestamp 1667941163
transform 1 0 4760 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_89
timestamp 1667941163
transform 1 0 5656 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_115
timestamp 1667941163
transform 1 0 7112 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1667941163
transform 1 0 8568 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1667941163
transform 1 0 8736 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_169
timestamp 1667941163
transform 1 0 10136 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_195
timestamp 1667941163
transform 1 0 11592 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_211
timestamp 1667941163
transform 1 0 12488 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1667941163
transform 1 0 12712 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_240
timestamp 1667941163
transform 1 0 14112 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_266
timestamp 1667941163
transform 1 0 15568 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_282
timestamp 1667941163
transform 1 0 16464 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_286
timestamp 1667941163
transform 1 0 16688 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_311
timestamp 1667941163
transform 1 0 18088 0 -1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_343
timestamp 1667941163
transform 1 0 19880 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_351
timestamp 1667941163
transform 1 0 20328 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_357
timestamp 1667941163
transform 1 0 20664 0 -1 22736
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_389
timestamp 1667941163
transform 1 0 22456 0 -1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_405
timestamp 1667941163
transform 1 0 23352 0 -1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_409
timestamp 1667941163
transform 1 0 23576 0 -1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1667941163
transform 1 0 24136 0 -1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_2
timestamp 1667941163
transform 1 0 784 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1667941163
transform 1 0 2576 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_37
timestamp 1667941163
transform 1 0 2744 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_53
timestamp 1667941163
transform 1 0 3640 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_79
timestamp 1667941163
transform 1 0 5096 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1667941163
transform 1 0 6552 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_108
timestamp 1667941163
transform 1 0 6720 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_124
timestamp 1667941163
transform 1 0 7616 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_126
timestamp 1667941163
transform 1 0 7728 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_151
timestamp 1667941163
transform 1 0 9128 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_167
timestamp 1667941163
transform 1 0 10024 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_175
timestamp 1667941163
transform 1 0 10472 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_179
timestamp 1667941163
transform 1 0 10696 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_204
timestamp 1667941163
transform 1 0 12096 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_230
timestamp 1667941163
transform 1 0 13552 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_246
timestamp 1667941163
transform 1 0 14448 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_250
timestamp 1667941163
transform 1 0 14672 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_275
timestamp 1667941163
transform 1 0 16072 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_301
timestamp 1667941163
transform 1 0 17528 0 1 22736
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_317
timestamp 1667941163
transform 1 0 18424 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1667941163
transform 1 0 18648 0 1 22736
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1667941163
transform 1 0 22232 0 1 22736
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1667941163
transform 1 0 22456 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_392
timestamp 1667941163
transform 1 0 22624 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_400
timestamp 1667941163
transform 1 0 23072 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_409
timestamp 1667941163
transform 1 0 23576 0 1 22736
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_419
timestamp 1667941163
transform 1 0 24136 0 1 22736
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_2
timestamp 1667941163
transform 1 0 784 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_18
timestamp 1667941163
transform 1 0 1680 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_44
timestamp 1667941163
transform 1 0 3136 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1667941163
transform 1 0 4592 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_73
timestamp 1667941163
transform 1 0 4760 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_75
timestamp 1667941163
transform 1 0 4872 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_100
timestamp 1667941163
transform 1 0 6272 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_126
timestamp 1667941163
transform 1 0 7728 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_144
timestamp 1667941163
transform 1 0 8736 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 10136 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_195
timestamp 1667941163
transform 1 0 11592 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_211
timestamp 1667941163
transform 1 0 12488 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_215
timestamp 1667941163
transform 1 0 12712 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_240
timestamp 1667941163
transform 1 0 14112 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_266
timestamp 1667941163
transform 1 0 15568 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_282
timestamp 1667941163
transform 1 0 16464 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1667941163
transform 1 0 16688 0 -1 23520
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1667941163
transform 1 0 20272 0 -1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1667941163
transform 1 0 20496 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_357
timestamp 1667941163
transform 1 0 20664 0 -1 23520
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_389
timestamp 1667941163
transform 1 0 22456 0 -1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_405
timestamp 1667941163
transform 1 0 23352 0 -1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_409
timestamp 1667941163
transform 1 0 23576 0 -1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_419
timestamp 1667941163
transform 1 0 24136 0 -1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_2
timestamp 1667941163
transform 1 0 784 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1667941163
transform 1 0 2576 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_37
timestamp 1667941163
transform 1 0 2744 0 1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_53
timestamp 1667941163
transform 1 0 3640 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_79
timestamp 1667941163
transform 1 0 5096 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1667941163
transform 1 0 6552 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_108
timestamp 1667941163
transform 1 0 6720 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_133
timestamp 1667941163
transform 1 0 8120 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_159
timestamp 1667941163
transform 1 0 9576 0 1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_175
timestamp 1667941163
transform 1 0 10472 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_179
timestamp 1667941163
transform 1 0 10696 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_204
timestamp 1667941163
transform 1 0 12096 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_230
timestamp 1667941163
transform 1 0 13552 0 1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_246
timestamp 1667941163
transform 1 0 14448 0 1 23520
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_250
timestamp 1667941163
transform 1 0 14672 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_275
timestamp 1667941163
transform 1 0 16072 0 1 23520
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_307
timestamp 1667941163
transform 1 0 17864 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_315
timestamp 1667941163
transform 1 0 18312 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1667941163
transform 1 0 18648 0 1 23520
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1667941163
transform 1 0 22232 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1667941163
transform 1 0 22456 0 1 23520
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_392
timestamp 1667941163
transform 1 0 22624 0 1 23520
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_408
timestamp 1667941163
transform 1 0 23520 0 1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_416
timestamp 1667941163
transform 1 0 23968 0 1 23520
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_2
timestamp 1667941163
transform 1 0 784 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_18
timestamp 1667941163
transform 1 0 1680 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_44
timestamp 1667941163
transform 1 0 3136 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1667941163
transform 1 0 4592 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_73
timestamp 1667941163
transform 1 0 4760 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_75
timestamp 1667941163
transform 1 0 4872 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_100
timestamp 1667941163
transform 1 0 6272 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_126
timestamp 1667941163
transform 1 0 7728 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_144
timestamp 1667941163
transform 1 0 8736 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 10136 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_195
timestamp 1667941163
transform 1 0 11592 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_211
timestamp 1667941163
transform 1 0 12488 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_215
timestamp 1667941163
transform 1 0 12712 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_240
timestamp 1667941163
transform 1 0 14112 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_266
timestamp 1667941163
transform 1 0 15568 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_282
timestamp 1667941163
transform 1 0 16464 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1667941163
transform 1 0 16688 0 -1 24304
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1667941163
transform 1 0 20272 0 -1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1667941163
transform 1 0 20496 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_357
timestamp 1667941163
transform 1 0 20664 0 -1 24304
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_389
timestamp 1667941163
transform 1 0 22456 0 -1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_405
timestamp 1667941163
transform 1 0 23352 0 -1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_409
timestamp 1667941163
transform 1 0 23576 0 -1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_419
timestamp 1667941163
transform 1 0 24136 0 -1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_2
timestamp 1667941163
transform 1 0 784 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1667941163
transform 1 0 2576 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_37
timestamp 1667941163
transform 1 0 2744 0 1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_53
timestamp 1667941163
transform 1 0 3640 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_79
timestamp 1667941163
transform 1 0 5096 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1667941163
transform 1 0 6552 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_108
timestamp 1667941163
transform 1 0 6720 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_133
timestamp 1667941163
transform 1 0 8120 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_159
timestamp 1667941163
transform 1 0 9576 0 1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_175
timestamp 1667941163
transform 1 0 10472 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_179
timestamp 1667941163
transform 1 0 10696 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_204
timestamp 1667941163
transform 1 0 12096 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_230
timestamp 1667941163
transform 1 0 13552 0 1 24304
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_246
timestamp 1667941163
transform 1 0 14448 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_250
timestamp 1667941163
transform 1 0 14672 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_275
timestamp 1667941163
transform 1 0 16072 0 1 24304
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_307
timestamp 1667941163
transform 1 0 17864 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_315
timestamp 1667941163
transform 1 0 18312 0 1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1667941163
transform 1 0 18648 0 1 24304
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1667941163
transform 1 0 22232 0 1 24304
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1667941163
transform 1 0 22456 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_392
timestamp 1667941163
transform 1 0 22624 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_400
timestamp 1667941163
transform 1 0 23072 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_409
timestamp 1667941163
transform 1 0 23576 0 1 24304
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_419
timestamp 1667941163
transform 1 0 24136 0 1 24304
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_2
timestamp 1667941163
transform 1 0 784 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_18
timestamp 1667941163
transform 1 0 1680 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_44
timestamp 1667941163
transform 1 0 3136 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1667941163
transform 1 0 4592 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_73
timestamp 1667941163
transform 1 0 4760 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_75
timestamp 1667941163
transform 1 0 4872 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_100
timestamp 1667941163
transform 1 0 6272 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_126
timestamp 1667941163
transform 1 0 7728 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_144
timestamp 1667941163
transform 1 0 8736 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_169
timestamp 1667941163
transform 1 0 10136 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_195
timestamp 1667941163
transform 1 0 11592 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_211
timestamp 1667941163
transform 1 0 12488 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_215
timestamp 1667941163
transform 1 0 12712 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_240
timestamp 1667941163
transform 1 0 14112 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_266
timestamp 1667941163
transform 1 0 15568 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_282
timestamp 1667941163
transform 1 0 16464 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1667941163
transform 1 0 16688 0 -1 25088
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1667941163
transform 1 0 20272 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1667941163
transform 1 0 20496 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_357
timestamp 1667941163
transform 1 0 20664 0 -1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_373
timestamp 1667941163
transform 1 0 21560 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_381
timestamp 1667941163
transform 1 0 22008 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_385
timestamp 1667941163
transform 1 0 22232 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_387
timestamp 1667941163
transform 1 0 22344 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_396
timestamp 1667941163
transform 1 0 22848 0 -1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_406
timestamp 1667941163
transform 1 0 23408 0 -1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_410
timestamp 1667941163
transform 1 0 23632 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_419
timestamp 1667941163
transform 1 0 24136 0 -1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_2
timestamp 1667941163
transform 1 0 784 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1667941163
transform 1 0 2576 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_37
timestamp 1667941163
transform 1 0 2744 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_65
timestamp 1667941163
transform 1 0 4312 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_91
timestamp 1667941163
transform 1 0 5768 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_99
timestamp 1667941163
transform 1 0 6216 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_103
timestamp 1667941163
transform 1 0 6440 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1667941163
transform 1 0 6552 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_108
timestamp 1667941163
transform 1 0 6720 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_133
timestamp 1667941163
transform 1 0 8120 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_159
timestamp 1667941163
transform 1 0 9576 0 1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_175
timestamp 1667941163
transform 1 0 10472 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_179
timestamp 1667941163
transform 1 0 10696 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_204
timestamp 1667941163
transform 1 0 12096 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_230
timestamp 1667941163
transform 1 0 13552 0 1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_246
timestamp 1667941163
transform 1 0 14448 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1667941163
transform 1 0 14672 0 1 25088
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1667941163
transform 1 0 18256 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1667941163
transform 1 0 18480 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_321
timestamp 1667941163
transform 1 0 18648 0 1 25088
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_353
timestamp 1667941163
transform 1 0 20440 0 1 25088
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_369
timestamp 1667941163
transform 1 0 21336 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_377
timestamp 1667941163
transform 1 0 21784 0 1 25088
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1667941163
transform 1 0 22456 0 1 25088
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_392
timestamp 1667941163
transform 1 0 22624 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_400
timestamp 1667941163
transform 1 0 23072 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_410
timestamp 1667941163
transform 1 0 23632 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_418
timestamp 1667941163
transform 1 0 24080 0 1 25088
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_2
timestamp 1667941163
transform 1 0 784 0 -1 25872
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_18
timestamp 1667941163
transform 1 0 1680 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_44
timestamp 1667941163
transform 1 0 3136 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1667941163
transform 1 0 4592 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_73
timestamp 1667941163
transform 1 0 4760 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_98
timestamp 1667941163
transform 1 0 6160 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_126
timestamp 1667941163
transform 1 0 7728 0 -1 25872
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_144
timestamp 1667941163
transform 1 0 8736 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 10136 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_195
timestamp 1667941163
transform 1 0 11592 0 -1 25872
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_211
timestamp 1667941163
transform 1 0 12488 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_215
timestamp 1667941163
transform 1 0 12712 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_240
timestamp 1667941163
transform 1 0 14112 0 -1 25872
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_272
timestamp 1667941163
transform 1 0 15904 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_280
timestamp 1667941163
transform 1 0 16352 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1667941163
transform 1 0 16688 0 -1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1667941163
transform 1 0 20272 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1667941163
transform 1 0 20496 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_357
timestamp 1667941163
transform 1 0 20664 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_365
timestamp 1667941163
transform 1 0 21112 0 -1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_369
timestamp 1667941163
transform 1 0 21336 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_371
timestamp 1667941163
transform 1 0 21448 0 -1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_380
timestamp 1667941163
transform 1 0 21952 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 22512 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_400
timestamp 1667941163
transform 1 0 23072 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_410
timestamp 1667941163
transform 1 0 23632 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_418
timestamp 1667941163
transform 1 0 24080 0 -1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_2
timestamp 1667941163
transform 1 0 784 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1667941163
transform 1 0 2576 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_37
timestamp 1667941163
transform 1 0 2744 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_65
timestamp 1667941163
transform 1 0 4312 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_91
timestamp 1667941163
transform 1 0 5768 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_99
timestamp 1667941163
transform 1 0 6216 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_103
timestamp 1667941163
transform 1 0 6440 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1667941163
transform 1 0 6552 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_108
timestamp 1667941163
transform 1 0 6720 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_133
timestamp 1667941163
transform 1 0 8120 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_159
timestamp 1667941163
transform 1 0 9576 0 1 25872
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_175
timestamp 1667941163
transform 1 0 10472 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_179
timestamp 1667941163
transform 1 0 10696 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_204
timestamp 1667941163
transform 1 0 12096 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_230
timestamp 1667941163
transform 1 0 13552 0 1 25872
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_246
timestamp 1667941163
transform 1 0 14448 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1667941163
transform 1 0 14672 0 1 25872
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1667941163
transform 1 0 18256 0 1 25872
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1667941163
transform 1 0 18480 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_321
timestamp 1667941163
transform 1 0 18648 0 1 25872
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_353
timestamp 1667941163
transform 1 0 20440 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_369
timestamp 1667941163
transform 1 0 21336 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_379
timestamp 1667941163
transform 1 0 21896 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1667941163
transform 1 0 22456 0 1 25872
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_392
timestamp 1667941163
transform 1 0 22624 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_400
timestamp 1667941163
transform 1 0 23072 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_410
timestamp 1667941163
transform 1 0 23632 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_418
timestamp 1667941163
transform 1 0 24080 0 1 25872
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_2
timestamp 1667941163
transform 1 0 784 0 -1 26656
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_18
timestamp 1667941163
transform 1 0 1680 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_44
timestamp 1667941163
transform 1 0 3136 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1667941163
transform 1 0 4592 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_73
timestamp 1667941163
transform 1 0 4760 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_98
timestamp 1667941163
transform 1 0 6160 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_124
timestamp 1667941163
transform 1 0 7616 0 -1 26656
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_140
timestamp 1667941163
transform 1 0 8512 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_144
timestamp 1667941163
transform 1 0 8736 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 10136 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_195
timestamp 1667941163
transform 1 0 11592 0 -1 26656
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_211
timestamp 1667941163
transform 1 0 12488 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1667941163
transform 1 0 12712 0 -1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1667941163
transform 1 0 16296 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1667941163
transform 1 0 16520 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1667941163
transform 1 0 16688 0 -1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1667941163
transform 1 0 20272 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1667941163
transform 1 0 20496 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_357
timestamp 1667941163
transform 1 0 20664 0 -1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_361
timestamp 1667941163
transform 1 0 20888 0 -1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_370
timestamp 1667941163
transform 1 0 21392 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_380
timestamp 1667941163
transform 1 0 21952 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 22512 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_400
timestamp 1667941163
transform 1 0 23072 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_410
timestamp 1667941163
transform 1 0 23632 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_418
timestamp 1667941163
transform 1 0 24080 0 -1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_2
timestamp 1667941163
transform 1 0 784 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1667941163
transform 1 0 2576 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_37
timestamp 1667941163
transform 1 0 2744 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_65
timestamp 1667941163
transform 1 0 4312 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_91
timestamp 1667941163
transform 1 0 5768 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_99
timestamp 1667941163
transform 1 0 6216 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_103
timestamp 1667941163
transform 1 0 6440 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1667941163
transform 1 0 6552 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_108
timestamp 1667941163
transform 1 0 6720 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_133
timestamp 1667941163
transform 1 0 8120 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_159
timestamp 1667941163
transform 1 0 9576 0 1 26656
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_175
timestamp 1667941163
transform 1 0 10472 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_179
timestamp 1667941163
transform 1 0 10696 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_204
timestamp 1667941163
transform 1 0 12096 0 1 26656
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_236
timestamp 1667941163
transform 1 0 13888 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_244
timestamp 1667941163
transform 1 0 14336 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1667941163
transform 1 0 14672 0 1 26656
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 18256 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1667941163
transform 1 0 18480 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_321
timestamp 1667941163
transform 1 0 18648 0 1 26656
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_337
timestamp 1667941163
transform 1 0 19544 0 1 26656
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_349
timestamp 1667941163
transform 1 0 20216 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_359
timestamp 1667941163
transform 1 0 20776 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_369
timestamp 1667941163
transform 1 0 21336 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 21896 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1667941163
transform 1 0 22456 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_392
timestamp 1667941163
transform 1 0 22624 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_401
timestamp 1667941163
transform 1 0 23128 0 1 26656
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_411
timestamp 1667941163
transform 1 0 23688 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_419
timestamp 1667941163
transform 1 0 24136 0 1 26656
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_2
timestamp 1667941163
transform 1 0 784 0 -1 27440
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_18
timestamp 1667941163
transform 1 0 1680 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_44
timestamp 1667941163
transform 1 0 3136 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1667941163
transform 1 0 4592 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_73
timestamp 1667941163
transform 1 0 4760 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_98
timestamp 1667941163
transform 1 0 6160 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_124
timestamp 1667941163
transform 1 0 7616 0 -1 27440
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_140
timestamp 1667941163
transform 1 0 8512 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_144
timestamp 1667941163
transform 1 0 8736 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_169
timestamp 1667941163
transform 1 0 10136 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_195
timestamp 1667941163
transform 1 0 11592 0 -1 27440
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_211
timestamp 1667941163
transform 1 0 12488 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1667941163
transform 1 0 12712 0 -1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1667941163
transform 1 0 16296 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1667941163
transform 1 0 16520 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1667941163
transform 1 0 16688 0 -1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1667941163
transform 1 0 20272 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1667941163
transform 1 0 20496 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_357
timestamp 1667941163
transform 1 0 20664 0 -1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_361
timestamp 1667941163
transform 1 0 20888 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_371
timestamp 1667941163
transform 1 0 21448 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_381
timestamp 1667941163
transform 1 0 22008 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_391
timestamp 1667941163
transform 1 0 22568 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_401
timestamp 1667941163
transform 1 0 23128 0 -1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_411
timestamp 1667941163
transform 1 0 23688 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_419
timestamp 1667941163
transform 1 0 24136 0 -1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_2
timestamp 1667941163
transform 1 0 784 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1667941163
transform 1 0 2576 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_37
timestamp 1667941163
transform 1 0 2744 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_65
timestamp 1667941163
transform 1 0 4312 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_91
timestamp 1667941163
transform 1 0 5768 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_99
timestamp 1667941163
transform 1 0 6216 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_103
timestamp 1667941163
transform 1 0 6440 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1667941163
transform 1 0 6552 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_108
timestamp 1667941163
transform 1 0 6720 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_133
timestamp 1667941163
transform 1 0 8120 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_159
timestamp 1667941163
transform 1 0 9576 0 1 27440
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_175
timestamp 1667941163
transform 1 0 10472 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_179
timestamp 1667941163
transform 1 0 10696 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_204
timestamp 1667941163
transform 1 0 12096 0 1 27440
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_236
timestamp 1667941163
transform 1 0 13888 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_244
timestamp 1667941163
transform 1 0 14336 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1667941163
transform 1 0 14672 0 1 27440
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1667941163
transform 1 0 18256 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1667941163
transform 1 0 18480 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_321
timestamp 1667941163
transform 1 0 18648 0 1 27440
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_353
timestamp 1667941163
transform 1 0 20440 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_369
timestamp 1667941163
transform 1 0 21336 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_379
timestamp 1667941163
transform 1 0 21896 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1667941163
transform 1 0 22456 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_392
timestamp 1667941163
transform 1 0 22624 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_396
timestamp 1667941163
transform 1 0 22848 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_405
timestamp 1667941163
transform 1 0 23352 0 1 27440
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_415
timestamp 1667941163
transform 1 0 23912 0 1 27440
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_419
timestamp 1667941163
transform 1 0 24136 0 1 27440
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_2
timestamp 1667941163
transform 1 0 784 0 -1 28224
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_18
timestamp 1667941163
transform 1 0 1680 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_44
timestamp 1667941163
transform 1 0 3136 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1667941163
transform 1 0 4592 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_73
timestamp 1667941163
transform 1 0 4760 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_98
timestamp 1667941163
transform 1 0 6160 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_124
timestamp 1667941163
transform 1 0 7616 0 -1 28224
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_140
timestamp 1667941163
transform 1 0 8512 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1667941163
transform 1 0 8736 0 -1 28224
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1667941163
transform 1 0 12320 0 -1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1667941163
transform 1 0 12544 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1667941163
transform 1 0 12712 0 -1 28224
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1667941163
transform 1 0 16296 0 -1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1667941163
transform 1 0 16520 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1667941163
transform 1 0 16688 0 -1 28224
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1667941163
transform 1 0 20272 0 -1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1667941163
transform 1 0 20496 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_357
timestamp 1667941163
transform 1 0 20664 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_365
timestamp 1667941163
transform 1 0 21112 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_367
timestamp 1667941163
transform 1 0 21224 0 -1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_376
timestamp 1667941163
transform 1 0 21728 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_386
timestamp 1667941163
transform 1 0 22288 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_396
timestamp 1667941163
transform 1 0 22848 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_406
timestamp 1667941163
transform 1 0 23408 0 -1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_416
timestamp 1667941163
transform 1 0 23968 0 -1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1667941163
transform 1 0 784 0 1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1667941163
transform 1 0 2576 0 1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_37
timestamp 1667941163
transform 1 0 2744 0 1 28224
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_53
timestamp 1667941163
transform 1 0 3640 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_81
timestamp 1667941163
transform 1 0 5208 0 1 28224
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_97
timestamp 1667941163
transform 1 0 6104 0 1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1667941163
transform 1 0 6552 0 1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1667941163
transform 1 0 6720 0 1 28224
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1667941163
transform 1 0 10304 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1667941163
transform 1 0 10528 0 1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1667941163
transform 1 0 10696 0 1 28224
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1667941163
transform 1 0 14280 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1667941163
transform 1 0 14504 0 1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1667941163
transform 1 0 14672 0 1 28224
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1667941163
transform 1 0 18256 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1667941163
transform 1 0 18480 0 1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_321
timestamp 1667941163
transform 1 0 18648 0 1 28224
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_353
timestamp 1667941163
transform 1 0 20440 0 1 28224
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_369
timestamp 1667941163
transform 1 0 21336 0 1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_377
timestamp 1667941163
transform 1 0 21784 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1667941163
transform 1 0 22456 0 1 28224
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_392
timestamp 1667941163
transform 1 0 22624 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_396
timestamp 1667941163
transform 1 0 22848 0 1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_406
timestamp 1667941163
transform 1 0 23408 0 1 28224
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_416
timestamp 1667941163
transform 1 0 23968 0 1 28224
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_2
timestamp 1667941163
transform 1 0 784 0 -1 29008
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_34
timestamp 1667941163
transform 1 0 2576 0 -1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_42
timestamp 1667941163
transform 1 0 3024 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1667941163
transform 1 0 4592 0 -1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_73
timestamp 1667941163
transform 1 0 4760 0 -1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_98
timestamp 1667941163
transform 1 0 6160 0 -1 29008
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_130
timestamp 1667941163
transform 1 0 7952 0 -1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_138
timestamp 1667941163
transform 1 0 8400 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1667941163
transform 1 0 8736 0 -1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1667941163
transform 1 0 12320 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1667941163
transform 1 0 12544 0 -1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1667941163
transform 1 0 12712 0 -1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1667941163
transform 1 0 16296 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1667941163
transform 1 0 16520 0 -1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1667941163
transform 1 0 16688 0 -1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1667941163
transform 1 0 20272 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1667941163
transform 1 0 20496 0 -1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_357
timestamp 1667941163
transform 1 0 20664 0 -1 29008
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_373
timestamp 1667941163
transform 1 0 21560 0 -1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_381
timestamp 1667941163
transform 1 0 22008 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_385
timestamp 1667941163
transform 1 0 22232 0 -1 29008
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_395
timestamp 1667941163
transform 1 0 22792 0 -1 29008
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_405
timestamp 1667941163
transform 1 0 23352 0 -1 29008
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_415
timestamp 1667941163
transform 1 0 23912 0 -1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_419
timestamp 1667941163
transform 1 0 24136 0 -1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_2
timestamp 1667941163
transform 1 0 784 0 1 29008
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_34
timestamp 1667941163
transform 1 0 2576 0 1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_37
timestamp 1667941163
transform 1 0 2744 0 1 29008
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_53
timestamp 1667941163
transform 1 0 3640 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_81
timestamp 1667941163
transform 1 0 5208 0 1 29008
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_97
timestamp 1667941163
transform 1 0 6104 0 1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1667941163
transform 1 0 6552 0 1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1667941163
transform 1 0 6720 0 1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1667941163
transform 1 0 10304 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1667941163
transform 1 0 10528 0 1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1667941163
transform 1 0 10696 0 1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1667941163
transform 1 0 14280 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1667941163
transform 1 0 14504 0 1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1667941163
transform 1 0 14672 0 1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1667941163
transform 1 0 18256 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1667941163
transform 1 0 18480 0 1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1667941163
transform 1 0 18648 0 1 29008
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1667941163
transform 1 0 22232 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1667941163
transform 1 0 22456 0 1 29008
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_392
timestamp 1667941163
transform 1 0 22624 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_396
timestamp 1667941163
transform 1 0 22848 0 1 29008
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_406
timestamp 1667941163
transform 1 0 23408 0 1 29008
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_416
timestamp 1667941163
transform 1 0 23968 0 1 29008
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_2
timestamp 1667941163
transform 1 0 784 0 -1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_66
timestamp 1667941163
transform 1 0 4368 0 -1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1667941163
transform 1 0 4592 0 -1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1667941163
transform 1 0 4760 0 -1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1667941163
transform 1 0 8344 0 -1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1667941163
transform 1 0 8568 0 -1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1667941163
transform 1 0 8736 0 -1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1667941163
transform 1 0 12320 0 -1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1667941163
transform 1 0 12544 0 -1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1667941163
transform 1 0 12712 0 -1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1667941163
transform 1 0 16296 0 -1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1667941163
transform 1 0 16520 0 -1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1667941163
transform 1 0 16688 0 -1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1667941163
transform 1 0 20272 0 -1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1667941163
transform 1 0 20496 0 -1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_357
timestamp 1667941163
transform 1 0 20664 0 -1 29792
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_389
timestamp 1667941163
transform 1 0 22456 0 -1 29792
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_397
timestamp 1667941163
transform 1 0 22904 0 -1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_401
timestamp 1667941163
transform 1 0 23128 0 -1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_410
timestamp 1667941163
transform 1 0 23632 0 -1 29792
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_418
timestamp 1667941163
transform 1 0 24080 0 -1 29792
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_2
timestamp 1667941163
transform 1 0 784 0 1 29792
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1667941163
transform 1 0 2576 0 1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1667941163
transform 1 0 2744 0 1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1667941163
transform 1 0 6328 0 1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1667941163
transform 1 0 6552 0 1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1667941163
transform 1 0 6720 0 1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1667941163
transform 1 0 10304 0 1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1667941163
transform 1 0 10528 0 1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1667941163
transform 1 0 10696 0 1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1667941163
transform 1 0 14280 0 1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1667941163
transform 1 0 14504 0 1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1667941163
transform 1 0 14672 0 1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1667941163
transform 1 0 18256 0 1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1667941163
transform 1 0 18480 0 1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1667941163
transform 1 0 18648 0 1 29792
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1667941163
transform 1 0 22232 0 1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1667941163
transform 1 0 22456 0 1 29792
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_392
timestamp 1667941163
transform 1 0 22624 0 1 29792
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_408
timestamp 1667941163
transform 1 0 23520 0 1 29792
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_416
timestamp 1667941163
transform 1 0 23968 0 1 29792
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_2
timestamp 1667941163
transform 1 0 784 0 -1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_66
timestamp 1667941163
transform 1 0 4368 0 -1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_70
timestamp 1667941163
transform 1 0 4592 0 -1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1667941163
transform 1 0 4760 0 -1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1667941163
transform 1 0 8344 0 -1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1667941163
transform 1 0 8568 0 -1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1667941163
transform 1 0 8736 0 -1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1667941163
transform 1 0 12320 0 -1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1667941163
transform 1 0 12544 0 -1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1667941163
transform 1 0 12712 0 -1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1667941163
transform 1 0 16296 0 -1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1667941163
transform 1 0 16520 0 -1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1667941163
transform 1 0 16688 0 -1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1667941163
transform 1 0 20272 0 -1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1667941163
transform 1 0 20496 0 -1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_357
timestamp 1667941163
transform 1 0 20664 0 -1 30576
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_389
timestamp 1667941163
transform 1 0 22456 0 -1 30576
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_405
timestamp 1667941163
transform 1 0 23352 0 -1 30576
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_413
timestamp 1667941163
transform 1 0 23800 0 -1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_417
timestamp 1667941163
transform 1 0 24024 0 -1 30576
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_419
timestamp 1667941163
transform 1 0 24136 0 -1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_2
timestamp 1667941163
transform 1 0 784 0 1 30576
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_34
timestamp 1667941163
transform 1 0 2576 0 1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1667941163
transform 1 0 2744 0 1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1667941163
transform 1 0 6328 0 1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1667941163
transform 1 0 6552 0 1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1667941163
transform 1 0 6720 0 1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1667941163
transform 1 0 10304 0 1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1667941163
transform 1 0 10528 0 1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1667941163
transform 1 0 10696 0 1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1667941163
transform 1 0 14280 0 1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1667941163
transform 1 0 14504 0 1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1667941163
transform 1 0 14672 0 1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1667941163
transform 1 0 18256 0 1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1667941163
transform 1 0 18480 0 1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1667941163
transform 1 0 18648 0 1 30576
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1667941163
transform 1 0 22232 0 1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1667941163
transform 1 0 22456 0 1 30576
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_392
timestamp 1667941163
transform 1 0 22624 0 1 30576
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_408
timestamp 1667941163
transform 1 0 23520 0 1 30576
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_416
timestamp 1667941163
transform 1 0 23968 0 1 30576
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_2
timestamp 1667941163
transform 1 0 784 0 -1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_66
timestamp 1667941163
transform 1 0 4368 0 -1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_70
timestamp 1667941163
transform 1 0 4592 0 -1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1667941163
transform 1 0 4760 0 -1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1667941163
transform 1 0 8344 0 -1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1667941163
transform 1 0 8568 0 -1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1667941163
transform 1 0 8736 0 -1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1667941163
transform 1 0 12320 0 -1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1667941163
transform 1 0 12544 0 -1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1667941163
transform 1 0 12712 0 -1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1667941163
transform 1 0 16296 0 -1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1667941163
transform 1 0 16520 0 -1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1667941163
transform 1 0 16688 0 -1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1667941163
transform 1 0 20272 0 -1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1667941163
transform 1 0 20496 0 -1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_357
timestamp 1667941163
transform 1 0 20664 0 -1 31360
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_389
timestamp 1667941163
transform 1 0 22456 0 -1 31360
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_405
timestamp 1667941163
transform 1 0 23352 0 -1 31360
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_413
timestamp 1667941163
transform 1 0 23800 0 -1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_417
timestamp 1667941163
transform 1 0 24024 0 -1 31360
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_419
timestamp 1667941163
transform 1 0 24136 0 -1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_2
timestamp 1667941163
transform 1 0 784 0 1 31360
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_34
timestamp 1667941163
transform 1 0 2576 0 1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1667941163
transform 1 0 2744 0 1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1667941163
transform 1 0 6328 0 1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1667941163
transform 1 0 6552 0 1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1667941163
transform 1 0 6720 0 1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1667941163
transform 1 0 10304 0 1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1667941163
transform 1 0 10528 0 1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1667941163
transform 1 0 10696 0 1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1667941163
transform 1 0 14280 0 1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1667941163
transform 1 0 14504 0 1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1667941163
transform 1 0 14672 0 1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1667941163
transform 1 0 18256 0 1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1667941163
transform 1 0 18480 0 1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1667941163
transform 1 0 18648 0 1 31360
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1667941163
transform 1 0 22232 0 1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1667941163
transform 1 0 22456 0 1 31360
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_392
timestamp 1667941163
transform 1 0 22624 0 1 31360
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_408
timestamp 1667941163
transform 1 0 23520 0 1 31360
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_416
timestamp 1667941163
transform 1 0 23968 0 1 31360
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_2
timestamp 1667941163
transform 1 0 784 0 -1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_66
timestamp 1667941163
transform 1 0 4368 0 -1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_70
timestamp 1667941163
transform 1 0 4592 0 -1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1667941163
transform 1 0 4760 0 -1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1667941163
transform 1 0 8344 0 -1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1667941163
transform 1 0 8568 0 -1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1667941163
transform 1 0 8736 0 -1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1667941163
transform 1 0 12320 0 -1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1667941163
transform 1 0 12544 0 -1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1667941163
transform 1 0 12712 0 -1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1667941163
transform 1 0 16296 0 -1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1667941163
transform 1 0 16520 0 -1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1667941163
transform 1 0 16688 0 -1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1667941163
transform 1 0 20272 0 -1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1667941163
transform 1 0 20496 0 -1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_357
timestamp 1667941163
transform 1 0 20664 0 -1 32144
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_389
timestamp 1667941163
transform 1 0 22456 0 -1 32144
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_405
timestamp 1667941163
transform 1 0 23352 0 -1 32144
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_413
timestamp 1667941163
transform 1 0 23800 0 -1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_417
timestamp 1667941163
transform 1 0 24024 0 -1 32144
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_419
timestamp 1667941163
transform 1 0 24136 0 -1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_2
timestamp 1667941163
transform 1 0 784 0 1 32144
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_34
timestamp 1667941163
transform 1 0 2576 0 1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1667941163
transform 1 0 2744 0 1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1667941163
transform 1 0 6328 0 1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1667941163
transform 1 0 6552 0 1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1667941163
transform 1 0 6720 0 1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1667941163
transform 1 0 10304 0 1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1667941163
transform 1 0 10528 0 1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1667941163
transform 1 0 10696 0 1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1667941163
transform 1 0 14280 0 1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1667941163
transform 1 0 14504 0 1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1667941163
transform 1 0 14672 0 1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1667941163
transform 1 0 18256 0 1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1667941163
transform 1 0 18480 0 1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1667941163
transform 1 0 18648 0 1 32144
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1667941163
transform 1 0 22232 0 1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1667941163
transform 1 0 22456 0 1 32144
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_392
timestamp 1667941163
transform 1 0 22624 0 1 32144
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_408
timestamp 1667941163
transform 1 0 23520 0 1 32144
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_416
timestamp 1667941163
transform 1 0 23968 0 1 32144
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_2
timestamp 1667941163
transform 1 0 784 0 -1 32928
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_66
timestamp 1667941163
transform 1 0 4368 0 -1 32928
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_70
timestamp 1667941163
transform 1 0 4592 0 -1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1667941163
transform 1 0 4760 0 -1 32928
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1667941163
transform 1 0 8344 0 -1 32928
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1667941163
transform 1 0 8568 0 -1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1667941163
transform 1 0 8736 0 -1 32928
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1667941163
transform 1 0 12320 0 -1 32928
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1667941163
transform 1 0 12544 0 -1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1667941163
transform 1 0 12712 0 -1 32928
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1667941163
transform 1 0 16296 0 -1 32928
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1667941163
transform 1 0 16520 0 -1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1667941163
transform 1 0 16688 0 -1 32928
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1667941163
transform 1 0 20272 0 -1 32928
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1667941163
transform 1 0 20496 0 -1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_357
timestamp 1667941163
transform 1 0 20664 0 -1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_389
timestamp 1667941163
transform 1 0 22456 0 -1 32928
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_405
timestamp 1667941163
transform 1 0 23352 0 -1 32928
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_413
timestamp 1667941163
transform 1 0 23800 0 -1 32928
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_417
timestamp 1667941163
transform 1 0 24024 0 -1 32928
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_419
timestamp 1667941163
transform 1 0 24136 0 -1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_2
timestamp 1667941163
transform 1 0 784 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_34
timestamp 1667941163
transform 1 0 2576 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_37
timestamp 1667941163
transform 1 0 2744 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_69
timestamp 1667941163
transform 1 0 4536 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_72
timestamp 1667941163
transform 1 0 4704 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_104
timestamp 1667941163
transform 1 0 6496 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_107
timestamp 1667941163
transform 1 0 6664 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_139
timestamp 1667941163
transform 1 0 8456 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_142
timestamp 1667941163
transform 1 0 8624 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_174
timestamp 1667941163
transform 1 0 10416 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_177
timestamp 1667941163
transform 1 0 10584 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_209
timestamp 1667941163
transform 1 0 12376 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_212
timestamp 1667941163
transform 1 0 12544 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_244
timestamp 1667941163
transform 1 0 14336 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_247
timestamp 1667941163
transform 1 0 14504 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_279
timestamp 1667941163
transform 1 0 16296 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_282
timestamp 1667941163
transform 1 0 16464 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_314
timestamp 1667941163
transform 1 0 18256 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_317
timestamp 1667941163
transform 1 0 18424 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_349
timestamp 1667941163
transform 1 0 20216 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_352
timestamp 1667941163
transform 1 0 20384 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_384
timestamp 1667941163
transform 1 0 22176 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_387
timestamp 1667941163
transform 1 0 22344 0 1 32928
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_419
timestamp 1667941163
transform 1 0 24136 0 1 32928
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 24304 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 24304 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 24304 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 24304 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 24304 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 24304 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 24304 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 24304 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 24304 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 24304 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 24304 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 24304 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 24304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 24304 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 24304 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 24304 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 24304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1667941163
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1667941163
transform -1 0 24304 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1667941163
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1667941163
transform -1 0 24304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1667941163
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1667941163
transform -1 0 24304 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1667941163
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1667941163
transform -1 0 24304 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1667941163
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1667941163
transform -1 0 24304 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1667941163
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1667941163
transform -1 0 24304 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1667941163
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1667941163
transform -1 0 24304 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1667941163
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1667941163
transform -1 0 24304 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1667941163
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1667941163
transform -1 0 24304 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1667941163
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1667941163
transform -1 0 24304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1667941163
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1667941163
transform -1 0 24304 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1667941163
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1667941163
transform -1 0 24304 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1667941163
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1667941163
transform -1 0 24304 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1667941163
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1667941163
transform -1 0 24304 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1667941163
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1667941163
transform -1 0 24304 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1667941163
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1667941163
transform -1 0 24304 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1667941163
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1667941163
transform -1 0 24304 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1667941163
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1667941163
transform -1 0 24304 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1667941163
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1667941163
transform -1 0 24304 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1667941163
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1667941163
transform -1 0 24304 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1667941163
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1667941163
transform -1 0 24304 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1667941163
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1667941163
transform -1 0 24304 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1667941163
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1667941163
transform -1 0 24304 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1667941163
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1667941163
transform -1 0 24304 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1667941163
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1667941163
transform -1 0 24304 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1667941163
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1667941163
transform -1 0 24304 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1667941163
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1667941163
transform -1 0 24304 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1667941163
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1667941163
transform -1 0 24304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1667941163
transform 1 0 672 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1667941163
transform -1 0 24304 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1667941163
transform 1 0 672 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1667941163
transform -1 0 24304 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1667941163
transform 1 0 672 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1667941163
transform -1 0 24304 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1667941163
transform 1 0 672 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1667941163
transform -1 0 24304 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1667941163
transform 1 0 672 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1667941163
transform -1 0 24304 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1667941163
transform 1 0 672 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1667941163
transform -1 0 24304 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1667941163
transform 1 0 672 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1667941163
transform -1 0 24304 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1667941163
transform 1 0 672 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1667941163
transform -1 0 24304 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1667941163
transform 1 0 672 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1667941163
transform -1 0 24304 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1667941163
transform 1 0 672 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1667941163
transform -1 0 24304 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1667941163
transform 1 0 672 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1667941163
transform -1 0 24304 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1667941163
transform 1 0 672 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1667941163
transform -1 0 24304 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1667941163
transform 1 0 672 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1667941163
transform -1 0 24304 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1667941163
transform 1 0 672 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1667941163
transform -1 0 24304 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1667941163
transform 1 0 672 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1667941163
transform -1 0 24304 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1667941163
transform 1 0 672 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1667941163
transform -1 0 24304 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1667941163
transform 1 0 672 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1667941163
transform -1 0 24304 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1667941163
transform 1 0 672 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1667941163
transform -1 0 24304 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1667941163
transform 1 0 672 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1667941163
transform -1 0 24304 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1667941163
transform 1 0 672 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1667941163
transform -1 0 24304 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1667941163
transform 1 0 672 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1667941163
transform -1 0 24304 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1667941163
transform 1 0 672 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1667941163
transform -1 0 24304 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1667941163
transform 1 0 672 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1667941163
transform -1 0 24304 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1667941163
transform 1 0 672 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1667941163
transform -1 0 24304 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1667941163
transform 1 0 672 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1667941163
transform -1 0 24304 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1667941163
transform 1 0 672 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1667941163
transform -1 0 24304 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1667941163
transform 1 0 672 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1667941163
transform -1 0 24304 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1667941163
transform 1 0 672 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1667941163
transform -1 0 24304 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1667941163
transform 1 0 672 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1667941163
transform -1 0 24304 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1667941163
transform 1 0 672 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1667941163
transform -1 0 24304 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1667941163
transform 1 0 672 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1667941163
transform -1 0 24304 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1667941163
transform 1 0 672 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1667941163
transform -1 0 24304 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1667941163
transform 1 0 672 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1667941163
transform -1 0 24304 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1667941163
transform 1 0 672 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1667941163
transform -1 0 24304 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1667941163
transform 1 0 672 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1667941163
transform -1 0 24304 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1667941163
transform 1 0 672 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1667941163
transform -1 0 24304 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 8512 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 10472 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 14392 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 16352 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 18312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 20272 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 22232 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 12600 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 16576 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 20552 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 10584 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 14560 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 18536 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 22512 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 12600 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 16576 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 20552 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 10584 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 14560 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 18536 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 22512 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 8624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 12600 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 16576 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 20552 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 10584 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 14560 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 18536 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 22512 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 8624 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 12600 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 16576 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 20552 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 10584 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 14560 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 18536 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 22512 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 8624 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 12600 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 16576 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 20552 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 10584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 14560 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 18536 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 22512 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 4648 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 12600 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 16576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 20552 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 6608 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 14560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 18536 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 22512 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 4648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 12600 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 16576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 20552 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 6608 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 14560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 18536 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 22512 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 4648 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 12600 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 16576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 20552 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 6608 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 14560 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 18536 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 22512 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 4648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 12600 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 16576 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 20552 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 6608 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 14560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 18536 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 22512 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 4648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 12600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 16576 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 20552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 6608 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 14560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 18536 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 22512 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 4648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 12600 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 16576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 20552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1667941163
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1667941163
transform 1 0 6608 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1667941163
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1667941163
transform 1 0 14560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1667941163
transform 1 0 18536 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1667941163
transform 1 0 22512 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1667941163
transform 1 0 4648 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1667941163
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1667941163
transform 1 0 12600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1667941163
transform 1 0 16576 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1667941163
transform 1 0 20552 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1667941163
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1667941163
transform 1 0 6608 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1667941163
transform 1 0 10584 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1667941163
transform 1 0 14560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1667941163
transform 1 0 18536 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1667941163
transform 1 0 22512 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1667941163
transform 1 0 4648 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1667941163
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1667941163
transform 1 0 12600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1667941163
transform 1 0 16576 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1667941163
transform 1 0 20552 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1667941163
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1667941163
transform 1 0 6608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1667941163
transform 1 0 10584 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1667941163
transform 1 0 14560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1667941163
transform 1 0 18536 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1667941163
transform 1 0 22512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1667941163
transform 1 0 4648 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1667941163
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1667941163
transform 1 0 12600 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1667941163
transform 1 0 16576 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1667941163
transform 1 0 20552 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1667941163
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1667941163
transform 1 0 6608 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1667941163
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1667941163
transform 1 0 14560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1667941163
transform 1 0 18536 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1667941163
transform 1 0 22512 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1667941163
transform 1 0 4648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1667941163
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1667941163
transform 1 0 12600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1667941163
transform 1 0 16576 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1667941163
transform 1 0 20552 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1667941163
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1667941163
transform 1 0 6608 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1667941163
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1667941163
transform 1 0 14560 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1667941163
transform 1 0 18536 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1667941163
transform 1 0 22512 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1667941163
transform 1 0 4648 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1667941163
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1667941163
transform 1 0 12600 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1667941163
transform 1 0 16576 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1667941163
transform 1 0 20552 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1667941163
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1667941163
transform 1 0 6608 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1667941163
transform 1 0 10584 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1667941163
transform 1 0 14560 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1667941163
transform 1 0 18536 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1667941163
transform 1 0 22512 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1667941163
transform 1 0 4648 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1667941163
transform 1 0 8624 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1667941163
transform 1 0 12600 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1667941163
transform 1 0 16576 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1667941163
transform 1 0 20552 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1667941163
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1667941163
transform 1 0 6608 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1667941163
transform 1 0 10584 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1667941163
transform 1 0 14560 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1667941163
transform 1 0 18536 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1667941163
transform 1 0 22512 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1667941163
transform 1 0 4648 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1667941163
transform 1 0 8624 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1667941163
transform 1 0 12600 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1667941163
transform 1 0 16576 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1667941163
transform 1 0 20552 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1667941163
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1667941163
transform 1 0 6608 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1667941163
transform 1 0 10584 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1667941163
transform 1 0 14560 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1667941163
transform 1 0 18536 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1667941163
transform 1 0 22512 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1667941163
transform 1 0 4648 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1667941163
transform 1 0 8624 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1667941163
transform 1 0 12600 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1667941163
transform 1 0 16576 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1667941163
transform 1 0 20552 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1667941163
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1667941163
transform 1 0 6608 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1667941163
transform 1 0 10584 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1667941163
transform 1 0 14560 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1667941163
transform 1 0 18536 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1667941163
transform 1 0 22512 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1667941163
transform 1 0 4648 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1667941163
transform 1 0 8624 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1667941163
transform 1 0 12600 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1667941163
transform 1 0 16576 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1667941163
transform 1 0 20552 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1667941163
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1667941163
transform 1 0 6608 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1667941163
transform 1 0 10584 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1667941163
transform 1 0 14560 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1667941163
transform 1 0 18536 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1667941163
transform 1 0 22512 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1667941163
transform 1 0 4648 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1667941163
transform 1 0 8624 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1667941163
transform 1 0 12600 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1667941163
transform 1 0 16576 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1667941163
transform 1 0 20552 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1667941163
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1667941163
transform 1 0 6608 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1667941163
transform 1 0 10584 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1667941163
transform 1 0 14560 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1667941163
transform 1 0 18536 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1667941163
transform 1 0 22512 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1667941163
transform 1 0 4648 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1667941163
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1667941163
transform 1 0 12600 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1667941163
transform 1 0 16576 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1667941163
transform 1 0 20552 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1667941163
transform 1 0 2632 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1667941163
transform 1 0 6608 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1667941163
transform 1 0 10584 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1667941163
transform 1 0 14560 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1667941163
transform 1 0 18536 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1667941163
transform 1 0 22512 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1667941163
transform 1 0 4648 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1667941163
transform 1 0 8624 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1667941163
transform 1 0 12600 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1667941163
transform 1 0 16576 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1667941163
transform 1 0 20552 0 -1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1667941163
transform 1 0 2632 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1667941163
transform 1 0 6608 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1667941163
transform 1 0 10584 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1667941163
transform 1 0 14560 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1667941163
transform 1 0 18536 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1667941163
transform 1 0 22512 0 1 19600
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1667941163
transform 1 0 4648 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1667941163
transform 1 0 8624 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1667941163
transform 1 0 12600 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1667941163
transform 1 0 16576 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1667941163
transform 1 0 20552 0 -1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1667941163
transform 1 0 2632 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1667941163
transform 1 0 6608 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1667941163
transform 1 0 10584 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1667941163
transform 1 0 14560 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1667941163
transform 1 0 18536 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1667941163
transform 1 0 22512 0 1 20384
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1667941163
transform 1 0 4648 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1667941163
transform 1 0 8624 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1667941163
transform 1 0 12600 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1667941163
transform 1 0 16576 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1667941163
transform 1 0 20552 0 -1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1667941163
transform 1 0 2632 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1667941163
transform 1 0 6608 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1667941163
transform 1 0 10584 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1667941163
transform 1 0 14560 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1667941163
transform 1 0 18536 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1667941163
transform 1 0 22512 0 1 21168
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1667941163
transform 1 0 4648 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1667941163
transform 1 0 8624 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1667941163
transform 1 0 12600 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1667941163
transform 1 0 16576 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1667941163
transform 1 0 20552 0 -1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1667941163
transform 1 0 2632 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1667941163
transform 1 0 6608 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1667941163
transform 1 0 10584 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1667941163
transform 1 0 14560 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1667941163
transform 1 0 18536 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1667941163
transform 1 0 22512 0 1 21952
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1667941163
transform 1 0 4648 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1667941163
transform 1 0 8624 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1667941163
transform 1 0 12600 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1667941163
transform 1 0 16576 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1667941163
transform 1 0 20552 0 -1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1667941163
transform 1 0 2632 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1667941163
transform 1 0 6608 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1667941163
transform 1 0 10584 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1667941163
transform 1 0 14560 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1667941163
transform 1 0 18536 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1667941163
transform 1 0 22512 0 1 22736
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1667941163
transform 1 0 4648 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1667941163
transform 1 0 8624 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1667941163
transform 1 0 12600 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1667941163
transform 1 0 16576 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1667941163
transform 1 0 20552 0 -1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1667941163
transform 1 0 2632 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1667941163
transform 1 0 6608 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1667941163
transform 1 0 10584 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1667941163
transform 1 0 14560 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1667941163
transform 1 0 18536 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1667941163
transform 1 0 22512 0 1 23520
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1667941163
transform 1 0 4648 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1667941163
transform 1 0 8624 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1667941163
transform 1 0 12600 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1667941163
transform 1 0 16576 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1667941163
transform 1 0 20552 0 -1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1667941163
transform 1 0 2632 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1667941163
transform 1 0 6608 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1667941163
transform 1 0 10584 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1667941163
transform 1 0 14560 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1667941163
transform 1 0 18536 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1667941163
transform 1 0 22512 0 1 24304
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1667941163
transform 1 0 4648 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1667941163
transform 1 0 8624 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1667941163
transform 1 0 12600 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1667941163
transform 1 0 16576 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1667941163
transform 1 0 20552 0 -1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1667941163
transform 1 0 2632 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1667941163
transform 1 0 6608 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1667941163
transform 1 0 10584 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1667941163
transform 1 0 14560 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1667941163
transform 1 0 18536 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1667941163
transform 1 0 22512 0 1 25088
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1667941163
transform 1 0 4648 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1667941163
transform 1 0 8624 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1667941163
transform 1 0 12600 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1667941163
transform 1 0 16576 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1667941163
transform 1 0 20552 0 -1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1667941163
transform 1 0 2632 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1667941163
transform 1 0 6608 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1667941163
transform 1 0 10584 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1667941163
transform 1 0 14560 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1667941163
transform 1 0 18536 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1667941163
transform 1 0 22512 0 1 25872
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1667941163
transform 1 0 4648 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1667941163
transform 1 0 8624 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1667941163
transform 1 0 12600 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1667941163
transform 1 0 16576 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1667941163
transform 1 0 20552 0 -1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1667941163
transform 1 0 2632 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1667941163
transform 1 0 6608 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1667941163
transform 1 0 10584 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1667941163
transform 1 0 14560 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1667941163
transform 1 0 18536 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1667941163
transform 1 0 22512 0 1 26656
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1667941163
transform 1 0 4648 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1667941163
transform 1 0 8624 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1667941163
transform 1 0 12600 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1667941163
transform 1 0 16576 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1667941163
transform 1 0 20552 0 -1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1667941163
transform 1 0 2632 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1667941163
transform 1 0 6608 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1667941163
transform 1 0 10584 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1667941163
transform 1 0 14560 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1667941163
transform 1 0 18536 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1667941163
transform 1 0 22512 0 1 27440
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1667941163
transform 1 0 4648 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1667941163
transform 1 0 8624 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1667941163
transform 1 0 12600 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1667941163
transform 1 0 16576 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1667941163
transform 1 0 20552 0 -1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1667941163
transform 1 0 2632 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1667941163
transform 1 0 6608 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1667941163
transform 1 0 10584 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1667941163
transform 1 0 14560 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1667941163
transform 1 0 18536 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1667941163
transform 1 0 22512 0 1 28224
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1667941163
transform 1 0 4648 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1667941163
transform 1 0 8624 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1667941163
transform 1 0 12600 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1667941163
transform 1 0 16576 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1667941163
transform 1 0 20552 0 -1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1667941163
transform 1 0 2632 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1667941163
transform 1 0 6608 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1667941163
transform 1 0 10584 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1667941163
transform 1 0 14560 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1667941163
transform 1 0 18536 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1667941163
transform 1 0 22512 0 1 29008
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1667941163
transform 1 0 4648 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1667941163
transform 1 0 8624 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1667941163
transform 1 0 12600 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1667941163
transform 1 0 16576 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1667941163
transform 1 0 20552 0 -1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1667941163
transform 1 0 2632 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1667941163
transform 1 0 6608 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1667941163
transform 1 0 10584 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1667941163
transform 1 0 14560 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1667941163
transform 1 0 18536 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1667941163
transform 1 0 22512 0 1 29792
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1667941163
transform 1 0 4648 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1667941163
transform 1 0 8624 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1667941163
transform 1 0 12600 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1667941163
transform 1 0 16576 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1667941163
transform 1 0 20552 0 -1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1667941163
transform 1 0 2632 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1667941163
transform 1 0 6608 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1667941163
transform 1 0 10584 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1667941163
transform 1 0 14560 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1667941163
transform 1 0 18536 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1667941163
transform 1 0 22512 0 1 30576
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1667941163
transform 1 0 4648 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1667941163
transform 1 0 8624 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1667941163
transform 1 0 12600 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1667941163
transform 1 0 16576 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1667941163
transform 1 0 20552 0 -1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1667941163
transform 1 0 2632 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1667941163
transform 1 0 6608 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1667941163
transform 1 0 10584 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1667941163
transform 1 0 14560 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1667941163
transform 1 0 18536 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1667941163
transform 1 0 22512 0 1 31360
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1667941163
transform 1 0 4648 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1667941163
transform 1 0 8624 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1667941163
transform 1 0 12600 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1667941163
transform 1 0 16576 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1667941163
transform 1 0 20552 0 -1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1667941163
transform 1 0 2632 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1667941163
transform 1 0 6608 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1667941163
transform 1 0 10584 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1667941163
transform 1 0 14560 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1667941163
transform 1 0 18536 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1667941163
transform 1 0 22512 0 1 32144
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1667941163
transform 1 0 4648 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1667941163
transform 1 0 8624 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1667941163
transform 1 0 12600 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1667941163
transform 1 0 16576 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1667941163
transform 1 0 20552 0 -1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1667941163
transform 1 0 2632 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1667941163
transform 1 0 4592 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1667941163
transform 1 0 6552 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1667941163
transform 1 0 8512 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1667941163
transform 1 0 10472 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1667941163
transform 1 0 12432 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1667941163
transform 1 0 14392 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1667941163
transform 1 0 16352 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1667941163
transform 1 0 18312 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1667941163
transform 1 0 20272 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1667941163
transform 1 0 22232 0 1 32928
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 15568 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 12544 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 16072 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 13048 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 18088 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 11088 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 12992 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 10528 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyp1
timestamp 1667941163
transform 1 0 7728 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 15568 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 12992 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 15568 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyp1
timestamp 1667941163
transform -1 0 16072 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 13048 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 12544 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 13552 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyp1
timestamp 1667941163
transform -1 0 14504 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 16072 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyp1
timestamp 1667941163
transform -1 0 14504 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 16072 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 13048 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 12544 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyp1
timestamp 1667941163
transform 1 0 7728 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[16\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[16\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[17\].u_series_gyn1
timestamp 1667941163
transform -1 0 14504 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[17\].u_series_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[18\].u_series_gyn1
timestamp 1667941163
transform -1 0 11088 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[18\].u_series_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[19\].u_series_gyn1
timestamp 1667941163
transform -1 0 15568 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[19\].u_series_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[20\].u_series_gyn1
timestamp 1667941163
transform -1 0 16072 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[20\].u_series_gyp1
timestamp 1667941163
transform -1 0 19544 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[21\].u_series_gyn1
timestamp 1667941163
transform -1 0 13048 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[21\].u_series_gyp1
timestamp 1667941163
transform -1 0 19544 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[22\].u_series_gyn1
timestamp 1667941163
transform -1 0 12544 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[22\].u_series_gyp1
timestamp 1667941163
transform 1 0 7224 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[23\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[23\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[24\].u_series_gyn1
timestamp 1667941163
transform -1 0 16072 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[24\].u_series_gyp1
timestamp 1667941163
transform -1 0 14112 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[25\].u_series_gyn1
timestamp 1667941163
transform -1 0 13552 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[25\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[26\].u_series_gyn1
timestamp 1667941163
transform -1 0 14504 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[26\].u_series_gyp1
timestamp 1667941163
transform -1 0 19544 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[27\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[27\].u_series_gyp1
timestamp 1667941163
transform -1 0 20048 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[28\].u_series_gyn1
timestamp 1667941163
transform -1 0 17528 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[28\].u_series_gyp1
timestamp 1667941163
transform -1 0 20048 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[29\].u_series_gyn1
timestamp 1667941163
transform -1 0 15568 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[29\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[30\].u_series_gyn1
timestamp 1667941163
transform -1 0 12544 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[30\].u_series_gyp1
timestamp 1667941163
transform -1 0 16072 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[31\].u_series_gyn1
timestamp 1667941163
transform -1 0 17528 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[31\].u_series_gyp1
timestamp 1667941163
transform -1 0 14112 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 6552 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 18088 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 12376 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 9072 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 8568 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 16072 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 19544 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 7112 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyp1
timestamp 1667941163
transform 1 0 3752 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 20048 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 18088 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 9072 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyp1
timestamp 1667941163
transform 1 0 5768 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 8568 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 9072 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyn1
timestamp 1667941163
transform 1 0 5768 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 8568 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 10416 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyp1
timestamp 1667941163
transform 1 0 5208 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 8288 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyp1
timestamp 1667941163
transform 1 0 5768 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 8288 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyp1
timestamp 1667941163
transform 1 0 5208 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 4144 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 3864 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 14448 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[0\].u_series_gyp1
timestamp 1667941163
transform 1 0 5208 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 12544 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 10528 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 11088 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 8568 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 15568 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[3\].u_series_gyp1
timestamp 1667941163
transform 1 0 5768 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 10528 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 19544 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 17528 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 22064 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 18088 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 12544 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 14448 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 13944 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[8\].u_series_gyp1
timestamp 1667941163
transform -1 0 11088 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 9072 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 14112 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[10\].u_series_gyp1
timestamp 1667941163
transform -1 0 20048 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 16072 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[11\].u_series_gyp1
timestamp 1667941163
transform -1 0 16072 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 19544 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[12\].u_series_gyp1
timestamp 1667941163
transform -1 0 17528 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 17528 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 18088 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[14\].u_series_gyp1
timestamp 1667941163
transform -1 0 21504 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 20048 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[15\].u_series_gyp1
timestamp 1667941163
transform -1 0 15568 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 8176 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 9688 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 6776 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 6832 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 8288 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 6776 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 6776 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 4704 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 9688 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 9744 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 6048 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 8176 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 4312 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_n
timestamp 1667941163
transform -1 0 9688 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_n
timestamp 1667941163
transform -1 0 6776 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_n
timestamp 1667941163
transform -1 0 9576 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_n
timestamp 1667941163
transform -1 0 9744 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[64\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[64\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[65\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[65\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[66\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[66\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[67\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[67\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[68\].u_shunt_n
timestamp 1667941163
transform -1 0 9688 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[68\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[69\].u_shunt_n
timestamp 1667941163
transform -1 0 6720 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[69\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[70\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[70\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[71\].u_shunt_n
timestamp 1667941163
transform -1 0 8288 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[71\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[72\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[72\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[73\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[73\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[74\].u_shunt_n
timestamp 1667941163
transform -1 0 8288 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[74\].u_shunt_p
timestamp 1667941163
transform -1 0 4704 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[75\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[75\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[76\].u_shunt_n
timestamp 1667941163
transform -1 0 8176 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[76\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[77\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[77\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[78\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[78\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[79\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[79\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[80\].u_shunt_n
timestamp 1667941163
transform -1 0 9744 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[80\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[81\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[81\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[82\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[82\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[83\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[83\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[84\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[84\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[85\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[85\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[86\].u_shunt_n
timestamp 1667941163
transform -1 0 9632 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[86\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[87\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[87\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[88\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[88\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[89\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[89\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[90\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[90\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[91\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[91\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[92\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[92\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[93\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[93\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[94\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[94\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[95\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[95\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[96\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[96\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[97\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[97\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[98\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[98\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[99\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[99\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[100\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[100\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[101\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[101\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[102\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[102\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[103\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[103\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[104\].u_shunt_n
timestamp 1667941163
transform -1 0 9632 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[104\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[105\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[105\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[106\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[106\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[107\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[107\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[108\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[108\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[109\].u_shunt_n
timestamp 1667941163
transform -1 0 8288 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[109\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[110\].u_shunt_n
timestamp 1667941163
transform -1 0 6272 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[110\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[111\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[111\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[112\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[112\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[113\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[113\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[114\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[114\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[115\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[115\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[116\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[116\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[117\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[117\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[118\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[118\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[119\].u_shunt_n
timestamp 1667941163
transform -1 0 8288 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[119\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[120\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[120\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[121\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[121\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[122\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[122\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[123\].u_shunt_n
timestamp 1667941163
transform -1 0 8232 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[123\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[124\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[124\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[125\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[125\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[126\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[126\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[127\].u_shunt_n
timestamp 1667941163
transform -1 0 8176 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[127\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 7728 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 6272 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 12096 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 7728 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[48\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[48\].u_shunt_p
timestamp 1667941163
transform -1 0 7728 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[49\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[49\].u_shunt_p
timestamp 1667941163
transform -1 0 6272 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[50\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[50\].u_shunt_p
timestamp 1667941163
transform -1 0 6272 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[51\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[51\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[52\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[52\].u_shunt_p
timestamp 1667941163
transform -1 0 7728 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[53\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[53\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[54\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[54\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[55\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[55\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[56\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[56\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[57\].u_shunt_n
timestamp 1667941163
transform -1 0 9128 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[57\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[58\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[58\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[59\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[59\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[60\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[60\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[61\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[61\].u_shunt_p
timestamp 1667941163
transform -1 0 7728 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[62\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[62\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[63\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[63\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 28224
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 6160 0 -1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 28224
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 28224
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 8120 0 1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 5768 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 7616 0 -1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 29008
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 4312 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 4312 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 6160 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 10136 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 5768 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 5768 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 5208 0 1 28224
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 4312 0 1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 5208 0 1 29008
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 5768 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 6160 0 -1 29008
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 4312 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 28224
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 5768 0 1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 6160 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 14112 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 21168
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 19600
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 18816
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 15568 0 -1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 13552 0 1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 23520
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 14112 0 -1 25872
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 11592 0 -1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 11592 0 -1 26656
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 15568 0 -1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 10136 0 -1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 24304
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 22736
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 20384
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 21952
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 12096 0 1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 13552 0 1 25088
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 9576 0 1 27440
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 3640 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 3640 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 4144 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 4144 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 3640 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g8\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 2184 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g8\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 2184 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 22456 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 23408 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 21336 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23128 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 21448 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 23912 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 23352 0 -1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 22456 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 23912 0 -1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 22512 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 22848 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 21952 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 20328 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 21896 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 23968 0 1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 22512 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 21896 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 20944 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 22456 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23128 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 22456 0 1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 23408 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 22008 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 22568 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 23408 0 1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 21896 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 23968 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23352 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 22848 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 23408 0 1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 22288 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 22456 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 21728 0 -1 28224
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 23688 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 23968 0 1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23632 0 1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 21336 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 22624 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 21952 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23632 0 1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 21336 0 1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 23688 0 -1 27440
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 22792 0 -1 29008
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23632 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 19768 0 1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 22624 0 -1 25872
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 23632 0 -1 29792
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 23632 0 -1 26656
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 23688 0 -1 25088
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 23128 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 23688 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 23688 0 1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 23128 0 1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 23688 0 -1 23520
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 23688 0 -1 24304
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 23688 0 -1 22736
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_n
timestamp 1667941163
transform 1 0 23688 0 -1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_p
timestamp 1667941163
transform 1 0 23688 0 1 19600
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 21112 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 21336 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 21112 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 21336 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 22680 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 19656 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 22456 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 22680 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 22456 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 20496 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 22680 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 21000 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 22792 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 22792 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn3
timestamp 1667941163
transform 1 0 22792 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 22792 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 22792 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp3
timestamp 1667941163
transform 1 0 22792 0 -1 7056
box -43 -43 1387 435
<< labels >>
flabel metal2 s 23240 34600 23296 35000 0 FreeSans 224 90 0 0 cap_series_gygyn
port 0 nsew signal bidirectional
flabel metal2 s 20160 34600 20216 35000 0 FreeSans 224 90 0 0 cap_series_gygyp
port 1 nsew signal bidirectional
flabel metal2 s 17080 34600 17136 35000 0 FreeSans 224 90 0 0 cap_series_gyn
port 2 nsew signal bidirectional
flabel metal2 s 14000 34600 14056 35000 0 FreeSans 224 90 0 0 cap_series_gyp
port 3 nsew signal bidirectional
flabel metal2 s 10920 34600 10976 35000 0 FreeSans 224 90 0 0 cap_shunt_gyn
port 4 nsew signal bidirectional
flabel metal2 s 7840 34600 7896 35000 0 FreeSans 224 90 0 0 cap_shunt_gyp
port 5 nsew signal bidirectional
flabel metal2 s 4760 34600 4816 35000 0 FreeSans 224 90 0 0 cap_shunt_n
port 6 nsew signal bidirectional
flabel metal2 s 1680 34600 1736 35000 0 FreeSans 224 90 0 0 cap_shunt_p
port 7 nsew signal bidirectional
flabel metal2 s 2072 0 2128 400 0 FreeSans 224 90 0 0 tune_series_gy[0]
port 8 nsew signal input
flabel metal2 s 6216 0 6272 400 0 FreeSans 224 90 0 0 tune_series_gy[1]
port 9 nsew signal input
flabel metal2 s 10360 0 10416 400 0 FreeSans 224 90 0 0 tune_series_gy[2]
port 10 nsew signal input
flabel metal2 s 14504 0 14560 400 0 FreeSans 224 90 0 0 tune_series_gy[3]
port 11 nsew signal input
flabel metal2 s 18648 0 18704 400 0 FreeSans 224 90 0 0 tune_series_gy[4]
port 12 nsew signal input
flabel metal2 s 22792 0 22848 400 0 FreeSans 224 90 0 0 tune_series_gy[5]
port 13 nsew signal input
flabel metal3 s 24600 1344 25000 1400 0 FreeSans 224 0 0 0 tune_series_gygy[0]
port 14 nsew signal input
flabel metal3 s 24600 4032 25000 4088 0 FreeSans 224 0 0 0 tune_series_gygy[1]
port 15 nsew signal input
flabel metal3 s 24600 6720 25000 6776 0 FreeSans 224 0 0 0 tune_series_gygy[2]
port 16 nsew signal input
flabel metal3 s 24600 9408 25000 9464 0 FreeSans 224 0 0 0 tune_series_gygy[3]
port 17 nsew signal input
flabel metal3 s 24600 12096 25000 12152 0 FreeSans 224 0 0 0 tune_series_gygy[4]
port 18 nsew signal input
flabel metal3 s 24600 14784 25000 14840 0 FreeSans 224 0 0 0 tune_series_gygy[5]
port 19 nsew signal input
flabel metal3 s 0 2184 400 2240 0 FreeSans 224 0 0 0 tune_shunt[0]
port 20 nsew signal input
flabel metal3 s 0 6552 400 6608 0 FreeSans 224 0 0 0 tune_shunt[1]
port 21 nsew signal input
flabel metal3 s 0 10920 400 10976 0 FreeSans 224 0 0 0 tune_shunt[2]
port 22 nsew signal input
flabel metal3 s 0 15288 400 15344 0 FreeSans 224 0 0 0 tune_shunt[3]
port 23 nsew signal input
flabel metal3 s 0 19656 400 19712 0 FreeSans 224 0 0 0 tune_shunt[4]
port 24 nsew signal input
flabel metal3 s 0 24024 400 24080 0 FreeSans 224 0 0 0 tune_shunt[5]
port 25 nsew signal input
flabel metal3 s 0 28392 400 28448 0 FreeSans 224 0 0 0 tune_shunt[6]
port 26 nsew signal input
flabel metal3 s 0 32760 400 32816 0 FreeSans 224 0 0 0 tune_shunt[7]
port 27 nsew signal input
flabel metal3 s 24600 17472 25000 17528 0 FreeSans 224 0 0 0 tune_shunt_gy[0]
port 28 nsew signal input
flabel metal3 s 24600 20160 25000 20216 0 FreeSans 224 0 0 0 tune_shunt_gy[1]
port 29 nsew signal input
flabel metal3 s 24600 22848 25000 22904 0 FreeSans 224 0 0 0 tune_shunt_gy[2]
port 30 nsew signal input
flabel metal3 s 24600 25536 25000 25592 0 FreeSans 224 0 0 0 tune_shunt_gy[3]
port 31 nsew signal input
flabel metal3 s 24600 28224 25000 28280 0 FreeSans 224 0 0 0 tune_shunt_gy[4]
port 32 nsew signal input
flabel metal3 s 24600 30912 25000 30968 0 FreeSans 224 0 0 0 tune_shunt_gy[5]
port 33 nsew signal input
flabel metal3 s 24600 33600 25000 33656 0 FreeSans 224 0 0 0 tune_shunt_gy[6]
port 34 nsew signal input
flabel metal4 s 2224 1538 2384 33350 0 FreeSans 640 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 17584 1538 17744 33350 0 FreeSans 640 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 9904 1538 10064 33350 0 FreeSans 640 90 0 0 vss
port 36 nsew ground bidirectional
rlabel metal1 12488 33320 12488 33320 0 vdd
rlabel metal1 12488 32928 12488 32928 0 vss
rlabel metal2 22932 4088 22932 4088 0 cap_series_gygyn
rlabel metal2 22876 14336 22876 14336 0 cap_series_gygyp
rlabel metal2 3836 1736 3836 1736 0 cap_series_gyn
rlabel metal2 3780 2380 3780 2380 0 cap_series_gyp
rlabel metal2 22708 26684 22708 26684 0 cap_shunt_gyn
rlabel metal2 23828 22540 23828 22540 0 cap_shunt_gyp
rlabel metal2 2128 2548 2128 2548 0 cap_shunt_n
rlabel metal2 1876 2968 1876 2968 0 cap_shunt_p
rlabel metal3 2492 1764 2492 1764 0 tune_series_gy[0]
rlabel metal2 6244 1463 6244 1463 0 tune_series_gy[1]
rlabel metal2 10388 1071 10388 1071 0 tune_series_gy[2]
rlabel metal2 11116 1904 11116 1904 0 tune_series_gy[3]
rlabel via2 15092 3724 15092 3724 0 tune_series_gy[4]
rlabel metal2 11788 2940 11788 2940 0 tune_series_gy[5]
rlabel metal2 24052 2744 24052 2744 0 tune_series_gygy[0]
rlabel metal3 24241 4060 24241 4060 0 tune_series_gygy[1]
rlabel metal2 24052 7196 24052 7196 0 tune_series_gygy[2]
rlabel metal3 19740 10052 19740 10052 0 tune_series_gygy[3]
rlabel metal3 24241 12124 24241 12124 0 tune_series_gygy[4]
rlabel metal2 24052 14560 24052 14560 0 tune_series_gygy[5]
rlabel metal2 924 2380 924 2380 0 tune_shunt[0]
rlabel metal2 1036 3920 1036 3920 0 tune_shunt[1]
rlabel metal3 1043 10948 1043 10948 0 tune_shunt[2]
rlabel metal3 1155 15316 1155 15316 0 tune_shunt[3]
rlabel metal2 15092 23324 15092 23324 0 tune_shunt[4]
rlabel metal3 1624 14700 1624 14700 0 tune_shunt[5]
rlabel metal2 1848 22540 1848 22540 0 tune_shunt[6]
rlabel metal2 3724 15484 3724 15484 0 tune_shunt[7]
rlabel metal2 24052 18452 24052 18452 0 tune_shunt_gy[0]
rlabel metal2 23520 22876 23520 22876 0 tune_shunt_gy[1]
rlabel metal2 24052 23492 24052 23492 0 tune_shunt_gy[2]
rlabel metal2 23324 25620 23324 25620 0 tune_shunt_gy[3]
rlabel metal2 23604 28868 23604 28868 0 tune_shunt_gy[4]
rlabel metal2 22764 27048 22764 27048 0 tune_shunt_gy[5]
rlabel metal2 22148 25116 22148 25116 0 tune_shunt_gy[6]
<< properties >>
string FIXED_BBOX 0 0 25000 35000
<< end >>
