magic
tech gf180mcuC
magscale 1 10
timestamp 1669999162
<< metal2 >>
rect 388000 -17191 397200 -17070
rect 388000 -17247 388146 -17191
rect 388202 -17247 388270 -17191
rect 388326 -17247 388394 -17191
rect 388450 -17247 388518 -17191
rect 388574 -17247 388642 -17191
rect 388698 -17247 388766 -17191
rect 388822 -17247 388890 -17191
rect 388946 -17247 389014 -17191
rect 389070 -17247 389138 -17191
rect 389194 -17247 389262 -17191
rect 389318 -17247 389386 -17191
rect 389442 -17247 389510 -17191
rect 389566 -17247 389634 -17191
rect 389690 -17247 389758 -17191
rect 389814 -17247 389882 -17191
rect 389938 -17247 390006 -17191
rect 390062 -17247 390130 -17191
rect 390186 -17247 390254 -17191
rect 390310 -17247 390378 -17191
rect 390434 -17247 390502 -17191
rect 390558 -17247 390626 -17191
rect 390682 -17247 390750 -17191
rect 390806 -17247 390874 -17191
rect 390930 -17247 390998 -17191
rect 391054 -17247 391122 -17191
rect 391178 -17247 391246 -17191
rect 391302 -17247 391370 -17191
rect 391426 -17247 391494 -17191
rect 391550 -17247 391618 -17191
rect 391674 -17247 391742 -17191
rect 391798 -17247 391866 -17191
rect 391922 -17247 391990 -17191
rect 392046 -17247 392114 -17191
rect 392170 -17247 392238 -17191
rect 392294 -17247 392362 -17191
rect 392418 -17247 392486 -17191
rect 392542 -17247 392610 -17191
rect 392666 -17247 392734 -17191
rect 392790 -17247 392858 -17191
rect 392914 -17247 392982 -17191
rect 393038 -17247 393106 -17191
rect 393162 -17247 393230 -17191
rect 393286 -17247 393354 -17191
rect 393410 -17247 393478 -17191
rect 393534 -17247 393602 -17191
rect 393658 -17247 393726 -17191
rect 393782 -17247 393850 -17191
rect 393906 -17247 393974 -17191
rect 394030 -17247 394098 -17191
rect 394154 -17247 394222 -17191
rect 394278 -17247 394346 -17191
rect 394402 -17247 394470 -17191
rect 394526 -17247 394594 -17191
rect 394650 -17247 394718 -17191
rect 394774 -17247 394842 -17191
rect 394898 -17247 394966 -17191
rect 395022 -17247 395090 -17191
rect 395146 -17247 395214 -17191
rect 395270 -17247 395338 -17191
rect 395394 -17247 395462 -17191
rect 395518 -17247 395586 -17191
rect 395642 -17247 395710 -17191
rect 395766 -17247 395898 -17191
rect 395954 -17247 396022 -17191
rect 396078 -17247 396146 -17191
rect 396202 -17247 396270 -17191
rect 396326 -17247 396394 -17191
rect 396450 -17247 396518 -17191
rect 396574 -17247 396642 -17191
rect 396698 -17247 396766 -17191
rect 396822 -17247 396890 -17191
rect 396946 -17247 397014 -17191
rect 397070 -17247 397200 -17191
rect 388000 -17315 397200 -17247
rect 388000 -17371 388146 -17315
rect 388202 -17371 388270 -17315
rect 388326 -17371 388394 -17315
rect 388450 -17371 388518 -17315
rect 388574 -17371 388642 -17315
rect 388698 -17371 388766 -17315
rect 388822 -17371 388890 -17315
rect 388946 -17371 389014 -17315
rect 389070 -17371 389138 -17315
rect 389194 -17371 389262 -17315
rect 389318 -17371 389386 -17315
rect 389442 -17371 389510 -17315
rect 389566 -17371 389634 -17315
rect 389690 -17371 389758 -17315
rect 389814 -17371 389882 -17315
rect 389938 -17371 390006 -17315
rect 390062 -17371 390130 -17315
rect 390186 -17371 390254 -17315
rect 390310 -17371 390378 -17315
rect 390434 -17371 390502 -17315
rect 390558 -17371 390626 -17315
rect 390682 -17371 390750 -17315
rect 390806 -17371 390874 -17315
rect 390930 -17371 390998 -17315
rect 391054 -17371 391122 -17315
rect 391178 -17371 391246 -17315
rect 391302 -17371 391370 -17315
rect 391426 -17371 391494 -17315
rect 391550 -17371 391618 -17315
rect 391674 -17371 391742 -17315
rect 391798 -17371 391866 -17315
rect 391922 -17371 391990 -17315
rect 392046 -17371 392114 -17315
rect 392170 -17371 392238 -17315
rect 392294 -17371 392362 -17315
rect 392418 -17371 392486 -17315
rect 392542 -17371 392610 -17315
rect 392666 -17371 392734 -17315
rect 392790 -17371 392858 -17315
rect 392914 -17371 392982 -17315
rect 393038 -17371 393106 -17315
rect 393162 -17371 393230 -17315
rect 393286 -17371 393354 -17315
rect 393410 -17371 393478 -17315
rect 393534 -17371 393602 -17315
rect 393658 -17371 393726 -17315
rect 393782 -17371 393850 -17315
rect 393906 -17371 393974 -17315
rect 394030 -17371 394098 -17315
rect 394154 -17371 394222 -17315
rect 394278 -17371 394346 -17315
rect 394402 -17371 394470 -17315
rect 394526 -17371 394594 -17315
rect 394650 -17371 394718 -17315
rect 394774 -17371 394842 -17315
rect 394898 -17371 394966 -17315
rect 395022 -17371 395090 -17315
rect 395146 -17371 395214 -17315
rect 395270 -17371 395338 -17315
rect 395394 -17371 395462 -17315
rect 395518 -17371 395586 -17315
rect 395642 -17371 395710 -17315
rect 395766 -17371 395898 -17315
rect 395954 -17371 396022 -17315
rect 396078 -17371 396146 -17315
rect 396202 -17371 396270 -17315
rect 396326 -17371 396394 -17315
rect 396450 -17371 396518 -17315
rect 396574 -17371 396642 -17315
rect 396698 -17371 396766 -17315
rect 396822 -17371 396890 -17315
rect 396946 -17371 397014 -17315
rect 397070 -17371 397200 -17315
rect 388000 -17439 397200 -17371
rect 388000 -17495 388146 -17439
rect 388202 -17495 388270 -17439
rect 388326 -17495 388394 -17439
rect 388450 -17495 388518 -17439
rect 388574 -17495 388642 -17439
rect 388698 -17495 388766 -17439
rect 388822 -17495 388890 -17439
rect 388946 -17495 389014 -17439
rect 389070 -17495 389138 -17439
rect 389194 -17495 389262 -17439
rect 389318 -17495 389386 -17439
rect 389442 -17495 389510 -17439
rect 389566 -17495 389634 -17439
rect 389690 -17495 389758 -17439
rect 389814 -17495 389882 -17439
rect 389938 -17495 390006 -17439
rect 390062 -17495 390130 -17439
rect 390186 -17495 390254 -17439
rect 390310 -17495 390378 -17439
rect 390434 -17495 390502 -17439
rect 390558 -17495 390626 -17439
rect 390682 -17495 390750 -17439
rect 390806 -17495 390874 -17439
rect 390930 -17495 390998 -17439
rect 391054 -17495 391122 -17439
rect 391178 -17495 391246 -17439
rect 391302 -17495 391370 -17439
rect 391426 -17495 391494 -17439
rect 391550 -17495 391618 -17439
rect 391674 -17495 391742 -17439
rect 391798 -17495 391866 -17439
rect 391922 -17495 391990 -17439
rect 392046 -17495 392114 -17439
rect 392170 -17495 392238 -17439
rect 392294 -17495 392362 -17439
rect 392418 -17495 392486 -17439
rect 392542 -17495 392610 -17439
rect 392666 -17495 392734 -17439
rect 392790 -17495 392858 -17439
rect 392914 -17495 392982 -17439
rect 393038 -17495 393106 -17439
rect 393162 -17495 393230 -17439
rect 393286 -17495 393354 -17439
rect 393410 -17495 393478 -17439
rect 393534 -17495 393602 -17439
rect 393658 -17495 393726 -17439
rect 393782 -17495 393850 -17439
rect 393906 -17495 393974 -17439
rect 394030 -17495 394098 -17439
rect 394154 -17495 394222 -17439
rect 394278 -17495 394346 -17439
rect 394402 -17495 394470 -17439
rect 394526 -17495 394594 -17439
rect 394650 -17495 394718 -17439
rect 394774 -17495 394842 -17439
rect 394898 -17495 394966 -17439
rect 395022 -17495 395090 -17439
rect 395146 -17495 395214 -17439
rect 395270 -17495 395338 -17439
rect 395394 -17495 395462 -17439
rect 395518 -17495 395586 -17439
rect 395642 -17495 395710 -17439
rect 395766 -17495 395898 -17439
rect 395954 -17495 396022 -17439
rect 396078 -17495 396146 -17439
rect 396202 -17495 396270 -17439
rect 396326 -17495 396394 -17439
rect 396450 -17495 396518 -17439
rect 396574 -17495 396642 -17439
rect 396698 -17495 396766 -17439
rect 396822 -17495 396890 -17439
rect 396946 -17495 397014 -17439
rect 397070 -17495 397200 -17439
rect 388000 -17563 397200 -17495
rect 388000 -17619 388146 -17563
rect 388202 -17619 388270 -17563
rect 388326 -17619 388394 -17563
rect 388450 -17619 388518 -17563
rect 388574 -17619 388642 -17563
rect 388698 -17619 388766 -17563
rect 388822 -17619 388890 -17563
rect 388946 -17619 389014 -17563
rect 389070 -17619 389138 -17563
rect 389194 -17619 389262 -17563
rect 389318 -17619 389386 -17563
rect 389442 -17619 389510 -17563
rect 389566 -17619 389634 -17563
rect 389690 -17619 389758 -17563
rect 389814 -17619 389882 -17563
rect 389938 -17619 390006 -17563
rect 390062 -17619 390130 -17563
rect 390186 -17619 390254 -17563
rect 390310 -17619 390378 -17563
rect 390434 -17619 390502 -17563
rect 390558 -17619 390626 -17563
rect 390682 -17619 390750 -17563
rect 390806 -17619 390874 -17563
rect 390930 -17619 390998 -17563
rect 391054 -17619 391122 -17563
rect 391178 -17619 391246 -17563
rect 391302 -17619 391370 -17563
rect 391426 -17619 391494 -17563
rect 391550 -17619 391618 -17563
rect 391674 -17619 391742 -17563
rect 391798 -17619 391866 -17563
rect 391922 -17619 391990 -17563
rect 392046 -17619 392114 -17563
rect 392170 -17619 392238 -17563
rect 392294 -17619 392362 -17563
rect 392418 -17619 392486 -17563
rect 392542 -17619 392610 -17563
rect 392666 -17619 392734 -17563
rect 392790 -17619 392858 -17563
rect 392914 -17619 392982 -17563
rect 393038 -17619 393106 -17563
rect 393162 -17619 393230 -17563
rect 393286 -17619 393354 -17563
rect 393410 -17619 393478 -17563
rect 393534 -17619 393602 -17563
rect 393658 -17619 393726 -17563
rect 393782 -17619 393850 -17563
rect 393906 -17619 393974 -17563
rect 394030 -17619 394098 -17563
rect 394154 -17619 394222 -17563
rect 394278 -17619 394346 -17563
rect 394402 -17619 394470 -17563
rect 394526 -17619 394594 -17563
rect 394650 -17619 394718 -17563
rect 394774 -17619 394842 -17563
rect 394898 -17619 394966 -17563
rect 395022 -17619 395090 -17563
rect 395146 -17619 395214 -17563
rect 395270 -17619 395338 -17563
rect 395394 -17619 395462 -17563
rect 395518 -17619 395586 -17563
rect 395642 -17619 395710 -17563
rect 395766 -17619 395898 -17563
rect 395954 -17619 396022 -17563
rect 396078 -17619 396146 -17563
rect 396202 -17619 396270 -17563
rect 396326 -17619 396394 -17563
rect 396450 -17619 396518 -17563
rect 396574 -17619 396642 -17563
rect 396698 -17619 396766 -17563
rect 396822 -17619 396890 -17563
rect 396946 -17619 397014 -17563
rect 397070 -17619 397200 -17563
rect 388000 -17740 397200 -17619
rect 388000 -17858 388800 -17740
rect 388000 -17914 388114 -17858
rect 388170 -17914 388238 -17858
rect 388294 -17914 388362 -17858
rect 388418 -17914 388486 -17858
rect 388542 -17914 388610 -17858
rect 388666 -17914 388800 -17858
rect 388000 -17982 388800 -17914
rect 388000 -18038 388114 -17982
rect 388170 -18038 388238 -17982
rect 388294 -18038 388362 -17982
rect 388418 -18038 388486 -17982
rect 388542 -18038 388610 -17982
rect 388666 -18038 388800 -17982
rect 388000 -18106 388800 -18038
rect 388000 -18162 388114 -18106
rect 388170 -18162 388238 -18106
rect 388294 -18162 388362 -18106
rect 388418 -18162 388486 -18106
rect 388542 -18162 388610 -18106
rect 388666 -18162 388800 -18106
rect 388000 -18230 388800 -18162
rect 388000 -18286 388114 -18230
rect 388170 -18286 388238 -18230
rect 388294 -18286 388362 -18230
rect 388418 -18286 388486 -18230
rect 388542 -18286 388610 -18230
rect 388666 -18286 388800 -18230
rect 388000 -18354 388800 -18286
rect 388000 -18410 388114 -18354
rect 388170 -18410 388238 -18354
rect 388294 -18410 388362 -18354
rect 388418 -18410 388486 -18354
rect 388542 -18410 388610 -18354
rect 388666 -18410 388800 -18354
rect 388000 -18478 388800 -18410
rect 388000 -18534 388114 -18478
rect 388170 -18534 388238 -18478
rect 388294 -18534 388362 -18478
rect 388418 -18534 388486 -18478
rect 388542 -18534 388610 -18478
rect 388666 -18534 388800 -18478
rect 388000 -18602 388800 -18534
rect 388000 -18658 388114 -18602
rect 388170 -18658 388238 -18602
rect 388294 -18658 388362 -18602
rect 388418 -18658 388486 -18602
rect 388542 -18658 388610 -18602
rect 388666 -18658 388800 -18602
rect 388000 -18726 388800 -18658
rect 388000 -18782 388114 -18726
rect 388170 -18782 388238 -18726
rect 388294 -18782 388362 -18726
rect 388418 -18782 388486 -18726
rect 388542 -18782 388610 -18726
rect 388666 -18782 388800 -18726
rect 388000 -18850 388800 -18782
rect 388000 -18906 388114 -18850
rect 388170 -18906 388238 -18850
rect 388294 -18906 388362 -18850
rect 388418 -18906 388486 -18850
rect 388542 -18906 388610 -18850
rect 388666 -18906 388800 -18850
rect 388000 -18974 388800 -18906
rect 388000 -19030 388114 -18974
rect 388170 -19030 388238 -18974
rect 388294 -19030 388362 -18974
rect 388418 -19030 388486 -18974
rect 388542 -19030 388610 -18974
rect 388666 -19030 388800 -18974
rect 388000 -19098 388800 -19030
rect 388000 -19154 388114 -19098
rect 388170 -19154 388238 -19098
rect 388294 -19154 388362 -19098
rect 388418 -19154 388486 -19098
rect 388542 -19154 388610 -19098
rect 388666 -19154 388800 -19098
rect 388000 -19222 388800 -19154
rect 388000 -19278 388114 -19222
rect 388170 -19278 388238 -19222
rect 388294 -19278 388362 -19222
rect 388418 -19278 388486 -19222
rect 388542 -19278 388610 -19222
rect 388666 -19278 388800 -19222
rect 388000 -19346 388800 -19278
rect 388000 -19402 388114 -19346
rect 388170 -19402 388238 -19346
rect 388294 -19402 388362 -19346
rect 388418 -19402 388486 -19346
rect 388542 -19402 388610 -19346
rect 388666 -19402 388800 -19346
rect 388000 -19470 388800 -19402
rect 388000 -19526 388114 -19470
rect 388170 -19526 388238 -19470
rect 388294 -19526 388362 -19470
rect 388418 -19526 388486 -19470
rect 388542 -19526 388610 -19470
rect 388666 -19526 388800 -19470
rect 388000 -19594 388800 -19526
rect 388000 -19650 388114 -19594
rect 388170 -19650 388238 -19594
rect 388294 -19650 388362 -19594
rect 388418 -19650 388486 -19594
rect 388542 -19650 388610 -19594
rect 388666 -19650 388800 -19594
rect 388000 -19718 388800 -19650
rect 388000 -19774 388114 -19718
rect 388170 -19774 388238 -19718
rect 388294 -19774 388362 -19718
rect 388418 -19774 388486 -19718
rect 388542 -19774 388610 -19718
rect 388666 -19774 388800 -19718
rect 388000 -19842 388800 -19774
rect 388000 -19898 388114 -19842
rect 388170 -19898 388238 -19842
rect 388294 -19898 388362 -19842
rect 388418 -19898 388486 -19842
rect 388542 -19898 388610 -19842
rect 388666 -19898 388800 -19842
rect 388000 -19966 388800 -19898
rect 388000 -20022 388114 -19966
rect 388170 -20022 388238 -19966
rect 388294 -20022 388362 -19966
rect 388418 -20022 388486 -19966
rect 388542 -20022 388610 -19966
rect 388666 -20022 388800 -19966
rect 388000 -20090 388800 -20022
rect 388000 -20146 388114 -20090
rect 388170 -20146 388238 -20090
rect 388294 -20146 388362 -20090
rect 388418 -20146 388486 -20090
rect 388542 -20146 388610 -20090
rect 388666 -20146 388800 -20090
rect 388000 -20214 388800 -20146
rect 388000 -20270 388114 -20214
rect 388170 -20270 388238 -20214
rect 388294 -20270 388362 -20214
rect 388418 -20270 388486 -20214
rect 388542 -20270 388610 -20214
rect 388666 -20270 388800 -20214
rect 388000 -20338 388800 -20270
rect 388000 -20394 388114 -20338
rect 388170 -20394 388238 -20338
rect 388294 -20394 388362 -20338
rect 388418 -20394 388486 -20338
rect 388542 -20394 388610 -20338
rect 388666 -20394 388800 -20338
rect 388000 -20462 388800 -20394
rect 388000 -20518 388114 -20462
rect 388170 -20518 388238 -20462
rect 388294 -20518 388362 -20462
rect 388418 -20518 388486 -20462
rect 388542 -20518 388610 -20462
rect 388666 -20518 388800 -20462
rect 388000 -20586 388800 -20518
rect 388000 -20642 388114 -20586
rect 388170 -20642 388238 -20586
rect 388294 -20642 388362 -20586
rect 388418 -20642 388486 -20586
rect 388542 -20642 388610 -20586
rect 388666 -20642 388800 -20586
rect 388000 -20710 388800 -20642
rect 388000 -20766 388114 -20710
rect 388170 -20766 388238 -20710
rect 388294 -20766 388362 -20710
rect 388418 -20766 388486 -20710
rect 388542 -20766 388610 -20710
rect 388666 -20766 388800 -20710
rect 388000 -20834 388800 -20766
rect 388000 -20890 388114 -20834
rect 388170 -20890 388238 -20834
rect 388294 -20890 388362 -20834
rect 388418 -20890 388486 -20834
rect 388542 -20890 388610 -20834
rect 388666 -20890 388800 -20834
rect 388000 -20958 388800 -20890
rect 388000 -21014 388114 -20958
rect 388170 -21014 388238 -20958
rect 388294 -21014 388362 -20958
rect 388418 -21014 388486 -20958
rect 388542 -21014 388610 -20958
rect 388666 -21014 388800 -20958
rect 388000 -21082 388800 -21014
rect 388000 -21138 388114 -21082
rect 388170 -21138 388238 -21082
rect 388294 -21138 388362 -21082
rect 388418 -21138 388486 -21082
rect 388542 -21138 388610 -21082
rect 388666 -21138 388800 -21082
rect 388000 -21206 388800 -21138
rect 388000 -21262 388114 -21206
rect 388170 -21262 388238 -21206
rect 388294 -21262 388362 -21206
rect 388418 -21262 388486 -21206
rect 388542 -21262 388610 -21206
rect 388666 -21262 388800 -21206
rect 388000 -21330 388800 -21262
rect 388000 -21386 388114 -21330
rect 388170 -21386 388238 -21330
rect 388294 -21386 388362 -21330
rect 388418 -21386 388486 -21330
rect 388542 -21386 388610 -21330
rect 388666 -21386 388800 -21330
rect 388000 -21454 388800 -21386
rect 388000 -21510 388114 -21454
rect 388170 -21510 388238 -21454
rect 388294 -21510 388362 -21454
rect 388418 -21510 388486 -21454
rect 388542 -21510 388610 -21454
rect 388666 -21510 388800 -21454
rect 388000 -21578 388800 -21510
rect 388000 -21634 388114 -21578
rect 388170 -21634 388238 -21578
rect 388294 -21634 388362 -21578
rect 388418 -21634 388486 -21578
rect 388542 -21634 388610 -21578
rect 388666 -21634 388800 -21578
rect 388000 -21702 388800 -21634
rect 388000 -21758 388114 -21702
rect 388170 -21758 388238 -21702
rect 388294 -21758 388362 -21702
rect 388418 -21758 388486 -21702
rect 388542 -21758 388610 -21702
rect 388666 -21758 388800 -21702
rect 388000 -21826 388800 -21758
rect 388000 -21882 388114 -21826
rect 388170 -21882 388238 -21826
rect 388294 -21882 388362 -21826
rect 388418 -21882 388486 -21826
rect 388542 -21882 388610 -21826
rect 388666 -21882 388800 -21826
rect 388000 -21950 388800 -21882
rect 388000 -22006 388114 -21950
rect 388170 -22006 388238 -21950
rect 388294 -22006 388362 -21950
rect 388418 -22006 388486 -21950
rect 388542 -22006 388610 -21950
rect 388666 -22006 388800 -21950
rect 388000 -22074 388800 -22006
rect 388000 -22130 388114 -22074
rect 388170 -22130 388238 -22074
rect 388294 -22130 388362 -22074
rect 388418 -22130 388486 -22074
rect 388542 -22130 388610 -22074
rect 388666 -22130 388800 -22074
rect 388000 -22198 388800 -22130
rect 388000 -22254 388114 -22198
rect 388170 -22254 388238 -22198
rect 388294 -22254 388362 -22198
rect 388418 -22254 388486 -22198
rect 388542 -22254 388610 -22198
rect 388666 -22254 388800 -22198
rect 388000 -22322 388800 -22254
rect 388000 -22378 388114 -22322
rect 388170 -22378 388238 -22322
rect 388294 -22378 388362 -22322
rect 388418 -22378 388486 -22322
rect 388542 -22378 388610 -22322
rect 388666 -22378 388800 -22322
rect 388000 -22446 388800 -22378
rect 388000 -22502 388114 -22446
rect 388170 -22502 388238 -22446
rect 388294 -22502 388362 -22446
rect 388418 -22502 388486 -22446
rect 388542 -22502 388610 -22446
rect 388666 -22502 388800 -22446
rect 388000 -22570 388800 -22502
rect 388000 -22626 388114 -22570
rect 388170 -22626 388238 -22570
rect 388294 -22626 388362 -22570
rect 388418 -22626 388486 -22570
rect 388542 -22626 388610 -22570
rect 388666 -22626 388800 -22570
rect 388000 -22694 388800 -22626
rect 388000 -22750 388114 -22694
rect 388170 -22750 388238 -22694
rect 388294 -22750 388362 -22694
rect 388418 -22750 388486 -22694
rect 388542 -22750 388610 -22694
rect 388666 -22750 388800 -22694
rect 388000 -22818 388800 -22750
rect 388000 -22874 388114 -22818
rect 388170 -22874 388238 -22818
rect 388294 -22874 388362 -22818
rect 388418 -22874 388486 -22818
rect 388542 -22874 388610 -22818
rect 388666 -22874 388800 -22818
rect 388000 -22942 388800 -22874
rect 388000 -22998 388114 -22942
rect 388170 -22998 388238 -22942
rect 388294 -22998 388362 -22942
rect 388418 -22998 388486 -22942
rect 388542 -22998 388610 -22942
rect 388666 -22998 388800 -22942
rect 388000 -23066 388800 -22998
rect 388000 -23122 388114 -23066
rect 388170 -23122 388238 -23066
rect 388294 -23122 388362 -23066
rect 388418 -23122 388486 -23066
rect 388542 -23122 388610 -23066
rect 388666 -23122 388800 -23066
rect 388000 -23190 388800 -23122
rect 388000 -23246 388114 -23190
rect 388170 -23246 388238 -23190
rect 388294 -23246 388362 -23190
rect 388418 -23246 388486 -23190
rect 388542 -23246 388610 -23190
rect 388666 -23246 388800 -23190
rect 388000 -23314 388800 -23246
rect 388000 -23370 388114 -23314
rect 388170 -23370 388238 -23314
rect 388294 -23370 388362 -23314
rect 388418 -23370 388486 -23314
rect 388542 -23370 388610 -23314
rect 388666 -23370 388800 -23314
rect 388000 -23438 388800 -23370
rect 388000 -23494 388114 -23438
rect 388170 -23494 388238 -23438
rect 388294 -23494 388362 -23438
rect 388418 -23494 388486 -23438
rect 388542 -23494 388610 -23438
rect 388666 -23494 388800 -23438
rect 388000 -23562 388800 -23494
rect 388000 -23618 388114 -23562
rect 388170 -23618 388238 -23562
rect 388294 -23618 388362 -23562
rect 388418 -23618 388486 -23562
rect 388542 -23618 388610 -23562
rect 388666 -23618 388800 -23562
rect 388000 -23686 388800 -23618
rect 388000 -23742 388114 -23686
rect 388170 -23742 388238 -23686
rect 388294 -23742 388362 -23686
rect 388418 -23742 388486 -23686
rect 388542 -23742 388610 -23686
rect 388666 -23742 388800 -23686
rect 388000 -23810 388800 -23742
rect 388000 -23866 388114 -23810
rect 388170 -23866 388238 -23810
rect 388294 -23866 388362 -23810
rect 388418 -23866 388486 -23810
rect 388542 -23866 388610 -23810
rect 388666 -23866 388800 -23810
rect 388000 -23934 388800 -23866
rect 388000 -23990 388114 -23934
rect 388170 -23990 388238 -23934
rect 388294 -23990 388362 -23934
rect 388418 -23990 388486 -23934
rect 388542 -23990 388610 -23934
rect 388666 -23990 388800 -23934
rect 388000 -24058 388800 -23990
rect 388000 -24114 388114 -24058
rect 388170 -24114 388238 -24058
rect 388294 -24114 388362 -24058
rect 388418 -24114 388486 -24058
rect 388542 -24114 388610 -24058
rect 388666 -24114 388800 -24058
rect 388000 -24182 388800 -24114
rect 388000 -24238 388114 -24182
rect 388170 -24238 388238 -24182
rect 388294 -24238 388362 -24182
rect 388418 -24238 388486 -24182
rect 388542 -24238 388610 -24182
rect 388666 -24238 388800 -24182
rect 388000 -24306 388800 -24238
rect 388000 -24362 388114 -24306
rect 388170 -24362 388238 -24306
rect 388294 -24362 388362 -24306
rect 388418 -24362 388486 -24306
rect 388542 -24362 388610 -24306
rect 388666 -24362 388800 -24306
rect 388000 -24430 388800 -24362
rect 388000 -24486 388114 -24430
rect 388170 -24486 388238 -24430
rect 388294 -24486 388362 -24430
rect 388418 -24486 388486 -24430
rect 388542 -24486 388610 -24430
rect 388666 -24486 388800 -24430
rect 388000 -24554 388800 -24486
rect 388000 -24610 388114 -24554
rect 388170 -24610 388238 -24554
rect 388294 -24610 388362 -24554
rect 388418 -24610 388486 -24554
rect 388542 -24610 388610 -24554
rect 388666 -24610 388800 -24554
rect 388000 -24678 388800 -24610
rect 388000 -24734 388114 -24678
rect 388170 -24734 388238 -24678
rect 388294 -24734 388362 -24678
rect 388418 -24734 388486 -24678
rect 388542 -24734 388610 -24678
rect 388666 -24734 388800 -24678
rect 388000 -24802 388800 -24734
rect 388000 -24858 388114 -24802
rect 388170 -24858 388238 -24802
rect 388294 -24858 388362 -24802
rect 388418 -24858 388486 -24802
rect 388542 -24858 388610 -24802
rect 388666 -24858 388800 -24802
rect 388000 -24926 388800 -24858
rect 388000 -24982 388114 -24926
rect 388170 -24982 388238 -24926
rect 388294 -24982 388362 -24926
rect 388418 -24982 388486 -24926
rect 388542 -24982 388610 -24926
rect 388666 -24982 388800 -24926
rect 388000 -25050 388800 -24982
rect 388000 -25106 388114 -25050
rect 388170 -25106 388238 -25050
rect 388294 -25106 388362 -25050
rect 388418 -25106 388486 -25050
rect 388542 -25106 388610 -25050
rect 388666 -25106 388800 -25050
rect 388000 -25174 388800 -25106
rect 388000 -25230 388114 -25174
rect 388170 -25230 388238 -25174
rect 388294 -25230 388362 -25174
rect 388418 -25230 388486 -25174
rect 388542 -25230 388610 -25174
rect 388666 -25230 388800 -25174
rect 388000 -25298 388800 -25230
rect 388000 -25354 388114 -25298
rect 388170 -25354 388238 -25298
rect 388294 -25354 388362 -25298
rect 388418 -25354 388486 -25298
rect 388542 -25354 388610 -25298
rect 388666 -25354 388800 -25298
rect 388000 -25422 388800 -25354
rect 388000 -25478 388114 -25422
rect 388170 -25478 388238 -25422
rect 388294 -25478 388362 -25422
rect 388418 -25478 388486 -25422
rect 388542 -25478 388610 -25422
rect 388666 -25478 388800 -25422
rect 388000 -25600 388800 -25478
rect 389068 -17950 389408 -17740
rect 389068 -18006 389141 -17950
rect 389197 -18006 389283 -17950
rect 389339 -18006 389408 -17950
rect 389068 -18092 389408 -18006
rect 389068 -18148 389141 -18092
rect 389197 -18148 389283 -18092
rect 389339 -18148 389408 -18092
rect 389068 -18234 389408 -18148
rect 389068 -18290 389141 -18234
rect 389197 -18290 389283 -18234
rect 389339 -18290 389408 -18234
rect 389068 -18376 389408 -18290
rect 389068 -18432 389141 -18376
rect 389197 -18432 389283 -18376
rect 389339 -18432 389408 -18376
rect 389068 -18518 389408 -18432
rect 389068 -18574 389141 -18518
rect 389197 -18574 389283 -18518
rect 389339 -18574 389408 -18518
rect 389068 -18660 389408 -18574
rect 389068 -18716 389141 -18660
rect 389197 -18716 389283 -18660
rect 389339 -18716 389408 -18660
rect 389068 -18802 389408 -18716
rect 389068 -18858 389141 -18802
rect 389197 -18858 389283 -18802
rect 389339 -18858 389408 -18802
rect 389068 -18944 389408 -18858
rect 389068 -19000 389141 -18944
rect 389197 -19000 389283 -18944
rect 389339 -19000 389408 -18944
rect 389068 -19086 389408 -19000
rect 389068 -19142 389141 -19086
rect 389197 -19142 389283 -19086
rect 389339 -19142 389408 -19086
rect 389068 -19228 389408 -19142
rect 389068 -19284 389141 -19228
rect 389197 -19284 389283 -19228
rect 389339 -19284 389408 -19228
rect 389068 -19370 389408 -19284
rect 389068 -19426 389141 -19370
rect 389197 -19426 389283 -19370
rect 389339 -19426 389408 -19370
rect 389068 -19512 389408 -19426
rect 389068 -19568 389141 -19512
rect 389197 -19568 389283 -19512
rect 389339 -19568 389408 -19512
rect 389068 -19654 389408 -19568
rect 389068 -19710 389141 -19654
rect 389197 -19710 389283 -19654
rect 389339 -19710 389408 -19654
rect 389068 -19796 389408 -19710
rect 389068 -19852 389141 -19796
rect 389197 -19852 389283 -19796
rect 389339 -19852 389408 -19796
rect 389068 -19938 389408 -19852
rect 389068 -19994 389141 -19938
rect 389197 -19994 389283 -19938
rect 389339 -19994 389408 -19938
rect 389068 -20080 389408 -19994
rect 389068 -20136 389141 -20080
rect 389197 -20136 389283 -20080
rect 389339 -20136 389408 -20080
rect 389068 -20222 389408 -20136
rect 389068 -20278 389141 -20222
rect 389197 -20278 389283 -20222
rect 389339 -20278 389408 -20222
rect 389068 -20364 389408 -20278
rect 389068 -20420 389141 -20364
rect 389197 -20420 389283 -20364
rect 389339 -20420 389408 -20364
rect 389068 -20506 389408 -20420
rect 389068 -20562 389141 -20506
rect 389197 -20562 389283 -20506
rect 389339 -20562 389408 -20506
rect 389068 -20648 389408 -20562
rect 389068 -20704 389141 -20648
rect 389197 -20704 389283 -20648
rect 389339 -20704 389408 -20648
rect 389068 -20790 389408 -20704
rect 389068 -20846 389141 -20790
rect 389197 -20846 389283 -20790
rect 389339 -20846 389408 -20790
rect 389068 -20932 389408 -20846
rect 389068 -20988 389141 -20932
rect 389197 -20988 389283 -20932
rect 389339 -20988 389408 -20932
rect 389068 -21074 389408 -20988
rect 389068 -21130 389141 -21074
rect 389197 -21130 389283 -21074
rect 389339 -21130 389408 -21074
rect 389068 -21216 389408 -21130
rect 389068 -21272 389141 -21216
rect 389197 -21272 389283 -21216
rect 389339 -21272 389408 -21216
rect 389068 -21358 389408 -21272
rect 389068 -21414 389141 -21358
rect 389197 -21414 389283 -21358
rect 389339 -21414 389408 -21358
rect 389068 -21500 389408 -21414
rect 389068 -21556 389141 -21500
rect 389197 -21556 389283 -21500
rect 389339 -21556 389408 -21500
rect 389068 -21642 389408 -21556
rect 389068 -21698 389141 -21642
rect 389197 -21698 389283 -21642
rect 389339 -21698 389408 -21642
rect 389068 -21784 389408 -21698
rect 389068 -21840 389141 -21784
rect 389197 -21840 389283 -21784
rect 389339 -21840 389408 -21784
rect 389068 -21926 389408 -21840
rect 389068 -21982 389141 -21926
rect 389197 -21982 389283 -21926
rect 389339 -21982 389408 -21926
rect 389068 -22068 389408 -21982
rect 389068 -22124 389141 -22068
rect 389197 -22124 389283 -22068
rect 389339 -22124 389408 -22068
rect 389068 -22210 389408 -22124
rect 389068 -22266 389141 -22210
rect 389197 -22266 389283 -22210
rect 389339 -22266 389408 -22210
rect 389068 -22352 389408 -22266
rect 389068 -22408 389141 -22352
rect 389197 -22408 389283 -22352
rect 389339 -22408 389408 -22352
rect 389068 -22494 389408 -22408
rect 389068 -22550 389141 -22494
rect 389197 -22550 389283 -22494
rect 389339 -22550 389408 -22494
rect 389068 -22636 389408 -22550
rect 389068 -22692 389141 -22636
rect 389197 -22692 389283 -22636
rect 389339 -22692 389408 -22636
rect 389068 -22778 389408 -22692
rect 389068 -22834 389141 -22778
rect 389197 -22834 389283 -22778
rect 389339 -22834 389408 -22778
rect 389068 -22920 389408 -22834
rect 389068 -22976 389141 -22920
rect 389197 -22976 389283 -22920
rect 389339 -22976 389408 -22920
rect 389068 -23062 389408 -22976
rect 389068 -23118 389141 -23062
rect 389197 -23118 389283 -23062
rect 389339 -23118 389408 -23062
rect 389068 -23204 389408 -23118
rect 389068 -23260 389141 -23204
rect 389197 -23260 389283 -23204
rect 389339 -23260 389408 -23204
rect 389068 -23346 389408 -23260
rect 389068 -23402 389141 -23346
rect 389197 -23402 389283 -23346
rect 389339 -23402 389408 -23346
rect 389068 -23488 389408 -23402
rect 389068 -23544 389141 -23488
rect 389197 -23544 389283 -23488
rect 389339 -23544 389408 -23488
rect 389068 -23630 389408 -23544
rect 389068 -23686 389141 -23630
rect 389197 -23686 389283 -23630
rect 389339 -23686 389408 -23630
rect 389068 -23772 389408 -23686
rect 389068 -23828 389141 -23772
rect 389197 -23828 389283 -23772
rect 389339 -23828 389408 -23772
rect 389068 -23914 389408 -23828
rect 389068 -23970 389141 -23914
rect 389197 -23970 389283 -23914
rect 389339 -23970 389408 -23914
rect 389068 -24056 389408 -23970
rect 389068 -24112 389141 -24056
rect 389197 -24112 389283 -24056
rect 389339 -24112 389408 -24056
rect 389068 -24198 389408 -24112
rect 389068 -24254 389141 -24198
rect 389197 -24254 389283 -24198
rect 389339 -24254 389408 -24198
rect 389068 -24340 389408 -24254
rect 389068 -24396 389141 -24340
rect 389197 -24396 389283 -24340
rect 389339 -24396 389408 -24340
rect 389068 -24482 389408 -24396
rect 389068 -24538 389141 -24482
rect 389197 -24538 389283 -24482
rect 389339 -24538 389408 -24482
rect 389068 -24624 389408 -24538
rect 389068 -24680 389141 -24624
rect 389197 -24680 389283 -24624
rect 389339 -24680 389408 -24624
rect 389068 -24766 389408 -24680
rect 389068 -24822 389141 -24766
rect 389197 -24822 389283 -24766
rect 389339 -24822 389408 -24766
rect 389068 -24908 389408 -24822
rect 389068 -24964 389141 -24908
rect 389197 -24964 389283 -24908
rect 389339 -24964 389408 -24908
rect 389068 -25050 389408 -24964
rect 389068 -25106 389141 -25050
rect 389197 -25106 389283 -25050
rect 389339 -25106 389408 -25050
rect 389068 -25192 389408 -25106
rect 389068 -25248 389141 -25192
rect 389197 -25248 389283 -25192
rect 389339 -25248 389408 -25192
rect 389068 -25334 389408 -25248
rect 389068 -25390 389141 -25334
rect 389197 -25390 389283 -25334
rect 389339 -25390 389408 -25334
rect 389068 -25476 389408 -25390
rect 389068 -25532 389141 -25476
rect 389197 -25532 389283 -25476
rect 389339 -25532 389408 -25476
rect 389068 -25600 389408 -25532
rect 389468 -17950 389808 -17740
rect 389468 -18006 389542 -17950
rect 389598 -18006 389684 -17950
rect 389740 -18006 389808 -17950
rect 389468 -18092 389808 -18006
rect 389468 -18148 389542 -18092
rect 389598 -18148 389684 -18092
rect 389740 -18148 389808 -18092
rect 389468 -18234 389808 -18148
rect 389468 -18290 389542 -18234
rect 389598 -18290 389684 -18234
rect 389740 -18290 389808 -18234
rect 389468 -18376 389808 -18290
rect 389468 -18432 389542 -18376
rect 389598 -18432 389684 -18376
rect 389740 -18432 389808 -18376
rect 389468 -18518 389808 -18432
rect 389468 -18574 389542 -18518
rect 389598 -18574 389684 -18518
rect 389740 -18574 389808 -18518
rect 389468 -18660 389808 -18574
rect 389468 -18716 389542 -18660
rect 389598 -18716 389684 -18660
rect 389740 -18716 389808 -18660
rect 389468 -18802 389808 -18716
rect 389468 -18858 389542 -18802
rect 389598 -18858 389684 -18802
rect 389740 -18858 389808 -18802
rect 389468 -18944 389808 -18858
rect 389468 -19000 389542 -18944
rect 389598 -19000 389684 -18944
rect 389740 -19000 389808 -18944
rect 389468 -19086 389808 -19000
rect 389468 -19142 389542 -19086
rect 389598 -19142 389684 -19086
rect 389740 -19142 389808 -19086
rect 389468 -19228 389808 -19142
rect 389468 -19284 389542 -19228
rect 389598 -19284 389684 -19228
rect 389740 -19284 389808 -19228
rect 389468 -19370 389808 -19284
rect 389468 -19426 389542 -19370
rect 389598 -19426 389684 -19370
rect 389740 -19426 389808 -19370
rect 389468 -19512 389808 -19426
rect 389468 -19568 389542 -19512
rect 389598 -19568 389684 -19512
rect 389740 -19568 389808 -19512
rect 389468 -19654 389808 -19568
rect 389468 -19710 389542 -19654
rect 389598 -19710 389684 -19654
rect 389740 -19710 389808 -19654
rect 389468 -19796 389808 -19710
rect 389468 -19852 389542 -19796
rect 389598 -19852 389684 -19796
rect 389740 -19852 389808 -19796
rect 389468 -19938 389808 -19852
rect 389468 -19994 389542 -19938
rect 389598 -19994 389684 -19938
rect 389740 -19994 389808 -19938
rect 389468 -20080 389808 -19994
rect 389468 -20136 389542 -20080
rect 389598 -20136 389684 -20080
rect 389740 -20136 389808 -20080
rect 389468 -20222 389808 -20136
rect 389468 -20278 389542 -20222
rect 389598 -20278 389684 -20222
rect 389740 -20278 389808 -20222
rect 389468 -20364 389808 -20278
rect 389468 -20420 389542 -20364
rect 389598 -20420 389684 -20364
rect 389740 -20420 389808 -20364
rect 389468 -20506 389808 -20420
rect 389468 -20562 389542 -20506
rect 389598 -20562 389684 -20506
rect 389740 -20562 389808 -20506
rect 389468 -20648 389808 -20562
rect 389468 -20704 389542 -20648
rect 389598 -20704 389684 -20648
rect 389740 -20704 389808 -20648
rect 389468 -20790 389808 -20704
rect 389468 -20846 389542 -20790
rect 389598 -20846 389684 -20790
rect 389740 -20846 389808 -20790
rect 389468 -20932 389808 -20846
rect 389468 -20988 389542 -20932
rect 389598 -20988 389684 -20932
rect 389740 -20988 389808 -20932
rect 389468 -21074 389808 -20988
rect 389468 -21130 389542 -21074
rect 389598 -21130 389684 -21074
rect 389740 -21130 389808 -21074
rect 389468 -21216 389808 -21130
rect 389468 -21272 389542 -21216
rect 389598 -21272 389684 -21216
rect 389740 -21272 389808 -21216
rect 389468 -21358 389808 -21272
rect 389468 -21414 389542 -21358
rect 389598 -21414 389684 -21358
rect 389740 -21414 389808 -21358
rect 389468 -21500 389808 -21414
rect 389468 -21556 389542 -21500
rect 389598 -21556 389684 -21500
rect 389740 -21556 389808 -21500
rect 389468 -21642 389808 -21556
rect 389468 -21698 389542 -21642
rect 389598 -21698 389684 -21642
rect 389740 -21698 389808 -21642
rect 389468 -21784 389808 -21698
rect 389468 -21840 389542 -21784
rect 389598 -21840 389684 -21784
rect 389740 -21840 389808 -21784
rect 389468 -21926 389808 -21840
rect 389468 -21982 389542 -21926
rect 389598 -21982 389684 -21926
rect 389740 -21982 389808 -21926
rect 389468 -22068 389808 -21982
rect 389468 -22124 389542 -22068
rect 389598 -22124 389684 -22068
rect 389740 -22124 389808 -22068
rect 389468 -22210 389808 -22124
rect 389468 -22266 389542 -22210
rect 389598 -22266 389684 -22210
rect 389740 -22266 389808 -22210
rect 389468 -22352 389808 -22266
rect 389468 -22408 389542 -22352
rect 389598 -22408 389684 -22352
rect 389740 -22408 389808 -22352
rect 389468 -22494 389808 -22408
rect 389468 -22550 389542 -22494
rect 389598 -22550 389684 -22494
rect 389740 -22550 389808 -22494
rect 389468 -22636 389808 -22550
rect 389468 -22692 389542 -22636
rect 389598 -22692 389684 -22636
rect 389740 -22692 389808 -22636
rect 389468 -22778 389808 -22692
rect 389468 -22834 389542 -22778
rect 389598 -22834 389684 -22778
rect 389740 -22834 389808 -22778
rect 389468 -22920 389808 -22834
rect 389468 -22976 389542 -22920
rect 389598 -22976 389684 -22920
rect 389740 -22976 389808 -22920
rect 389468 -23062 389808 -22976
rect 389468 -23118 389542 -23062
rect 389598 -23118 389684 -23062
rect 389740 -23118 389808 -23062
rect 389468 -23204 389808 -23118
rect 389468 -23260 389542 -23204
rect 389598 -23260 389684 -23204
rect 389740 -23260 389808 -23204
rect 389468 -23346 389808 -23260
rect 389468 -23402 389542 -23346
rect 389598 -23402 389684 -23346
rect 389740 -23402 389808 -23346
rect 389468 -23488 389808 -23402
rect 389468 -23544 389542 -23488
rect 389598 -23544 389684 -23488
rect 389740 -23544 389808 -23488
rect 389468 -23630 389808 -23544
rect 389468 -23686 389542 -23630
rect 389598 -23686 389684 -23630
rect 389740 -23686 389808 -23630
rect 389468 -23772 389808 -23686
rect 389468 -23828 389542 -23772
rect 389598 -23828 389684 -23772
rect 389740 -23828 389808 -23772
rect 389468 -23914 389808 -23828
rect 389468 -23970 389542 -23914
rect 389598 -23970 389684 -23914
rect 389740 -23970 389808 -23914
rect 389468 -24056 389808 -23970
rect 389468 -24112 389542 -24056
rect 389598 -24112 389684 -24056
rect 389740 -24112 389808 -24056
rect 389468 -24198 389808 -24112
rect 389468 -24254 389542 -24198
rect 389598 -24254 389684 -24198
rect 389740 -24254 389808 -24198
rect 389468 -24340 389808 -24254
rect 389468 -24396 389542 -24340
rect 389598 -24396 389684 -24340
rect 389740 -24396 389808 -24340
rect 389468 -24482 389808 -24396
rect 389468 -24538 389542 -24482
rect 389598 -24538 389684 -24482
rect 389740 -24538 389808 -24482
rect 389468 -24624 389808 -24538
rect 389468 -24680 389542 -24624
rect 389598 -24680 389684 -24624
rect 389740 -24680 389808 -24624
rect 389468 -24766 389808 -24680
rect 389468 -24822 389542 -24766
rect 389598 -24822 389684 -24766
rect 389740 -24822 389808 -24766
rect 389468 -24908 389808 -24822
rect 389468 -24964 389542 -24908
rect 389598 -24964 389684 -24908
rect 389740 -24964 389808 -24908
rect 389468 -25050 389808 -24964
rect 389468 -25106 389542 -25050
rect 389598 -25106 389684 -25050
rect 389740 -25106 389808 -25050
rect 389468 -25192 389808 -25106
rect 389468 -25248 389542 -25192
rect 389598 -25248 389684 -25192
rect 389740 -25248 389808 -25192
rect 389468 -25334 389808 -25248
rect 389468 -25390 389542 -25334
rect 389598 -25390 389684 -25334
rect 389740 -25390 389808 -25334
rect 389468 -25476 389808 -25390
rect 389468 -25532 389542 -25476
rect 389598 -25532 389684 -25476
rect 389740 -25532 389808 -25476
rect 389468 -25600 389808 -25532
rect 389868 -17950 390208 -17740
rect 389868 -18006 389942 -17950
rect 389998 -18006 390084 -17950
rect 390140 -18006 390208 -17950
rect 389868 -18092 390208 -18006
rect 389868 -18148 389942 -18092
rect 389998 -18148 390084 -18092
rect 390140 -18148 390208 -18092
rect 389868 -18234 390208 -18148
rect 389868 -18290 389942 -18234
rect 389998 -18290 390084 -18234
rect 390140 -18290 390208 -18234
rect 389868 -18376 390208 -18290
rect 389868 -18432 389942 -18376
rect 389998 -18432 390084 -18376
rect 390140 -18432 390208 -18376
rect 389868 -18518 390208 -18432
rect 389868 -18574 389942 -18518
rect 389998 -18574 390084 -18518
rect 390140 -18574 390208 -18518
rect 389868 -18660 390208 -18574
rect 389868 -18716 389942 -18660
rect 389998 -18716 390084 -18660
rect 390140 -18716 390208 -18660
rect 389868 -18802 390208 -18716
rect 389868 -18858 389942 -18802
rect 389998 -18858 390084 -18802
rect 390140 -18858 390208 -18802
rect 389868 -18944 390208 -18858
rect 389868 -19000 389942 -18944
rect 389998 -19000 390084 -18944
rect 390140 -19000 390208 -18944
rect 389868 -19086 390208 -19000
rect 389868 -19142 389942 -19086
rect 389998 -19142 390084 -19086
rect 390140 -19142 390208 -19086
rect 389868 -19228 390208 -19142
rect 389868 -19284 389942 -19228
rect 389998 -19284 390084 -19228
rect 390140 -19284 390208 -19228
rect 389868 -19370 390208 -19284
rect 389868 -19426 389942 -19370
rect 389998 -19426 390084 -19370
rect 390140 -19426 390208 -19370
rect 389868 -19512 390208 -19426
rect 389868 -19568 389942 -19512
rect 389998 -19568 390084 -19512
rect 390140 -19568 390208 -19512
rect 389868 -19654 390208 -19568
rect 389868 -19710 389942 -19654
rect 389998 -19710 390084 -19654
rect 390140 -19710 390208 -19654
rect 389868 -19796 390208 -19710
rect 389868 -19852 389942 -19796
rect 389998 -19852 390084 -19796
rect 390140 -19852 390208 -19796
rect 389868 -19938 390208 -19852
rect 389868 -19994 389942 -19938
rect 389998 -19994 390084 -19938
rect 390140 -19994 390208 -19938
rect 389868 -20080 390208 -19994
rect 389868 -20136 389942 -20080
rect 389998 -20136 390084 -20080
rect 390140 -20136 390208 -20080
rect 389868 -20222 390208 -20136
rect 389868 -20278 389942 -20222
rect 389998 -20278 390084 -20222
rect 390140 -20278 390208 -20222
rect 389868 -20364 390208 -20278
rect 389868 -20420 389942 -20364
rect 389998 -20420 390084 -20364
rect 390140 -20420 390208 -20364
rect 389868 -20506 390208 -20420
rect 389868 -20562 389942 -20506
rect 389998 -20562 390084 -20506
rect 390140 -20562 390208 -20506
rect 389868 -20648 390208 -20562
rect 389868 -20704 389942 -20648
rect 389998 -20704 390084 -20648
rect 390140 -20704 390208 -20648
rect 389868 -20790 390208 -20704
rect 389868 -20846 389942 -20790
rect 389998 -20846 390084 -20790
rect 390140 -20846 390208 -20790
rect 389868 -20932 390208 -20846
rect 389868 -20988 389942 -20932
rect 389998 -20988 390084 -20932
rect 390140 -20988 390208 -20932
rect 389868 -21074 390208 -20988
rect 389868 -21130 389942 -21074
rect 389998 -21130 390084 -21074
rect 390140 -21130 390208 -21074
rect 389868 -21216 390208 -21130
rect 389868 -21272 389942 -21216
rect 389998 -21272 390084 -21216
rect 390140 -21272 390208 -21216
rect 389868 -21358 390208 -21272
rect 389868 -21414 389942 -21358
rect 389998 -21414 390084 -21358
rect 390140 -21414 390208 -21358
rect 389868 -21500 390208 -21414
rect 389868 -21556 389942 -21500
rect 389998 -21556 390084 -21500
rect 390140 -21556 390208 -21500
rect 389868 -21642 390208 -21556
rect 389868 -21698 389942 -21642
rect 389998 -21698 390084 -21642
rect 390140 -21698 390208 -21642
rect 389868 -21784 390208 -21698
rect 389868 -21840 389942 -21784
rect 389998 -21840 390084 -21784
rect 390140 -21840 390208 -21784
rect 389868 -21926 390208 -21840
rect 389868 -21982 389942 -21926
rect 389998 -21982 390084 -21926
rect 390140 -21982 390208 -21926
rect 389868 -22068 390208 -21982
rect 389868 -22124 389942 -22068
rect 389998 -22124 390084 -22068
rect 390140 -22124 390208 -22068
rect 389868 -22210 390208 -22124
rect 389868 -22266 389942 -22210
rect 389998 -22266 390084 -22210
rect 390140 -22266 390208 -22210
rect 389868 -22352 390208 -22266
rect 389868 -22408 389942 -22352
rect 389998 -22408 390084 -22352
rect 390140 -22408 390208 -22352
rect 389868 -22494 390208 -22408
rect 389868 -22550 389942 -22494
rect 389998 -22550 390084 -22494
rect 390140 -22550 390208 -22494
rect 389868 -22636 390208 -22550
rect 389868 -22692 389942 -22636
rect 389998 -22692 390084 -22636
rect 390140 -22692 390208 -22636
rect 389868 -22778 390208 -22692
rect 389868 -22834 389942 -22778
rect 389998 -22834 390084 -22778
rect 390140 -22834 390208 -22778
rect 389868 -22920 390208 -22834
rect 389868 -22976 389942 -22920
rect 389998 -22976 390084 -22920
rect 390140 -22976 390208 -22920
rect 389868 -23062 390208 -22976
rect 389868 -23118 389942 -23062
rect 389998 -23118 390084 -23062
rect 390140 -23118 390208 -23062
rect 389868 -23204 390208 -23118
rect 389868 -23260 389942 -23204
rect 389998 -23260 390084 -23204
rect 390140 -23260 390208 -23204
rect 389868 -23346 390208 -23260
rect 389868 -23402 389942 -23346
rect 389998 -23402 390084 -23346
rect 390140 -23402 390208 -23346
rect 389868 -23488 390208 -23402
rect 389868 -23544 389942 -23488
rect 389998 -23544 390084 -23488
rect 390140 -23544 390208 -23488
rect 389868 -23630 390208 -23544
rect 389868 -23686 389942 -23630
rect 389998 -23686 390084 -23630
rect 390140 -23686 390208 -23630
rect 389868 -23772 390208 -23686
rect 389868 -23828 389942 -23772
rect 389998 -23828 390084 -23772
rect 390140 -23828 390208 -23772
rect 389868 -23914 390208 -23828
rect 389868 -23970 389942 -23914
rect 389998 -23970 390084 -23914
rect 390140 -23970 390208 -23914
rect 389868 -24056 390208 -23970
rect 389868 -24112 389942 -24056
rect 389998 -24112 390084 -24056
rect 390140 -24112 390208 -24056
rect 389868 -24198 390208 -24112
rect 389868 -24254 389942 -24198
rect 389998 -24254 390084 -24198
rect 390140 -24254 390208 -24198
rect 389868 -24340 390208 -24254
rect 389868 -24396 389942 -24340
rect 389998 -24396 390084 -24340
rect 390140 -24396 390208 -24340
rect 389868 -24482 390208 -24396
rect 389868 -24538 389942 -24482
rect 389998 -24538 390084 -24482
rect 390140 -24538 390208 -24482
rect 389868 -24624 390208 -24538
rect 389868 -24680 389942 -24624
rect 389998 -24680 390084 -24624
rect 390140 -24680 390208 -24624
rect 389868 -24766 390208 -24680
rect 389868 -24822 389942 -24766
rect 389998 -24822 390084 -24766
rect 390140 -24822 390208 -24766
rect 389868 -24908 390208 -24822
rect 389868 -24964 389942 -24908
rect 389998 -24964 390084 -24908
rect 390140 -24964 390208 -24908
rect 389868 -25050 390208 -24964
rect 389868 -25106 389942 -25050
rect 389998 -25106 390084 -25050
rect 390140 -25106 390208 -25050
rect 389868 -25192 390208 -25106
rect 389868 -25248 389942 -25192
rect 389998 -25248 390084 -25192
rect 390140 -25248 390208 -25192
rect 389868 -25334 390208 -25248
rect 389868 -25390 389942 -25334
rect 389998 -25390 390084 -25334
rect 390140 -25390 390208 -25334
rect 389868 -25476 390208 -25390
rect 389868 -25532 389942 -25476
rect 389998 -25532 390084 -25476
rect 390140 -25532 390208 -25476
rect 389868 -25600 390208 -25532
rect 390268 -17950 390608 -17740
rect 390268 -18006 390339 -17950
rect 390395 -18006 390481 -17950
rect 390537 -18006 390608 -17950
rect 390268 -18092 390608 -18006
rect 390268 -18148 390339 -18092
rect 390395 -18148 390481 -18092
rect 390537 -18148 390608 -18092
rect 390268 -18234 390608 -18148
rect 390268 -18290 390339 -18234
rect 390395 -18290 390481 -18234
rect 390537 -18290 390608 -18234
rect 390268 -18376 390608 -18290
rect 390268 -18432 390339 -18376
rect 390395 -18432 390481 -18376
rect 390537 -18432 390608 -18376
rect 390268 -18518 390608 -18432
rect 390268 -18574 390339 -18518
rect 390395 -18574 390481 -18518
rect 390537 -18574 390608 -18518
rect 390268 -18660 390608 -18574
rect 390268 -18716 390339 -18660
rect 390395 -18716 390481 -18660
rect 390537 -18716 390608 -18660
rect 390268 -18802 390608 -18716
rect 390268 -18858 390339 -18802
rect 390395 -18858 390481 -18802
rect 390537 -18858 390608 -18802
rect 390268 -18944 390608 -18858
rect 390268 -19000 390339 -18944
rect 390395 -19000 390481 -18944
rect 390537 -19000 390608 -18944
rect 390268 -19086 390608 -19000
rect 390268 -19142 390339 -19086
rect 390395 -19142 390481 -19086
rect 390537 -19142 390608 -19086
rect 390268 -19228 390608 -19142
rect 390268 -19284 390339 -19228
rect 390395 -19284 390481 -19228
rect 390537 -19284 390608 -19228
rect 390268 -19370 390608 -19284
rect 390268 -19426 390339 -19370
rect 390395 -19426 390481 -19370
rect 390537 -19426 390608 -19370
rect 390268 -19512 390608 -19426
rect 390268 -19568 390339 -19512
rect 390395 -19568 390481 -19512
rect 390537 -19568 390608 -19512
rect 390268 -19654 390608 -19568
rect 390268 -19710 390339 -19654
rect 390395 -19710 390481 -19654
rect 390537 -19710 390608 -19654
rect 390268 -19796 390608 -19710
rect 390268 -19852 390339 -19796
rect 390395 -19852 390481 -19796
rect 390537 -19852 390608 -19796
rect 390268 -19938 390608 -19852
rect 390268 -19994 390339 -19938
rect 390395 -19994 390481 -19938
rect 390537 -19994 390608 -19938
rect 390268 -20080 390608 -19994
rect 390268 -20136 390339 -20080
rect 390395 -20136 390481 -20080
rect 390537 -20136 390608 -20080
rect 390268 -20222 390608 -20136
rect 390268 -20278 390339 -20222
rect 390395 -20278 390481 -20222
rect 390537 -20278 390608 -20222
rect 390268 -20364 390608 -20278
rect 390268 -20420 390339 -20364
rect 390395 -20420 390481 -20364
rect 390537 -20420 390608 -20364
rect 390268 -20506 390608 -20420
rect 390268 -20562 390339 -20506
rect 390395 -20562 390481 -20506
rect 390537 -20562 390608 -20506
rect 390268 -20648 390608 -20562
rect 390268 -20704 390339 -20648
rect 390395 -20704 390481 -20648
rect 390537 -20704 390608 -20648
rect 390268 -20790 390608 -20704
rect 390268 -20846 390339 -20790
rect 390395 -20846 390481 -20790
rect 390537 -20846 390608 -20790
rect 390268 -20932 390608 -20846
rect 390268 -20988 390339 -20932
rect 390395 -20988 390481 -20932
rect 390537 -20988 390608 -20932
rect 390268 -21074 390608 -20988
rect 390268 -21130 390339 -21074
rect 390395 -21130 390481 -21074
rect 390537 -21130 390608 -21074
rect 390268 -21216 390608 -21130
rect 390268 -21272 390339 -21216
rect 390395 -21272 390481 -21216
rect 390537 -21272 390608 -21216
rect 390268 -21358 390608 -21272
rect 390268 -21414 390339 -21358
rect 390395 -21414 390481 -21358
rect 390537 -21414 390608 -21358
rect 390268 -21500 390608 -21414
rect 390268 -21556 390339 -21500
rect 390395 -21556 390481 -21500
rect 390537 -21556 390608 -21500
rect 390268 -21642 390608 -21556
rect 390268 -21698 390339 -21642
rect 390395 -21698 390481 -21642
rect 390537 -21698 390608 -21642
rect 390268 -21784 390608 -21698
rect 390268 -21840 390339 -21784
rect 390395 -21840 390481 -21784
rect 390537 -21840 390608 -21784
rect 390268 -21926 390608 -21840
rect 390268 -21982 390339 -21926
rect 390395 -21982 390481 -21926
rect 390537 -21982 390608 -21926
rect 390268 -22068 390608 -21982
rect 390268 -22124 390339 -22068
rect 390395 -22124 390481 -22068
rect 390537 -22124 390608 -22068
rect 390268 -22210 390608 -22124
rect 390268 -22266 390339 -22210
rect 390395 -22266 390481 -22210
rect 390537 -22266 390608 -22210
rect 390268 -22352 390608 -22266
rect 390268 -22408 390339 -22352
rect 390395 -22408 390481 -22352
rect 390537 -22408 390608 -22352
rect 390268 -22494 390608 -22408
rect 390268 -22550 390339 -22494
rect 390395 -22550 390481 -22494
rect 390537 -22550 390608 -22494
rect 390268 -22636 390608 -22550
rect 390268 -22692 390339 -22636
rect 390395 -22692 390481 -22636
rect 390537 -22692 390608 -22636
rect 390268 -22778 390608 -22692
rect 390268 -22834 390339 -22778
rect 390395 -22834 390481 -22778
rect 390537 -22834 390608 -22778
rect 390268 -22920 390608 -22834
rect 390268 -22976 390339 -22920
rect 390395 -22976 390481 -22920
rect 390537 -22976 390608 -22920
rect 390268 -23062 390608 -22976
rect 390268 -23118 390339 -23062
rect 390395 -23118 390481 -23062
rect 390537 -23118 390608 -23062
rect 390268 -23204 390608 -23118
rect 390268 -23260 390339 -23204
rect 390395 -23260 390481 -23204
rect 390537 -23260 390608 -23204
rect 390268 -23346 390608 -23260
rect 390268 -23402 390339 -23346
rect 390395 -23402 390481 -23346
rect 390537 -23402 390608 -23346
rect 390268 -23488 390608 -23402
rect 390268 -23544 390339 -23488
rect 390395 -23544 390481 -23488
rect 390537 -23544 390608 -23488
rect 390268 -23630 390608 -23544
rect 390268 -23686 390339 -23630
rect 390395 -23686 390481 -23630
rect 390537 -23686 390608 -23630
rect 390268 -23772 390608 -23686
rect 390268 -23828 390339 -23772
rect 390395 -23828 390481 -23772
rect 390537 -23828 390608 -23772
rect 390268 -23914 390608 -23828
rect 390268 -23970 390339 -23914
rect 390395 -23970 390481 -23914
rect 390537 -23970 390608 -23914
rect 390268 -24056 390608 -23970
rect 390268 -24112 390339 -24056
rect 390395 -24112 390481 -24056
rect 390537 -24112 390608 -24056
rect 390268 -24198 390608 -24112
rect 390268 -24254 390339 -24198
rect 390395 -24254 390481 -24198
rect 390537 -24254 390608 -24198
rect 390268 -24340 390608 -24254
rect 390268 -24396 390339 -24340
rect 390395 -24396 390481 -24340
rect 390537 -24396 390608 -24340
rect 390268 -24482 390608 -24396
rect 390268 -24538 390339 -24482
rect 390395 -24538 390481 -24482
rect 390537 -24538 390608 -24482
rect 390268 -24624 390608 -24538
rect 390268 -24680 390339 -24624
rect 390395 -24680 390481 -24624
rect 390537 -24680 390608 -24624
rect 390268 -24766 390608 -24680
rect 390268 -24822 390339 -24766
rect 390395 -24822 390481 -24766
rect 390537 -24822 390608 -24766
rect 390268 -24908 390608 -24822
rect 390268 -24964 390339 -24908
rect 390395 -24964 390481 -24908
rect 390537 -24964 390608 -24908
rect 390268 -25050 390608 -24964
rect 390268 -25106 390339 -25050
rect 390395 -25106 390481 -25050
rect 390537 -25106 390608 -25050
rect 390268 -25192 390608 -25106
rect 390268 -25248 390339 -25192
rect 390395 -25248 390481 -25192
rect 390537 -25248 390608 -25192
rect 390268 -25334 390608 -25248
rect 390268 -25390 390339 -25334
rect 390395 -25390 390481 -25334
rect 390537 -25390 390608 -25334
rect 390268 -25476 390608 -25390
rect 390268 -25532 390339 -25476
rect 390395 -25532 390481 -25476
rect 390537 -25532 390608 -25476
rect 390268 -25600 390608 -25532
rect 390668 -17950 391008 -17740
rect 390668 -18006 390736 -17950
rect 390792 -18006 390878 -17950
rect 390934 -18006 391008 -17950
rect 390668 -18092 391008 -18006
rect 390668 -18148 390736 -18092
rect 390792 -18148 390878 -18092
rect 390934 -18148 391008 -18092
rect 390668 -18234 391008 -18148
rect 390668 -18290 390736 -18234
rect 390792 -18290 390878 -18234
rect 390934 -18290 391008 -18234
rect 390668 -18376 391008 -18290
rect 390668 -18432 390736 -18376
rect 390792 -18432 390878 -18376
rect 390934 -18432 391008 -18376
rect 390668 -18518 391008 -18432
rect 390668 -18574 390736 -18518
rect 390792 -18574 390878 -18518
rect 390934 -18574 391008 -18518
rect 390668 -18660 391008 -18574
rect 390668 -18716 390736 -18660
rect 390792 -18716 390878 -18660
rect 390934 -18716 391008 -18660
rect 390668 -18802 391008 -18716
rect 390668 -18858 390736 -18802
rect 390792 -18858 390878 -18802
rect 390934 -18858 391008 -18802
rect 390668 -18944 391008 -18858
rect 390668 -19000 390736 -18944
rect 390792 -19000 390878 -18944
rect 390934 -19000 391008 -18944
rect 390668 -19086 391008 -19000
rect 390668 -19142 390736 -19086
rect 390792 -19142 390878 -19086
rect 390934 -19142 391008 -19086
rect 390668 -19228 391008 -19142
rect 390668 -19284 390736 -19228
rect 390792 -19284 390878 -19228
rect 390934 -19284 391008 -19228
rect 390668 -19370 391008 -19284
rect 390668 -19426 390736 -19370
rect 390792 -19426 390878 -19370
rect 390934 -19426 391008 -19370
rect 390668 -19512 391008 -19426
rect 390668 -19568 390736 -19512
rect 390792 -19568 390878 -19512
rect 390934 -19568 391008 -19512
rect 390668 -19654 391008 -19568
rect 390668 -19710 390736 -19654
rect 390792 -19710 390878 -19654
rect 390934 -19710 391008 -19654
rect 390668 -19796 391008 -19710
rect 390668 -19852 390736 -19796
rect 390792 -19852 390878 -19796
rect 390934 -19852 391008 -19796
rect 390668 -19938 391008 -19852
rect 390668 -19994 390736 -19938
rect 390792 -19994 390878 -19938
rect 390934 -19994 391008 -19938
rect 390668 -20080 391008 -19994
rect 390668 -20136 390736 -20080
rect 390792 -20136 390878 -20080
rect 390934 -20136 391008 -20080
rect 390668 -20222 391008 -20136
rect 390668 -20278 390736 -20222
rect 390792 -20278 390878 -20222
rect 390934 -20278 391008 -20222
rect 390668 -20364 391008 -20278
rect 390668 -20420 390736 -20364
rect 390792 -20420 390878 -20364
rect 390934 -20420 391008 -20364
rect 390668 -20506 391008 -20420
rect 390668 -20562 390736 -20506
rect 390792 -20562 390878 -20506
rect 390934 -20562 391008 -20506
rect 390668 -20648 391008 -20562
rect 390668 -20704 390736 -20648
rect 390792 -20704 390878 -20648
rect 390934 -20704 391008 -20648
rect 390668 -20790 391008 -20704
rect 390668 -20846 390736 -20790
rect 390792 -20846 390878 -20790
rect 390934 -20846 391008 -20790
rect 390668 -20932 391008 -20846
rect 390668 -20988 390736 -20932
rect 390792 -20988 390878 -20932
rect 390934 -20988 391008 -20932
rect 390668 -21074 391008 -20988
rect 390668 -21130 390736 -21074
rect 390792 -21130 390878 -21074
rect 390934 -21130 391008 -21074
rect 390668 -21216 391008 -21130
rect 390668 -21272 390736 -21216
rect 390792 -21272 390878 -21216
rect 390934 -21272 391008 -21216
rect 390668 -21358 391008 -21272
rect 390668 -21414 390736 -21358
rect 390792 -21414 390878 -21358
rect 390934 -21414 391008 -21358
rect 390668 -21500 391008 -21414
rect 390668 -21556 390736 -21500
rect 390792 -21556 390878 -21500
rect 390934 -21556 391008 -21500
rect 390668 -21642 391008 -21556
rect 390668 -21698 390736 -21642
rect 390792 -21698 390878 -21642
rect 390934 -21698 391008 -21642
rect 390668 -21784 391008 -21698
rect 390668 -21840 390736 -21784
rect 390792 -21840 390878 -21784
rect 390934 -21840 391008 -21784
rect 390668 -21926 391008 -21840
rect 390668 -21982 390736 -21926
rect 390792 -21982 390878 -21926
rect 390934 -21982 391008 -21926
rect 390668 -22068 391008 -21982
rect 390668 -22124 390736 -22068
rect 390792 -22124 390878 -22068
rect 390934 -22124 391008 -22068
rect 390668 -22210 391008 -22124
rect 390668 -22266 390736 -22210
rect 390792 -22266 390878 -22210
rect 390934 -22266 391008 -22210
rect 390668 -22352 391008 -22266
rect 390668 -22408 390736 -22352
rect 390792 -22408 390878 -22352
rect 390934 -22408 391008 -22352
rect 390668 -22494 391008 -22408
rect 390668 -22550 390736 -22494
rect 390792 -22550 390878 -22494
rect 390934 -22550 391008 -22494
rect 390668 -22636 391008 -22550
rect 390668 -22692 390736 -22636
rect 390792 -22692 390878 -22636
rect 390934 -22692 391008 -22636
rect 390668 -22778 391008 -22692
rect 390668 -22834 390736 -22778
rect 390792 -22834 390878 -22778
rect 390934 -22834 391008 -22778
rect 390668 -22920 391008 -22834
rect 390668 -22976 390736 -22920
rect 390792 -22976 390878 -22920
rect 390934 -22976 391008 -22920
rect 390668 -23062 391008 -22976
rect 390668 -23118 390736 -23062
rect 390792 -23118 390878 -23062
rect 390934 -23118 391008 -23062
rect 390668 -23204 391008 -23118
rect 390668 -23260 390736 -23204
rect 390792 -23260 390878 -23204
rect 390934 -23260 391008 -23204
rect 390668 -23346 391008 -23260
rect 390668 -23402 390736 -23346
rect 390792 -23402 390878 -23346
rect 390934 -23402 391008 -23346
rect 390668 -23488 391008 -23402
rect 390668 -23544 390736 -23488
rect 390792 -23544 390878 -23488
rect 390934 -23544 391008 -23488
rect 390668 -23630 391008 -23544
rect 390668 -23686 390736 -23630
rect 390792 -23686 390878 -23630
rect 390934 -23686 391008 -23630
rect 390668 -23772 391008 -23686
rect 390668 -23828 390736 -23772
rect 390792 -23828 390878 -23772
rect 390934 -23828 391008 -23772
rect 390668 -23914 391008 -23828
rect 390668 -23970 390736 -23914
rect 390792 -23970 390878 -23914
rect 390934 -23970 391008 -23914
rect 390668 -24056 391008 -23970
rect 390668 -24112 390736 -24056
rect 390792 -24112 390878 -24056
rect 390934 -24112 391008 -24056
rect 390668 -24198 391008 -24112
rect 390668 -24254 390736 -24198
rect 390792 -24254 390878 -24198
rect 390934 -24254 391008 -24198
rect 390668 -24340 391008 -24254
rect 390668 -24396 390736 -24340
rect 390792 -24396 390878 -24340
rect 390934 -24396 391008 -24340
rect 390668 -24482 391008 -24396
rect 390668 -24538 390736 -24482
rect 390792 -24538 390878 -24482
rect 390934 -24538 391008 -24482
rect 390668 -24624 391008 -24538
rect 390668 -24680 390736 -24624
rect 390792 -24680 390878 -24624
rect 390934 -24680 391008 -24624
rect 390668 -24766 391008 -24680
rect 390668 -24822 390736 -24766
rect 390792 -24822 390878 -24766
rect 390934 -24822 391008 -24766
rect 390668 -24908 391008 -24822
rect 390668 -24964 390736 -24908
rect 390792 -24964 390878 -24908
rect 390934 -24964 391008 -24908
rect 390668 -25050 391008 -24964
rect 390668 -25106 390736 -25050
rect 390792 -25106 390878 -25050
rect 390934 -25106 391008 -25050
rect 390668 -25192 391008 -25106
rect 390668 -25248 390736 -25192
rect 390792 -25248 390878 -25192
rect 390934 -25248 391008 -25192
rect 390668 -25334 391008 -25248
rect 390668 -25390 390736 -25334
rect 390792 -25390 390878 -25334
rect 390934 -25390 391008 -25334
rect 390668 -25476 391008 -25390
rect 390668 -25532 390736 -25476
rect 390792 -25532 390878 -25476
rect 390934 -25532 391008 -25476
rect 390668 -25600 391008 -25532
rect 391068 -17950 391408 -17740
rect 391068 -18006 391140 -17950
rect 391196 -18006 391282 -17950
rect 391338 -18006 391408 -17950
rect 391068 -18092 391408 -18006
rect 391068 -18148 391140 -18092
rect 391196 -18148 391282 -18092
rect 391338 -18148 391408 -18092
rect 391068 -18234 391408 -18148
rect 391068 -18290 391140 -18234
rect 391196 -18290 391282 -18234
rect 391338 -18290 391408 -18234
rect 391068 -18376 391408 -18290
rect 391068 -18432 391140 -18376
rect 391196 -18432 391282 -18376
rect 391338 -18432 391408 -18376
rect 391068 -18518 391408 -18432
rect 391068 -18574 391140 -18518
rect 391196 -18574 391282 -18518
rect 391338 -18574 391408 -18518
rect 391068 -18660 391408 -18574
rect 391068 -18716 391140 -18660
rect 391196 -18716 391282 -18660
rect 391338 -18716 391408 -18660
rect 391068 -18802 391408 -18716
rect 391068 -18858 391140 -18802
rect 391196 -18858 391282 -18802
rect 391338 -18858 391408 -18802
rect 391068 -18944 391408 -18858
rect 391068 -19000 391140 -18944
rect 391196 -19000 391282 -18944
rect 391338 -19000 391408 -18944
rect 391068 -19086 391408 -19000
rect 391068 -19142 391140 -19086
rect 391196 -19142 391282 -19086
rect 391338 -19142 391408 -19086
rect 391068 -19228 391408 -19142
rect 391068 -19284 391140 -19228
rect 391196 -19284 391282 -19228
rect 391338 -19284 391408 -19228
rect 391068 -19370 391408 -19284
rect 391068 -19426 391140 -19370
rect 391196 -19426 391282 -19370
rect 391338 -19426 391408 -19370
rect 391068 -19512 391408 -19426
rect 391068 -19568 391140 -19512
rect 391196 -19568 391282 -19512
rect 391338 -19568 391408 -19512
rect 391068 -19654 391408 -19568
rect 391068 -19710 391140 -19654
rect 391196 -19710 391282 -19654
rect 391338 -19710 391408 -19654
rect 391068 -19796 391408 -19710
rect 391068 -19852 391140 -19796
rect 391196 -19852 391282 -19796
rect 391338 -19852 391408 -19796
rect 391068 -19938 391408 -19852
rect 391068 -19994 391140 -19938
rect 391196 -19994 391282 -19938
rect 391338 -19994 391408 -19938
rect 391068 -20080 391408 -19994
rect 391068 -20136 391140 -20080
rect 391196 -20136 391282 -20080
rect 391338 -20136 391408 -20080
rect 391068 -20222 391408 -20136
rect 391068 -20278 391140 -20222
rect 391196 -20278 391282 -20222
rect 391338 -20278 391408 -20222
rect 391068 -20364 391408 -20278
rect 391068 -20420 391140 -20364
rect 391196 -20420 391282 -20364
rect 391338 -20420 391408 -20364
rect 391068 -20506 391408 -20420
rect 391068 -20562 391140 -20506
rect 391196 -20562 391282 -20506
rect 391338 -20562 391408 -20506
rect 391068 -20648 391408 -20562
rect 391068 -20704 391140 -20648
rect 391196 -20704 391282 -20648
rect 391338 -20704 391408 -20648
rect 391068 -20790 391408 -20704
rect 391068 -20846 391140 -20790
rect 391196 -20846 391282 -20790
rect 391338 -20846 391408 -20790
rect 391068 -20932 391408 -20846
rect 391068 -20988 391140 -20932
rect 391196 -20988 391282 -20932
rect 391338 -20988 391408 -20932
rect 391068 -21074 391408 -20988
rect 391068 -21130 391140 -21074
rect 391196 -21130 391282 -21074
rect 391338 -21130 391408 -21074
rect 391068 -21216 391408 -21130
rect 391068 -21272 391140 -21216
rect 391196 -21272 391282 -21216
rect 391338 -21272 391408 -21216
rect 391068 -21358 391408 -21272
rect 391068 -21414 391140 -21358
rect 391196 -21414 391282 -21358
rect 391338 -21414 391408 -21358
rect 391068 -21500 391408 -21414
rect 391068 -21556 391140 -21500
rect 391196 -21556 391282 -21500
rect 391338 -21556 391408 -21500
rect 391068 -21642 391408 -21556
rect 391068 -21698 391140 -21642
rect 391196 -21698 391282 -21642
rect 391338 -21698 391408 -21642
rect 391068 -21784 391408 -21698
rect 391068 -21840 391140 -21784
rect 391196 -21840 391282 -21784
rect 391338 -21840 391408 -21784
rect 391068 -21926 391408 -21840
rect 391068 -21982 391140 -21926
rect 391196 -21982 391282 -21926
rect 391338 -21982 391408 -21926
rect 391068 -22068 391408 -21982
rect 391068 -22124 391140 -22068
rect 391196 -22124 391282 -22068
rect 391338 -22124 391408 -22068
rect 391068 -22210 391408 -22124
rect 391068 -22266 391140 -22210
rect 391196 -22266 391282 -22210
rect 391338 -22266 391408 -22210
rect 391068 -22352 391408 -22266
rect 391068 -22408 391140 -22352
rect 391196 -22408 391282 -22352
rect 391338 -22408 391408 -22352
rect 391068 -22494 391408 -22408
rect 391068 -22550 391140 -22494
rect 391196 -22550 391282 -22494
rect 391338 -22550 391408 -22494
rect 391068 -22636 391408 -22550
rect 391068 -22692 391140 -22636
rect 391196 -22692 391282 -22636
rect 391338 -22692 391408 -22636
rect 391068 -22778 391408 -22692
rect 391068 -22834 391140 -22778
rect 391196 -22834 391282 -22778
rect 391338 -22834 391408 -22778
rect 391068 -22920 391408 -22834
rect 391068 -22976 391140 -22920
rect 391196 -22976 391282 -22920
rect 391338 -22976 391408 -22920
rect 391068 -23062 391408 -22976
rect 391068 -23118 391140 -23062
rect 391196 -23118 391282 -23062
rect 391338 -23118 391408 -23062
rect 391068 -23204 391408 -23118
rect 391068 -23260 391140 -23204
rect 391196 -23260 391282 -23204
rect 391338 -23260 391408 -23204
rect 391068 -23346 391408 -23260
rect 391068 -23402 391140 -23346
rect 391196 -23402 391282 -23346
rect 391338 -23402 391408 -23346
rect 391068 -23488 391408 -23402
rect 391068 -23544 391140 -23488
rect 391196 -23544 391282 -23488
rect 391338 -23544 391408 -23488
rect 391068 -23630 391408 -23544
rect 391068 -23686 391140 -23630
rect 391196 -23686 391282 -23630
rect 391338 -23686 391408 -23630
rect 391068 -23772 391408 -23686
rect 391068 -23828 391140 -23772
rect 391196 -23828 391282 -23772
rect 391338 -23828 391408 -23772
rect 391068 -23914 391408 -23828
rect 391068 -23970 391140 -23914
rect 391196 -23970 391282 -23914
rect 391338 -23970 391408 -23914
rect 391068 -24056 391408 -23970
rect 391068 -24112 391140 -24056
rect 391196 -24112 391282 -24056
rect 391338 -24112 391408 -24056
rect 391068 -24198 391408 -24112
rect 391068 -24254 391140 -24198
rect 391196 -24254 391282 -24198
rect 391338 -24254 391408 -24198
rect 391068 -24340 391408 -24254
rect 391068 -24396 391140 -24340
rect 391196 -24396 391282 -24340
rect 391338 -24396 391408 -24340
rect 391068 -24482 391408 -24396
rect 391068 -24538 391140 -24482
rect 391196 -24538 391282 -24482
rect 391338 -24538 391408 -24482
rect 391068 -24624 391408 -24538
rect 391068 -24680 391140 -24624
rect 391196 -24680 391282 -24624
rect 391338 -24680 391408 -24624
rect 391068 -24766 391408 -24680
rect 391068 -24822 391140 -24766
rect 391196 -24822 391282 -24766
rect 391338 -24822 391408 -24766
rect 391068 -24908 391408 -24822
rect 391068 -24964 391140 -24908
rect 391196 -24964 391282 -24908
rect 391338 -24964 391408 -24908
rect 391068 -25050 391408 -24964
rect 391068 -25106 391140 -25050
rect 391196 -25106 391282 -25050
rect 391338 -25106 391408 -25050
rect 391068 -25192 391408 -25106
rect 391068 -25248 391140 -25192
rect 391196 -25248 391282 -25192
rect 391338 -25248 391408 -25192
rect 391068 -25334 391408 -25248
rect 391068 -25390 391140 -25334
rect 391196 -25390 391282 -25334
rect 391338 -25390 391408 -25334
rect 391068 -25476 391408 -25390
rect 391068 -25532 391140 -25476
rect 391196 -25532 391282 -25476
rect 391338 -25532 391408 -25476
rect 391068 -25600 391408 -25532
rect 391468 -17950 391808 -17740
rect 391468 -18006 391536 -17950
rect 391592 -18006 391678 -17950
rect 391734 -18006 391808 -17950
rect 391468 -18092 391808 -18006
rect 391468 -18148 391536 -18092
rect 391592 -18148 391678 -18092
rect 391734 -18148 391808 -18092
rect 391468 -18234 391808 -18148
rect 391468 -18290 391536 -18234
rect 391592 -18290 391678 -18234
rect 391734 -18290 391808 -18234
rect 391468 -18376 391808 -18290
rect 391468 -18432 391536 -18376
rect 391592 -18432 391678 -18376
rect 391734 -18432 391808 -18376
rect 391468 -18518 391808 -18432
rect 391468 -18574 391536 -18518
rect 391592 -18574 391678 -18518
rect 391734 -18574 391808 -18518
rect 391468 -18660 391808 -18574
rect 391468 -18716 391536 -18660
rect 391592 -18716 391678 -18660
rect 391734 -18716 391808 -18660
rect 391468 -18802 391808 -18716
rect 391468 -18858 391536 -18802
rect 391592 -18858 391678 -18802
rect 391734 -18858 391808 -18802
rect 391468 -18944 391808 -18858
rect 391468 -19000 391536 -18944
rect 391592 -19000 391678 -18944
rect 391734 -19000 391808 -18944
rect 391468 -19086 391808 -19000
rect 391468 -19142 391536 -19086
rect 391592 -19142 391678 -19086
rect 391734 -19142 391808 -19086
rect 391468 -19228 391808 -19142
rect 391468 -19284 391536 -19228
rect 391592 -19284 391678 -19228
rect 391734 -19284 391808 -19228
rect 391468 -19370 391808 -19284
rect 391468 -19426 391536 -19370
rect 391592 -19426 391678 -19370
rect 391734 -19426 391808 -19370
rect 391468 -19512 391808 -19426
rect 391468 -19568 391536 -19512
rect 391592 -19568 391678 -19512
rect 391734 -19568 391808 -19512
rect 391468 -19654 391808 -19568
rect 391468 -19710 391536 -19654
rect 391592 -19710 391678 -19654
rect 391734 -19710 391808 -19654
rect 391468 -19796 391808 -19710
rect 391468 -19852 391536 -19796
rect 391592 -19852 391678 -19796
rect 391734 -19852 391808 -19796
rect 391468 -19938 391808 -19852
rect 391468 -19994 391536 -19938
rect 391592 -19994 391678 -19938
rect 391734 -19994 391808 -19938
rect 391468 -20080 391808 -19994
rect 391468 -20136 391536 -20080
rect 391592 -20136 391678 -20080
rect 391734 -20136 391808 -20080
rect 391468 -20222 391808 -20136
rect 391468 -20278 391536 -20222
rect 391592 -20278 391678 -20222
rect 391734 -20278 391808 -20222
rect 391468 -20364 391808 -20278
rect 391468 -20420 391536 -20364
rect 391592 -20420 391678 -20364
rect 391734 -20420 391808 -20364
rect 391468 -20506 391808 -20420
rect 391468 -20562 391536 -20506
rect 391592 -20562 391678 -20506
rect 391734 -20562 391808 -20506
rect 391468 -20648 391808 -20562
rect 391468 -20704 391536 -20648
rect 391592 -20704 391678 -20648
rect 391734 -20704 391808 -20648
rect 391468 -20790 391808 -20704
rect 391468 -20846 391536 -20790
rect 391592 -20846 391678 -20790
rect 391734 -20846 391808 -20790
rect 391468 -20932 391808 -20846
rect 391468 -20988 391536 -20932
rect 391592 -20988 391678 -20932
rect 391734 -20988 391808 -20932
rect 391468 -21074 391808 -20988
rect 391468 -21130 391536 -21074
rect 391592 -21130 391678 -21074
rect 391734 -21130 391808 -21074
rect 391468 -21216 391808 -21130
rect 391468 -21272 391536 -21216
rect 391592 -21272 391678 -21216
rect 391734 -21272 391808 -21216
rect 391468 -21358 391808 -21272
rect 391468 -21414 391536 -21358
rect 391592 -21414 391678 -21358
rect 391734 -21414 391808 -21358
rect 391468 -21500 391808 -21414
rect 391468 -21556 391536 -21500
rect 391592 -21556 391678 -21500
rect 391734 -21556 391808 -21500
rect 391468 -21642 391808 -21556
rect 391468 -21698 391536 -21642
rect 391592 -21698 391678 -21642
rect 391734 -21698 391808 -21642
rect 391468 -21784 391808 -21698
rect 391468 -21840 391536 -21784
rect 391592 -21840 391678 -21784
rect 391734 -21840 391808 -21784
rect 391468 -21926 391808 -21840
rect 391468 -21982 391536 -21926
rect 391592 -21982 391678 -21926
rect 391734 -21982 391808 -21926
rect 391468 -22068 391808 -21982
rect 391468 -22124 391536 -22068
rect 391592 -22124 391678 -22068
rect 391734 -22124 391808 -22068
rect 391468 -22210 391808 -22124
rect 391468 -22266 391536 -22210
rect 391592 -22266 391678 -22210
rect 391734 -22266 391808 -22210
rect 391468 -22352 391808 -22266
rect 391468 -22408 391536 -22352
rect 391592 -22408 391678 -22352
rect 391734 -22408 391808 -22352
rect 391468 -22494 391808 -22408
rect 391468 -22550 391536 -22494
rect 391592 -22550 391678 -22494
rect 391734 -22550 391808 -22494
rect 391468 -22636 391808 -22550
rect 391468 -22692 391536 -22636
rect 391592 -22692 391678 -22636
rect 391734 -22692 391808 -22636
rect 391468 -22778 391808 -22692
rect 391468 -22834 391536 -22778
rect 391592 -22834 391678 -22778
rect 391734 -22834 391808 -22778
rect 391468 -22920 391808 -22834
rect 391468 -22976 391536 -22920
rect 391592 -22976 391678 -22920
rect 391734 -22976 391808 -22920
rect 391468 -23062 391808 -22976
rect 391468 -23118 391536 -23062
rect 391592 -23118 391678 -23062
rect 391734 -23118 391808 -23062
rect 391468 -23204 391808 -23118
rect 391468 -23260 391536 -23204
rect 391592 -23260 391678 -23204
rect 391734 -23260 391808 -23204
rect 391468 -23346 391808 -23260
rect 391468 -23402 391536 -23346
rect 391592 -23402 391678 -23346
rect 391734 -23402 391808 -23346
rect 391468 -23488 391808 -23402
rect 391468 -23544 391536 -23488
rect 391592 -23544 391678 -23488
rect 391734 -23544 391808 -23488
rect 391468 -23630 391808 -23544
rect 391468 -23686 391536 -23630
rect 391592 -23686 391678 -23630
rect 391734 -23686 391808 -23630
rect 391468 -23772 391808 -23686
rect 391468 -23828 391536 -23772
rect 391592 -23828 391678 -23772
rect 391734 -23828 391808 -23772
rect 391468 -23914 391808 -23828
rect 391468 -23970 391536 -23914
rect 391592 -23970 391678 -23914
rect 391734 -23970 391808 -23914
rect 391468 -24056 391808 -23970
rect 391468 -24112 391536 -24056
rect 391592 -24112 391678 -24056
rect 391734 -24112 391808 -24056
rect 391468 -24198 391808 -24112
rect 391468 -24254 391536 -24198
rect 391592 -24254 391678 -24198
rect 391734 -24254 391808 -24198
rect 391468 -24340 391808 -24254
rect 391468 -24396 391536 -24340
rect 391592 -24396 391678 -24340
rect 391734 -24396 391808 -24340
rect 391468 -24482 391808 -24396
rect 391468 -24538 391536 -24482
rect 391592 -24538 391678 -24482
rect 391734 -24538 391808 -24482
rect 391468 -24624 391808 -24538
rect 391468 -24680 391536 -24624
rect 391592 -24680 391678 -24624
rect 391734 -24680 391808 -24624
rect 391468 -24766 391808 -24680
rect 391468 -24822 391536 -24766
rect 391592 -24822 391678 -24766
rect 391734 -24822 391808 -24766
rect 391468 -24908 391808 -24822
rect 391468 -24964 391536 -24908
rect 391592 -24964 391678 -24908
rect 391734 -24964 391808 -24908
rect 391468 -25050 391808 -24964
rect 391468 -25106 391536 -25050
rect 391592 -25106 391678 -25050
rect 391734 -25106 391808 -25050
rect 391468 -25192 391808 -25106
rect 391468 -25248 391536 -25192
rect 391592 -25248 391678 -25192
rect 391734 -25248 391808 -25192
rect 391468 -25334 391808 -25248
rect 391468 -25390 391536 -25334
rect 391592 -25390 391678 -25334
rect 391734 -25390 391808 -25334
rect 391468 -25476 391808 -25390
rect 391468 -25532 391536 -25476
rect 391592 -25532 391678 -25476
rect 391734 -25532 391808 -25476
rect 391468 -25600 391808 -25532
rect 391868 -17950 392208 -17740
rect 391868 -18006 391936 -17950
rect 391992 -18006 392078 -17950
rect 392134 -18006 392208 -17950
rect 391868 -18092 392208 -18006
rect 391868 -18148 391936 -18092
rect 391992 -18148 392078 -18092
rect 392134 -18148 392208 -18092
rect 391868 -18234 392208 -18148
rect 391868 -18290 391936 -18234
rect 391992 -18290 392078 -18234
rect 392134 -18290 392208 -18234
rect 391868 -18376 392208 -18290
rect 391868 -18432 391936 -18376
rect 391992 -18432 392078 -18376
rect 392134 -18432 392208 -18376
rect 391868 -18518 392208 -18432
rect 391868 -18574 391936 -18518
rect 391992 -18574 392078 -18518
rect 392134 -18574 392208 -18518
rect 391868 -18660 392208 -18574
rect 391868 -18716 391936 -18660
rect 391992 -18716 392078 -18660
rect 392134 -18716 392208 -18660
rect 391868 -18802 392208 -18716
rect 391868 -18858 391936 -18802
rect 391992 -18858 392078 -18802
rect 392134 -18858 392208 -18802
rect 391868 -18944 392208 -18858
rect 391868 -19000 391936 -18944
rect 391992 -19000 392078 -18944
rect 392134 -19000 392208 -18944
rect 391868 -19086 392208 -19000
rect 391868 -19142 391936 -19086
rect 391992 -19142 392078 -19086
rect 392134 -19142 392208 -19086
rect 391868 -19228 392208 -19142
rect 391868 -19284 391936 -19228
rect 391992 -19284 392078 -19228
rect 392134 -19284 392208 -19228
rect 391868 -19370 392208 -19284
rect 391868 -19426 391936 -19370
rect 391992 -19426 392078 -19370
rect 392134 -19426 392208 -19370
rect 391868 -19512 392208 -19426
rect 391868 -19568 391936 -19512
rect 391992 -19568 392078 -19512
rect 392134 -19568 392208 -19512
rect 391868 -19654 392208 -19568
rect 391868 -19710 391936 -19654
rect 391992 -19710 392078 -19654
rect 392134 -19710 392208 -19654
rect 391868 -19796 392208 -19710
rect 391868 -19852 391936 -19796
rect 391992 -19852 392078 -19796
rect 392134 -19852 392208 -19796
rect 391868 -19938 392208 -19852
rect 391868 -19994 391936 -19938
rect 391992 -19994 392078 -19938
rect 392134 -19994 392208 -19938
rect 391868 -20080 392208 -19994
rect 391868 -20136 391936 -20080
rect 391992 -20136 392078 -20080
rect 392134 -20136 392208 -20080
rect 391868 -20222 392208 -20136
rect 391868 -20278 391936 -20222
rect 391992 -20278 392078 -20222
rect 392134 -20278 392208 -20222
rect 391868 -20364 392208 -20278
rect 391868 -20420 391936 -20364
rect 391992 -20420 392078 -20364
rect 392134 -20420 392208 -20364
rect 391868 -20506 392208 -20420
rect 391868 -20562 391936 -20506
rect 391992 -20562 392078 -20506
rect 392134 -20562 392208 -20506
rect 391868 -20648 392208 -20562
rect 391868 -20704 391936 -20648
rect 391992 -20704 392078 -20648
rect 392134 -20704 392208 -20648
rect 391868 -20790 392208 -20704
rect 391868 -20846 391936 -20790
rect 391992 -20846 392078 -20790
rect 392134 -20846 392208 -20790
rect 391868 -20932 392208 -20846
rect 391868 -20988 391936 -20932
rect 391992 -20988 392078 -20932
rect 392134 -20988 392208 -20932
rect 391868 -21074 392208 -20988
rect 391868 -21130 391936 -21074
rect 391992 -21130 392078 -21074
rect 392134 -21130 392208 -21074
rect 391868 -21216 392208 -21130
rect 391868 -21272 391936 -21216
rect 391992 -21272 392078 -21216
rect 392134 -21272 392208 -21216
rect 391868 -21358 392208 -21272
rect 391868 -21414 391936 -21358
rect 391992 -21414 392078 -21358
rect 392134 -21414 392208 -21358
rect 391868 -21500 392208 -21414
rect 391868 -21556 391936 -21500
rect 391992 -21556 392078 -21500
rect 392134 -21556 392208 -21500
rect 391868 -21642 392208 -21556
rect 391868 -21698 391936 -21642
rect 391992 -21698 392078 -21642
rect 392134 -21698 392208 -21642
rect 391868 -21784 392208 -21698
rect 391868 -21840 391936 -21784
rect 391992 -21840 392078 -21784
rect 392134 -21840 392208 -21784
rect 391868 -21926 392208 -21840
rect 391868 -21982 391936 -21926
rect 391992 -21982 392078 -21926
rect 392134 -21982 392208 -21926
rect 391868 -22068 392208 -21982
rect 391868 -22124 391936 -22068
rect 391992 -22124 392078 -22068
rect 392134 -22124 392208 -22068
rect 391868 -22210 392208 -22124
rect 391868 -22266 391936 -22210
rect 391992 -22266 392078 -22210
rect 392134 -22266 392208 -22210
rect 391868 -22352 392208 -22266
rect 391868 -22408 391936 -22352
rect 391992 -22408 392078 -22352
rect 392134 -22408 392208 -22352
rect 391868 -22494 392208 -22408
rect 391868 -22550 391936 -22494
rect 391992 -22550 392078 -22494
rect 392134 -22550 392208 -22494
rect 391868 -22636 392208 -22550
rect 391868 -22692 391936 -22636
rect 391992 -22692 392078 -22636
rect 392134 -22692 392208 -22636
rect 391868 -22778 392208 -22692
rect 391868 -22834 391936 -22778
rect 391992 -22834 392078 -22778
rect 392134 -22834 392208 -22778
rect 391868 -22920 392208 -22834
rect 391868 -22976 391936 -22920
rect 391992 -22976 392078 -22920
rect 392134 -22976 392208 -22920
rect 391868 -23062 392208 -22976
rect 391868 -23118 391936 -23062
rect 391992 -23118 392078 -23062
rect 392134 -23118 392208 -23062
rect 391868 -23204 392208 -23118
rect 391868 -23260 391936 -23204
rect 391992 -23260 392078 -23204
rect 392134 -23260 392208 -23204
rect 391868 -23346 392208 -23260
rect 391868 -23402 391936 -23346
rect 391992 -23402 392078 -23346
rect 392134 -23402 392208 -23346
rect 391868 -23488 392208 -23402
rect 391868 -23544 391936 -23488
rect 391992 -23544 392078 -23488
rect 392134 -23544 392208 -23488
rect 391868 -23630 392208 -23544
rect 391868 -23686 391936 -23630
rect 391992 -23686 392078 -23630
rect 392134 -23686 392208 -23630
rect 391868 -23772 392208 -23686
rect 391868 -23828 391936 -23772
rect 391992 -23828 392078 -23772
rect 392134 -23828 392208 -23772
rect 391868 -23914 392208 -23828
rect 391868 -23970 391936 -23914
rect 391992 -23970 392078 -23914
rect 392134 -23970 392208 -23914
rect 391868 -24056 392208 -23970
rect 391868 -24112 391936 -24056
rect 391992 -24112 392078 -24056
rect 392134 -24112 392208 -24056
rect 391868 -24198 392208 -24112
rect 391868 -24254 391936 -24198
rect 391992 -24254 392078 -24198
rect 392134 -24254 392208 -24198
rect 391868 -24340 392208 -24254
rect 391868 -24396 391936 -24340
rect 391992 -24396 392078 -24340
rect 392134 -24396 392208 -24340
rect 391868 -24482 392208 -24396
rect 391868 -24538 391936 -24482
rect 391992 -24538 392078 -24482
rect 392134 -24538 392208 -24482
rect 391868 -24624 392208 -24538
rect 391868 -24680 391936 -24624
rect 391992 -24680 392078 -24624
rect 392134 -24680 392208 -24624
rect 391868 -24766 392208 -24680
rect 391868 -24822 391936 -24766
rect 391992 -24822 392078 -24766
rect 392134 -24822 392208 -24766
rect 391868 -24908 392208 -24822
rect 391868 -24964 391936 -24908
rect 391992 -24964 392078 -24908
rect 392134 -24964 392208 -24908
rect 391868 -25050 392208 -24964
rect 391868 -25106 391936 -25050
rect 391992 -25106 392078 -25050
rect 392134 -25106 392208 -25050
rect 391868 -25192 392208 -25106
rect 391868 -25248 391936 -25192
rect 391992 -25248 392078 -25192
rect 392134 -25248 392208 -25192
rect 391868 -25334 392208 -25248
rect 391868 -25390 391936 -25334
rect 391992 -25390 392078 -25334
rect 392134 -25390 392208 -25334
rect 391868 -25476 392208 -25390
rect 391868 -25532 391936 -25476
rect 391992 -25532 392078 -25476
rect 392134 -25532 392208 -25476
rect 391868 -25600 392208 -25532
rect 392268 -17950 392608 -17740
rect 392268 -18006 392333 -17950
rect 392389 -18006 392475 -17950
rect 392531 -18006 392608 -17950
rect 392268 -18092 392608 -18006
rect 392268 -18148 392333 -18092
rect 392389 -18148 392475 -18092
rect 392531 -18148 392608 -18092
rect 392268 -18234 392608 -18148
rect 392268 -18290 392333 -18234
rect 392389 -18290 392475 -18234
rect 392531 -18290 392608 -18234
rect 392268 -18376 392608 -18290
rect 392268 -18432 392333 -18376
rect 392389 -18432 392475 -18376
rect 392531 -18432 392608 -18376
rect 392268 -18518 392608 -18432
rect 392268 -18574 392333 -18518
rect 392389 -18574 392475 -18518
rect 392531 -18574 392608 -18518
rect 392268 -18660 392608 -18574
rect 392268 -18716 392333 -18660
rect 392389 -18716 392475 -18660
rect 392531 -18716 392608 -18660
rect 392268 -18802 392608 -18716
rect 392268 -18858 392333 -18802
rect 392389 -18858 392475 -18802
rect 392531 -18858 392608 -18802
rect 392268 -18944 392608 -18858
rect 392268 -19000 392333 -18944
rect 392389 -19000 392475 -18944
rect 392531 -19000 392608 -18944
rect 392268 -19086 392608 -19000
rect 392268 -19142 392333 -19086
rect 392389 -19142 392475 -19086
rect 392531 -19142 392608 -19086
rect 392268 -19228 392608 -19142
rect 392268 -19284 392333 -19228
rect 392389 -19284 392475 -19228
rect 392531 -19284 392608 -19228
rect 392268 -19370 392608 -19284
rect 392268 -19426 392333 -19370
rect 392389 -19426 392475 -19370
rect 392531 -19426 392608 -19370
rect 392268 -19512 392608 -19426
rect 392268 -19568 392333 -19512
rect 392389 -19568 392475 -19512
rect 392531 -19568 392608 -19512
rect 392268 -19654 392608 -19568
rect 392268 -19710 392333 -19654
rect 392389 -19710 392475 -19654
rect 392531 -19710 392608 -19654
rect 392268 -19796 392608 -19710
rect 392268 -19852 392333 -19796
rect 392389 -19852 392475 -19796
rect 392531 -19852 392608 -19796
rect 392268 -19938 392608 -19852
rect 392268 -19994 392333 -19938
rect 392389 -19994 392475 -19938
rect 392531 -19994 392608 -19938
rect 392268 -20080 392608 -19994
rect 392268 -20136 392333 -20080
rect 392389 -20136 392475 -20080
rect 392531 -20136 392608 -20080
rect 392268 -20222 392608 -20136
rect 392268 -20278 392333 -20222
rect 392389 -20278 392475 -20222
rect 392531 -20278 392608 -20222
rect 392268 -20364 392608 -20278
rect 392268 -20420 392333 -20364
rect 392389 -20420 392475 -20364
rect 392531 -20420 392608 -20364
rect 392268 -20506 392608 -20420
rect 392268 -20562 392333 -20506
rect 392389 -20562 392475 -20506
rect 392531 -20562 392608 -20506
rect 392268 -20648 392608 -20562
rect 392268 -20704 392333 -20648
rect 392389 -20704 392475 -20648
rect 392531 -20704 392608 -20648
rect 392268 -20790 392608 -20704
rect 392268 -20846 392333 -20790
rect 392389 -20846 392475 -20790
rect 392531 -20846 392608 -20790
rect 392268 -20932 392608 -20846
rect 392268 -20988 392333 -20932
rect 392389 -20988 392475 -20932
rect 392531 -20988 392608 -20932
rect 392268 -21074 392608 -20988
rect 392268 -21130 392333 -21074
rect 392389 -21130 392475 -21074
rect 392531 -21130 392608 -21074
rect 392268 -21216 392608 -21130
rect 392268 -21272 392333 -21216
rect 392389 -21272 392475 -21216
rect 392531 -21272 392608 -21216
rect 392268 -21358 392608 -21272
rect 392268 -21414 392333 -21358
rect 392389 -21414 392475 -21358
rect 392531 -21414 392608 -21358
rect 392268 -21500 392608 -21414
rect 392268 -21556 392333 -21500
rect 392389 -21556 392475 -21500
rect 392531 -21556 392608 -21500
rect 392268 -21642 392608 -21556
rect 392268 -21698 392333 -21642
rect 392389 -21698 392475 -21642
rect 392531 -21698 392608 -21642
rect 392268 -21784 392608 -21698
rect 392268 -21840 392333 -21784
rect 392389 -21840 392475 -21784
rect 392531 -21840 392608 -21784
rect 392268 -21926 392608 -21840
rect 392268 -21982 392333 -21926
rect 392389 -21982 392475 -21926
rect 392531 -21982 392608 -21926
rect 392268 -22068 392608 -21982
rect 392268 -22124 392333 -22068
rect 392389 -22124 392475 -22068
rect 392531 -22124 392608 -22068
rect 392268 -22210 392608 -22124
rect 392268 -22266 392333 -22210
rect 392389 -22266 392475 -22210
rect 392531 -22266 392608 -22210
rect 392268 -22352 392608 -22266
rect 392268 -22408 392333 -22352
rect 392389 -22408 392475 -22352
rect 392531 -22408 392608 -22352
rect 392268 -22494 392608 -22408
rect 392268 -22550 392333 -22494
rect 392389 -22550 392475 -22494
rect 392531 -22550 392608 -22494
rect 392268 -22636 392608 -22550
rect 392268 -22692 392333 -22636
rect 392389 -22692 392475 -22636
rect 392531 -22692 392608 -22636
rect 392268 -22778 392608 -22692
rect 392268 -22834 392333 -22778
rect 392389 -22834 392475 -22778
rect 392531 -22834 392608 -22778
rect 392268 -22920 392608 -22834
rect 392268 -22976 392333 -22920
rect 392389 -22976 392475 -22920
rect 392531 -22976 392608 -22920
rect 392268 -23062 392608 -22976
rect 392268 -23118 392333 -23062
rect 392389 -23118 392475 -23062
rect 392531 -23118 392608 -23062
rect 392268 -23204 392608 -23118
rect 392268 -23260 392333 -23204
rect 392389 -23260 392475 -23204
rect 392531 -23260 392608 -23204
rect 392268 -23346 392608 -23260
rect 392268 -23402 392333 -23346
rect 392389 -23402 392475 -23346
rect 392531 -23402 392608 -23346
rect 392268 -23488 392608 -23402
rect 392268 -23544 392333 -23488
rect 392389 -23544 392475 -23488
rect 392531 -23544 392608 -23488
rect 392268 -23630 392608 -23544
rect 392268 -23686 392333 -23630
rect 392389 -23686 392475 -23630
rect 392531 -23686 392608 -23630
rect 392268 -23772 392608 -23686
rect 392268 -23828 392333 -23772
rect 392389 -23828 392475 -23772
rect 392531 -23828 392608 -23772
rect 392268 -23914 392608 -23828
rect 392268 -23970 392333 -23914
rect 392389 -23970 392475 -23914
rect 392531 -23970 392608 -23914
rect 392268 -24056 392608 -23970
rect 392268 -24112 392333 -24056
rect 392389 -24112 392475 -24056
rect 392531 -24112 392608 -24056
rect 392268 -24198 392608 -24112
rect 392268 -24254 392333 -24198
rect 392389 -24254 392475 -24198
rect 392531 -24254 392608 -24198
rect 392268 -24340 392608 -24254
rect 392268 -24396 392333 -24340
rect 392389 -24396 392475 -24340
rect 392531 -24396 392608 -24340
rect 392268 -24482 392608 -24396
rect 392268 -24538 392333 -24482
rect 392389 -24538 392475 -24482
rect 392531 -24538 392608 -24482
rect 392268 -24624 392608 -24538
rect 392268 -24680 392333 -24624
rect 392389 -24680 392475 -24624
rect 392531 -24680 392608 -24624
rect 392268 -24766 392608 -24680
rect 392268 -24822 392333 -24766
rect 392389 -24822 392475 -24766
rect 392531 -24822 392608 -24766
rect 392268 -24908 392608 -24822
rect 392268 -24964 392333 -24908
rect 392389 -24964 392475 -24908
rect 392531 -24964 392608 -24908
rect 392268 -25050 392608 -24964
rect 392268 -25106 392333 -25050
rect 392389 -25106 392475 -25050
rect 392531 -25106 392608 -25050
rect 392268 -25192 392608 -25106
rect 392268 -25248 392333 -25192
rect 392389 -25248 392475 -25192
rect 392531 -25248 392608 -25192
rect 392268 -25334 392608 -25248
rect 392268 -25390 392333 -25334
rect 392389 -25390 392475 -25334
rect 392531 -25390 392608 -25334
rect 392268 -25476 392608 -25390
rect 392268 -25532 392333 -25476
rect 392389 -25532 392475 -25476
rect 392531 -25532 392608 -25476
rect 392268 -25600 392608 -25532
rect 392668 -17950 393008 -17740
rect 392668 -18006 392738 -17950
rect 392794 -18006 392880 -17950
rect 392936 -18006 393008 -17950
rect 392668 -18092 393008 -18006
rect 392668 -18148 392738 -18092
rect 392794 -18148 392880 -18092
rect 392936 -18148 393008 -18092
rect 392668 -18234 393008 -18148
rect 392668 -18290 392738 -18234
rect 392794 -18290 392880 -18234
rect 392936 -18290 393008 -18234
rect 392668 -18376 393008 -18290
rect 392668 -18432 392738 -18376
rect 392794 -18432 392880 -18376
rect 392936 -18432 393008 -18376
rect 392668 -18518 393008 -18432
rect 392668 -18574 392738 -18518
rect 392794 -18574 392880 -18518
rect 392936 -18574 393008 -18518
rect 392668 -18660 393008 -18574
rect 392668 -18716 392738 -18660
rect 392794 -18716 392880 -18660
rect 392936 -18716 393008 -18660
rect 392668 -18802 393008 -18716
rect 392668 -18858 392738 -18802
rect 392794 -18858 392880 -18802
rect 392936 -18858 393008 -18802
rect 392668 -18944 393008 -18858
rect 392668 -19000 392738 -18944
rect 392794 -19000 392880 -18944
rect 392936 -19000 393008 -18944
rect 392668 -19086 393008 -19000
rect 392668 -19142 392738 -19086
rect 392794 -19142 392880 -19086
rect 392936 -19142 393008 -19086
rect 392668 -19228 393008 -19142
rect 392668 -19284 392738 -19228
rect 392794 -19284 392880 -19228
rect 392936 -19284 393008 -19228
rect 392668 -19370 393008 -19284
rect 392668 -19426 392738 -19370
rect 392794 -19426 392880 -19370
rect 392936 -19426 393008 -19370
rect 392668 -19512 393008 -19426
rect 392668 -19568 392738 -19512
rect 392794 -19568 392880 -19512
rect 392936 -19568 393008 -19512
rect 392668 -19654 393008 -19568
rect 392668 -19710 392738 -19654
rect 392794 -19710 392880 -19654
rect 392936 -19710 393008 -19654
rect 392668 -19796 393008 -19710
rect 392668 -19852 392738 -19796
rect 392794 -19852 392880 -19796
rect 392936 -19852 393008 -19796
rect 392668 -19938 393008 -19852
rect 392668 -19994 392738 -19938
rect 392794 -19994 392880 -19938
rect 392936 -19994 393008 -19938
rect 392668 -20080 393008 -19994
rect 392668 -20136 392738 -20080
rect 392794 -20136 392880 -20080
rect 392936 -20136 393008 -20080
rect 392668 -20222 393008 -20136
rect 392668 -20278 392738 -20222
rect 392794 -20278 392880 -20222
rect 392936 -20278 393008 -20222
rect 392668 -20364 393008 -20278
rect 392668 -20420 392738 -20364
rect 392794 -20420 392880 -20364
rect 392936 -20420 393008 -20364
rect 392668 -20506 393008 -20420
rect 392668 -20562 392738 -20506
rect 392794 -20562 392880 -20506
rect 392936 -20562 393008 -20506
rect 392668 -20648 393008 -20562
rect 392668 -20704 392738 -20648
rect 392794 -20704 392880 -20648
rect 392936 -20704 393008 -20648
rect 392668 -20790 393008 -20704
rect 392668 -20846 392738 -20790
rect 392794 -20846 392880 -20790
rect 392936 -20846 393008 -20790
rect 392668 -20932 393008 -20846
rect 392668 -20988 392738 -20932
rect 392794 -20988 392880 -20932
rect 392936 -20988 393008 -20932
rect 392668 -21074 393008 -20988
rect 392668 -21130 392738 -21074
rect 392794 -21130 392880 -21074
rect 392936 -21130 393008 -21074
rect 392668 -21216 393008 -21130
rect 392668 -21272 392738 -21216
rect 392794 -21272 392880 -21216
rect 392936 -21272 393008 -21216
rect 392668 -21358 393008 -21272
rect 392668 -21414 392738 -21358
rect 392794 -21414 392880 -21358
rect 392936 -21414 393008 -21358
rect 392668 -21500 393008 -21414
rect 392668 -21556 392738 -21500
rect 392794 -21556 392880 -21500
rect 392936 -21556 393008 -21500
rect 392668 -21642 393008 -21556
rect 392668 -21698 392738 -21642
rect 392794 -21698 392880 -21642
rect 392936 -21698 393008 -21642
rect 392668 -21784 393008 -21698
rect 392668 -21840 392738 -21784
rect 392794 -21840 392880 -21784
rect 392936 -21840 393008 -21784
rect 392668 -21926 393008 -21840
rect 392668 -21982 392738 -21926
rect 392794 -21982 392880 -21926
rect 392936 -21982 393008 -21926
rect 392668 -22068 393008 -21982
rect 392668 -22124 392738 -22068
rect 392794 -22124 392880 -22068
rect 392936 -22124 393008 -22068
rect 392668 -22210 393008 -22124
rect 392668 -22266 392738 -22210
rect 392794 -22266 392880 -22210
rect 392936 -22266 393008 -22210
rect 392668 -22352 393008 -22266
rect 392668 -22408 392738 -22352
rect 392794 -22408 392880 -22352
rect 392936 -22408 393008 -22352
rect 392668 -22494 393008 -22408
rect 392668 -22550 392738 -22494
rect 392794 -22550 392880 -22494
rect 392936 -22550 393008 -22494
rect 392668 -22636 393008 -22550
rect 392668 -22692 392738 -22636
rect 392794 -22692 392880 -22636
rect 392936 -22692 393008 -22636
rect 392668 -22778 393008 -22692
rect 392668 -22834 392738 -22778
rect 392794 -22834 392880 -22778
rect 392936 -22834 393008 -22778
rect 392668 -22920 393008 -22834
rect 392668 -22976 392738 -22920
rect 392794 -22976 392880 -22920
rect 392936 -22976 393008 -22920
rect 392668 -23062 393008 -22976
rect 392668 -23118 392738 -23062
rect 392794 -23118 392880 -23062
rect 392936 -23118 393008 -23062
rect 392668 -23204 393008 -23118
rect 392668 -23260 392738 -23204
rect 392794 -23260 392880 -23204
rect 392936 -23260 393008 -23204
rect 392668 -23346 393008 -23260
rect 392668 -23402 392738 -23346
rect 392794 -23402 392880 -23346
rect 392936 -23402 393008 -23346
rect 392668 -23488 393008 -23402
rect 392668 -23544 392738 -23488
rect 392794 -23544 392880 -23488
rect 392936 -23544 393008 -23488
rect 392668 -23630 393008 -23544
rect 392668 -23686 392738 -23630
rect 392794 -23686 392880 -23630
rect 392936 -23686 393008 -23630
rect 392668 -23772 393008 -23686
rect 392668 -23828 392738 -23772
rect 392794 -23828 392880 -23772
rect 392936 -23828 393008 -23772
rect 392668 -23914 393008 -23828
rect 392668 -23970 392738 -23914
rect 392794 -23970 392880 -23914
rect 392936 -23970 393008 -23914
rect 392668 -24056 393008 -23970
rect 392668 -24112 392738 -24056
rect 392794 -24112 392880 -24056
rect 392936 -24112 393008 -24056
rect 392668 -24198 393008 -24112
rect 392668 -24254 392738 -24198
rect 392794 -24254 392880 -24198
rect 392936 -24254 393008 -24198
rect 392668 -24340 393008 -24254
rect 392668 -24396 392738 -24340
rect 392794 -24396 392880 -24340
rect 392936 -24396 393008 -24340
rect 392668 -24482 393008 -24396
rect 392668 -24538 392738 -24482
rect 392794 -24538 392880 -24482
rect 392936 -24538 393008 -24482
rect 392668 -24624 393008 -24538
rect 392668 -24680 392738 -24624
rect 392794 -24680 392880 -24624
rect 392936 -24680 393008 -24624
rect 392668 -24766 393008 -24680
rect 392668 -24822 392738 -24766
rect 392794 -24822 392880 -24766
rect 392936 -24822 393008 -24766
rect 392668 -24908 393008 -24822
rect 392668 -24964 392738 -24908
rect 392794 -24964 392880 -24908
rect 392936 -24964 393008 -24908
rect 392668 -25050 393008 -24964
rect 392668 -25106 392738 -25050
rect 392794 -25106 392880 -25050
rect 392936 -25106 393008 -25050
rect 392668 -25192 393008 -25106
rect 392668 -25248 392738 -25192
rect 392794 -25248 392880 -25192
rect 392936 -25248 393008 -25192
rect 392668 -25334 393008 -25248
rect 392668 -25390 392738 -25334
rect 392794 -25390 392880 -25334
rect 392936 -25390 393008 -25334
rect 392668 -25476 393008 -25390
rect 392668 -25532 392738 -25476
rect 392794 -25532 392880 -25476
rect 392936 -25532 393008 -25476
rect 392668 -25600 393008 -25532
rect 393068 -17950 393408 -17740
rect 393068 -18006 393138 -17950
rect 393194 -18006 393280 -17950
rect 393336 -18006 393408 -17950
rect 393068 -18092 393408 -18006
rect 393068 -18148 393138 -18092
rect 393194 -18148 393280 -18092
rect 393336 -18148 393408 -18092
rect 393068 -18234 393408 -18148
rect 393068 -18290 393138 -18234
rect 393194 -18290 393280 -18234
rect 393336 -18290 393408 -18234
rect 393068 -18376 393408 -18290
rect 393068 -18432 393138 -18376
rect 393194 -18432 393280 -18376
rect 393336 -18432 393408 -18376
rect 393068 -18518 393408 -18432
rect 393068 -18574 393138 -18518
rect 393194 -18574 393280 -18518
rect 393336 -18574 393408 -18518
rect 393068 -18660 393408 -18574
rect 393068 -18716 393138 -18660
rect 393194 -18716 393280 -18660
rect 393336 -18716 393408 -18660
rect 393068 -18802 393408 -18716
rect 393068 -18858 393138 -18802
rect 393194 -18858 393280 -18802
rect 393336 -18858 393408 -18802
rect 393068 -18944 393408 -18858
rect 393068 -19000 393138 -18944
rect 393194 -19000 393280 -18944
rect 393336 -19000 393408 -18944
rect 393068 -19086 393408 -19000
rect 393068 -19142 393138 -19086
rect 393194 -19142 393280 -19086
rect 393336 -19142 393408 -19086
rect 393068 -19228 393408 -19142
rect 393068 -19284 393138 -19228
rect 393194 -19284 393280 -19228
rect 393336 -19284 393408 -19228
rect 393068 -19370 393408 -19284
rect 393068 -19426 393138 -19370
rect 393194 -19426 393280 -19370
rect 393336 -19426 393408 -19370
rect 393068 -19512 393408 -19426
rect 393068 -19568 393138 -19512
rect 393194 -19568 393280 -19512
rect 393336 -19568 393408 -19512
rect 393068 -19654 393408 -19568
rect 393068 -19710 393138 -19654
rect 393194 -19710 393280 -19654
rect 393336 -19710 393408 -19654
rect 393068 -19796 393408 -19710
rect 393068 -19852 393138 -19796
rect 393194 -19852 393280 -19796
rect 393336 -19852 393408 -19796
rect 393068 -19938 393408 -19852
rect 393068 -19994 393138 -19938
rect 393194 -19994 393280 -19938
rect 393336 -19994 393408 -19938
rect 393068 -20080 393408 -19994
rect 393068 -20136 393138 -20080
rect 393194 -20136 393280 -20080
rect 393336 -20136 393408 -20080
rect 393068 -20222 393408 -20136
rect 393068 -20278 393138 -20222
rect 393194 -20278 393280 -20222
rect 393336 -20278 393408 -20222
rect 393068 -20364 393408 -20278
rect 393068 -20420 393138 -20364
rect 393194 -20420 393280 -20364
rect 393336 -20420 393408 -20364
rect 393068 -20506 393408 -20420
rect 393068 -20562 393138 -20506
rect 393194 -20562 393280 -20506
rect 393336 -20562 393408 -20506
rect 393068 -20648 393408 -20562
rect 393068 -20704 393138 -20648
rect 393194 -20704 393280 -20648
rect 393336 -20704 393408 -20648
rect 393068 -20790 393408 -20704
rect 393068 -20846 393138 -20790
rect 393194 -20846 393280 -20790
rect 393336 -20846 393408 -20790
rect 393068 -20932 393408 -20846
rect 393068 -20988 393138 -20932
rect 393194 -20988 393280 -20932
rect 393336 -20988 393408 -20932
rect 393068 -21074 393408 -20988
rect 393068 -21130 393138 -21074
rect 393194 -21130 393280 -21074
rect 393336 -21130 393408 -21074
rect 393068 -21216 393408 -21130
rect 393068 -21272 393138 -21216
rect 393194 -21272 393280 -21216
rect 393336 -21272 393408 -21216
rect 393068 -21358 393408 -21272
rect 393068 -21414 393138 -21358
rect 393194 -21414 393280 -21358
rect 393336 -21414 393408 -21358
rect 393068 -21500 393408 -21414
rect 393068 -21556 393138 -21500
rect 393194 -21556 393280 -21500
rect 393336 -21556 393408 -21500
rect 393068 -21642 393408 -21556
rect 393068 -21698 393138 -21642
rect 393194 -21698 393280 -21642
rect 393336 -21698 393408 -21642
rect 393068 -21784 393408 -21698
rect 393068 -21840 393138 -21784
rect 393194 -21840 393280 -21784
rect 393336 -21840 393408 -21784
rect 393068 -21926 393408 -21840
rect 393068 -21982 393138 -21926
rect 393194 -21982 393280 -21926
rect 393336 -21982 393408 -21926
rect 393068 -22068 393408 -21982
rect 393068 -22124 393138 -22068
rect 393194 -22124 393280 -22068
rect 393336 -22124 393408 -22068
rect 393068 -22210 393408 -22124
rect 393068 -22266 393138 -22210
rect 393194 -22266 393280 -22210
rect 393336 -22266 393408 -22210
rect 393068 -22352 393408 -22266
rect 393068 -22408 393138 -22352
rect 393194 -22408 393280 -22352
rect 393336 -22408 393408 -22352
rect 393068 -22494 393408 -22408
rect 393068 -22550 393138 -22494
rect 393194 -22550 393280 -22494
rect 393336 -22550 393408 -22494
rect 393068 -22636 393408 -22550
rect 393068 -22692 393138 -22636
rect 393194 -22692 393280 -22636
rect 393336 -22692 393408 -22636
rect 393068 -22778 393408 -22692
rect 393068 -22834 393138 -22778
rect 393194 -22834 393280 -22778
rect 393336 -22834 393408 -22778
rect 393068 -22920 393408 -22834
rect 393068 -22976 393138 -22920
rect 393194 -22976 393280 -22920
rect 393336 -22976 393408 -22920
rect 393068 -23062 393408 -22976
rect 393068 -23118 393138 -23062
rect 393194 -23118 393280 -23062
rect 393336 -23118 393408 -23062
rect 393068 -23204 393408 -23118
rect 393068 -23260 393138 -23204
rect 393194 -23260 393280 -23204
rect 393336 -23260 393408 -23204
rect 393068 -23346 393408 -23260
rect 393068 -23402 393138 -23346
rect 393194 -23402 393280 -23346
rect 393336 -23402 393408 -23346
rect 393068 -23488 393408 -23402
rect 393068 -23544 393138 -23488
rect 393194 -23544 393280 -23488
rect 393336 -23544 393408 -23488
rect 393068 -23630 393408 -23544
rect 393068 -23686 393138 -23630
rect 393194 -23686 393280 -23630
rect 393336 -23686 393408 -23630
rect 393068 -23772 393408 -23686
rect 393068 -23828 393138 -23772
rect 393194 -23828 393280 -23772
rect 393336 -23828 393408 -23772
rect 393068 -23914 393408 -23828
rect 393068 -23970 393138 -23914
rect 393194 -23970 393280 -23914
rect 393336 -23970 393408 -23914
rect 393068 -24056 393408 -23970
rect 393068 -24112 393138 -24056
rect 393194 -24112 393280 -24056
rect 393336 -24112 393408 -24056
rect 393068 -24198 393408 -24112
rect 393068 -24254 393138 -24198
rect 393194 -24254 393280 -24198
rect 393336 -24254 393408 -24198
rect 393068 -24340 393408 -24254
rect 393068 -24396 393138 -24340
rect 393194 -24396 393280 -24340
rect 393336 -24396 393408 -24340
rect 393068 -24482 393408 -24396
rect 393068 -24538 393138 -24482
rect 393194 -24538 393280 -24482
rect 393336 -24538 393408 -24482
rect 393068 -24624 393408 -24538
rect 393068 -24680 393138 -24624
rect 393194 -24680 393280 -24624
rect 393336 -24680 393408 -24624
rect 393068 -24766 393408 -24680
rect 393068 -24822 393138 -24766
rect 393194 -24822 393280 -24766
rect 393336 -24822 393408 -24766
rect 393068 -24908 393408 -24822
rect 393068 -24964 393138 -24908
rect 393194 -24964 393280 -24908
rect 393336 -24964 393408 -24908
rect 393068 -25050 393408 -24964
rect 393068 -25106 393138 -25050
rect 393194 -25106 393280 -25050
rect 393336 -25106 393408 -25050
rect 393068 -25192 393408 -25106
rect 393068 -25248 393138 -25192
rect 393194 -25248 393280 -25192
rect 393336 -25248 393408 -25192
rect 393068 -25334 393408 -25248
rect 393068 -25390 393138 -25334
rect 393194 -25390 393280 -25334
rect 393336 -25390 393408 -25334
rect 393068 -25476 393408 -25390
rect 393068 -25532 393138 -25476
rect 393194 -25532 393280 -25476
rect 393336 -25532 393408 -25476
rect 393068 -25600 393408 -25532
rect 393468 -17950 393808 -17740
rect 393468 -18006 393543 -17950
rect 393599 -18006 393685 -17950
rect 393741 -18006 393808 -17950
rect 393468 -18092 393808 -18006
rect 393468 -18148 393543 -18092
rect 393599 -18148 393685 -18092
rect 393741 -18148 393808 -18092
rect 393468 -18234 393808 -18148
rect 393468 -18290 393543 -18234
rect 393599 -18290 393685 -18234
rect 393741 -18290 393808 -18234
rect 393468 -18376 393808 -18290
rect 393468 -18432 393543 -18376
rect 393599 -18432 393685 -18376
rect 393741 -18432 393808 -18376
rect 393468 -18518 393808 -18432
rect 393468 -18574 393543 -18518
rect 393599 -18574 393685 -18518
rect 393741 -18574 393808 -18518
rect 393468 -18660 393808 -18574
rect 393468 -18716 393543 -18660
rect 393599 -18716 393685 -18660
rect 393741 -18716 393808 -18660
rect 393468 -18802 393808 -18716
rect 393468 -18858 393543 -18802
rect 393599 -18858 393685 -18802
rect 393741 -18858 393808 -18802
rect 393468 -18944 393808 -18858
rect 393468 -19000 393543 -18944
rect 393599 -19000 393685 -18944
rect 393741 -19000 393808 -18944
rect 393468 -19086 393808 -19000
rect 393468 -19142 393543 -19086
rect 393599 -19142 393685 -19086
rect 393741 -19142 393808 -19086
rect 393468 -19228 393808 -19142
rect 393468 -19284 393543 -19228
rect 393599 -19284 393685 -19228
rect 393741 -19284 393808 -19228
rect 393468 -19370 393808 -19284
rect 393468 -19426 393543 -19370
rect 393599 -19426 393685 -19370
rect 393741 -19426 393808 -19370
rect 393468 -19512 393808 -19426
rect 393468 -19568 393543 -19512
rect 393599 -19568 393685 -19512
rect 393741 -19568 393808 -19512
rect 393468 -19654 393808 -19568
rect 393468 -19710 393543 -19654
rect 393599 -19710 393685 -19654
rect 393741 -19710 393808 -19654
rect 393468 -19796 393808 -19710
rect 393468 -19852 393543 -19796
rect 393599 -19852 393685 -19796
rect 393741 -19852 393808 -19796
rect 393468 -19938 393808 -19852
rect 393468 -19994 393543 -19938
rect 393599 -19994 393685 -19938
rect 393741 -19994 393808 -19938
rect 393468 -20080 393808 -19994
rect 393468 -20136 393543 -20080
rect 393599 -20136 393685 -20080
rect 393741 -20136 393808 -20080
rect 393468 -20222 393808 -20136
rect 393468 -20278 393543 -20222
rect 393599 -20278 393685 -20222
rect 393741 -20278 393808 -20222
rect 393468 -20364 393808 -20278
rect 393468 -20420 393543 -20364
rect 393599 -20420 393685 -20364
rect 393741 -20420 393808 -20364
rect 393468 -20506 393808 -20420
rect 393468 -20562 393543 -20506
rect 393599 -20562 393685 -20506
rect 393741 -20562 393808 -20506
rect 393468 -20648 393808 -20562
rect 393468 -20704 393543 -20648
rect 393599 -20704 393685 -20648
rect 393741 -20704 393808 -20648
rect 393468 -20790 393808 -20704
rect 393468 -20846 393543 -20790
rect 393599 -20846 393685 -20790
rect 393741 -20846 393808 -20790
rect 393468 -20932 393808 -20846
rect 393468 -20988 393543 -20932
rect 393599 -20988 393685 -20932
rect 393741 -20988 393808 -20932
rect 393468 -21074 393808 -20988
rect 393468 -21130 393543 -21074
rect 393599 -21130 393685 -21074
rect 393741 -21130 393808 -21074
rect 393468 -21216 393808 -21130
rect 393468 -21272 393543 -21216
rect 393599 -21272 393685 -21216
rect 393741 -21272 393808 -21216
rect 393468 -21358 393808 -21272
rect 393468 -21414 393543 -21358
rect 393599 -21414 393685 -21358
rect 393741 -21414 393808 -21358
rect 393468 -21500 393808 -21414
rect 393468 -21556 393543 -21500
rect 393599 -21556 393685 -21500
rect 393741 -21556 393808 -21500
rect 393468 -21642 393808 -21556
rect 393468 -21698 393543 -21642
rect 393599 -21698 393685 -21642
rect 393741 -21698 393808 -21642
rect 393468 -21784 393808 -21698
rect 393468 -21840 393543 -21784
rect 393599 -21840 393685 -21784
rect 393741 -21840 393808 -21784
rect 393468 -21926 393808 -21840
rect 393468 -21982 393543 -21926
rect 393599 -21982 393685 -21926
rect 393741 -21982 393808 -21926
rect 393468 -22068 393808 -21982
rect 393468 -22124 393543 -22068
rect 393599 -22124 393685 -22068
rect 393741 -22124 393808 -22068
rect 393468 -22210 393808 -22124
rect 393468 -22266 393543 -22210
rect 393599 -22266 393685 -22210
rect 393741 -22266 393808 -22210
rect 393468 -22352 393808 -22266
rect 393468 -22408 393543 -22352
rect 393599 -22408 393685 -22352
rect 393741 -22408 393808 -22352
rect 393468 -22494 393808 -22408
rect 393468 -22550 393543 -22494
rect 393599 -22550 393685 -22494
rect 393741 -22550 393808 -22494
rect 393468 -22636 393808 -22550
rect 393468 -22692 393543 -22636
rect 393599 -22692 393685 -22636
rect 393741 -22692 393808 -22636
rect 393468 -22778 393808 -22692
rect 393468 -22834 393543 -22778
rect 393599 -22834 393685 -22778
rect 393741 -22834 393808 -22778
rect 393468 -22920 393808 -22834
rect 393468 -22976 393543 -22920
rect 393599 -22976 393685 -22920
rect 393741 -22976 393808 -22920
rect 393468 -23062 393808 -22976
rect 393468 -23118 393543 -23062
rect 393599 -23118 393685 -23062
rect 393741 -23118 393808 -23062
rect 393468 -23204 393808 -23118
rect 393468 -23260 393543 -23204
rect 393599 -23260 393685 -23204
rect 393741 -23260 393808 -23204
rect 393468 -23346 393808 -23260
rect 393468 -23402 393543 -23346
rect 393599 -23402 393685 -23346
rect 393741 -23402 393808 -23346
rect 393468 -23488 393808 -23402
rect 393468 -23544 393543 -23488
rect 393599 -23544 393685 -23488
rect 393741 -23544 393808 -23488
rect 393468 -23630 393808 -23544
rect 393468 -23686 393543 -23630
rect 393599 -23686 393685 -23630
rect 393741 -23686 393808 -23630
rect 393468 -23772 393808 -23686
rect 393468 -23828 393543 -23772
rect 393599 -23828 393685 -23772
rect 393741 -23828 393808 -23772
rect 393468 -23914 393808 -23828
rect 393468 -23970 393543 -23914
rect 393599 -23970 393685 -23914
rect 393741 -23970 393808 -23914
rect 393468 -24056 393808 -23970
rect 393468 -24112 393543 -24056
rect 393599 -24112 393685 -24056
rect 393741 -24112 393808 -24056
rect 393468 -24198 393808 -24112
rect 393468 -24254 393543 -24198
rect 393599 -24254 393685 -24198
rect 393741 -24254 393808 -24198
rect 393468 -24340 393808 -24254
rect 393468 -24396 393543 -24340
rect 393599 -24396 393685 -24340
rect 393741 -24396 393808 -24340
rect 393468 -24482 393808 -24396
rect 393468 -24538 393543 -24482
rect 393599 -24538 393685 -24482
rect 393741 -24538 393808 -24482
rect 393468 -24624 393808 -24538
rect 393468 -24680 393543 -24624
rect 393599 -24680 393685 -24624
rect 393741 -24680 393808 -24624
rect 393468 -24766 393808 -24680
rect 393468 -24822 393543 -24766
rect 393599 -24822 393685 -24766
rect 393741 -24822 393808 -24766
rect 393468 -24908 393808 -24822
rect 393468 -24964 393543 -24908
rect 393599 -24964 393685 -24908
rect 393741 -24964 393808 -24908
rect 393468 -25050 393808 -24964
rect 393468 -25106 393543 -25050
rect 393599 -25106 393685 -25050
rect 393741 -25106 393808 -25050
rect 393468 -25192 393808 -25106
rect 393468 -25248 393543 -25192
rect 393599 -25248 393685 -25192
rect 393741 -25248 393808 -25192
rect 393468 -25334 393808 -25248
rect 393468 -25390 393543 -25334
rect 393599 -25390 393685 -25334
rect 393741 -25390 393808 -25334
rect 393468 -25476 393808 -25390
rect 393468 -25532 393543 -25476
rect 393599 -25532 393685 -25476
rect 393741 -25532 393808 -25476
rect 393468 -25600 393808 -25532
rect 393868 -17950 394208 -17740
rect 393868 -18006 393940 -17950
rect 393996 -18006 394082 -17950
rect 394138 -18006 394208 -17950
rect 393868 -18092 394208 -18006
rect 393868 -18148 393940 -18092
rect 393996 -18148 394082 -18092
rect 394138 -18148 394208 -18092
rect 393868 -18234 394208 -18148
rect 393868 -18290 393940 -18234
rect 393996 -18290 394082 -18234
rect 394138 -18290 394208 -18234
rect 393868 -18376 394208 -18290
rect 393868 -18432 393940 -18376
rect 393996 -18432 394082 -18376
rect 394138 -18432 394208 -18376
rect 393868 -18518 394208 -18432
rect 393868 -18574 393940 -18518
rect 393996 -18574 394082 -18518
rect 394138 -18574 394208 -18518
rect 393868 -18660 394208 -18574
rect 393868 -18716 393940 -18660
rect 393996 -18716 394082 -18660
rect 394138 -18716 394208 -18660
rect 393868 -18802 394208 -18716
rect 393868 -18858 393940 -18802
rect 393996 -18858 394082 -18802
rect 394138 -18858 394208 -18802
rect 393868 -18944 394208 -18858
rect 393868 -19000 393940 -18944
rect 393996 -19000 394082 -18944
rect 394138 -19000 394208 -18944
rect 393868 -19086 394208 -19000
rect 393868 -19142 393940 -19086
rect 393996 -19142 394082 -19086
rect 394138 -19142 394208 -19086
rect 393868 -19228 394208 -19142
rect 393868 -19284 393940 -19228
rect 393996 -19284 394082 -19228
rect 394138 -19284 394208 -19228
rect 393868 -19370 394208 -19284
rect 393868 -19426 393940 -19370
rect 393996 -19426 394082 -19370
rect 394138 -19426 394208 -19370
rect 393868 -19512 394208 -19426
rect 393868 -19568 393940 -19512
rect 393996 -19568 394082 -19512
rect 394138 -19568 394208 -19512
rect 393868 -19654 394208 -19568
rect 393868 -19710 393940 -19654
rect 393996 -19710 394082 -19654
rect 394138 -19710 394208 -19654
rect 393868 -19796 394208 -19710
rect 393868 -19852 393940 -19796
rect 393996 -19852 394082 -19796
rect 394138 -19852 394208 -19796
rect 393868 -19938 394208 -19852
rect 393868 -19994 393940 -19938
rect 393996 -19994 394082 -19938
rect 394138 -19994 394208 -19938
rect 393868 -20080 394208 -19994
rect 393868 -20136 393940 -20080
rect 393996 -20136 394082 -20080
rect 394138 -20136 394208 -20080
rect 393868 -20222 394208 -20136
rect 393868 -20278 393940 -20222
rect 393996 -20278 394082 -20222
rect 394138 -20278 394208 -20222
rect 393868 -20364 394208 -20278
rect 393868 -20420 393940 -20364
rect 393996 -20420 394082 -20364
rect 394138 -20420 394208 -20364
rect 393868 -20506 394208 -20420
rect 393868 -20562 393940 -20506
rect 393996 -20562 394082 -20506
rect 394138 -20562 394208 -20506
rect 393868 -20648 394208 -20562
rect 393868 -20704 393940 -20648
rect 393996 -20704 394082 -20648
rect 394138 -20704 394208 -20648
rect 393868 -20790 394208 -20704
rect 393868 -20846 393940 -20790
rect 393996 -20846 394082 -20790
rect 394138 -20846 394208 -20790
rect 393868 -20932 394208 -20846
rect 393868 -20988 393940 -20932
rect 393996 -20988 394082 -20932
rect 394138 -20988 394208 -20932
rect 393868 -21074 394208 -20988
rect 393868 -21130 393940 -21074
rect 393996 -21130 394082 -21074
rect 394138 -21130 394208 -21074
rect 393868 -21216 394208 -21130
rect 393868 -21272 393940 -21216
rect 393996 -21272 394082 -21216
rect 394138 -21272 394208 -21216
rect 393868 -21358 394208 -21272
rect 393868 -21414 393940 -21358
rect 393996 -21414 394082 -21358
rect 394138 -21414 394208 -21358
rect 393868 -21500 394208 -21414
rect 393868 -21556 393940 -21500
rect 393996 -21556 394082 -21500
rect 394138 -21556 394208 -21500
rect 393868 -21642 394208 -21556
rect 393868 -21698 393940 -21642
rect 393996 -21698 394082 -21642
rect 394138 -21698 394208 -21642
rect 393868 -21784 394208 -21698
rect 393868 -21840 393940 -21784
rect 393996 -21840 394082 -21784
rect 394138 -21840 394208 -21784
rect 393868 -21926 394208 -21840
rect 393868 -21982 393940 -21926
rect 393996 -21982 394082 -21926
rect 394138 -21982 394208 -21926
rect 393868 -22068 394208 -21982
rect 393868 -22124 393940 -22068
rect 393996 -22124 394082 -22068
rect 394138 -22124 394208 -22068
rect 393868 -22210 394208 -22124
rect 393868 -22266 393940 -22210
rect 393996 -22266 394082 -22210
rect 394138 -22266 394208 -22210
rect 393868 -22352 394208 -22266
rect 393868 -22408 393940 -22352
rect 393996 -22408 394082 -22352
rect 394138 -22408 394208 -22352
rect 393868 -22494 394208 -22408
rect 393868 -22550 393940 -22494
rect 393996 -22550 394082 -22494
rect 394138 -22550 394208 -22494
rect 393868 -22636 394208 -22550
rect 393868 -22692 393940 -22636
rect 393996 -22692 394082 -22636
rect 394138 -22692 394208 -22636
rect 393868 -22778 394208 -22692
rect 393868 -22834 393940 -22778
rect 393996 -22834 394082 -22778
rect 394138 -22834 394208 -22778
rect 393868 -22920 394208 -22834
rect 393868 -22976 393940 -22920
rect 393996 -22976 394082 -22920
rect 394138 -22976 394208 -22920
rect 393868 -23062 394208 -22976
rect 393868 -23118 393940 -23062
rect 393996 -23118 394082 -23062
rect 394138 -23118 394208 -23062
rect 393868 -23204 394208 -23118
rect 393868 -23260 393940 -23204
rect 393996 -23260 394082 -23204
rect 394138 -23260 394208 -23204
rect 393868 -23346 394208 -23260
rect 393868 -23402 393940 -23346
rect 393996 -23402 394082 -23346
rect 394138 -23402 394208 -23346
rect 393868 -23488 394208 -23402
rect 393868 -23544 393940 -23488
rect 393996 -23544 394082 -23488
rect 394138 -23544 394208 -23488
rect 393868 -23630 394208 -23544
rect 393868 -23686 393940 -23630
rect 393996 -23686 394082 -23630
rect 394138 -23686 394208 -23630
rect 393868 -23772 394208 -23686
rect 393868 -23828 393940 -23772
rect 393996 -23828 394082 -23772
rect 394138 -23828 394208 -23772
rect 393868 -23914 394208 -23828
rect 393868 -23970 393940 -23914
rect 393996 -23970 394082 -23914
rect 394138 -23970 394208 -23914
rect 393868 -24056 394208 -23970
rect 393868 -24112 393940 -24056
rect 393996 -24112 394082 -24056
rect 394138 -24112 394208 -24056
rect 393868 -24198 394208 -24112
rect 393868 -24254 393940 -24198
rect 393996 -24254 394082 -24198
rect 394138 -24254 394208 -24198
rect 393868 -24340 394208 -24254
rect 393868 -24396 393940 -24340
rect 393996 -24396 394082 -24340
rect 394138 -24396 394208 -24340
rect 393868 -24482 394208 -24396
rect 393868 -24538 393940 -24482
rect 393996 -24538 394082 -24482
rect 394138 -24538 394208 -24482
rect 393868 -24624 394208 -24538
rect 393868 -24680 393940 -24624
rect 393996 -24680 394082 -24624
rect 394138 -24680 394208 -24624
rect 393868 -24766 394208 -24680
rect 393868 -24822 393940 -24766
rect 393996 -24822 394082 -24766
rect 394138 -24822 394208 -24766
rect 393868 -24908 394208 -24822
rect 393868 -24964 393940 -24908
rect 393996 -24964 394082 -24908
rect 394138 -24964 394208 -24908
rect 393868 -25050 394208 -24964
rect 393868 -25106 393940 -25050
rect 393996 -25106 394082 -25050
rect 394138 -25106 394208 -25050
rect 393868 -25192 394208 -25106
rect 393868 -25248 393940 -25192
rect 393996 -25248 394082 -25192
rect 394138 -25248 394208 -25192
rect 393868 -25334 394208 -25248
rect 393868 -25390 393940 -25334
rect 393996 -25390 394082 -25334
rect 394138 -25390 394208 -25334
rect 393868 -25476 394208 -25390
rect 393868 -25532 393940 -25476
rect 393996 -25532 394082 -25476
rect 394138 -25532 394208 -25476
rect 393868 -25600 394208 -25532
rect 394268 -17950 394608 -17740
rect 394268 -18006 394337 -17950
rect 394393 -18006 394479 -17950
rect 394535 -18006 394608 -17950
rect 394268 -18092 394608 -18006
rect 394268 -18148 394337 -18092
rect 394393 -18148 394479 -18092
rect 394535 -18148 394608 -18092
rect 394268 -18234 394608 -18148
rect 394268 -18290 394337 -18234
rect 394393 -18290 394479 -18234
rect 394535 -18290 394608 -18234
rect 394268 -18376 394608 -18290
rect 394268 -18432 394337 -18376
rect 394393 -18432 394479 -18376
rect 394535 -18432 394608 -18376
rect 394268 -18518 394608 -18432
rect 394268 -18574 394337 -18518
rect 394393 -18574 394479 -18518
rect 394535 -18574 394608 -18518
rect 394268 -18660 394608 -18574
rect 394268 -18716 394337 -18660
rect 394393 -18716 394479 -18660
rect 394535 -18716 394608 -18660
rect 394268 -18802 394608 -18716
rect 394268 -18858 394337 -18802
rect 394393 -18858 394479 -18802
rect 394535 -18858 394608 -18802
rect 394268 -18944 394608 -18858
rect 394268 -19000 394337 -18944
rect 394393 -19000 394479 -18944
rect 394535 -19000 394608 -18944
rect 394268 -19086 394608 -19000
rect 394268 -19142 394337 -19086
rect 394393 -19142 394479 -19086
rect 394535 -19142 394608 -19086
rect 394268 -19228 394608 -19142
rect 394268 -19284 394337 -19228
rect 394393 -19284 394479 -19228
rect 394535 -19284 394608 -19228
rect 394268 -19370 394608 -19284
rect 394268 -19426 394337 -19370
rect 394393 -19426 394479 -19370
rect 394535 -19426 394608 -19370
rect 394268 -19512 394608 -19426
rect 394268 -19568 394337 -19512
rect 394393 -19568 394479 -19512
rect 394535 -19568 394608 -19512
rect 394268 -19654 394608 -19568
rect 394268 -19710 394337 -19654
rect 394393 -19710 394479 -19654
rect 394535 -19710 394608 -19654
rect 394268 -19796 394608 -19710
rect 394268 -19852 394337 -19796
rect 394393 -19852 394479 -19796
rect 394535 -19852 394608 -19796
rect 394268 -19938 394608 -19852
rect 394268 -19994 394337 -19938
rect 394393 -19994 394479 -19938
rect 394535 -19994 394608 -19938
rect 394268 -20080 394608 -19994
rect 394268 -20136 394337 -20080
rect 394393 -20136 394479 -20080
rect 394535 -20136 394608 -20080
rect 394268 -20222 394608 -20136
rect 394268 -20278 394337 -20222
rect 394393 -20278 394479 -20222
rect 394535 -20278 394608 -20222
rect 394268 -20364 394608 -20278
rect 394268 -20420 394337 -20364
rect 394393 -20420 394479 -20364
rect 394535 -20420 394608 -20364
rect 394268 -20506 394608 -20420
rect 394268 -20562 394337 -20506
rect 394393 -20562 394479 -20506
rect 394535 -20562 394608 -20506
rect 394268 -20648 394608 -20562
rect 394268 -20704 394337 -20648
rect 394393 -20704 394479 -20648
rect 394535 -20704 394608 -20648
rect 394268 -20790 394608 -20704
rect 394268 -20846 394337 -20790
rect 394393 -20846 394479 -20790
rect 394535 -20846 394608 -20790
rect 394268 -20932 394608 -20846
rect 394268 -20988 394337 -20932
rect 394393 -20988 394479 -20932
rect 394535 -20988 394608 -20932
rect 394268 -21074 394608 -20988
rect 394268 -21130 394337 -21074
rect 394393 -21130 394479 -21074
rect 394535 -21130 394608 -21074
rect 394268 -21216 394608 -21130
rect 394268 -21272 394337 -21216
rect 394393 -21272 394479 -21216
rect 394535 -21272 394608 -21216
rect 394268 -21358 394608 -21272
rect 394268 -21414 394337 -21358
rect 394393 -21414 394479 -21358
rect 394535 -21414 394608 -21358
rect 394268 -21500 394608 -21414
rect 394268 -21556 394337 -21500
rect 394393 -21556 394479 -21500
rect 394535 -21556 394608 -21500
rect 394268 -21642 394608 -21556
rect 394268 -21698 394337 -21642
rect 394393 -21698 394479 -21642
rect 394535 -21698 394608 -21642
rect 394268 -21784 394608 -21698
rect 394268 -21840 394337 -21784
rect 394393 -21840 394479 -21784
rect 394535 -21840 394608 -21784
rect 394268 -21926 394608 -21840
rect 394268 -21982 394337 -21926
rect 394393 -21982 394479 -21926
rect 394535 -21982 394608 -21926
rect 394268 -22068 394608 -21982
rect 394268 -22124 394337 -22068
rect 394393 -22124 394479 -22068
rect 394535 -22124 394608 -22068
rect 394268 -22210 394608 -22124
rect 394268 -22266 394337 -22210
rect 394393 -22266 394479 -22210
rect 394535 -22266 394608 -22210
rect 394268 -22352 394608 -22266
rect 394268 -22408 394337 -22352
rect 394393 -22408 394479 -22352
rect 394535 -22408 394608 -22352
rect 394268 -22494 394608 -22408
rect 394268 -22550 394337 -22494
rect 394393 -22550 394479 -22494
rect 394535 -22550 394608 -22494
rect 394268 -22636 394608 -22550
rect 394268 -22692 394337 -22636
rect 394393 -22692 394479 -22636
rect 394535 -22692 394608 -22636
rect 394268 -22778 394608 -22692
rect 394268 -22834 394337 -22778
rect 394393 -22834 394479 -22778
rect 394535 -22834 394608 -22778
rect 394268 -22920 394608 -22834
rect 394268 -22976 394337 -22920
rect 394393 -22976 394479 -22920
rect 394535 -22976 394608 -22920
rect 394268 -23062 394608 -22976
rect 394268 -23118 394337 -23062
rect 394393 -23118 394479 -23062
rect 394535 -23118 394608 -23062
rect 394268 -23204 394608 -23118
rect 394268 -23260 394337 -23204
rect 394393 -23260 394479 -23204
rect 394535 -23260 394608 -23204
rect 394268 -23346 394608 -23260
rect 394268 -23402 394337 -23346
rect 394393 -23402 394479 -23346
rect 394535 -23402 394608 -23346
rect 394268 -23488 394608 -23402
rect 394268 -23544 394337 -23488
rect 394393 -23544 394479 -23488
rect 394535 -23544 394608 -23488
rect 394268 -23630 394608 -23544
rect 394268 -23686 394337 -23630
rect 394393 -23686 394479 -23630
rect 394535 -23686 394608 -23630
rect 394268 -23772 394608 -23686
rect 394268 -23828 394337 -23772
rect 394393 -23828 394479 -23772
rect 394535 -23828 394608 -23772
rect 394268 -23914 394608 -23828
rect 394268 -23970 394337 -23914
rect 394393 -23970 394479 -23914
rect 394535 -23970 394608 -23914
rect 394268 -24056 394608 -23970
rect 394268 -24112 394337 -24056
rect 394393 -24112 394479 -24056
rect 394535 -24112 394608 -24056
rect 394268 -24198 394608 -24112
rect 394268 -24254 394337 -24198
rect 394393 -24254 394479 -24198
rect 394535 -24254 394608 -24198
rect 394268 -24340 394608 -24254
rect 394268 -24396 394337 -24340
rect 394393 -24396 394479 -24340
rect 394535 -24396 394608 -24340
rect 394268 -24482 394608 -24396
rect 394268 -24538 394337 -24482
rect 394393 -24538 394479 -24482
rect 394535 -24538 394608 -24482
rect 394268 -24624 394608 -24538
rect 394268 -24680 394337 -24624
rect 394393 -24680 394479 -24624
rect 394535 -24680 394608 -24624
rect 394268 -24766 394608 -24680
rect 394268 -24822 394337 -24766
rect 394393 -24822 394479 -24766
rect 394535 -24822 394608 -24766
rect 394268 -24908 394608 -24822
rect 394268 -24964 394337 -24908
rect 394393 -24964 394479 -24908
rect 394535 -24964 394608 -24908
rect 394268 -25050 394608 -24964
rect 394268 -25106 394337 -25050
rect 394393 -25106 394479 -25050
rect 394535 -25106 394608 -25050
rect 394268 -25192 394608 -25106
rect 394268 -25248 394337 -25192
rect 394393 -25248 394479 -25192
rect 394535 -25248 394608 -25192
rect 394268 -25334 394608 -25248
rect 394268 -25390 394337 -25334
rect 394393 -25390 394479 -25334
rect 394535 -25390 394608 -25334
rect 394268 -25476 394608 -25390
rect 394268 -25532 394337 -25476
rect 394393 -25532 394479 -25476
rect 394535 -25532 394608 -25476
rect 394268 -25600 394608 -25532
rect 394668 -17950 395008 -17740
rect 394668 -18006 394740 -17950
rect 394796 -18006 394882 -17950
rect 394938 -18006 395008 -17950
rect 394668 -18092 395008 -18006
rect 394668 -18148 394740 -18092
rect 394796 -18148 394882 -18092
rect 394938 -18148 395008 -18092
rect 394668 -18234 395008 -18148
rect 394668 -18290 394740 -18234
rect 394796 -18290 394882 -18234
rect 394938 -18290 395008 -18234
rect 394668 -18376 395008 -18290
rect 394668 -18432 394740 -18376
rect 394796 -18432 394882 -18376
rect 394938 -18432 395008 -18376
rect 394668 -18518 395008 -18432
rect 394668 -18574 394740 -18518
rect 394796 -18574 394882 -18518
rect 394938 -18574 395008 -18518
rect 394668 -18660 395008 -18574
rect 394668 -18716 394740 -18660
rect 394796 -18716 394882 -18660
rect 394938 -18716 395008 -18660
rect 394668 -18802 395008 -18716
rect 394668 -18858 394740 -18802
rect 394796 -18858 394882 -18802
rect 394938 -18858 395008 -18802
rect 394668 -18944 395008 -18858
rect 394668 -19000 394740 -18944
rect 394796 -19000 394882 -18944
rect 394938 -19000 395008 -18944
rect 394668 -19086 395008 -19000
rect 394668 -19142 394740 -19086
rect 394796 -19142 394882 -19086
rect 394938 -19142 395008 -19086
rect 394668 -19228 395008 -19142
rect 394668 -19284 394740 -19228
rect 394796 -19284 394882 -19228
rect 394938 -19284 395008 -19228
rect 394668 -19370 395008 -19284
rect 394668 -19426 394740 -19370
rect 394796 -19426 394882 -19370
rect 394938 -19426 395008 -19370
rect 394668 -19512 395008 -19426
rect 394668 -19568 394740 -19512
rect 394796 -19568 394882 -19512
rect 394938 -19568 395008 -19512
rect 394668 -19654 395008 -19568
rect 394668 -19710 394740 -19654
rect 394796 -19710 394882 -19654
rect 394938 -19710 395008 -19654
rect 394668 -19796 395008 -19710
rect 394668 -19852 394740 -19796
rect 394796 -19852 394882 -19796
rect 394938 -19852 395008 -19796
rect 394668 -19938 395008 -19852
rect 394668 -19994 394740 -19938
rect 394796 -19994 394882 -19938
rect 394938 -19994 395008 -19938
rect 394668 -20080 395008 -19994
rect 394668 -20136 394740 -20080
rect 394796 -20136 394882 -20080
rect 394938 -20136 395008 -20080
rect 394668 -20222 395008 -20136
rect 394668 -20278 394740 -20222
rect 394796 -20278 394882 -20222
rect 394938 -20278 395008 -20222
rect 394668 -20364 395008 -20278
rect 394668 -20420 394740 -20364
rect 394796 -20420 394882 -20364
rect 394938 -20420 395008 -20364
rect 394668 -20506 395008 -20420
rect 394668 -20562 394740 -20506
rect 394796 -20562 394882 -20506
rect 394938 -20562 395008 -20506
rect 394668 -20648 395008 -20562
rect 394668 -20704 394740 -20648
rect 394796 -20704 394882 -20648
rect 394938 -20704 395008 -20648
rect 394668 -20790 395008 -20704
rect 394668 -20846 394740 -20790
rect 394796 -20846 394882 -20790
rect 394938 -20846 395008 -20790
rect 394668 -20932 395008 -20846
rect 394668 -20988 394740 -20932
rect 394796 -20988 394882 -20932
rect 394938 -20988 395008 -20932
rect 394668 -21074 395008 -20988
rect 394668 -21130 394740 -21074
rect 394796 -21130 394882 -21074
rect 394938 -21130 395008 -21074
rect 394668 -21216 395008 -21130
rect 394668 -21272 394740 -21216
rect 394796 -21272 394882 -21216
rect 394938 -21272 395008 -21216
rect 394668 -21358 395008 -21272
rect 394668 -21414 394740 -21358
rect 394796 -21414 394882 -21358
rect 394938 -21414 395008 -21358
rect 394668 -21500 395008 -21414
rect 394668 -21556 394740 -21500
rect 394796 -21556 394882 -21500
rect 394938 -21556 395008 -21500
rect 394668 -21642 395008 -21556
rect 394668 -21698 394740 -21642
rect 394796 -21698 394882 -21642
rect 394938 -21698 395008 -21642
rect 394668 -21784 395008 -21698
rect 394668 -21840 394740 -21784
rect 394796 -21840 394882 -21784
rect 394938 -21840 395008 -21784
rect 394668 -21926 395008 -21840
rect 394668 -21982 394740 -21926
rect 394796 -21982 394882 -21926
rect 394938 -21982 395008 -21926
rect 394668 -22068 395008 -21982
rect 394668 -22124 394740 -22068
rect 394796 -22124 394882 -22068
rect 394938 -22124 395008 -22068
rect 394668 -22210 395008 -22124
rect 394668 -22266 394740 -22210
rect 394796 -22266 394882 -22210
rect 394938 -22266 395008 -22210
rect 394668 -22352 395008 -22266
rect 394668 -22408 394740 -22352
rect 394796 -22408 394882 -22352
rect 394938 -22408 395008 -22352
rect 394668 -22494 395008 -22408
rect 394668 -22550 394740 -22494
rect 394796 -22550 394882 -22494
rect 394938 -22550 395008 -22494
rect 394668 -22636 395008 -22550
rect 394668 -22692 394740 -22636
rect 394796 -22692 394882 -22636
rect 394938 -22692 395008 -22636
rect 394668 -22778 395008 -22692
rect 394668 -22834 394740 -22778
rect 394796 -22834 394882 -22778
rect 394938 -22834 395008 -22778
rect 394668 -22920 395008 -22834
rect 394668 -22976 394740 -22920
rect 394796 -22976 394882 -22920
rect 394938 -22976 395008 -22920
rect 394668 -23062 395008 -22976
rect 394668 -23118 394740 -23062
rect 394796 -23118 394882 -23062
rect 394938 -23118 395008 -23062
rect 394668 -23204 395008 -23118
rect 394668 -23260 394740 -23204
rect 394796 -23260 394882 -23204
rect 394938 -23260 395008 -23204
rect 394668 -23346 395008 -23260
rect 394668 -23402 394740 -23346
rect 394796 -23402 394882 -23346
rect 394938 -23402 395008 -23346
rect 394668 -23488 395008 -23402
rect 394668 -23544 394740 -23488
rect 394796 -23544 394882 -23488
rect 394938 -23544 395008 -23488
rect 394668 -23630 395008 -23544
rect 394668 -23686 394740 -23630
rect 394796 -23686 394882 -23630
rect 394938 -23686 395008 -23630
rect 394668 -23772 395008 -23686
rect 394668 -23828 394740 -23772
rect 394796 -23828 394882 -23772
rect 394938 -23828 395008 -23772
rect 394668 -23914 395008 -23828
rect 394668 -23970 394740 -23914
rect 394796 -23970 394882 -23914
rect 394938 -23970 395008 -23914
rect 394668 -24056 395008 -23970
rect 394668 -24112 394740 -24056
rect 394796 -24112 394882 -24056
rect 394938 -24112 395008 -24056
rect 394668 -24198 395008 -24112
rect 394668 -24254 394740 -24198
rect 394796 -24254 394882 -24198
rect 394938 -24254 395008 -24198
rect 394668 -24340 395008 -24254
rect 394668 -24396 394740 -24340
rect 394796 -24396 394882 -24340
rect 394938 -24396 395008 -24340
rect 394668 -24482 395008 -24396
rect 394668 -24538 394740 -24482
rect 394796 -24538 394882 -24482
rect 394938 -24538 395008 -24482
rect 394668 -24624 395008 -24538
rect 394668 -24680 394740 -24624
rect 394796 -24680 394882 -24624
rect 394938 -24680 395008 -24624
rect 394668 -24766 395008 -24680
rect 394668 -24822 394740 -24766
rect 394796 -24822 394882 -24766
rect 394938 -24822 395008 -24766
rect 394668 -24908 395008 -24822
rect 394668 -24964 394740 -24908
rect 394796 -24964 394882 -24908
rect 394938 -24964 395008 -24908
rect 394668 -25050 395008 -24964
rect 394668 -25106 394740 -25050
rect 394796 -25106 394882 -25050
rect 394938 -25106 395008 -25050
rect 394668 -25192 395008 -25106
rect 394668 -25248 394740 -25192
rect 394796 -25248 394882 -25192
rect 394938 -25248 395008 -25192
rect 394668 -25334 395008 -25248
rect 394668 -25390 394740 -25334
rect 394796 -25390 394882 -25334
rect 394938 -25390 395008 -25334
rect 394668 -25476 395008 -25390
rect 394668 -25532 394740 -25476
rect 394796 -25532 394882 -25476
rect 394938 -25532 395008 -25476
rect 394668 -25600 395008 -25532
rect 395068 -17950 395408 -17740
rect 395068 -18006 395142 -17950
rect 395198 -18006 395284 -17950
rect 395340 -18006 395408 -17950
rect 395068 -18092 395408 -18006
rect 395068 -18148 395142 -18092
rect 395198 -18148 395284 -18092
rect 395340 -18148 395408 -18092
rect 395068 -18234 395408 -18148
rect 395068 -18290 395142 -18234
rect 395198 -18290 395284 -18234
rect 395340 -18290 395408 -18234
rect 395068 -18376 395408 -18290
rect 395068 -18432 395142 -18376
rect 395198 -18432 395284 -18376
rect 395340 -18432 395408 -18376
rect 395068 -18518 395408 -18432
rect 395068 -18574 395142 -18518
rect 395198 -18574 395284 -18518
rect 395340 -18574 395408 -18518
rect 395068 -18660 395408 -18574
rect 395068 -18716 395142 -18660
rect 395198 -18716 395284 -18660
rect 395340 -18716 395408 -18660
rect 395068 -18802 395408 -18716
rect 395068 -18858 395142 -18802
rect 395198 -18858 395284 -18802
rect 395340 -18858 395408 -18802
rect 395068 -18944 395408 -18858
rect 395068 -19000 395142 -18944
rect 395198 -19000 395284 -18944
rect 395340 -19000 395408 -18944
rect 395068 -19086 395408 -19000
rect 395068 -19142 395142 -19086
rect 395198 -19142 395284 -19086
rect 395340 -19142 395408 -19086
rect 395068 -19228 395408 -19142
rect 395068 -19284 395142 -19228
rect 395198 -19284 395284 -19228
rect 395340 -19284 395408 -19228
rect 395068 -19370 395408 -19284
rect 395068 -19426 395142 -19370
rect 395198 -19426 395284 -19370
rect 395340 -19426 395408 -19370
rect 395068 -19512 395408 -19426
rect 395068 -19568 395142 -19512
rect 395198 -19568 395284 -19512
rect 395340 -19568 395408 -19512
rect 395068 -19654 395408 -19568
rect 395068 -19710 395142 -19654
rect 395198 -19710 395284 -19654
rect 395340 -19710 395408 -19654
rect 395068 -19796 395408 -19710
rect 395068 -19852 395142 -19796
rect 395198 -19852 395284 -19796
rect 395340 -19852 395408 -19796
rect 395068 -19938 395408 -19852
rect 395068 -19994 395142 -19938
rect 395198 -19994 395284 -19938
rect 395340 -19994 395408 -19938
rect 395068 -20080 395408 -19994
rect 395068 -20136 395142 -20080
rect 395198 -20136 395284 -20080
rect 395340 -20136 395408 -20080
rect 395068 -20222 395408 -20136
rect 395068 -20278 395142 -20222
rect 395198 -20278 395284 -20222
rect 395340 -20278 395408 -20222
rect 395068 -20364 395408 -20278
rect 395068 -20420 395142 -20364
rect 395198 -20420 395284 -20364
rect 395340 -20420 395408 -20364
rect 395068 -20506 395408 -20420
rect 395068 -20562 395142 -20506
rect 395198 -20562 395284 -20506
rect 395340 -20562 395408 -20506
rect 395068 -20648 395408 -20562
rect 395068 -20704 395142 -20648
rect 395198 -20704 395284 -20648
rect 395340 -20704 395408 -20648
rect 395068 -20790 395408 -20704
rect 395068 -20846 395142 -20790
rect 395198 -20846 395284 -20790
rect 395340 -20846 395408 -20790
rect 395068 -20932 395408 -20846
rect 395068 -20988 395142 -20932
rect 395198 -20988 395284 -20932
rect 395340 -20988 395408 -20932
rect 395068 -21074 395408 -20988
rect 395068 -21130 395142 -21074
rect 395198 -21130 395284 -21074
rect 395340 -21130 395408 -21074
rect 395068 -21216 395408 -21130
rect 395068 -21272 395142 -21216
rect 395198 -21272 395284 -21216
rect 395340 -21272 395408 -21216
rect 395068 -21358 395408 -21272
rect 395068 -21414 395142 -21358
rect 395198 -21414 395284 -21358
rect 395340 -21414 395408 -21358
rect 395068 -21500 395408 -21414
rect 395068 -21556 395142 -21500
rect 395198 -21556 395284 -21500
rect 395340 -21556 395408 -21500
rect 395068 -21642 395408 -21556
rect 395068 -21698 395142 -21642
rect 395198 -21698 395284 -21642
rect 395340 -21698 395408 -21642
rect 395068 -21784 395408 -21698
rect 395068 -21840 395142 -21784
rect 395198 -21840 395284 -21784
rect 395340 -21840 395408 -21784
rect 395068 -21926 395408 -21840
rect 395068 -21982 395142 -21926
rect 395198 -21982 395284 -21926
rect 395340 -21982 395408 -21926
rect 395068 -22068 395408 -21982
rect 395068 -22124 395142 -22068
rect 395198 -22124 395284 -22068
rect 395340 -22124 395408 -22068
rect 395068 -22210 395408 -22124
rect 395068 -22266 395142 -22210
rect 395198 -22266 395284 -22210
rect 395340 -22266 395408 -22210
rect 395068 -22352 395408 -22266
rect 395068 -22408 395142 -22352
rect 395198 -22408 395284 -22352
rect 395340 -22408 395408 -22352
rect 395068 -22494 395408 -22408
rect 395068 -22550 395142 -22494
rect 395198 -22550 395284 -22494
rect 395340 -22550 395408 -22494
rect 395068 -22636 395408 -22550
rect 395068 -22692 395142 -22636
rect 395198 -22692 395284 -22636
rect 395340 -22692 395408 -22636
rect 395068 -22778 395408 -22692
rect 395068 -22834 395142 -22778
rect 395198 -22834 395284 -22778
rect 395340 -22834 395408 -22778
rect 395068 -22920 395408 -22834
rect 395068 -22976 395142 -22920
rect 395198 -22976 395284 -22920
rect 395340 -22976 395408 -22920
rect 395068 -23062 395408 -22976
rect 395068 -23118 395142 -23062
rect 395198 -23118 395284 -23062
rect 395340 -23118 395408 -23062
rect 395068 -23204 395408 -23118
rect 395068 -23260 395142 -23204
rect 395198 -23260 395284 -23204
rect 395340 -23260 395408 -23204
rect 395068 -23346 395408 -23260
rect 395068 -23402 395142 -23346
rect 395198 -23402 395284 -23346
rect 395340 -23402 395408 -23346
rect 395068 -23488 395408 -23402
rect 395068 -23544 395142 -23488
rect 395198 -23544 395284 -23488
rect 395340 -23544 395408 -23488
rect 395068 -23630 395408 -23544
rect 395068 -23686 395142 -23630
rect 395198 -23686 395284 -23630
rect 395340 -23686 395408 -23630
rect 395068 -23772 395408 -23686
rect 395068 -23828 395142 -23772
rect 395198 -23828 395284 -23772
rect 395340 -23828 395408 -23772
rect 395068 -23914 395408 -23828
rect 395068 -23970 395142 -23914
rect 395198 -23970 395284 -23914
rect 395340 -23970 395408 -23914
rect 395068 -24056 395408 -23970
rect 395068 -24112 395142 -24056
rect 395198 -24112 395284 -24056
rect 395340 -24112 395408 -24056
rect 395068 -24198 395408 -24112
rect 395068 -24254 395142 -24198
rect 395198 -24254 395284 -24198
rect 395340 -24254 395408 -24198
rect 395068 -24340 395408 -24254
rect 395068 -24396 395142 -24340
rect 395198 -24396 395284 -24340
rect 395340 -24396 395408 -24340
rect 395068 -24482 395408 -24396
rect 395068 -24538 395142 -24482
rect 395198 -24538 395284 -24482
rect 395340 -24538 395408 -24482
rect 395068 -24624 395408 -24538
rect 395068 -24680 395142 -24624
rect 395198 -24680 395284 -24624
rect 395340 -24680 395408 -24624
rect 395068 -24766 395408 -24680
rect 395068 -24822 395142 -24766
rect 395198 -24822 395284 -24766
rect 395340 -24822 395408 -24766
rect 395068 -24908 395408 -24822
rect 395068 -24964 395142 -24908
rect 395198 -24964 395284 -24908
rect 395340 -24964 395408 -24908
rect 395068 -25050 395408 -24964
rect 395068 -25106 395142 -25050
rect 395198 -25106 395284 -25050
rect 395340 -25106 395408 -25050
rect 395068 -25192 395408 -25106
rect 395068 -25248 395142 -25192
rect 395198 -25248 395284 -25192
rect 395340 -25248 395408 -25192
rect 395068 -25334 395408 -25248
rect 395068 -25390 395142 -25334
rect 395198 -25390 395284 -25334
rect 395340 -25390 395408 -25334
rect 395068 -25476 395408 -25390
rect 395068 -25532 395142 -25476
rect 395198 -25532 395284 -25476
rect 395340 -25532 395408 -25476
rect 395068 -25600 395408 -25532
rect 395468 -17950 395808 -17740
rect 395468 -18006 395545 -17950
rect 395601 -18006 395687 -17950
rect 395743 -18006 395808 -17950
rect 395468 -18092 395808 -18006
rect 395468 -18148 395545 -18092
rect 395601 -18148 395687 -18092
rect 395743 -18148 395808 -18092
rect 395468 -18234 395808 -18148
rect 395468 -18290 395545 -18234
rect 395601 -18290 395687 -18234
rect 395743 -18290 395808 -18234
rect 395468 -18376 395808 -18290
rect 395468 -18432 395545 -18376
rect 395601 -18432 395687 -18376
rect 395743 -18432 395808 -18376
rect 395468 -18518 395808 -18432
rect 395468 -18574 395545 -18518
rect 395601 -18574 395687 -18518
rect 395743 -18574 395808 -18518
rect 395468 -18660 395808 -18574
rect 395468 -18716 395545 -18660
rect 395601 -18716 395687 -18660
rect 395743 -18716 395808 -18660
rect 395468 -18802 395808 -18716
rect 395468 -18858 395545 -18802
rect 395601 -18858 395687 -18802
rect 395743 -18858 395808 -18802
rect 395468 -18944 395808 -18858
rect 395468 -19000 395545 -18944
rect 395601 -19000 395687 -18944
rect 395743 -19000 395808 -18944
rect 395468 -19086 395808 -19000
rect 395468 -19142 395545 -19086
rect 395601 -19142 395687 -19086
rect 395743 -19142 395808 -19086
rect 395468 -19228 395808 -19142
rect 395468 -19284 395545 -19228
rect 395601 -19284 395687 -19228
rect 395743 -19284 395808 -19228
rect 395468 -19370 395808 -19284
rect 395468 -19426 395545 -19370
rect 395601 -19426 395687 -19370
rect 395743 -19426 395808 -19370
rect 395468 -19512 395808 -19426
rect 395468 -19568 395545 -19512
rect 395601 -19568 395687 -19512
rect 395743 -19568 395808 -19512
rect 395468 -19654 395808 -19568
rect 395468 -19710 395545 -19654
rect 395601 -19710 395687 -19654
rect 395743 -19710 395808 -19654
rect 395468 -19796 395808 -19710
rect 395468 -19852 395545 -19796
rect 395601 -19852 395687 -19796
rect 395743 -19852 395808 -19796
rect 395468 -19938 395808 -19852
rect 395468 -19994 395545 -19938
rect 395601 -19994 395687 -19938
rect 395743 -19994 395808 -19938
rect 395468 -20080 395808 -19994
rect 395468 -20136 395545 -20080
rect 395601 -20136 395687 -20080
rect 395743 -20136 395808 -20080
rect 395468 -20222 395808 -20136
rect 395468 -20278 395545 -20222
rect 395601 -20278 395687 -20222
rect 395743 -20278 395808 -20222
rect 395468 -20364 395808 -20278
rect 395468 -20420 395545 -20364
rect 395601 -20420 395687 -20364
rect 395743 -20420 395808 -20364
rect 395468 -20506 395808 -20420
rect 395468 -20562 395545 -20506
rect 395601 -20562 395687 -20506
rect 395743 -20562 395808 -20506
rect 395468 -20648 395808 -20562
rect 395468 -20704 395545 -20648
rect 395601 -20704 395687 -20648
rect 395743 -20704 395808 -20648
rect 395468 -20790 395808 -20704
rect 395468 -20846 395545 -20790
rect 395601 -20846 395687 -20790
rect 395743 -20846 395808 -20790
rect 395468 -20932 395808 -20846
rect 395468 -20988 395545 -20932
rect 395601 -20988 395687 -20932
rect 395743 -20988 395808 -20932
rect 395468 -21074 395808 -20988
rect 395468 -21130 395545 -21074
rect 395601 -21130 395687 -21074
rect 395743 -21130 395808 -21074
rect 395468 -21216 395808 -21130
rect 395468 -21272 395545 -21216
rect 395601 -21272 395687 -21216
rect 395743 -21272 395808 -21216
rect 395468 -21358 395808 -21272
rect 395468 -21414 395545 -21358
rect 395601 -21414 395687 -21358
rect 395743 -21414 395808 -21358
rect 395468 -21500 395808 -21414
rect 395468 -21556 395545 -21500
rect 395601 -21556 395687 -21500
rect 395743 -21556 395808 -21500
rect 395468 -21642 395808 -21556
rect 395468 -21698 395545 -21642
rect 395601 -21698 395687 -21642
rect 395743 -21698 395808 -21642
rect 395468 -21784 395808 -21698
rect 395468 -21840 395545 -21784
rect 395601 -21840 395687 -21784
rect 395743 -21840 395808 -21784
rect 395468 -21926 395808 -21840
rect 395468 -21982 395545 -21926
rect 395601 -21982 395687 -21926
rect 395743 -21982 395808 -21926
rect 395468 -22068 395808 -21982
rect 395468 -22124 395545 -22068
rect 395601 -22124 395687 -22068
rect 395743 -22124 395808 -22068
rect 395468 -22210 395808 -22124
rect 395468 -22266 395545 -22210
rect 395601 -22266 395687 -22210
rect 395743 -22266 395808 -22210
rect 395468 -22352 395808 -22266
rect 395468 -22408 395545 -22352
rect 395601 -22408 395687 -22352
rect 395743 -22408 395808 -22352
rect 395468 -22494 395808 -22408
rect 395468 -22550 395545 -22494
rect 395601 -22550 395687 -22494
rect 395743 -22550 395808 -22494
rect 395468 -22636 395808 -22550
rect 395468 -22692 395545 -22636
rect 395601 -22692 395687 -22636
rect 395743 -22692 395808 -22636
rect 395468 -22778 395808 -22692
rect 395468 -22834 395545 -22778
rect 395601 -22834 395687 -22778
rect 395743 -22834 395808 -22778
rect 395468 -22920 395808 -22834
rect 395468 -22976 395545 -22920
rect 395601 -22976 395687 -22920
rect 395743 -22976 395808 -22920
rect 395468 -23062 395808 -22976
rect 395468 -23118 395545 -23062
rect 395601 -23118 395687 -23062
rect 395743 -23118 395808 -23062
rect 395468 -23204 395808 -23118
rect 395468 -23260 395545 -23204
rect 395601 -23260 395687 -23204
rect 395743 -23260 395808 -23204
rect 395468 -23346 395808 -23260
rect 395468 -23402 395545 -23346
rect 395601 -23402 395687 -23346
rect 395743 -23402 395808 -23346
rect 395468 -23488 395808 -23402
rect 395468 -23544 395545 -23488
rect 395601 -23544 395687 -23488
rect 395743 -23544 395808 -23488
rect 395468 -23630 395808 -23544
rect 395468 -23686 395545 -23630
rect 395601 -23686 395687 -23630
rect 395743 -23686 395808 -23630
rect 395468 -23772 395808 -23686
rect 395468 -23828 395545 -23772
rect 395601 -23828 395687 -23772
rect 395743 -23828 395808 -23772
rect 395468 -23914 395808 -23828
rect 395468 -23970 395545 -23914
rect 395601 -23970 395687 -23914
rect 395743 -23970 395808 -23914
rect 395468 -24056 395808 -23970
rect 395468 -24112 395545 -24056
rect 395601 -24112 395687 -24056
rect 395743 -24112 395808 -24056
rect 395468 -24198 395808 -24112
rect 395468 -24254 395545 -24198
rect 395601 -24254 395687 -24198
rect 395743 -24254 395808 -24198
rect 395468 -24340 395808 -24254
rect 395468 -24396 395545 -24340
rect 395601 -24396 395687 -24340
rect 395743 -24396 395808 -24340
rect 395468 -24482 395808 -24396
rect 395468 -24538 395545 -24482
rect 395601 -24538 395687 -24482
rect 395743 -24538 395808 -24482
rect 395468 -24624 395808 -24538
rect 395468 -24680 395545 -24624
rect 395601 -24680 395687 -24624
rect 395743 -24680 395808 -24624
rect 395468 -24766 395808 -24680
rect 395468 -24822 395545 -24766
rect 395601 -24822 395687 -24766
rect 395743 -24822 395808 -24766
rect 395468 -24908 395808 -24822
rect 395468 -24964 395545 -24908
rect 395601 -24964 395687 -24908
rect 395743 -24964 395808 -24908
rect 395468 -25050 395808 -24964
rect 395468 -25106 395545 -25050
rect 395601 -25106 395687 -25050
rect 395743 -25106 395808 -25050
rect 395468 -25192 395808 -25106
rect 395468 -25248 395545 -25192
rect 395601 -25248 395687 -25192
rect 395743 -25248 395808 -25192
rect 395468 -25334 395808 -25248
rect 395468 -25390 395545 -25334
rect 395601 -25390 395687 -25334
rect 395743 -25390 395808 -25334
rect 395468 -25476 395808 -25390
rect 395468 -25532 395545 -25476
rect 395601 -25532 395687 -25476
rect 395743 -25532 395808 -25476
rect 395468 -25600 395808 -25532
rect 395868 -17950 396208 -17740
rect 395868 -18006 395941 -17950
rect 395997 -18006 396083 -17950
rect 396139 -18006 396208 -17950
rect 395868 -18092 396208 -18006
rect 395868 -18148 395941 -18092
rect 395997 -18148 396083 -18092
rect 396139 -18148 396208 -18092
rect 395868 -18234 396208 -18148
rect 395868 -18290 395941 -18234
rect 395997 -18290 396083 -18234
rect 396139 -18290 396208 -18234
rect 395868 -18376 396208 -18290
rect 395868 -18432 395941 -18376
rect 395997 -18432 396083 -18376
rect 396139 -18432 396208 -18376
rect 395868 -18518 396208 -18432
rect 395868 -18574 395941 -18518
rect 395997 -18574 396083 -18518
rect 396139 -18574 396208 -18518
rect 395868 -18660 396208 -18574
rect 395868 -18716 395941 -18660
rect 395997 -18716 396083 -18660
rect 396139 -18716 396208 -18660
rect 395868 -18802 396208 -18716
rect 395868 -18858 395941 -18802
rect 395997 -18858 396083 -18802
rect 396139 -18858 396208 -18802
rect 395868 -18944 396208 -18858
rect 395868 -19000 395941 -18944
rect 395997 -19000 396083 -18944
rect 396139 -19000 396208 -18944
rect 395868 -19086 396208 -19000
rect 395868 -19142 395941 -19086
rect 395997 -19142 396083 -19086
rect 396139 -19142 396208 -19086
rect 395868 -19228 396208 -19142
rect 395868 -19284 395941 -19228
rect 395997 -19284 396083 -19228
rect 396139 -19284 396208 -19228
rect 395868 -19370 396208 -19284
rect 395868 -19426 395941 -19370
rect 395997 -19426 396083 -19370
rect 396139 -19426 396208 -19370
rect 395868 -19512 396208 -19426
rect 395868 -19568 395941 -19512
rect 395997 -19568 396083 -19512
rect 396139 -19568 396208 -19512
rect 395868 -19654 396208 -19568
rect 395868 -19710 395941 -19654
rect 395997 -19710 396083 -19654
rect 396139 -19710 396208 -19654
rect 395868 -19796 396208 -19710
rect 395868 -19852 395941 -19796
rect 395997 -19852 396083 -19796
rect 396139 -19852 396208 -19796
rect 395868 -19938 396208 -19852
rect 395868 -19994 395941 -19938
rect 395997 -19994 396083 -19938
rect 396139 -19994 396208 -19938
rect 395868 -20080 396208 -19994
rect 395868 -20136 395941 -20080
rect 395997 -20136 396083 -20080
rect 396139 -20136 396208 -20080
rect 395868 -20222 396208 -20136
rect 395868 -20278 395941 -20222
rect 395997 -20278 396083 -20222
rect 396139 -20278 396208 -20222
rect 395868 -20364 396208 -20278
rect 395868 -20420 395941 -20364
rect 395997 -20420 396083 -20364
rect 396139 -20420 396208 -20364
rect 395868 -20506 396208 -20420
rect 395868 -20562 395941 -20506
rect 395997 -20562 396083 -20506
rect 396139 -20562 396208 -20506
rect 395868 -20648 396208 -20562
rect 395868 -20704 395941 -20648
rect 395997 -20704 396083 -20648
rect 396139 -20704 396208 -20648
rect 395868 -20790 396208 -20704
rect 395868 -20846 395941 -20790
rect 395997 -20846 396083 -20790
rect 396139 -20846 396208 -20790
rect 395868 -20932 396208 -20846
rect 395868 -20988 395941 -20932
rect 395997 -20988 396083 -20932
rect 396139 -20988 396208 -20932
rect 395868 -21074 396208 -20988
rect 395868 -21130 395941 -21074
rect 395997 -21130 396083 -21074
rect 396139 -21130 396208 -21074
rect 395868 -21216 396208 -21130
rect 395868 -21272 395941 -21216
rect 395997 -21272 396083 -21216
rect 396139 -21272 396208 -21216
rect 395868 -21358 396208 -21272
rect 395868 -21414 395941 -21358
rect 395997 -21414 396083 -21358
rect 396139 -21414 396208 -21358
rect 395868 -21500 396208 -21414
rect 395868 -21556 395941 -21500
rect 395997 -21556 396083 -21500
rect 396139 -21556 396208 -21500
rect 395868 -21642 396208 -21556
rect 395868 -21698 395941 -21642
rect 395997 -21698 396083 -21642
rect 396139 -21698 396208 -21642
rect 395868 -21784 396208 -21698
rect 395868 -21840 395941 -21784
rect 395997 -21840 396083 -21784
rect 396139 -21840 396208 -21784
rect 395868 -21926 396208 -21840
rect 395868 -21982 395941 -21926
rect 395997 -21982 396083 -21926
rect 396139 -21982 396208 -21926
rect 395868 -22068 396208 -21982
rect 395868 -22124 395941 -22068
rect 395997 -22124 396083 -22068
rect 396139 -22124 396208 -22068
rect 395868 -22210 396208 -22124
rect 395868 -22266 395941 -22210
rect 395997 -22266 396083 -22210
rect 396139 -22266 396208 -22210
rect 395868 -22352 396208 -22266
rect 395868 -22408 395941 -22352
rect 395997 -22408 396083 -22352
rect 396139 -22408 396208 -22352
rect 395868 -22494 396208 -22408
rect 395868 -22550 395941 -22494
rect 395997 -22550 396083 -22494
rect 396139 -22550 396208 -22494
rect 395868 -22636 396208 -22550
rect 395868 -22692 395941 -22636
rect 395997 -22692 396083 -22636
rect 396139 -22692 396208 -22636
rect 395868 -22778 396208 -22692
rect 395868 -22834 395941 -22778
rect 395997 -22834 396083 -22778
rect 396139 -22834 396208 -22778
rect 395868 -22920 396208 -22834
rect 395868 -22976 395941 -22920
rect 395997 -22976 396083 -22920
rect 396139 -22976 396208 -22920
rect 395868 -23062 396208 -22976
rect 395868 -23118 395941 -23062
rect 395997 -23118 396083 -23062
rect 396139 -23118 396208 -23062
rect 395868 -23204 396208 -23118
rect 395868 -23260 395941 -23204
rect 395997 -23260 396083 -23204
rect 396139 -23260 396208 -23204
rect 395868 -23346 396208 -23260
rect 395868 -23402 395941 -23346
rect 395997 -23402 396083 -23346
rect 396139 -23402 396208 -23346
rect 395868 -23488 396208 -23402
rect 395868 -23544 395941 -23488
rect 395997 -23544 396083 -23488
rect 396139 -23544 396208 -23488
rect 395868 -23630 396208 -23544
rect 395868 -23686 395941 -23630
rect 395997 -23686 396083 -23630
rect 396139 -23686 396208 -23630
rect 395868 -23772 396208 -23686
rect 395868 -23828 395941 -23772
rect 395997 -23828 396083 -23772
rect 396139 -23828 396208 -23772
rect 395868 -23914 396208 -23828
rect 395868 -23970 395941 -23914
rect 395997 -23970 396083 -23914
rect 396139 -23970 396208 -23914
rect 395868 -24056 396208 -23970
rect 395868 -24112 395941 -24056
rect 395997 -24112 396083 -24056
rect 396139 -24112 396208 -24056
rect 395868 -24198 396208 -24112
rect 395868 -24254 395941 -24198
rect 395997 -24254 396083 -24198
rect 396139 -24254 396208 -24198
rect 395868 -24340 396208 -24254
rect 395868 -24396 395941 -24340
rect 395997 -24396 396083 -24340
rect 396139 -24396 396208 -24340
rect 395868 -24482 396208 -24396
rect 395868 -24538 395941 -24482
rect 395997 -24538 396083 -24482
rect 396139 -24538 396208 -24482
rect 395868 -24624 396208 -24538
rect 395868 -24680 395941 -24624
rect 395997 -24680 396083 -24624
rect 396139 -24680 396208 -24624
rect 395868 -24766 396208 -24680
rect 395868 -24822 395941 -24766
rect 395997 -24822 396083 -24766
rect 396139 -24822 396208 -24766
rect 395868 -24908 396208 -24822
rect 395868 -24964 395941 -24908
rect 395997 -24964 396083 -24908
rect 396139 -24964 396208 -24908
rect 395868 -25050 396208 -24964
rect 395868 -25106 395941 -25050
rect 395997 -25106 396083 -25050
rect 396139 -25106 396208 -25050
rect 395868 -25192 396208 -25106
rect 395868 -25248 395941 -25192
rect 395997 -25248 396083 -25192
rect 396139 -25248 396208 -25192
rect 395868 -25334 396208 -25248
rect 395868 -25390 395941 -25334
rect 395997 -25390 396083 -25334
rect 396139 -25390 396208 -25334
rect 395868 -25476 396208 -25390
rect 395868 -25532 395941 -25476
rect 395997 -25532 396083 -25476
rect 396139 -25532 396208 -25476
rect 395868 -25600 396208 -25532
rect 396400 -17858 397200 -17740
rect 396400 -17914 396526 -17858
rect 396582 -17914 396650 -17858
rect 396706 -17914 396774 -17858
rect 396830 -17914 396898 -17858
rect 396954 -17914 397022 -17858
rect 397078 -17914 397200 -17858
rect 396400 -17982 397200 -17914
rect 396400 -18038 396526 -17982
rect 396582 -18038 396650 -17982
rect 396706 -18038 396774 -17982
rect 396830 -18038 396898 -17982
rect 396954 -18038 397022 -17982
rect 397078 -18038 397200 -17982
rect 396400 -18106 397200 -18038
rect 396400 -18162 396526 -18106
rect 396582 -18162 396650 -18106
rect 396706 -18162 396774 -18106
rect 396830 -18162 396898 -18106
rect 396954 -18162 397022 -18106
rect 397078 -18162 397200 -18106
rect 396400 -18230 397200 -18162
rect 396400 -18286 396526 -18230
rect 396582 -18286 396650 -18230
rect 396706 -18286 396774 -18230
rect 396830 -18286 396898 -18230
rect 396954 -18286 397022 -18230
rect 397078 -18286 397200 -18230
rect 396400 -18354 397200 -18286
rect 396400 -18410 396526 -18354
rect 396582 -18410 396650 -18354
rect 396706 -18410 396774 -18354
rect 396830 -18410 396898 -18354
rect 396954 -18410 397022 -18354
rect 397078 -18410 397200 -18354
rect 396400 -18478 397200 -18410
rect 396400 -18534 396526 -18478
rect 396582 -18534 396650 -18478
rect 396706 -18534 396774 -18478
rect 396830 -18534 396898 -18478
rect 396954 -18534 397022 -18478
rect 397078 -18534 397200 -18478
rect 396400 -18602 397200 -18534
rect 396400 -18658 396526 -18602
rect 396582 -18658 396650 -18602
rect 396706 -18658 396774 -18602
rect 396830 -18658 396898 -18602
rect 396954 -18658 397022 -18602
rect 397078 -18658 397200 -18602
rect 396400 -18726 397200 -18658
rect 396400 -18782 396526 -18726
rect 396582 -18782 396650 -18726
rect 396706 -18782 396774 -18726
rect 396830 -18782 396898 -18726
rect 396954 -18782 397022 -18726
rect 397078 -18782 397200 -18726
rect 396400 -18850 397200 -18782
rect 396400 -18906 396526 -18850
rect 396582 -18906 396650 -18850
rect 396706 -18906 396774 -18850
rect 396830 -18906 396898 -18850
rect 396954 -18906 397022 -18850
rect 397078 -18906 397200 -18850
rect 396400 -18974 397200 -18906
rect 396400 -19030 396526 -18974
rect 396582 -19030 396650 -18974
rect 396706 -19030 396774 -18974
rect 396830 -19030 396898 -18974
rect 396954 -19030 397022 -18974
rect 397078 -19030 397200 -18974
rect 396400 -19098 397200 -19030
rect 396400 -19154 396526 -19098
rect 396582 -19154 396650 -19098
rect 396706 -19154 396774 -19098
rect 396830 -19154 396898 -19098
rect 396954 -19154 397022 -19098
rect 397078 -19154 397200 -19098
rect 396400 -19222 397200 -19154
rect 396400 -19278 396526 -19222
rect 396582 -19278 396650 -19222
rect 396706 -19278 396774 -19222
rect 396830 -19278 396898 -19222
rect 396954 -19278 397022 -19222
rect 397078 -19278 397200 -19222
rect 396400 -19346 397200 -19278
rect 396400 -19402 396526 -19346
rect 396582 -19402 396650 -19346
rect 396706 -19402 396774 -19346
rect 396830 -19402 396898 -19346
rect 396954 -19402 397022 -19346
rect 397078 -19402 397200 -19346
rect 396400 -19470 397200 -19402
rect 396400 -19526 396526 -19470
rect 396582 -19526 396650 -19470
rect 396706 -19526 396774 -19470
rect 396830 -19526 396898 -19470
rect 396954 -19526 397022 -19470
rect 397078 -19526 397200 -19470
rect 396400 -19594 397200 -19526
rect 396400 -19650 396526 -19594
rect 396582 -19650 396650 -19594
rect 396706 -19650 396774 -19594
rect 396830 -19650 396898 -19594
rect 396954 -19650 397022 -19594
rect 397078 -19650 397200 -19594
rect 396400 -19718 397200 -19650
rect 396400 -19774 396526 -19718
rect 396582 -19774 396650 -19718
rect 396706 -19774 396774 -19718
rect 396830 -19774 396898 -19718
rect 396954 -19774 397022 -19718
rect 397078 -19774 397200 -19718
rect 396400 -19842 397200 -19774
rect 396400 -19898 396526 -19842
rect 396582 -19898 396650 -19842
rect 396706 -19898 396774 -19842
rect 396830 -19898 396898 -19842
rect 396954 -19898 397022 -19842
rect 397078 -19898 397200 -19842
rect 396400 -19966 397200 -19898
rect 396400 -20022 396526 -19966
rect 396582 -20022 396650 -19966
rect 396706 -20022 396774 -19966
rect 396830 -20022 396898 -19966
rect 396954 -20022 397022 -19966
rect 397078 -20022 397200 -19966
rect 396400 -20090 397200 -20022
rect 396400 -20146 396526 -20090
rect 396582 -20146 396650 -20090
rect 396706 -20146 396774 -20090
rect 396830 -20146 396898 -20090
rect 396954 -20146 397022 -20090
rect 397078 -20146 397200 -20090
rect 396400 -20214 397200 -20146
rect 396400 -20270 396526 -20214
rect 396582 -20270 396650 -20214
rect 396706 -20270 396774 -20214
rect 396830 -20270 396898 -20214
rect 396954 -20270 397022 -20214
rect 397078 -20270 397200 -20214
rect 396400 -20338 397200 -20270
rect 396400 -20394 396526 -20338
rect 396582 -20394 396650 -20338
rect 396706 -20394 396774 -20338
rect 396830 -20394 396898 -20338
rect 396954 -20394 397022 -20338
rect 397078 -20394 397200 -20338
rect 396400 -20462 397200 -20394
rect 396400 -20518 396526 -20462
rect 396582 -20518 396650 -20462
rect 396706 -20518 396774 -20462
rect 396830 -20518 396898 -20462
rect 396954 -20518 397022 -20462
rect 397078 -20518 397200 -20462
rect 396400 -20586 397200 -20518
rect 396400 -20642 396526 -20586
rect 396582 -20642 396650 -20586
rect 396706 -20642 396774 -20586
rect 396830 -20642 396898 -20586
rect 396954 -20642 397022 -20586
rect 397078 -20642 397200 -20586
rect 396400 -20710 397200 -20642
rect 396400 -20766 396526 -20710
rect 396582 -20766 396650 -20710
rect 396706 -20766 396774 -20710
rect 396830 -20766 396898 -20710
rect 396954 -20766 397022 -20710
rect 397078 -20766 397200 -20710
rect 396400 -20834 397200 -20766
rect 396400 -20890 396526 -20834
rect 396582 -20890 396650 -20834
rect 396706 -20890 396774 -20834
rect 396830 -20890 396898 -20834
rect 396954 -20890 397022 -20834
rect 397078 -20890 397200 -20834
rect 396400 -20958 397200 -20890
rect 396400 -21014 396526 -20958
rect 396582 -21014 396650 -20958
rect 396706 -21014 396774 -20958
rect 396830 -21014 396898 -20958
rect 396954 -21014 397022 -20958
rect 397078 -21014 397200 -20958
rect 396400 -21082 397200 -21014
rect 396400 -21138 396526 -21082
rect 396582 -21138 396650 -21082
rect 396706 -21138 396774 -21082
rect 396830 -21138 396898 -21082
rect 396954 -21138 397022 -21082
rect 397078 -21138 397200 -21082
rect 396400 -21206 397200 -21138
rect 396400 -21262 396526 -21206
rect 396582 -21262 396650 -21206
rect 396706 -21262 396774 -21206
rect 396830 -21262 396898 -21206
rect 396954 -21262 397022 -21206
rect 397078 -21262 397200 -21206
rect 396400 -21330 397200 -21262
rect 396400 -21386 396526 -21330
rect 396582 -21386 396650 -21330
rect 396706 -21386 396774 -21330
rect 396830 -21386 396898 -21330
rect 396954 -21386 397022 -21330
rect 397078 -21386 397200 -21330
rect 396400 -21454 397200 -21386
rect 396400 -21510 396526 -21454
rect 396582 -21510 396650 -21454
rect 396706 -21510 396774 -21454
rect 396830 -21510 396898 -21454
rect 396954 -21510 397022 -21454
rect 397078 -21510 397200 -21454
rect 396400 -21578 397200 -21510
rect 396400 -21634 396526 -21578
rect 396582 -21634 396650 -21578
rect 396706 -21634 396774 -21578
rect 396830 -21634 396898 -21578
rect 396954 -21634 397022 -21578
rect 397078 -21634 397200 -21578
rect 396400 -21702 397200 -21634
rect 396400 -21758 396526 -21702
rect 396582 -21758 396650 -21702
rect 396706 -21758 396774 -21702
rect 396830 -21758 396898 -21702
rect 396954 -21758 397022 -21702
rect 397078 -21758 397200 -21702
rect 396400 -21826 397200 -21758
rect 396400 -21882 396526 -21826
rect 396582 -21882 396650 -21826
rect 396706 -21882 396774 -21826
rect 396830 -21882 396898 -21826
rect 396954 -21882 397022 -21826
rect 397078 -21882 397200 -21826
rect 396400 -21950 397200 -21882
rect 396400 -22006 396526 -21950
rect 396582 -22006 396650 -21950
rect 396706 -22006 396774 -21950
rect 396830 -22006 396898 -21950
rect 396954 -22006 397022 -21950
rect 397078 -22006 397200 -21950
rect 396400 -22074 397200 -22006
rect 396400 -22130 396526 -22074
rect 396582 -22130 396650 -22074
rect 396706 -22130 396774 -22074
rect 396830 -22130 396898 -22074
rect 396954 -22130 397022 -22074
rect 397078 -22130 397200 -22074
rect 396400 -22198 397200 -22130
rect 396400 -22254 396526 -22198
rect 396582 -22254 396650 -22198
rect 396706 -22254 396774 -22198
rect 396830 -22254 396898 -22198
rect 396954 -22254 397022 -22198
rect 397078 -22254 397200 -22198
rect 396400 -22322 397200 -22254
rect 396400 -22378 396526 -22322
rect 396582 -22378 396650 -22322
rect 396706 -22378 396774 -22322
rect 396830 -22378 396898 -22322
rect 396954 -22378 397022 -22322
rect 397078 -22378 397200 -22322
rect 396400 -22446 397200 -22378
rect 396400 -22502 396526 -22446
rect 396582 -22502 396650 -22446
rect 396706 -22502 396774 -22446
rect 396830 -22502 396898 -22446
rect 396954 -22502 397022 -22446
rect 397078 -22502 397200 -22446
rect 396400 -22570 397200 -22502
rect 396400 -22626 396526 -22570
rect 396582 -22626 396650 -22570
rect 396706 -22626 396774 -22570
rect 396830 -22626 396898 -22570
rect 396954 -22626 397022 -22570
rect 397078 -22626 397200 -22570
rect 396400 -22694 397200 -22626
rect 396400 -22750 396526 -22694
rect 396582 -22750 396650 -22694
rect 396706 -22750 396774 -22694
rect 396830 -22750 396898 -22694
rect 396954 -22750 397022 -22694
rect 397078 -22750 397200 -22694
rect 396400 -22818 397200 -22750
rect 396400 -22874 396526 -22818
rect 396582 -22874 396650 -22818
rect 396706 -22874 396774 -22818
rect 396830 -22874 396898 -22818
rect 396954 -22874 397022 -22818
rect 397078 -22874 397200 -22818
rect 396400 -22942 397200 -22874
rect 396400 -22998 396526 -22942
rect 396582 -22998 396650 -22942
rect 396706 -22998 396774 -22942
rect 396830 -22998 396898 -22942
rect 396954 -22998 397022 -22942
rect 397078 -22998 397200 -22942
rect 396400 -23066 397200 -22998
rect 396400 -23122 396526 -23066
rect 396582 -23122 396650 -23066
rect 396706 -23122 396774 -23066
rect 396830 -23122 396898 -23066
rect 396954 -23122 397022 -23066
rect 397078 -23122 397200 -23066
rect 396400 -23190 397200 -23122
rect 396400 -23246 396526 -23190
rect 396582 -23246 396650 -23190
rect 396706 -23246 396774 -23190
rect 396830 -23246 396898 -23190
rect 396954 -23246 397022 -23190
rect 397078 -23246 397200 -23190
rect 396400 -23314 397200 -23246
rect 396400 -23370 396526 -23314
rect 396582 -23370 396650 -23314
rect 396706 -23370 396774 -23314
rect 396830 -23370 396898 -23314
rect 396954 -23370 397022 -23314
rect 397078 -23370 397200 -23314
rect 396400 -23438 397200 -23370
rect 396400 -23494 396526 -23438
rect 396582 -23494 396650 -23438
rect 396706 -23494 396774 -23438
rect 396830 -23494 396898 -23438
rect 396954 -23494 397022 -23438
rect 397078 -23494 397200 -23438
rect 396400 -23562 397200 -23494
rect 396400 -23618 396526 -23562
rect 396582 -23618 396650 -23562
rect 396706 -23618 396774 -23562
rect 396830 -23618 396898 -23562
rect 396954 -23618 397022 -23562
rect 397078 -23618 397200 -23562
rect 396400 -23686 397200 -23618
rect 396400 -23742 396526 -23686
rect 396582 -23742 396650 -23686
rect 396706 -23742 396774 -23686
rect 396830 -23742 396898 -23686
rect 396954 -23742 397022 -23686
rect 397078 -23742 397200 -23686
rect 396400 -23810 397200 -23742
rect 396400 -23866 396526 -23810
rect 396582 -23866 396650 -23810
rect 396706 -23866 396774 -23810
rect 396830 -23866 396898 -23810
rect 396954 -23866 397022 -23810
rect 397078 -23866 397200 -23810
rect 396400 -23934 397200 -23866
rect 396400 -23990 396526 -23934
rect 396582 -23990 396650 -23934
rect 396706 -23990 396774 -23934
rect 396830 -23990 396898 -23934
rect 396954 -23990 397022 -23934
rect 397078 -23990 397200 -23934
rect 396400 -24058 397200 -23990
rect 396400 -24114 396526 -24058
rect 396582 -24114 396650 -24058
rect 396706 -24114 396774 -24058
rect 396830 -24114 396898 -24058
rect 396954 -24114 397022 -24058
rect 397078 -24114 397200 -24058
rect 396400 -24182 397200 -24114
rect 396400 -24238 396526 -24182
rect 396582 -24238 396650 -24182
rect 396706 -24238 396774 -24182
rect 396830 -24238 396898 -24182
rect 396954 -24238 397022 -24182
rect 397078 -24238 397200 -24182
rect 396400 -24306 397200 -24238
rect 396400 -24362 396526 -24306
rect 396582 -24362 396650 -24306
rect 396706 -24362 396774 -24306
rect 396830 -24362 396898 -24306
rect 396954 -24362 397022 -24306
rect 397078 -24362 397200 -24306
rect 396400 -24430 397200 -24362
rect 396400 -24486 396526 -24430
rect 396582 -24486 396650 -24430
rect 396706 -24486 396774 -24430
rect 396830 -24486 396898 -24430
rect 396954 -24486 397022 -24430
rect 397078 -24486 397200 -24430
rect 396400 -24554 397200 -24486
rect 396400 -24610 396526 -24554
rect 396582 -24610 396650 -24554
rect 396706 -24610 396774 -24554
rect 396830 -24610 396898 -24554
rect 396954 -24610 397022 -24554
rect 397078 -24610 397200 -24554
rect 396400 -24678 397200 -24610
rect 396400 -24734 396526 -24678
rect 396582 -24734 396650 -24678
rect 396706 -24734 396774 -24678
rect 396830 -24734 396898 -24678
rect 396954 -24734 397022 -24678
rect 397078 -24734 397200 -24678
rect 396400 -24802 397200 -24734
rect 396400 -24858 396526 -24802
rect 396582 -24858 396650 -24802
rect 396706 -24858 396774 -24802
rect 396830 -24858 396898 -24802
rect 396954 -24858 397022 -24802
rect 397078 -24858 397200 -24802
rect 396400 -24926 397200 -24858
rect 396400 -24982 396526 -24926
rect 396582 -24982 396650 -24926
rect 396706 -24982 396774 -24926
rect 396830 -24982 396898 -24926
rect 396954 -24982 397022 -24926
rect 397078 -24982 397200 -24926
rect 396400 -25050 397200 -24982
rect 396400 -25106 396526 -25050
rect 396582 -25106 396650 -25050
rect 396706 -25106 396774 -25050
rect 396830 -25106 396898 -25050
rect 396954 -25106 397022 -25050
rect 397078 -25106 397200 -25050
rect 396400 -25174 397200 -25106
rect 396400 -25230 396526 -25174
rect 396582 -25230 396650 -25174
rect 396706 -25230 396774 -25174
rect 396830 -25230 396898 -25174
rect 396954 -25230 397022 -25174
rect 397078 -25230 397200 -25174
rect 396400 -25298 397200 -25230
rect 396400 -25354 396526 -25298
rect 396582 -25354 396650 -25298
rect 396706 -25354 396774 -25298
rect 396830 -25354 396898 -25298
rect 396954 -25354 397022 -25298
rect 397078 -25354 397200 -25298
rect 396400 -25422 397200 -25354
rect 396400 -25478 396526 -25422
rect 396582 -25478 396650 -25422
rect 396706 -25478 396774 -25422
rect 396830 -25478 396898 -25422
rect 396954 -25478 397022 -25422
rect 397078 -25478 397200 -25422
rect 396400 -25600 397200 -25478
rect 388000 -25721 397200 -25600
rect 388000 -25777 388146 -25721
rect 388202 -25777 388270 -25721
rect 388326 -25777 388394 -25721
rect 388450 -25777 388518 -25721
rect 388574 -25777 388642 -25721
rect 388698 -25777 388766 -25721
rect 388822 -25777 388890 -25721
rect 388946 -25777 389014 -25721
rect 389070 -25777 389138 -25721
rect 389194 -25777 389262 -25721
rect 389318 -25777 389386 -25721
rect 389442 -25777 389510 -25721
rect 389566 -25777 389634 -25721
rect 389690 -25777 389758 -25721
rect 389814 -25777 389882 -25721
rect 389938 -25777 390006 -25721
rect 390062 -25777 390130 -25721
rect 390186 -25777 390254 -25721
rect 390310 -25777 390378 -25721
rect 390434 -25777 390502 -25721
rect 390558 -25777 390626 -25721
rect 390682 -25777 390750 -25721
rect 390806 -25777 390874 -25721
rect 390930 -25777 390998 -25721
rect 391054 -25777 391122 -25721
rect 391178 -25777 391246 -25721
rect 391302 -25777 391370 -25721
rect 391426 -25777 391494 -25721
rect 391550 -25777 391618 -25721
rect 391674 -25777 391742 -25721
rect 391798 -25777 391866 -25721
rect 391922 -25777 391990 -25721
rect 392046 -25777 392114 -25721
rect 392170 -25777 392238 -25721
rect 392294 -25777 392362 -25721
rect 392418 -25777 392486 -25721
rect 392542 -25777 392610 -25721
rect 392666 -25777 392734 -25721
rect 392790 -25777 392858 -25721
rect 392914 -25777 392982 -25721
rect 393038 -25777 393106 -25721
rect 393162 -25777 393230 -25721
rect 393286 -25777 393354 -25721
rect 393410 -25777 393478 -25721
rect 393534 -25777 393602 -25721
rect 393658 -25777 393726 -25721
rect 393782 -25777 393850 -25721
rect 393906 -25777 393974 -25721
rect 394030 -25777 394098 -25721
rect 394154 -25777 394222 -25721
rect 394278 -25777 394346 -25721
rect 394402 -25777 394470 -25721
rect 394526 -25777 394594 -25721
rect 394650 -25777 394718 -25721
rect 394774 -25777 394842 -25721
rect 394898 -25777 394966 -25721
rect 395022 -25777 395090 -25721
rect 395146 -25777 395214 -25721
rect 395270 -25777 395338 -25721
rect 395394 -25777 395462 -25721
rect 395518 -25777 395586 -25721
rect 395642 -25777 395710 -25721
rect 395766 -25777 395898 -25721
rect 395954 -25777 396022 -25721
rect 396078 -25777 396146 -25721
rect 396202 -25777 396270 -25721
rect 396326 -25777 396394 -25721
rect 396450 -25777 396518 -25721
rect 396574 -25777 396642 -25721
rect 396698 -25777 396766 -25721
rect 396822 -25777 396890 -25721
rect 396946 -25777 397014 -25721
rect 397070 -25777 397200 -25721
rect 388000 -25845 397200 -25777
rect 388000 -25901 388146 -25845
rect 388202 -25901 388270 -25845
rect 388326 -25901 388394 -25845
rect 388450 -25901 388518 -25845
rect 388574 -25901 388642 -25845
rect 388698 -25901 388766 -25845
rect 388822 -25901 388890 -25845
rect 388946 -25901 389014 -25845
rect 389070 -25901 389138 -25845
rect 389194 -25901 389262 -25845
rect 389318 -25901 389386 -25845
rect 389442 -25901 389510 -25845
rect 389566 -25901 389634 -25845
rect 389690 -25901 389758 -25845
rect 389814 -25901 389882 -25845
rect 389938 -25901 390006 -25845
rect 390062 -25901 390130 -25845
rect 390186 -25901 390254 -25845
rect 390310 -25901 390378 -25845
rect 390434 -25901 390502 -25845
rect 390558 -25901 390626 -25845
rect 390682 -25901 390750 -25845
rect 390806 -25901 390874 -25845
rect 390930 -25901 390998 -25845
rect 391054 -25901 391122 -25845
rect 391178 -25901 391246 -25845
rect 391302 -25901 391370 -25845
rect 391426 -25901 391494 -25845
rect 391550 -25901 391618 -25845
rect 391674 -25901 391742 -25845
rect 391798 -25901 391866 -25845
rect 391922 -25901 391990 -25845
rect 392046 -25901 392114 -25845
rect 392170 -25901 392238 -25845
rect 392294 -25901 392362 -25845
rect 392418 -25901 392486 -25845
rect 392542 -25901 392610 -25845
rect 392666 -25901 392734 -25845
rect 392790 -25901 392858 -25845
rect 392914 -25901 392982 -25845
rect 393038 -25901 393106 -25845
rect 393162 -25901 393230 -25845
rect 393286 -25901 393354 -25845
rect 393410 -25901 393478 -25845
rect 393534 -25901 393602 -25845
rect 393658 -25901 393726 -25845
rect 393782 -25901 393850 -25845
rect 393906 -25901 393974 -25845
rect 394030 -25901 394098 -25845
rect 394154 -25901 394222 -25845
rect 394278 -25901 394346 -25845
rect 394402 -25901 394470 -25845
rect 394526 -25901 394594 -25845
rect 394650 -25901 394718 -25845
rect 394774 -25901 394842 -25845
rect 394898 -25901 394966 -25845
rect 395022 -25901 395090 -25845
rect 395146 -25901 395214 -25845
rect 395270 -25901 395338 -25845
rect 395394 -25901 395462 -25845
rect 395518 -25901 395586 -25845
rect 395642 -25901 395710 -25845
rect 395766 -25901 395898 -25845
rect 395954 -25901 396022 -25845
rect 396078 -25901 396146 -25845
rect 396202 -25901 396270 -25845
rect 396326 -25901 396394 -25845
rect 396450 -25901 396518 -25845
rect 396574 -25901 396642 -25845
rect 396698 -25901 396766 -25845
rect 396822 -25901 396890 -25845
rect 396946 -25901 397014 -25845
rect 397070 -25901 397200 -25845
rect 388000 -25969 397200 -25901
rect 388000 -26025 388146 -25969
rect 388202 -26025 388270 -25969
rect 388326 -26025 388394 -25969
rect 388450 -26025 388518 -25969
rect 388574 -26025 388642 -25969
rect 388698 -26025 388766 -25969
rect 388822 -26025 388890 -25969
rect 388946 -26025 389014 -25969
rect 389070 -26025 389138 -25969
rect 389194 -26025 389262 -25969
rect 389318 -26025 389386 -25969
rect 389442 -26025 389510 -25969
rect 389566 -26025 389634 -25969
rect 389690 -26025 389758 -25969
rect 389814 -26025 389882 -25969
rect 389938 -26025 390006 -25969
rect 390062 -26025 390130 -25969
rect 390186 -26025 390254 -25969
rect 390310 -26025 390378 -25969
rect 390434 -26025 390502 -25969
rect 390558 -26025 390626 -25969
rect 390682 -26025 390750 -25969
rect 390806 -26025 390874 -25969
rect 390930 -26025 390998 -25969
rect 391054 -26025 391122 -25969
rect 391178 -26025 391246 -25969
rect 391302 -26025 391370 -25969
rect 391426 -26025 391494 -25969
rect 391550 -26025 391618 -25969
rect 391674 -26025 391742 -25969
rect 391798 -26025 391866 -25969
rect 391922 -26025 391990 -25969
rect 392046 -26025 392114 -25969
rect 392170 -26025 392238 -25969
rect 392294 -26025 392362 -25969
rect 392418 -26025 392486 -25969
rect 392542 -26025 392610 -25969
rect 392666 -26025 392734 -25969
rect 392790 -26025 392858 -25969
rect 392914 -26025 392982 -25969
rect 393038 -26025 393106 -25969
rect 393162 -26025 393230 -25969
rect 393286 -26025 393354 -25969
rect 393410 -26025 393478 -25969
rect 393534 -26025 393602 -25969
rect 393658 -26025 393726 -25969
rect 393782 -26025 393850 -25969
rect 393906 -26025 393974 -25969
rect 394030 -26025 394098 -25969
rect 394154 -26025 394222 -25969
rect 394278 -26025 394346 -25969
rect 394402 -26025 394470 -25969
rect 394526 -26025 394594 -25969
rect 394650 -26025 394718 -25969
rect 394774 -26025 394842 -25969
rect 394898 -26025 394966 -25969
rect 395022 -26025 395090 -25969
rect 395146 -26025 395214 -25969
rect 395270 -26025 395338 -25969
rect 395394 -26025 395462 -25969
rect 395518 -26025 395586 -25969
rect 395642 -26025 395710 -25969
rect 395766 -26025 395898 -25969
rect 395954 -26025 396022 -25969
rect 396078 -26025 396146 -25969
rect 396202 -26025 396270 -25969
rect 396326 -26025 396394 -25969
rect 396450 -26025 396518 -25969
rect 396574 -26025 396642 -25969
rect 396698 -26025 396766 -25969
rect 396822 -26025 396890 -25969
rect 396946 -26025 397014 -25969
rect 397070 -26025 397200 -25969
rect 388000 -26093 397200 -26025
rect 388000 -26149 388146 -26093
rect 388202 -26149 388270 -26093
rect 388326 -26149 388394 -26093
rect 388450 -26149 388518 -26093
rect 388574 -26149 388642 -26093
rect 388698 -26149 388766 -26093
rect 388822 -26149 388890 -26093
rect 388946 -26149 389014 -26093
rect 389070 -26149 389138 -26093
rect 389194 -26149 389262 -26093
rect 389318 -26149 389386 -26093
rect 389442 -26149 389510 -26093
rect 389566 -26149 389634 -26093
rect 389690 -26149 389758 -26093
rect 389814 -26149 389882 -26093
rect 389938 -26149 390006 -26093
rect 390062 -26149 390130 -26093
rect 390186 -26149 390254 -26093
rect 390310 -26149 390378 -26093
rect 390434 -26149 390502 -26093
rect 390558 -26149 390626 -26093
rect 390682 -26149 390750 -26093
rect 390806 -26149 390874 -26093
rect 390930 -26149 390998 -26093
rect 391054 -26149 391122 -26093
rect 391178 -26149 391246 -26093
rect 391302 -26149 391370 -26093
rect 391426 -26149 391494 -26093
rect 391550 -26149 391618 -26093
rect 391674 -26149 391742 -26093
rect 391798 -26149 391866 -26093
rect 391922 -26149 391990 -26093
rect 392046 -26149 392114 -26093
rect 392170 -26149 392238 -26093
rect 392294 -26149 392362 -26093
rect 392418 -26149 392486 -26093
rect 392542 -26149 392610 -26093
rect 392666 -26149 392734 -26093
rect 392790 -26149 392858 -26093
rect 392914 -26149 392982 -26093
rect 393038 -26149 393106 -26093
rect 393162 -26149 393230 -26093
rect 393286 -26149 393354 -26093
rect 393410 -26149 393478 -26093
rect 393534 -26149 393602 -26093
rect 393658 -26149 393726 -26093
rect 393782 -26149 393850 -26093
rect 393906 -26149 393974 -26093
rect 394030 -26149 394098 -26093
rect 394154 -26149 394222 -26093
rect 394278 -26149 394346 -26093
rect 394402 -26149 394470 -26093
rect 394526 -26149 394594 -26093
rect 394650 -26149 394718 -26093
rect 394774 -26149 394842 -26093
rect 394898 -26149 394966 -26093
rect 395022 -26149 395090 -26093
rect 395146 -26149 395214 -26093
rect 395270 -26149 395338 -26093
rect 395394 -26149 395462 -26093
rect 395518 -26149 395586 -26093
rect 395642 -26149 395710 -26093
rect 395766 -26149 395898 -26093
rect 395954 -26149 396022 -26093
rect 396078 -26149 396146 -26093
rect 396202 -26149 396270 -26093
rect 396326 -26149 396394 -26093
rect 396450 -26149 396518 -26093
rect 396574 -26149 396642 -26093
rect 396698 -26149 396766 -26093
rect 396822 -26149 396890 -26093
rect 396946 -26149 397014 -26093
rect 397070 -26149 397200 -26093
rect 388000 -26270 397200 -26149
<< via2 >>
rect 388146 -17247 388202 -17191
rect 388270 -17247 388326 -17191
rect 388394 -17247 388450 -17191
rect 388518 -17247 388574 -17191
rect 388642 -17247 388698 -17191
rect 388766 -17247 388822 -17191
rect 388890 -17247 388946 -17191
rect 389014 -17247 389070 -17191
rect 389138 -17247 389194 -17191
rect 389262 -17247 389318 -17191
rect 389386 -17247 389442 -17191
rect 389510 -17247 389566 -17191
rect 389634 -17247 389690 -17191
rect 389758 -17247 389814 -17191
rect 389882 -17247 389938 -17191
rect 390006 -17247 390062 -17191
rect 390130 -17247 390186 -17191
rect 390254 -17247 390310 -17191
rect 390378 -17247 390434 -17191
rect 390502 -17247 390558 -17191
rect 390626 -17247 390682 -17191
rect 390750 -17247 390806 -17191
rect 390874 -17247 390930 -17191
rect 390998 -17247 391054 -17191
rect 391122 -17247 391178 -17191
rect 391246 -17247 391302 -17191
rect 391370 -17247 391426 -17191
rect 391494 -17247 391550 -17191
rect 391618 -17247 391674 -17191
rect 391742 -17247 391798 -17191
rect 391866 -17247 391922 -17191
rect 391990 -17247 392046 -17191
rect 392114 -17247 392170 -17191
rect 392238 -17247 392294 -17191
rect 392362 -17247 392418 -17191
rect 392486 -17247 392542 -17191
rect 392610 -17247 392666 -17191
rect 392734 -17247 392790 -17191
rect 392858 -17247 392914 -17191
rect 392982 -17247 393038 -17191
rect 393106 -17247 393162 -17191
rect 393230 -17247 393286 -17191
rect 393354 -17247 393410 -17191
rect 393478 -17247 393534 -17191
rect 393602 -17247 393658 -17191
rect 393726 -17247 393782 -17191
rect 393850 -17247 393906 -17191
rect 393974 -17247 394030 -17191
rect 394098 -17247 394154 -17191
rect 394222 -17247 394278 -17191
rect 394346 -17247 394402 -17191
rect 394470 -17247 394526 -17191
rect 394594 -17247 394650 -17191
rect 394718 -17247 394774 -17191
rect 394842 -17247 394898 -17191
rect 394966 -17247 395022 -17191
rect 395090 -17247 395146 -17191
rect 395214 -17247 395270 -17191
rect 395338 -17247 395394 -17191
rect 395462 -17247 395518 -17191
rect 395586 -17247 395642 -17191
rect 395710 -17247 395766 -17191
rect 395898 -17247 395954 -17191
rect 396022 -17247 396078 -17191
rect 396146 -17247 396202 -17191
rect 396270 -17247 396326 -17191
rect 396394 -17247 396450 -17191
rect 396518 -17247 396574 -17191
rect 396642 -17247 396698 -17191
rect 396766 -17247 396822 -17191
rect 396890 -17247 396946 -17191
rect 397014 -17247 397070 -17191
rect 388146 -17371 388202 -17315
rect 388270 -17371 388326 -17315
rect 388394 -17371 388450 -17315
rect 388518 -17371 388574 -17315
rect 388642 -17371 388698 -17315
rect 388766 -17371 388822 -17315
rect 388890 -17371 388946 -17315
rect 389014 -17371 389070 -17315
rect 389138 -17371 389194 -17315
rect 389262 -17371 389318 -17315
rect 389386 -17371 389442 -17315
rect 389510 -17371 389566 -17315
rect 389634 -17371 389690 -17315
rect 389758 -17371 389814 -17315
rect 389882 -17371 389938 -17315
rect 390006 -17371 390062 -17315
rect 390130 -17371 390186 -17315
rect 390254 -17371 390310 -17315
rect 390378 -17371 390434 -17315
rect 390502 -17371 390558 -17315
rect 390626 -17371 390682 -17315
rect 390750 -17371 390806 -17315
rect 390874 -17371 390930 -17315
rect 390998 -17371 391054 -17315
rect 391122 -17371 391178 -17315
rect 391246 -17371 391302 -17315
rect 391370 -17371 391426 -17315
rect 391494 -17371 391550 -17315
rect 391618 -17371 391674 -17315
rect 391742 -17371 391798 -17315
rect 391866 -17371 391922 -17315
rect 391990 -17371 392046 -17315
rect 392114 -17371 392170 -17315
rect 392238 -17371 392294 -17315
rect 392362 -17371 392418 -17315
rect 392486 -17371 392542 -17315
rect 392610 -17371 392666 -17315
rect 392734 -17371 392790 -17315
rect 392858 -17371 392914 -17315
rect 392982 -17371 393038 -17315
rect 393106 -17371 393162 -17315
rect 393230 -17371 393286 -17315
rect 393354 -17371 393410 -17315
rect 393478 -17371 393534 -17315
rect 393602 -17371 393658 -17315
rect 393726 -17371 393782 -17315
rect 393850 -17371 393906 -17315
rect 393974 -17371 394030 -17315
rect 394098 -17371 394154 -17315
rect 394222 -17371 394278 -17315
rect 394346 -17371 394402 -17315
rect 394470 -17371 394526 -17315
rect 394594 -17371 394650 -17315
rect 394718 -17371 394774 -17315
rect 394842 -17371 394898 -17315
rect 394966 -17371 395022 -17315
rect 395090 -17371 395146 -17315
rect 395214 -17371 395270 -17315
rect 395338 -17371 395394 -17315
rect 395462 -17371 395518 -17315
rect 395586 -17371 395642 -17315
rect 395710 -17371 395766 -17315
rect 395898 -17371 395954 -17315
rect 396022 -17371 396078 -17315
rect 396146 -17371 396202 -17315
rect 396270 -17371 396326 -17315
rect 396394 -17371 396450 -17315
rect 396518 -17371 396574 -17315
rect 396642 -17371 396698 -17315
rect 396766 -17371 396822 -17315
rect 396890 -17371 396946 -17315
rect 397014 -17371 397070 -17315
rect 388146 -17495 388202 -17439
rect 388270 -17495 388326 -17439
rect 388394 -17495 388450 -17439
rect 388518 -17495 388574 -17439
rect 388642 -17495 388698 -17439
rect 388766 -17495 388822 -17439
rect 388890 -17495 388946 -17439
rect 389014 -17495 389070 -17439
rect 389138 -17495 389194 -17439
rect 389262 -17495 389318 -17439
rect 389386 -17495 389442 -17439
rect 389510 -17495 389566 -17439
rect 389634 -17495 389690 -17439
rect 389758 -17495 389814 -17439
rect 389882 -17495 389938 -17439
rect 390006 -17495 390062 -17439
rect 390130 -17495 390186 -17439
rect 390254 -17495 390310 -17439
rect 390378 -17495 390434 -17439
rect 390502 -17495 390558 -17439
rect 390626 -17495 390682 -17439
rect 390750 -17495 390806 -17439
rect 390874 -17495 390930 -17439
rect 390998 -17495 391054 -17439
rect 391122 -17495 391178 -17439
rect 391246 -17495 391302 -17439
rect 391370 -17495 391426 -17439
rect 391494 -17495 391550 -17439
rect 391618 -17495 391674 -17439
rect 391742 -17495 391798 -17439
rect 391866 -17495 391922 -17439
rect 391990 -17495 392046 -17439
rect 392114 -17495 392170 -17439
rect 392238 -17495 392294 -17439
rect 392362 -17495 392418 -17439
rect 392486 -17495 392542 -17439
rect 392610 -17495 392666 -17439
rect 392734 -17495 392790 -17439
rect 392858 -17495 392914 -17439
rect 392982 -17495 393038 -17439
rect 393106 -17495 393162 -17439
rect 393230 -17495 393286 -17439
rect 393354 -17495 393410 -17439
rect 393478 -17495 393534 -17439
rect 393602 -17495 393658 -17439
rect 393726 -17495 393782 -17439
rect 393850 -17495 393906 -17439
rect 393974 -17495 394030 -17439
rect 394098 -17495 394154 -17439
rect 394222 -17495 394278 -17439
rect 394346 -17495 394402 -17439
rect 394470 -17495 394526 -17439
rect 394594 -17495 394650 -17439
rect 394718 -17495 394774 -17439
rect 394842 -17495 394898 -17439
rect 394966 -17495 395022 -17439
rect 395090 -17495 395146 -17439
rect 395214 -17495 395270 -17439
rect 395338 -17495 395394 -17439
rect 395462 -17495 395518 -17439
rect 395586 -17495 395642 -17439
rect 395710 -17495 395766 -17439
rect 395898 -17495 395954 -17439
rect 396022 -17495 396078 -17439
rect 396146 -17495 396202 -17439
rect 396270 -17495 396326 -17439
rect 396394 -17495 396450 -17439
rect 396518 -17495 396574 -17439
rect 396642 -17495 396698 -17439
rect 396766 -17495 396822 -17439
rect 396890 -17495 396946 -17439
rect 397014 -17495 397070 -17439
rect 388146 -17619 388202 -17563
rect 388270 -17619 388326 -17563
rect 388394 -17619 388450 -17563
rect 388518 -17619 388574 -17563
rect 388642 -17619 388698 -17563
rect 388766 -17619 388822 -17563
rect 388890 -17619 388946 -17563
rect 389014 -17619 389070 -17563
rect 389138 -17619 389194 -17563
rect 389262 -17619 389318 -17563
rect 389386 -17619 389442 -17563
rect 389510 -17619 389566 -17563
rect 389634 -17619 389690 -17563
rect 389758 -17619 389814 -17563
rect 389882 -17619 389938 -17563
rect 390006 -17619 390062 -17563
rect 390130 -17619 390186 -17563
rect 390254 -17619 390310 -17563
rect 390378 -17619 390434 -17563
rect 390502 -17619 390558 -17563
rect 390626 -17619 390682 -17563
rect 390750 -17619 390806 -17563
rect 390874 -17619 390930 -17563
rect 390998 -17619 391054 -17563
rect 391122 -17619 391178 -17563
rect 391246 -17619 391302 -17563
rect 391370 -17619 391426 -17563
rect 391494 -17619 391550 -17563
rect 391618 -17619 391674 -17563
rect 391742 -17619 391798 -17563
rect 391866 -17619 391922 -17563
rect 391990 -17619 392046 -17563
rect 392114 -17619 392170 -17563
rect 392238 -17619 392294 -17563
rect 392362 -17619 392418 -17563
rect 392486 -17619 392542 -17563
rect 392610 -17619 392666 -17563
rect 392734 -17619 392790 -17563
rect 392858 -17619 392914 -17563
rect 392982 -17619 393038 -17563
rect 393106 -17619 393162 -17563
rect 393230 -17619 393286 -17563
rect 393354 -17619 393410 -17563
rect 393478 -17619 393534 -17563
rect 393602 -17619 393658 -17563
rect 393726 -17619 393782 -17563
rect 393850 -17619 393906 -17563
rect 393974 -17619 394030 -17563
rect 394098 -17619 394154 -17563
rect 394222 -17619 394278 -17563
rect 394346 -17619 394402 -17563
rect 394470 -17619 394526 -17563
rect 394594 -17619 394650 -17563
rect 394718 -17619 394774 -17563
rect 394842 -17619 394898 -17563
rect 394966 -17619 395022 -17563
rect 395090 -17619 395146 -17563
rect 395214 -17619 395270 -17563
rect 395338 -17619 395394 -17563
rect 395462 -17619 395518 -17563
rect 395586 -17619 395642 -17563
rect 395710 -17619 395766 -17563
rect 395898 -17619 395954 -17563
rect 396022 -17619 396078 -17563
rect 396146 -17619 396202 -17563
rect 396270 -17619 396326 -17563
rect 396394 -17619 396450 -17563
rect 396518 -17619 396574 -17563
rect 396642 -17619 396698 -17563
rect 396766 -17619 396822 -17563
rect 396890 -17619 396946 -17563
rect 397014 -17619 397070 -17563
rect 388114 -17914 388170 -17858
rect 388238 -17914 388294 -17858
rect 388362 -17914 388418 -17858
rect 388486 -17914 388542 -17858
rect 388610 -17914 388666 -17858
rect 388114 -18038 388170 -17982
rect 388238 -18038 388294 -17982
rect 388362 -18038 388418 -17982
rect 388486 -18038 388542 -17982
rect 388610 -18038 388666 -17982
rect 388114 -18162 388170 -18106
rect 388238 -18162 388294 -18106
rect 388362 -18162 388418 -18106
rect 388486 -18162 388542 -18106
rect 388610 -18162 388666 -18106
rect 388114 -18286 388170 -18230
rect 388238 -18286 388294 -18230
rect 388362 -18286 388418 -18230
rect 388486 -18286 388542 -18230
rect 388610 -18286 388666 -18230
rect 388114 -18410 388170 -18354
rect 388238 -18410 388294 -18354
rect 388362 -18410 388418 -18354
rect 388486 -18410 388542 -18354
rect 388610 -18410 388666 -18354
rect 388114 -18534 388170 -18478
rect 388238 -18534 388294 -18478
rect 388362 -18534 388418 -18478
rect 388486 -18534 388542 -18478
rect 388610 -18534 388666 -18478
rect 388114 -18658 388170 -18602
rect 388238 -18658 388294 -18602
rect 388362 -18658 388418 -18602
rect 388486 -18658 388542 -18602
rect 388610 -18658 388666 -18602
rect 388114 -18782 388170 -18726
rect 388238 -18782 388294 -18726
rect 388362 -18782 388418 -18726
rect 388486 -18782 388542 -18726
rect 388610 -18782 388666 -18726
rect 388114 -18906 388170 -18850
rect 388238 -18906 388294 -18850
rect 388362 -18906 388418 -18850
rect 388486 -18906 388542 -18850
rect 388610 -18906 388666 -18850
rect 388114 -19030 388170 -18974
rect 388238 -19030 388294 -18974
rect 388362 -19030 388418 -18974
rect 388486 -19030 388542 -18974
rect 388610 -19030 388666 -18974
rect 388114 -19154 388170 -19098
rect 388238 -19154 388294 -19098
rect 388362 -19154 388418 -19098
rect 388486 -19154 388542 -19098
rect 388610 -19154 388666 -19098
rect 388114 -19278 388170 -19222
rect 388238 -19278 388294 -19222
rect 388362 -19278 388418 -19222
rect 388486 -19278 388542 -19222
rect 388610 -19278 388666 -19222
rect 388114 -19402 388170 -19346
rect 388238 -19402 388294 -19346
rect 388362 -19402 388418 -19346
rect 388486 -19402 388542 -19346
rect 388610 -19402 388666 -19346
rect 388114 -19526 388170 -19470
rect 388238 -19526 388294 -19470
rect 388362 -19526 388418 -19470
rect 388486 -19526 388542 -19470
rect 388610 -19526 388666 -19470
rect 388114 -19650 388170 -19594
rect 388238 -19650 388294 -19594
rect 388362 -19650 388418 -19594
rect 388486 -19650 388542 -19594
rect 388610 -19650 388666 -19594
rect 388114 -19774 388170 -19718
rect 388238 -19774 388294 -19718
rect 388362 -19774 388418 -19718
rect 388486 -19774 388542 -19718
rect 388610 -19774 388666 -19718
rect 388114 -19898 388170 -19842
rect 388238 -19898 388294 -19842
rect 388362 -19898 388418 -19842
rect 388486 -19898 388542 -19842
rect 388610 -19898 388666 -19842
rect 388114 -20022 388170 -19966
rect 388238 -20022 388294 -19966
rect 388362 -20022 388418 -19966
rect 388486 -20022 388542 -19966
rect 388610 -20022 388666 -19966
rect 388114 -20146 388170 -20090
rect 388238 -20146 388294 -20090
rect 388362 -20146 388418 -20090
rect 388486 -20146 388542 -20090
rect 388610 -20146 388666 -20090
rect 388114 -20270 388170 -20214
rect 388238 -20270 388294 -20214
rect 388362 -20270 388418 -20214
rect 388486 -20270 388542 -20214
rect 388610 -20270 388666 -20214
rect 388114 -20394 388170 -20338
rect 388238 -20394 388294 -20338
rect 388362 -20394 388418 -20338
rect 388486 -20394 388542 -20338
rect 388610 -20394 388666 -20338
rect 388114 -20518 388170 -20462
rect 388238 -20518 388294 -20462
rect 388362 -20518 388418 -20462
rect 388486 -20518 388542 -20462
rect 388610 -20518 388666 -20462
rect 388114 -20642 388170 -20586
rect 388238 -20642 388294 -20586
rect 388362 -20642 388418 -20586
rect 388486 -20642 388542 -20586
rect 388610 -20642 388666 -20586
rect 388114 -20766 388170 -20710
rect 388238 -20766 388294 -20710
rect 388362 -20766 388418 -20710
rect 388486 -20766 388542 -20710
rect 388610 -20766 388666 -20710
rect 388114 -20890 388170 -20834
rect 388238 -20890 388294 -20834
rect 388362 -20890 388418 -20834
rect 388486 -20890 388542 -20834
rect 388610 -20890 388666 -20834
rect 388114 -21014 388170 -20958
rect 388238 -21014 388294 -20958
rect 388362 -21014 388418 -20958
rect 388486 -21014 388542 -20958
rect 388610 -21014 388666 -20958
rect 388114 -21138 388170 -21082
rect 388238 -21138 388294 -21082
rect 388362 -21138 388418 -21082
rect 388486 -21138 388542 -21082
rect 388610 -21138 388666 -21082
rect 388114 -21262 388170 -21206
rect 388238 -21262 388294 -21206
rect 388362 -21262 388418 -21206
rect 388486 -21262 388542 -21206
rect 388610 -21262 388666 -21206
rect 388114 -21386 388170 -21330
rect 388238 -21386 388294 -21330
rect 388362 -21386 388418 -21330
rect 388486 -21386 388542 -21330
rect 388610 -21386 388666 -21330
rect 388114 -21510 388170 -21454
rect 388238 -21510 388294 -21454
rect 388362 -21510 388418 -21454
rect 388486 -21510 388542 -21454
rect 388610 -21510 388666 -21454
rect 388114 -21634 388170 -21578
rect 388238 -21634 388294 -21578
rect 388362 -21634 388418 -21578
rect 388486 -21634 388542 -21578
rect 388610 -21634 388666 -21578
rect 388114 -21758 388170 -21702
rect 388238 -21758 388294 -21702
rect 388362 -21758 388418 -21702
rect 388486 -21758 388542 -21702
rect 388610 -21758 388666 -21702
rect 388114 -21882 388170 -21826
rect 388238 -21882 388294 -21826
rect 388362 -21882 388418 -21826
rect 388486 -21882 388542 -21826
rect 388610 -21882 388666 -21826
rect 388114 -22006 388170 -21950
rect 388238 -22006 388294 -21950
rect 388362 -22006 388418 -21950
rect 388486 -22006 388542 -21950
rect 388610 -22006 388666 -21950
rect 388114 -22130 388170 -22074
rect 388238 -22130 388294 -22074
rect 388362 -22130 388418 -22074
rect 388486 -22130 388542 -22074
rect 388610 -22130 388666 -22074
rect 388114 -22254 388170 -22198
rect 388238 -22254 388294 -22198
rect 388362 -22254 388418 -22198
rect 388486 -22254 388542 -22198
rect 388610 -22254 388666 -22198
rect 388114 -22378 388170 -22322
rect 388238 -22378 388294 -22322
rect 388362 -22378 388418 -22322
rect 388486 -22378 388542 -22322
rect 388610 -22378 388666 -22322
rect 388114 -22502 388170 -22446
rect 388238 -22502 388294 -22446
rect 388362 -22502 388418 -22446
rect 388486 -22502 388542 -22446
rect 388610 -22502 388666 -22446
rect 388114 -22626 388170 -22570
rect 388238 -22626 388294 -22570
rect 388362 -22626 388418 -22570
rect 388486 -22626 388542 -22570
rect 388610 -22626 388666 -22570
rect 388114 -22750 388170 -22694
rect 388238 -22750 388294 -22694
rect 388362 -22750 388418 -22694
rect 388486 -22750 388542 -22694
rect 388610 -22750 388666 -22694
rect 388114 -22874 388170 -22818
rect 388238 -22874 388294 -22818
rect 388362 -22874 388418 -22818
rect 388486 -22874 388542 -22818
rect 388610 -22874 388666 -22818
rect 388114 -22998 388170 -22942
rect 388238 -22998 388294 -22942
rect 388362 -22998 388418 -22942
rect 388486 -22998 388542 -22942
rect 388610 -22998 388666 -22942
rect 388114 -23122 388170 -23066
rect 388238 -23122 388294 -23066
rect 388362 -23122 388418 -23066
rect 388486 -23122 388542 -23066
rect 388610 -23122 388666 -23066
rect 388114 -23246 388170 -23190
rect 388238 -23246 388294 -23190
rect 388362 -23246 388418 -23190
rect 388486 -23246 388542 -23190
rect 388610 -23246 388666 -23190
rect 388114 -23370 388170 -23314
rect 388238 -23370 388294 -23314
rect 388362 -23370 388418 -23314
rect 388486 -23370 388542 -23314
rect 388610 -23370 388666 -23314
rect 388114 -23494 388170 -23438
rect 388238 -23494 388294 -23438
rect 388362 -23494 388418 -23438
rect 388486 -23494 388542 -23438
rect 388610 -23494 388666 -23438
rect 388114 -23618 388170 -23562
rect 388238 -23618 388294 -23562
rect 388362 -23618 388418 -23562
rect 388486 -23618 388542 -23562
rect 388610 -23618 388666 -23562
rect 388114 -23742 388170 -23686
rect 388238 -23742 388294 -23686
rect 388362 -23742 388418 -23686
rect 388486 -23742 388542 -23686
rect 388610 -23742 388666 -23686
rect 388114 -23866 388170 -23810
rect 388238 -23866 388294 -23810
rect 388362 -23866 388418 -23810
rect 388486 -23866 388542 -23810
rect 388610 -23866 388666 -23810
rect 388114 -23990 388170 -23934
rect 388238 -23990 388294 -23934
rect 388362 -23990 388418 -23934
rect 388486 -23990 388542 -23934
rect 388610 -23990 388666 -23934
rect 388114 -24114 388170 -24058
rect 388238 -24114 388294 -24058
rect 388362 -24114 388418 -24058
rect 388486 -24114 388542 -24058
rect 388610 -24114 388666 -24058
rect 388114 -24238 388170 -24182
rect 388238 -24238 388294 -24182
rect 388362 -24238 388418 -24182
rect 388486 -24238 388542 -24182
rect 388610 -24238 388666 -24182
rect 388114 -24362 388170 -24306
rect 388238 -24362 388294 -24306
rect 388362 -24362 388418 -24306
rect 388486 -24362 388542 -24306
rect 388610 -24362 388666 -24306
rect 388114 -24486 388170 -24430
rect 388238 -24486 388294 -24430
rect 388362 -24486 388418 -24430
rect 388486 -24486 388542 -24430
rect 388610 -24486 388666 -24430
rect 388114 -24610 388170 -24554
rect 388238 -24610 388294 -24554
rect 388362 -24610 388418 -24554
rect 388486 -24610 388542 -24554
rect 388610 -24610 388666 -24554
rect 388114 -24734 388170 -24678
rect 388238 -24734 388294 -24678
rect 388362 -24734 388418 -24678
rect 388486 -24734 388542 -24678
rect 388610 -24734 388666 -24678
rect 388114 -24858 388170 -24802
rect 388238 -24858 388294 -24802
rect 388362 -24858 388418 -24802
rect 388486 -24858 388542 -24802
rect 388610 -24858 388666 -24802
rect 388114 -24982 388170 -24926
rect 388238 -24982 388294 -24926
rect 388362 -24982 388418 -24926
rect 388486 -24982 388542 -24926
rect 388610 -24982 388666 -24926
rect 388114 -25106 388170 -25050
rect 388238 -25106 388294 -25050
rect 388362 -25106 388418 -25050
rect 388486 -25106 388542 -25050
rect 388610 -25106 388666 -25050
rect 388114 -25230 388170 -25174
rect 388238 -25230 388294 -25174
rect 388362 -25230 388418 -25174
rect 388486 -25230 388542 -25174
rect 388610 -25230 388666 -25174
rect 388114 -25354 388170 -25298
rect 388238 -25354 388294 -25298
rect 388362 -25354 388418 -25298
rect 388486 -25354 388542 -25298
rect 388610 -25354 388666 -25298
rect 388114 -25478 388170 -25422
rect 388238 -25478 388294 -25422
rect 388362 -25478 388418 -25422
rect 388486 -25478 388542 -25422
rect 388610 -25478 388666 -25422
rect 389141 -18006 389197 -17950
rect 389283 -18006 389339 -17950
rect 389141 -18148 389197 -18092
rect 389283 -18148 389339 -18092
rect 389141 -18290 389197 -18234
rect 389283 -18290 389339 -18234
rect 389141 -18432 389197 -18376
rect 389283 -18432 389339 -18376
rect 389141 -18574 389197 -18518
rect 389283 -18574 389339 -18518
rect 389141 -18716 389197 -18660
rect 389283 -18716 389339 -18660
rect 389141 -18858 389197 -18802
rect 389283 -18858 389339 -18802
rect 389141 -19000 389197 -18944
rect 389283 -19000 389339 -18944
rect 389141 -19142 389197 -19086
rect 389283 -19142 389339 -19086
rect 389141 -19284 389197 -19228
rect 389283 -19284 389339 -19228
rect 389141 -19426 389197 -19370
rect 389283 -19426 389339 -19370
rect 389141 -19568 389197 -19512
rect 389283 -19568 389339 -19512
rect 389141 -19710 389197 -19654
rect 389283 -19710 389339 -19654
rect 389141 -19852 389197 -19796
rect 389283 -19852 389339 -19796
rect 389141 -19994 389197 -19938
rect 389283 -19994 389339 -19938
rect 389141 -20136 389197 -20080
rect 389283 -20136 389339 -20080
rect 389141 -20278 389197 -20222
rect 389283 -20278 389339 -20222
rect 389141 -20420 389197 -20364
rect 389283 -20420 389339 -20364
rect 389141 -20562 389197 -20506
rect 389283 -20562 389339 -20506
rect 389141 -20704 389197 -20648
rect 389283 -20704 389339 -20648
rect 389141 -20846 389197 -20790
rect 389283 -20846 389339 -20790
rect 389141 -20988 389197 -20932
rect 389283 -20988 389339 -20932
rect 389141 -21130 389197 -21074
rect 389283 -21130 389339 -21074
rect 389141 -21272 389197 -21216
rect 389283 -21272 389339 -21216
rect 389141 -21414 389197 -21358
rect 389283 -21414 389339 -21358
rect 389141 -21556 389197 -21500
rect 389283 -21556 389339 -21500
rect 389141 -21698 389197 -21642
rect 389283 -21698 389339 -21642
rect 389141 -21840 389197 -21784
rect 389283 -21840 389339 -21784
rect 389141 -21982 389197 -21926
rect 389283 -21982 389339 -21926
rect 389141 -22124 389197 -22068
rect 389283 -22124 389339 -22068
rect 389141 -22266 389197 -22210
rect 389283 -22266 389339 -22210
rect 389141 -22408 389197 -22352
rect 389283 -22408 389339 -22352
rect 389141 -22550 389197 -22494
rect 389283 -22550 389339 -22494
rect 389141 -22692 389197 -22636
rect 389283 -22692 389339 -22636
rect 389141 -22834 389197 -22778
rect 389283 -22834 389339 -22778
rect 389141 -22976 389197 -22920
rect 389283 -22976 389339 -22920
rect 389141 -23118 389197 -23062
rect 389283 -23118 389339 -23062
rect 389141 -23260 389197 -23204
rect 389283 -23260 389339 -23204
rect 389141 -23402 389197 -23346
rect 389283 -23402 389339 -23346
rect 389141 -23544 389197 -23488
rect 389283 -23544 389339 -23488
rect 389141 -23686 389197 -23630
rect 389283 -23686 389339 -23630
rect 389141 -23828 389197 -23772
rect 389283 -23828 389339 -23772
rect 389141 -23970 389197 -23914
rect 389283 -23970 389339 -23914
rect 389141 -24112 389197 -24056
rect 389283 -24112 389339 -24056
rect 389141 -24254 389197 -24198
rect 389283 -24254 389339 -24198
rect 389141 -24396 389197 -24340
rect 389283 -24396 389339 -24340
rect 389141 -24538 389197 -24482
rect 389283 -24538 389339 -24482
rect 389141 -24680 389197 -24624
rect 389283 -24680 389339 -24624
rect 389141 -24822 389197 -24766
rect 389283 -24822 389339 -24766
rect 389141 -24964 389197 -24908
rect 389283 -24964 389339 -24908
rect 389141 -25106 389197 -25050
rect 389283 -25106 389339 -25050
rect 389141 -25248 389197 -25192
rect 389283 -25248 389339 -25192
rect 389141 -25390 389197 -25334
rect 389283 -25390 389339 -25334
rect 389141 -25532 389197 -25476
rect 389283 -25532 389339 -25476
rect 389542 -18006 389598 -17950
rect 389684 -18006 389740 -17950
rect 389542 -18148 389598 -18092
rect 389684 -18148 389740 -18092
rect 389542 -18290 389598 -18234
rect 389684 -18290 389740 -18234
rect 389542 -18432 389598 -18376
rect 389684 -18432 389740 -18376
rect 389542 -18574 389598 -18518
rect 389684 -18574 389740 -18518
rect 389542 -18716 389598 -18660
rect 389684 -18716 389740 -18660
rect 389542 -18858 389598 -18802
rect 389684 -18858 389740 -18802
rect 389542 -19000 389598 -18944
rect 389684 -19000 389740 -18944
rect 389542 -19142 389598 -19086
rect 389684 -19142 389740 -19086
rect 389542 -19284 389598 -19228
rect 389684 -19284 389740 -19228
rect 389542 -19426 389598 -19370
rect 389684 -19426 389740 -19370
rect 389542 -19568 389598 -19512
rect 389684 -19568 389740 -19512
rect 389542 -19710 389598 -19654
rect 389684 -19710 389740 -19654
rect 389542 -19852 389598 -19796
rect 389684 -19852 389740 -19796
rect 389542 -19994 389598 -19938
rect 389684 -19994 389740 -19938
rect 389542 -20136 389598 -20080
rect 389684 -20136 389740 -20080
rect 389542 -20278 389598 -20222
rect 389684 -20278 389740 -20222
rect 389542 -20420 389598 -20364
rect 389684 -20420 389740 -20364
rect 389542 -20562 389598 -20506
rect 389684 -20562 389740 -20506
rect 389542 -20704 389598 -20648
rect 389684 -20704 389740 -20648
rect 389542 -20846 389598 -20790
rect 389684 -20846 389740 -20790
rect 389542 -20988 389598 -20932
rect 389684 -20988 389740 -20932
rect 389542 -21130 389598 -21074
rect 389684 -21130 389740 -21074
rect 389542 -21272 389598 -21216
rect 389684 -21272 389740 -21216
rect 389542 -21414 389598 -21358
rect 389684 -21414 389740 -21358
rect 389542 -21556 389598 -21500
rect 389684 -21556 389740 -21500
rect 389542 -21698 389598 -21642
rect 389684 -21698 389740 -21642
rect 389542 -21840 389598 -21784
rect 389684 -21840 389740 -21784
rect 389542 -21982 389598 -21926
rect 389684 -21982 389740 -21926
rect 389542 -22124 389598 -22068
rect 389684 -22124 389740 -22068
rect 389542 -22266 389598 -22210
rect 389684 -22266 389740 -22210
rect 389542 -22408 389598 -22352
rect 389684 -22408 389740 -22352
rect 389542 -22550 389598 -22494
rect 389684 -22550 389740 -22494
rect 389542 -22692 389598 -22636
rect 389684 -22692 389740 -22636
rect 389542 -22834 389598 -22778
rect 389684 -22834 389740 -22778
rect 389542 -22976 389598 -22920
rect 389684 -22976 389740 -22920
rect 389542 -23118 389598 -23062
rect 389684 -23118 389740 -23062
rect 389542 -23260 389598 -23204
rect 389684 -23260 389740 -23204
rect 389542 -23402 389598 -23346
rect 389684 -23402 389740 -23346
rect 389542 -23544 389598 -23488
rect 389684 -23544 389740 -23488
rect 389542 -23686 389598 -23630
rect 389684 -23686 389740 -23630
rect 389542 -23828 389598 -23772
rect 389684 -23828 389740 -23772
rect 389542 -23970 389598 -23914
rect 389684 -23970 389740 -23914
rect 389542 -24112 389598 -24056
rect 389684 -24112 389740 -24056
rect 389542 -24254 389598 -24198
rect 389684 -24254 389740 -24198
rect 389542 -24396 389598 -24340
rect 389684 -24396 389740 -24340
rect 389542 -24538 389598 -24482
rect 389684 -24538 389740 -24482
rect 389542 -24680 389598 -24624
rect 389684 -24680 389740 -24624
rect 389542 -24822 389598 -24766
rect 389684 -24822 389740 -24766
rect 389542 -24964 389598 -24908
rect 389684 -24964 389740 -24908
rect 389542 -25106 389598 -25050
rect 389684 -25106 389740 -25050
rect 389542 -25248 389598 -25192
rect 389684 -25248 389740 -25192
rect 389542 -25390 389598 -25334
rect 389684 -25390 389740 -25334
rect 389542 -25532 389598 -25476
rect 389684 -25532 389740 -25476
rect 389942 -18006 389998 -17950
rect 390084 -18006 390140 -17950
rect 389942 -18148 389998 -18092
rect 390084 -18148 390140 -18092
rect 389942 -18290 389998 -18234
rect 390084 -18290 390140 -18234
rect 389942 -18432 389998 -18376
rect 390084 -18432 390140 -18376
rect 389942 -18574 389998 -18518
rect 390084 -18574 390140 -18518
rect 389942 -18716 389998 -18660
rect 390084 -18716 390140 -18660
rect 389942 -18858 389998 -18802
rect 390084 -18858 390140 -18802
rect 389942 -19000 389998 -18944
rect 390084 -19000 390140 -18944
rect 389942 -19142 389998 -19086
rect 390084 -19142 390140 -19086
rect 389942 -19284 389998 -19228
rect 390084 -19284 390140 -19228
rect 389942 -19426 389998 -19370
rect 390084 -19426 390140 -19370
rect 389942 -19568 389998 -19512
rect 390084 -19568 390140 -19512
rect 389942 -19710 389998 -19654
rect 390084 -19710 390140 -19654
rect 389942 -19852 389998 -19796
rect 390084 -19852 390140 -19796
rect 389942 -19994 389998 -19938
rect 390084 -19994 390140 -19938
rect 389942 -20136 389998 -20080
rect 390084 -20136 390140 -20080
rect 389942 -20278 389998 -20222
rect 390084 -20278 390140 -20222
rect 389942 -20420 389998 -20364
rect 390084 -20420 390140 -20364
rect 389942 -20562 389998 -20506
rect 390084 -20562 390140 -20506
rect 389942 -20704 389998 -20648
rect 390084 -20704 390140 -20648
rect 389942 -20846 389998 -20790
rect 390084 -20846 390140 -20790
rect 389942 -20988 389998 -20932
rect 390084 -20988 390140 -20932
rect 389942 -21130 389998 -21074
rect 390084 -21130 390140 -21074
rect 389942 -21272 389998 -21216
rect 390084 -21272 390140 -21216
rect 389942 -21414 389998 -21358
rect 390084 -21414 390140 -21358
rect 389942 -21556 389998 -21500
rect 390084 -21556 390140 -21500
rect 389942 -21698 389998 -21642
rect 390084 -21698 390140 -21642
rect 389942 -21840 389998 -21784
rect 390084 -21840 390140 -21784
rect 389942 -21982 389998 -21926
rect 390084 -21982 390140 -21926
rect 389942 -22124 389998 -22068
rect 390084 -22124 390140 -22068
rect 389942 -22266 389998 -22210
rect 390084 -22266 390140 -22210
rect 389942 -22408 389998 -22352
rect 390084 -22408 390140 -22352
rect 389942 -22550 389998 -22494
rect 390084 -22550 390140 -22494
rect 389942 -22692 389998 -22636
rect 390084 -22692 390140 -22636
rect 389942 -22834 389998 -22778
rect 390084 -22834 390140 -22778
rect 389942 -22976 389998 -22920
rect 390084 -22976 390140 -22920
rect 389942 -23118 389998 -23062
rect 390084 -23118 390140 -23062
rect 389942 -23260 389998 -23204
rect 390084 -23260 390140 -23204
rect 389942 -23402 389998 -23346
rect 390084 -23402 390140 -23346
rect 389942 -23544 389998 -23488
rect 390084 -23544 390140 -23488
rect 389942 -23686 389998 -23630
rect 390084 -23686 390140 -23630
rect 389942 -23828 389998 -23772
rect 390084 -23828 390140 -23772
rect 389942 -23970 389998 -23914
rect 390084 -23970 390140 -23914
rect 389942 -24112 389998 -24056
rect 390084 -24112 390140 -24056
rect 389942 -24254 389998 -24198
rect 390084 -24254 390140 -24198
rect 389942 -24396 389998 -24340
rect 390084 -24396 390140 -24340
rect 389942 -24538 389998 -24482
rect 390084 -24538 390140 -24482
rect 389942 -24680 389998 -24624
rect 390084 -24680 390140 -24624
rect 389942 -24822 389998 -24766
rect 390084 -24822 390140 -24766
rect 389942 -24964 389998 -24908
rect 390084 -24964 390140 -24908
rect 389942 -25106 389998 -25050
rect 390084 -25106 390140 -25050
rect 389942 -25248 389998 -25192
rect 390084 -25248 390140 -25192
rect 389942 -25390 389998 -25334
rect 390084 -25390 390140 -25334
rect 389942 -25532 389998 -25476
rect 390084 -25532 390140 -25476
rect 390339 -18006 390395 -17950
rect 390481 -18006 390537 -17950
rect 390339 -18148 390395 -18092
rect 390481 -18148 390537 -18092
rect 390339 -18290 390395 -18234
rect 390481 -18290 390537 -18234
rect 390339 -18432 390395 -18376
rect 390481 -18432 390537 -18376
rect 390339 -18574 390395 -18518
rect 390481 -18574 390537 -18518
rect 390339 -18716 390395 -18660
rect 390481 -18716 390537 -18660
rect 390339 -18858 390395 -18802
rect 390481 -18858 390537 -18802
rect 390339 -19000 390395 -18944
rect 390481 -19000 390537 -18944
rect 390339 -19142 390395 -19086
rect 390481 -19142 390537 -19086
rect 390339 -19284 390395 -19228
rect 390481 -19284 390537 -19228
rect 390339 -19426 390395 -19370
rect 390481 -19426 390537 -19370
rect 390339 -19568 390395 -19512
rect 390481 -19568 390537 -19512
rect 390339 -19710 390395 -19654
rect 390481 -19710 390537 -19654
rect 390339 -19852 390395 -19796
rect 390481 -19852 390537 -19796
rect 390339 -19994 390395 -19938
rect 390481 -19994 390537 -19938
rect 390339 -20136 390395 -20080
rect 390481 -20136 390537 -20080
rect 390339 -20278 390395 -20222
rect 390481 -20278 390537 -20222
rect 390339 -20420 390395 -20364
rect 390481 -20420 390537 -20364
rect 390339 -20562 390395 -20506
rect 390481 -20562 390537 -20506
rect 390339 -20704 390395 -20648
rect 390481 -20704 390537 -20648
rect 390339 -20846 390395 -20790
rect 390481 -20846 390537 -20790
rect 390339 -20988 390395 -20932
rect 390481 -20988 390537 -20932
rect 390339 -21130 390395 -21074
rect 390481 -21130 390537 -21074
rect 390339 -21272 390395 -21216
rect 390481 -21272 390537 -21216
rect 390339 -21414 390395 -21358
rect 390481 -21414 390537 -21358
rect 390339 -21556 390395 -21500
rect 390481 -21556 390537 -21500
rect 390339 -21698 390395 -21642
rect 390481 -21698 390537 -21642
rect 390339 -21840 390395 -21784
rect 390481 -21840 390537 -21784
rect 390339 -21982 390395 -21926
rect 390481 -21982 390537 -21926
rect 390339 -22124 390395 -22068
rect 390481 -22124 390537 -22068
rect 390339 -22266 390395 -22210
rect 390481 -22266 390537 -22210
rect 390339 -22408 390395 -22352
rect 390481 -22408 390537 -22352
rect 390339 -22550 390395 -22494
rect 390481 -22550 390537 -22494
rect 390339 -22692 390395 -22636
rect 390481 -22692 390537 -22636
rect 390339 -22834 390395 -22778
rect 390481 -22834 390537 -22778
rect 390339 -22976 390395 -22920
rect 390481 -22976 390537 -22920
rect 390339 -23118 390395 -23062
rect 390481 -23118 390537 -23062
rect 390339 -23260 390395 -23204
rect 390481 -23260 390537 -23204
rect 390339 -23402 390395 -23346
rect 390481 -23402 390537 -23346
rect 390339 -23544 390395 -23488
rect 390481 -23544 390537 -23488
rect 390339 -23686 390395 -23630
rect 390481 -23686 390537 -23630
rect 390339 -23828 390395 -23772
rect 390481 -23828 390537 -23772
rect 390339 -23970 390395 -23914
rect 390481 -23970 390537 -23914
rect 390339 -24112 390395 -24056
rect 390481 -24112 390537 -24056
rect 390339 -24254 390395 -24198
rect 390481 -24254 390537 -24198
rect 390339 -24396 390395 -24340
rect 390481 -24396 390537 -24340
rect 390339 -24538 390395 -24482
rect 390481 -24538 390537 -24482
rect 390339 -24680 390395 -24624
rect 390481 -24680 390537 -24624
rect 390339 -24822 390395 -24766
rect 390481 -24822 390537 -24766
rect 390339 -24964 390395 -24908
rect 390481 -24964 390537 -24908
rect 390339 -25106 390395 -25050
rect 390481 -25106 390537 -25050
rect 390339 -25248 390395 -25192
rect 390481 -25248 390537 -25192
rect 390339 -25390 390395 -25334
rect 390481 -25390 390537 -25334
rect 390339 -25532 390395 -25476
rect 390481 -25532 390537 -25476
rect 390736 -18006 390792 -17950
rect 390878 -18006 390934 -17950
rect 390736 -18148 390792 -18092
rect 390878 -18148 390934 -18092
rect 390736 -18290 390792 -18234
rect 390878 -18290 390934 -18234
rect 390736 -18432 390792 -18376
rect 390878 -18432 390934 -18376
rect 390736 -18574 390792 -18518
rect 390878 -18574 390934 -18518
rect 390736 -18716 390792 -18660
rect 390878 -18716 390934 -18660
rect 390736 -18858 390792 -18802
rect 390878 -18858 390934 -18802
rect 390736 -19000 390792 -18944
rect 390878 -19000 390934 -18944
rect 390736 -19142 390792 -19086
rect 390878 -19142 390934 -19086
rect 390736 -19284 390792 -19228
rect 390878 -19284 390934 -19228
rect 390736 -19426 390792 -19370
rect 390878 -19426 390934 -19370
rect 390736 -19568 390792 -19512
rect 390878 -19568 390934 -19512
rect 390736 -19710 390792 -19654
rect 390878 -19710 390934 -19654
rect 390736 -19852 390792 -19796
rect 390878 -19852 390934 -19796
rect 390736 -19994 390792 -19938
rect 390878 -19994 390934 -19938
rect 390736 -20136 390792 -20080
rect 390878 -20136 390934 -20080
rect 390736 -20278 390792 -20222
rect 390878 -20278 390934 -20222
rect 390736 -20420 390792 -20364
rect 390878 -20420 390934 -20364
rect 390736 -20562 390792 -20506
rect 390878 -20562 390934 -20506
rect 390736 -20704 390792 -20648
rect 390878 -20704 390934 -20648
rect 390736 -20846 390792 -20790
rect 390878 -20846 390934 -20790
rect 390736 -20988 390792 -20932
rect 390878 -20988 390934 -20932
rect 390736 -21130 390792 -21074
rect 390878 -21130 390934 -21074
rect 390736 -21272 390792 -21216
rect 390878 -21272 390934 -21216
rect 390736 -21414 390792 -21358
rect 390878 -21414 390934 -21358
rect 390736 -21556 390792 -21500
rect 390878 -21556 390934 -21500
rect 390736 -21698 390792 -21642
rect 390878 -21698 390934 -21642
rect 390736 -21840 390792 -21784
rect 390878 -21840 390934 -21784
rect 390736 -21982 390792 -21926
rect 390878 -21982 390934 -21926
rect 390736 -22124 390792 -22068
rect 390878 -22124 390934 -22068
rect 390736 -22266 390792 -22210
rect 390878 -22266 390934 -22210
rect 390736 -22408 390792 -22352
rect 390878 -22408 390934 -22352
rect 390736 -22550 390792 -22494
rect 390878 -22550 390934 -22494
rect 390736 -22692 390792 -22636
rect 390878 -22692 390934 -22636
rect 390736 -22834 390792 -22778
rect 390878 -22834 390934 -22778
rect 390736 -22976 390792 -22920
rect 390878 -22976 390934 -22920
rect 390736 -23118 390792 -23062
rect 390878 -23118 390934 -23062
rect 390736 -23260 390792 -23204
rect 390878 -23260 390934 -23204
rect 390736 -23402 390792 -23346
rect 390878 -23402 390934 -23346
rect 390736 -23544 390792 -23488
rect 390878 -23544 390934 -23488
rect 390736 -23686 390792 -23630
rect 390878 -23686 390934 -23630
rect 390736 -23828 390792 -23772
rect 390878 -23828 390934 -23772
rect 390736 -23970 390792 -23914
rect 390878 -23970 390934 -23914
rect 390736 -24112 390792 -24056
rect 390878 -24112 390934 -24056
rect 390736 -24254 390792 -24198
rect 390878 -24254 390934 -24198
rect 390736 -24396 390792 -24340
rect 390878 -24396 390934 -24340
rect 390736 -24538 390792 -24482
rect 390878 -24538 390934 -24482
rect 390736 -24680 390792 -24624
rect 390878 -24680 390934 -24624
rect 390736 -24822 390792 -24766
rect 390878 -24822 390934 -24766
rect 390736 -24964 390792 -24908
rect 390878 -24964 390934 -24908
rect 390736 -25106 390792 -25050
rect 390878 -25106 390934 -25050
rect 390736 -25248 390792 -25192
rect 390878 -25248 390934 -25192
rect 390736 -25390 390792 -25334
rect 390878 -25390 390934 -25334
rect 390736 -25532 390792 -25476
rect 390878 -25532 390934 -25476
rect 391140 -18006 391196 -17950
rect 391282 -18006 391338 -17950
rect 391140 -18148 391196 -18092
rect 391282 -18148 391338 -18092
rect 391140 -18290 391196 -18234
rect 391282 -18290 391338 -18234
rect 391140 -18432 391196 -18376
rect 391282 -18432 391338 -18376
rect 391140 -18574 391196 -18518
rect 391282 -18574 391338 -18518
rect 391140 -18716 391196 -18660
rect 391282 -18716 391338 -18660
rect 391140 -18858 391196 -18802
rect 391282 -18858 391338 -18802
rect 391140 -19000 391196 -18944
rect 391282 -19000 391338 -18944
rect 391140 -19142 391196 -19086
rect 391282 -19142 391338 -19086
rect 391140 -19284 391196 -19228
rect 391282 -19284 391338 -19228
rect 391140 -19426 391196 -19370
rect 391282 -19426 391338 -19370
rect 391140 -19568 391196 -19512
rect 391282 -19568 391338 -19512
rect 391140 -19710 391196 -19654
rect 391282 -19710 391338 -19654
rect 391140 -19852 391196 -19796
rect 391282 -19852 391338 -19796
rect 391140 -19994 391196 -19938
rect 391282 -19994 391338 -19938
rect 391140 -20136 391196 -20080
rect 391282 -20136 391338 -20080
rect 391140 -20278 391196 -20222
rect 391282 -20278 391338 -20222
rect 391140 -20420 391196 -20364
rect 391282 -20420 391338 -20364
rect 391140 -20562 391196 -20506
rect 391282 -20562 391338 -20506
rect 391140 -20704 391196 -20648
rect 391282 -20704 391338 -20648
rect 391140 -20846 391196 -20790
rect 391282 -20846 391338 -20790
rect 391140 -20988 391196 -20932
rect 391282 -20988 391338 -20932
rect 391140 -21130 391196 -21074
rect 391282 -21130 391338 -21074
rect 391140 -21272 391196 -21216
rect 391282 -21272 391338 -21216
rect 391140 -21414 391196 -21358
rect 391282 -21414 391338 -21358
rect 391140 -21556 391196 -21500
rect 391282 -21556 391338 -21500
rect 391140 -21698 391196 -21642
rect 391282 -21698 391338 -21642
rect 391140 -21840 391196 -21784
rect 391282 -21840 391338 -21784
rect 391140 -21982 391196 -21926
rect 391282 -21982 391338 -21926
rect 391140 -22124 391196 -22068
rect 391282 -22124 391338 -22068
rect 391140 -22266 391196 -22210
rect 391282 -22266 391338 -22210
rect 391140 -22408 391196 -22352
rect 391282 -22408 391338 -22352
rect 391140 -22550 391196 -22494
rect 391282 -22550 391338 -22494
rect 391140 -22692 391196 -22636
rect 391282 -22692 391338 -22636
rect 391140 -22834 391196 -22778
rect 391282 -22834 391338 -22778
rect 391140 -22976 391196 -22920
rect 391282 -22976 391338 -22920
rect 391140 -23118 391196 -23062
rect 391282 -23118 391338 -23062
rect 391140 -23260 391196 -23204
rect 391282 -23260 391338 -23204
rect 391140 -23402 391196 -23346
rect 391282 -23402 391338 -23346
rect 391140 -23544 391196 -23488
rect 391282 -23544 391338 -23488
rect 391140 -23686 391196 -23630
rect 391282 -23686 391338 -23630
rect 391140 -23828 391196 -23772
rect 391282 -23828 391338 -23772
rect 391140 -23970 391196 -23914
rect 391282 -23970 391338 -23914
rect 391140 -24112 391196 -24056
rect 391282 -24112 391338 -24056
rect 391140 -24254 391196 -24198
rect 391282 -24254 391338 -24198
rect 391140 -24396 391196 -24340
rect 391282 -24396 391338 -24340
rect 391140 -24538 391196 -24482
rect 391282 -24538 391338 -24482
rect 391140 -24680 391196 -24624
rect 391282 -24680 391338 -24624
rect 391140 -24822 391196 -24766
rect 391282 -24822 391338 -24766
rect 391140 -24964 391196 -24908
rect 391282 -24964 391338 -24908
rect 391140 -25106 391196 -25050
rect 391282 -25106 391338 -25050
rect 391140 -25248 391196 -25192
rect 391282 -25248 391338 -25192
rect 391140 -25390 391196 -25334
rect 391282 -25390 391338 -25334
rect 391140 -25532 391196 -25476
rect 391282 -25532 391338 -25476
rect 391536 -18006 391592 -17950
rect 391678 -18006 391734 -17950
rect 391536 -18148 391592 -18092
rect 391678 -18148 391734 -18092
rect 391536 -18290 391592 -18234
rect 391678 -18290 391734 -18234
rect 391536 -18432 391592 -18376
rect 391678 -18432 391734 -18376
rect 391536 -18574 391592 -18518
rect 391678 -18574 391734 -18518
rect 391536 -18716 391592 -18660
rect 391678 -18716 391734 -18660
rect 391536 -18858 391592 -18802
rect 391678 -18858 391734 -18802
rect 391536 -19000 391592 -18944
rect 391678 -19000 391734 -18944
rect 391536 -19142 391592 -19086
rect 391678 -19142 391734 -19086
rect 391536 -19284 391592 -19228
rect 391678 -19284 391734 -19228
rect 391536 -19426 391592 -19370
rect 391678 -19426 391734 -19370
rect 391536 -19568 391592 -19512
rect 391678 -19568 391734 -19512
rect 391536 -19710 391592 -19654
rect 391678 -19710 391734 -19654
rect 391536 -19852 391592 -19796
rect 391678 -19852 391734 -19796
rect 391536 -19994 391592 -19938
rect 391678 -19994 391734 -19938
rect 391536 -20136 391592 -20080
rect 391678 -20136 391734 -20080
rect 391536 -20278 391592 -20222
rect 391678 -20278 391734 -20222
rect 391536 -20420 391592 -20364
rect 391678 -20420 391734 -20364
rect 391536 -20562 391592 -20506
rect 391678 -20562 391734 -20506
rect 391536 -20704 391592 -20648
rect 391678 -20704 391734 -20648
rect 391536 -20846 391592 -20790
rect 391678 -20846 391734 -20790
rect 391536 -20988 391592 -20932
rect 391678 -20988 391734 -20932
rect 391536 -21130 391592 -21074
rect 391678 -21130 391734 -21074
rect 391536 -21272 391592 -21216
rect 391678 -21272 391734 -21216
rect 391536 -21414 391592 -21358
rect 391678 -21414 391734 -21358
rect 391536 -21556 391592 -21500
rect 391678 -21556 391734 -21500
rect 391536 -21698 391592 -21642
rect 391678 -21698 391734 -21642
rect 391536 -21840 391592 -21784
rect 391678 -21840 391734 -21784
rect 391536 -21982 391592 -21926
rect 391678 -21982 391734 -21926
rect 391536 -22124 391592 -22068
rect 391678 -22124 391734 -22068
rect 391536 -22266 391592 -22210
rect 391678 -22266 391734 -22210
rect 391536 -22408 391592 -22352
rect 391678 -22408 391734 -22352
rect 391536 -22550 391592 -22494
rect 391678 -22550 391734 -22494
rect 391536 -22692 391592 -22636
rect 391678 -22692 391734 -22636
rect 391536 -22834 391592 -22778
rect 391678 -22834 391734 -22778
rect 391536 -22976 391592 -22920
rect 391678 -22976 391734 -22920
rect 391536 -23118 391592 -23062
rect 391678 -23118 391734 -23062
rect 391536 -23260 391592 -23204
rect 391678 -23260 391734 -23204
rect 391536 -23402 391592 -23346
rect 391678 -23402 391734 -23346
rect 391536 -23544 391592 -23488
rect 391678 -23544 391734 -23488
rect 391536 -23686 391592 -23630
rect 391678 -23686 391734 -23630
rect 391536 -23828 391592 -23772
rect 391678 -23828 391734 -23772
rect 391536 -23970 391592 -23914
rect 391678 -23970 391734 -23914
rect 391536 -24112 391592 -24056
rect 391678 -24112 391734 -24056
rect 391536 -24254 391592 -24198
rect 391678 -24254 391734 -24198
rect 391536 -24396 391592 -24340
rect 391678 -24396 391734 -24340
rect 391536 -24538 391592 -24482
rect 391678 -24538 391734 -24482
rect 391536 -24680 391592 -24624
rect 391678 -24680 391734 -24624
rect 391536 -24822 391592 -24766
rect 391678 -24822 391734 -24766
rect 391536 -24964 391592 -24908
rect 391678 -24964 391734 -24908
rect 391536 -25106 391592 -25050
rect 391678 -25106 391734 -25050
rect 391536 -25248 391592 -25192
rect 391678 -25248 391734 -25192
rect 391536 -25390 391592 -25334
rect 391678 -25390 391734 -25334
rect 391536 -25532 391592 -25476
rect 391678 -25532 391734 -25476
rect 391936 -18006 391992 -17950
rect 392078 -18006 392134 -17950
rect 391936 -18148 391992 -18092
rect 392078 -18148 392134 -18092
rect 391936 -18290 391992 -18234
rect 392078 -18290 392134 -18234
rect 391936 -18432 391992 -18376
rect 392078 -18432 392134 -18376
rect 391936 -18574 391992 -18518
rect 392078 -18574 392134 -18518
rect 391936 -18716 391992 -18660
rect 392078 -18716 392134 -18660
rect 391936 -18858 391992 -18802
rect 392078 -18858 392134 -18802
rect 391936 -19000 391992 -18944
rect 392078 -19000 392134 -18944
rect 391936 -19142 391992 -19086
rect 392078 -19142 392134 -19086
rect 391936 -19284 391992 -19228
rect 392078 -19284 392134 -19228
rect 391936 -19426 391992 -19370
rect 392078 -19426 392134 -19370
rect 391936 -19568 391992 -19512
rect 392078 -19568 392134 -19512
rect 391936 -19710 391992 -19654
rect 392078 -19710 392134 -19654
rect 391936 -19852 391992 -19796
rect 392078 -19852 392134 -19796
rect 391936 -19994 391992 -19938
rect 392078 -19994 392134 -19938
rect 391936 -20136 391992 -20080
rect 392078 -20136 392134 -20080
rect 391936 -20278 391992 -20222
rect 392078 -20278 392134 -20222
rect 391936 -20420 391992 -20364
rect 392078 -20420 392134 -20364
rect 391936 -20562 391992 -20506
rect 392078 -20562 392134 -20506
rect 391936 -20704 391992 -20648
rect 392078 -20704 392134 -20648
rect 391936 -20846 391992 -20790
rect 392078 -20846 392134 -20790
rect 391936 -20988 391992 -20932
rect 392078 -20988 392134 -20932
rect 391936 -21130 391992 -21074
rect 392078 -21130 392134 -21074
rect 391936 -21272 391992 -21216
rect 392078 -21272 392134 -21216
rect 391936 -21414 391992 -21358
rect 392078 -21414 392134 -21358
rect 391936 -21556 391992 -21500
rect 392078 -21556 392134 -21500
rect 391936 -21698 391992 -21642
rect 392078 -21698 392134 -21642
rect 391936 -21840 391992 -21784
rect 392078 -21840 392134 -21784
rect 391936 -21982 391992 -21926
rect 392078 -21982 392134 -21926
rect 391936 -22124 391992 -22068
rect 392078 -22124 392134 -22068
rect 391936 -22266 391992 -22210
rect 392078 -22266 392134 -22210
rect 391936 -22408 391992 -22352
rect 392078 -22408 392134 -22352
rect 391936 -22550 391992 -22494
rect 392078 -22550 392134 -22494
rect 391936 -22692 391992 -22636
rect 392078 -22692 392134 -22636
rect 391936 -22834 391992 -22778
rect 392078 -22834 392134 -22778
rect 391936 -22976 391992 -22920
rect 392078 -22976 392134 -22920
rect 391936 -23118 391992 -23062
rect 392078 -23118 392134 -23062
rect 391936 -23260 391992 -23204
rect 392078 -23260 392134 -23204
rect 391936 -23402 391992 -23346
rect 392078 -23402 392134 -23346
rect 391936 -23544 391992 -23488
rect 392078 -23544 392134 -23488
rect 391936 -23686 391992 -23630
rect 392078 -23686 392134 -23630
rect 391936 -23828 391992 -23772
rect 392078 -23828 392134 -23772
rect 391936 -23970 391992 -23914
rect 392078 -23970 392134 -23914
rect 391936 -24112 391992 -24056
rect 392078 -24112 392134 -24056
rect 391936 -24254 391992 -24198
rect 392078 -24254 392134 -24198
rect 391936 -24396 391992 -24340
rect 392078 -24396 392134 -24340
rect 391936 -24538 391992 -24482
rect 392078 -24538 392134 -24482
rect 391936 -24680 391992 -24624
rect 392078 -24680 392134 -24624
rect 391936 -24822 391992 -24766
rect 392078 -24822 392134 -24766
rect 391936 -24964 391992 -24908
rect 392078 -24964 392134 -24908
rect 391936 -25106 391992 -25050
rect 392078 -25106 392134 -25050
rect 391936 -25248 391992 -25192
rect 392078 -25248 392134 -25192
rect 391936 -25390 391992 -25334
rect 392078 -25390 392134 -25334
rect 391936 -25532 391992 -25476
rect 392078 -25532 392134 -25476
rect 392333 -18006 392389 -17950
rect 392475 -18006 392531 -17950
rect 392333 -18148 392389 -18092
rect 392475 -18148 392531 -18092
rect 392333 -18290 392389 -18234
rect 392475 -18290 392531 -18234
rect 392333 -18432 392389 -18376
rect 392475 -18432 392531 -18376
rect 392333 -18574 392389 -18518
rect 392475 -18574 392531 -18518
rect 392333 -18716 392389 -18660
rect 392475 -18716 392531 -18660
rect 392333 -18858 392389 -18802
rect 392475 -18858 392531 -18802
rect 392333 -19000 392389 -18944
rect 392475 -19000 392531 -18944
rect 392333 -19142 392389 -19086
rect 392475 -19142 392531 -19086
rect 392333 -19284 392389 -19228
rect 392475 -19284 392531 -19228
rect 392333 -19426 392389 -19370
rect 392475 -19426 392531 -19370
rect 392333 -19568 392389 -19512
rect 392475 -19568 392531 -19512
rect 392333 -19710 392389 -19654
rect 392475 -19710 392531 -19654
rect 392333 -19852 392389 -19796
rect 392475 -19852 392531 -19796
rect 392333 -19994 392389 -19938
rect 392475 -19994 392531 -19938
rect 392333 -20136 392389 -20080
rect 392475 -20136 392531 -20080
rect 392333 -20278 392389 -20222
rect 392475 -20278 392531 -20222
rect 392333 -20420 392389 -20364
rect 392475 -20420 392531 -20364
rect 392333 -20562 392389 -20506
rect 392475 -20562 392531 -20506
rect 392333 -20704 392389 -20648
rect 392475 -20704 392531 -20648
rect 392333 -20846 392389 -20790
rect 392475 -20846 392531 -20790
rect 392333 -20988 392389 -20932
rect 392475 -20988 392531 -20932
rect 392333 -21130 392389 -21074
rect 392475 -21130 392531 -21074
rect 392333 -21272 392389 -21216
rect 392475 -21272 392531 -21216
rect 392333 -21414 392389 -21358
rect 392475 -21414 392531 -21358
rect 392333 -21556 392389 -21500
rect 392475 -21556 392531 -21500
rect 392333 -21698 392389 -21642
rect 392475 -21698 392531 -21642
rect 392333 -21840 392389 -21784
rect 392475 -21840 392531 -21784
rect 392333 -21982 392389 -21926
rect 392475 -21982 392531 -21926
rect 392333 -22124 392389 -22068
rect 392475 -22124 392531 -22068
rect 392333 -22266 392389 -22210
rect 392475 -22266 392531 -22210
rect 392333 -22408 392389 -22352
rect 392475 -22408 392531 -22352
rect 392333 -22550 392389 -22494
rect 392475 -22550 392531 -22494
rect 392333 -22692 392389 -22636
rect 392475 -22692 392531 -22636
rect 392333 -22834 392389 -22778
rect 392475 -22834 392531 -22778
rect 392333 -22976 392389 -22920
rect 392475 -22976 392531 -22920
rect 392333 -23118 392389 -23062
rect 392475 -23118 392531 -23062
rect 392333 -23260 392389 -23204
rect 392475 -23260 392531 -23204
rect 392333 -23402 392389 -23346
rect 392475 -23402 392531 -23346
rect 392333 -23544 392389 -23488
rect 392475 -23544 392531 -23488
rect 392333 -23686 392389 -23630
rect 392475 -23686 392531 -23630
rect 392333 -23828 392389 -23772
rect 392475 -23828 392531 -23772
rect 392333 -23970 392389 -23914
rect 392475 -23970 392531 -23914
rect 392333 -24112 392389 -24056
rect 392475 -24112 392531 -24056
rect 392333 -24254 392389 -24198
rect 392475 -24254 392531 -24198
rect 392333 -24396 392389 -24340
rect 392475 -24396 392531 -24340
rect 392333 -24538 392389 -24482
rect 392475 -24538 392531 -24482
rect 392333 -24680 392389 -24624
rect 392475 -24680 392531 -24624
rect 392333 -24822 392389 -24766
rect 392475 -24822 392531 -24766
rect 392333 -24964 392389 -24908
rect 392475 -24964 392531 -24908
rect 392333 -25106 392389 -25050
rect 392475 -25106 392531 -25050
rect 392333 -25248 392389 -25192
rect 392475 -25248 392531 -25192
rect 392333 -25390 392389 -25334
rect 392475 -25390 392531 -25334
rect 392333 -25532 392389 -25476
rect 392475 -25532 392531 -25476
rect 392738 -18006 392794 -17950
rect 392880 -18006 392936 -17950
rect 392738 -18148 392794 -18092
rect 392880 -18148 392936 -18092
rect 392738 -18290 392794 -18234
rect 392880 -18290 392936 -18234
rect 392738 -18432 392794 -18376
rect 392880 -18432 392936 -18376
rect 392738 -18574 392794 -18518
rect 392880 -18574 392936 -18518
rect 392738 -18716 392794 -18660
rect 392880 -18716 392936 -18660
rect 392738 -18858 392794 -18802
rect 392880 -18858 392936 -18802
rect 392738 -19000 392794 -18944
rect 392880 -19000 392936 -18944
rect 392738 -19142 392794 -19086
rect 392880 -19142 392936 -19086
rect 392738 -19284 392794 -19228
rect 392880 -19284 392936 -19228
rect 392738 -19426 392794 -19370
rect 392880 -19426 392936 -19370
rect 392738 -19568 392794 -19512
rect 392880 -19568 392936 -19512
rect 392738 -19710 392794 -19654
rect 392880 -19710 392936 -19654
rect 392738 -19852 392794 -19796
rect 392880 -19852 392936 -19796
rect 392738 -19994 392794 -19938
rect 392880 -19994 392936 -19938
rect 392738 -20136 392794 -20080
rect 392880 -20136 392936 -20080
rect 392738 -20278 392794 -20222
rect 392880 -20278 392936 -20222
rect 392738 -20420 392794 -20364
rect 392880 -20420 392936 -20364
rect 392738 -20562 392794 -20506
rect 392880 -20562 392936 -20506
rect 392738 -20704 392794 -20648
rect 392880 -20704 392936 -20648
rect 392738 -20846 392794 -20790
rect 392880 -20846 392936 -20790
rect 392738 -20988 392794 -20932
rect 392880 -20988 392936 -20932
rect 392738 -21130 392794 -21074
rect 392880 -21130 392936 -21074
rect 392738 -21272 392794 -21216
rect 392880 -21272 392936 -21216
rect 392738 -21414 392794 -21358
rect 392880 -21414 392936 -21358
rect 392738 -21556 392794 -21500
rect 392880 -21556 392936 -21500
rect 392738 -21698 392794 -21642
rect 392880 -21698 392936 -21642
rect 392738 -21840 392794 -21784
rect 392880 -21840 392936 -21784
rect 392738 -21982 392794 -21926
rect 392880 -21982 392936 -21926
rect 392738 -22124 392794 -22068
rect 392880 -22124 392936 -22068
rect 392738 -22266 392794 -22210
rect 392880 -22266 392936 -22210
rect 392738 -22408 392794 -22352
rect 392880 -22408 392936 -22352
rect 392738 -22550 392794 -22494
rect 392880 -22550 392936 -22494
rect 392738 -22692 392794 -22636
rect 392880 -22692 392936 -22636
rect 392738 -22834 392794 -22778
rect 392880 -22834 392936 -22778
rect 392738 -22976 392794 -22920
rect 392880 -22976 392936 -22920
rect 392738 -23118 392794 -23062
rect 392880 -23118 392936 -23062
rect 392738 -23260 392794 -23204
rect 392880 -23260 392936 -23204
rect 392738 -23402 392794 -23346
rect 392880 -23402 392936 -23346
rect 392738 -23544 392794 -23488
rect 392880 -23544 392936 -23488
rect 392738 -23686 392794 -23630
rect 392880 -23686 392936 -23630
rect 392738 -23828 392794 -23772
rect 392880 -23828 392936 -23772
rect 392738 -23970 392794 -23914
rect 392880 -23970 392936 -23914
rect 392738 -24112 392794 -24056
rect 392880 -24112 392936 -24056
rect 392738 -24254 392794 -24198
rect 392880 -24254 392936 -24198
rect 392738 -24396 392794 -24340
rect 392880 -24396 392936 -24340
rect 392738 -24538 392794 -24482
rect 392880 -24538 392936 -24482
rect 392738 -24680 392794 -24624
rect 392880 -24680 392936 -24624
rect 392738 -24822 392794 -24766
rect 392880 -24822 392936 -24766
rect 392738 -24964 392794 -24908
rect 392880 -24964 392936 -24908
rect 392738 -25106 392794 -25050
rect 392880 -25106 392936 -25050
rect 392738 -25248 392794 -25192
rect 392880 -25248 392936 -25192
rect 392738 -25390 392794 -25334
rect 392880 -25390 392936 -25334
rect 392738 -25532 392794 -25476
rect 392880 -25532 392936 -25476
rect 393138 -18006 393194 -17950
rect 393280 -18006 393336 -17950
rect 393138 -18148 393194 -18092
rect 393280 -18148 393336 -18092
rect 393138 -18290 393194 -18234
rect 393280 -18290 393336 -18234
rect 393138 -18432 393194 -18376
rect 393280 -18432 393336 -18376
rect 393138 -18574 393194 -18518
rect 393280 -18574 393336 -18518
rect 393138 -18716 393194 -18660
rect 393280 -18716 393336 -18660
rect 393138 -18858 393194 -18802
rect 393280 -18858 393336 -18802
rect 393138 -19000 393194 -18944
rect 393280 -19000 393336 -18944
rect 393138 -19142 393194 -19086
rect 393280 -19142 393336 -19086
rect 393138 -19284 393194 -19228
rect 393280 -19284 393336 -19228
rect 393138 -19426 393194 -19370
rect 393280 -19426 393336 -19370
rect 393138 -19568 393194 -19512
rect 393280 -19568 393336 -19512
rect 393138 -19710 393194 -19654
rect 393280 -19710 393336 -19654
rect 393138 -19852 393194 -19796
rect 393280 -19852 393336 -19796
rect 393138 -19994 393194 -19938
rect 393280 -19994 393336 -19938
rect 393138 -20136 393194 -20080
rect 393280 -20136 393336 -20080
rect 393138 -20278 393194 -20222
rect 393280 -20278 393336 -20222
rect 393138 -20420 393194 -20364
rect 393280 -20420 393336 -20364
rect 393138 -20562 393194 -20506
rect 393280 -20562 393336 -20506
rect 393138 -20704 393194 -20648
rect 393280 -20704 393336 -20648
rect 393138 -20846 393194 -20790
rect 393280 -20846 393336 -20790
rect 393138 -20988 393194 -20932
rect 393280 -20988 393336 -20932
rect 393138 -21130 393194 -21074
rect 393280 -21130 393336 -21074
rect 393138 -21272 393194 -21216
rect 393280 -21272 393336 -21216
rect 393138 -21414 393194 -21358
rect 393280 -21414 393336 -21358
rect 393138 -21556 393194 -21500
rect 393280 -21556 393336 -21500
rect 393138 -21698 393194 -21642
rect 393280 -21698 393336 -21642
rect 393138 -21840 393194 -21784
rect 393280 -21840 393336 -21784
rect 393138 -21982 393194 -21926
rect 393280 -21982 393336 -21926
rect 393138 -22124 393194 -22068
rect 393280 -22124 393336 -22068
rect 393138 -22266 393194 -22210
rect 393280 -22266 393336 -22210
rect 393138 -22408 393194 -22352
rect 393280 -22408 393336 -22352
rect 393138 -22550 393194 -22494
rect 393280 -22550 393336 -22494
rect 393138 -22692 393194 -22636
rect 393280 -22692 393336 -22636
rect 393138 -22834 393194 -22778
rect 393280 -22834 393336 -22778
rect 393138 -22976 393194 -22920
rect 393280 -22976 393336 -22920
rect 393138 -23118 393194 -23062
rect 393280 -23118 393336 -23062
rect 393138 -23260 393194 -23204
rect 393280 -23260 393336 -23204
rect 393138 -23402 393194 -23346
rect 393280 -23402 393336 -23346
rect 393138 -23544 393194 -23488
rect 393280 -23544 393336 -23488
rect 393138 -23686 393194 -23630
rect 393280 -23686 393336 -23630
rect 393138 -23828 393194 -23772
rect 393280 -23828 393336 -23772
rect 393138 -23970 393194 -23914
rect 393280 -23970 393336 -23914
rect 393138 -24112 393194 -24056
rect 393280 -24112 393336 -24056
rect 393138 -24254 393194 -24198
rect 393280 -24254 393336 -24198
rect 393138 -24396 393194 -24340
rect 393280 -24396 393336 -24340
rect 393138 -24538 393194 -24482
rect 393280 -24538 393336 -24482
rect 393138 -24680 393194 -24624
rect 393280 -24680 393336 -24624
rect 393138 -24822 393194 -24766
rect 393280 -24822 393336 -24766
rect 393138 -24964 393194 -24908
rect 393280 -24964 393336 -24908
rect 393138 -25106 393194 -25050
rect 393280 -25106 393336 -25050
rect 393138 -25248 393194 -25192
rect 393280 -25248 393336 -25192
rect 393138 -25390 393194 -25334
rect 393280 -25390 393336 -25334
rect 393138 -25532 393194 -25476
rect 393280 -25532 393336 -25476
rect 393543 -18006 393599 -17950
rect 393685 -18006 393741 -17950
rect 393543 -18148 393599 -18092
rect 393685 -18148 393741 -18092
rect 393543 -18290 393599 -18234
rect 393685 -18290 393741 -18234
rect 393543 -18432 393599 -18376
rect 393685 -18432 393741 -18376
rect 393543 -18574 393599 -18518
rect 393685 -18574 393741 -18518
rect 393543 -18716 393599 -18660
rect 393685 -18716 393741 -18660
rect 393543 -18858 393599 -18802
rect 393685 -18858 393741 -18802
rect 393543 -19000 393599 -18944
rect 393685 -19000 393741 -18944
rect 393543 -19142 393599 -19086
rect 393685 -19142 393741 -19086
rect 393543 -19284 393599 -19228
rect 393685 -19284 393741 -19228
rect 393543 -19426 393599 -19370
rect 393685 -19426 393741 -19370
rect 393543 -19568 393599 -19512
rect 393685 -19568 393741 -19512
rect 393543 -19710 393599 -19654
rect 393685 -19710 393741 -19654
rect 393543 -19852 393599 -19796
rect 393685 -19852 393741 -19796
rect 393543 -19994 393599 -19938
rect 393685 -19994 393741 -19938
rect 393543 -20136 393599 -20080
rect 393685 -20136 393741 -20080
rect 393543 -20278 393599 -20222
rect 393685 -20278 393741 -20222
rect 393543 -20420 393599 -20364
rect 393685 -20420 393741 -20364
rect 393543 -20562 393599 -20506
rect 393685 -20562 393741 -20506
rect 393543 -20704 393599 -20648
rect 393685 -20704 393741 -20648
rect 393543 -20846 393599 -20790
rect 393685 -20846 393741 -20790
rect 393543 -20988 393599 -20932
rect 393685 -20988 393741 -20932
rect 393543 -21130 393599 -21074
rect 393685 -21130 393741 -21074
rect 393543 -21272 393599 -21216
rect 393685 -21272 393741 -21216
rect 393543 -21414 393599 -21358
rect 393685 -21414 393741 -21358
rect 393543 -21556 393599 -21500
rect 393685 -21556 393741 -21500
rect 393543 -21698 393599 -21642
rect 393685 -21698 393741 -21642
rect 393543 -21840 393599 -21784
rect 393685 -21840 393741 -21784
rect 393543 -21982 393599 -21926
rect 393685 -21982 393741 -21926
rect 393543 -22124 393599 -22068
rect 393685 -22124 393741 -22068
rect 393543 -22266 393599 -22210
rect 393685 -22266 393741 -22210
rect 393543 -22408 393599 -22352
rect 393685 -22408 393741 -22352
rect 393543 -22550 393599 -22494
rect 393685 -22550 393741 -22494
rect 393543 -22692 393599 -22636
rect 393685 -22692 393741 -22636
rect 393543 -22834 393599 -22778
rect 393685 -22834 393741 -22778
rect 393543 -22976 393599 -22920
rect 393685 -22976 393741 -22920
rect 393543 -23118 393599 -23062
rect 393685 -23118 393741 -23062
rect 393543 -23260 393599 -23204
rect 393685 -23260 393741 -23204
rect 393543 -23402 393599 -23346
rect 393685 -23402 393741 -23346
rect 393543 -23544 393599 -23488
rect 393685 -23544 393741 -23488
rect 393543 -23686 393599 -23630
rect 393685 -23686 393741 -23630
rect 393543 -23828 393599 -23772
rect 393685 -23828 393741 -23772
rect 393543 -23970 393599 -23914
rect 393685 -23970 393741 -23914
rect 393543 -24112 393599 -24056
rect 393685 -24112 393741 -24056
rect 393543 -24254 393599 -24198
rect 393685 -24254 393741 -24198
rect 393543 -24396 393599 -24340
rect 393685 -24396 393741 -24340
rect 393543 -24538 393599 -24482
rect 393685 -24538 393741 -24482
rect 393543 -24680 393599 -24624
rect 393685 -24680 393741 -24624
rect 393543 -24822 393599 -24766
rect 393685 -24822 393741 -24766
rect 393543 -24964 393599 -24908
rect 393685 -24964 393741 -24908
rect 393543 -25106 393599 -25050
rect 393685 -25106 393741 -25050
rect 393543 -25248 393599 -25192
rect 393685 -25248 393741 -25192
rect 393543 -25390 393599 -25334
rect 393685 -25390 393741 -25334
rect 393543 -25532 393599 -25476
rect 393685 -25532 393741 -25476
rect 393940 -18006 393996 -17950
rect 394082 -18006 394138 -17950
rect 393940 -18148 393996 -18092
rect 394082 -18148 394138 -18092
rect 393940 -18290 393996 -18234
rect 394082 -18290 394138 -18234
rect 393940 -18432 393996 -18376
rect 394082 -18432 394138 -18376
rect 393940 -18574 393996 -18518
rect 394082 -18574 394138 -18518
rect 393940 -18716 393996 -18660
rect 394082 -18716 394138 -18660
rect 393940 -18858 393996 -18802
rect 394082 -18858 394138 -18802
rect 393940 -19000 393996 -18944
rect 394082 -19000 394138 -18944
rect 393940 -19142 393996 -19086
rect 394082 -19142 394138 -19086
rect 393940 -19284 393996 -19228
rect 394082 -19284 394138 -19228
rect 393940 -19426 393996 -19370
rect 394082 -19426 394138 -19370
rect 393940 -19568 393996 -19512
rect 394082 -19568 394138 -19512
rect 393940 -19710 393996 -19654
rect 394082 -19710 394138 -19654
rect 393940 -19852 393996 -19796
rect 394082 -19852 394138 -19796
rect 393940 -19994 393996 -19938
rect 394082 -19994 394138 -19938
rect 393940 -20136 393996 -20080
rect 394082 -20136 394138 -20080
rect 393940 -20278 393996 -20222
rect 394082 -20278 394138 -20222
rect 393940 -20420 393996 -20364
rect 394082 -20420 394138 -20364
rect 393940 -20562 393996 -20506
rect 394082 -20562 394138 -20506
rect 393940 -20704 393996 -20648
rect 394082 -20704 394138 -20648
rect 393940 -20846 393996 -20790
rect 394082 -20846 394138 -20790
rect 393940 -20988 393996 -20932
rect 394082 -20988 394138 -20932
rect 393940 -21130 393996 -21074
rect 394082 -21130 394138 -21074
rect 393940 -21272 393996 -21216
rect 394082 -21272 394138 -21216
rect 393940 -21414 393996 -21358
rect 394082 -21414 394138 -21358
rect 393940 -21556 393996 -21500
rect 394082 -21556 394138 -21500
rect 393940 -21698 393996 -21642
rect 394082 -21698 394138 -21642
rect 393940 -21840 393996 -21784
rect 394082 -21840 394138 -21784
rect 393940 -21982 393996 -21926
rect 394082 -21982 394138 -21926
rect 393940 -22124 393996 -22068
rect 394082 -22124 394138 -22068
rect 393940 -22266 393996 -22210
rect 394082 -22266 394138 -22210
rect 393940 -22408 393996 -22352
rect 394082 -22408 394138 -22352
rect 393940 -22550 393996 -22494
rect 394082 -22550 394138 -22494
rect 393940 -22692 393996 -22636
rect 394082 -22692 394138 -22636
rect 393940 -22834 393996 -22778
rect 394082 -22834 394138 -22778
rect 393940 -22976 393996 -22920
rect 394082 -22976 394138 -22920
rect 393940 -23118 393996 -23062
rect 394082 -23118 394138 -23062
rect 393940 -23260 393996 -23204
rect 394082 -23260 394138 -23204
rect 393940 -23402 393996 -23346
rect 394082 -23402 394138 -23346
rect 393940 -23544 393996 -23488
rect 394082 -23544 394138 -23488
rect 393940 -23686 393996 -23630
rect 394082 -23686 394138 -23630
rect 393940 -23828 393996 -23772
rect 394082 -23828 394138 -23772
rect 393940 -23970 393996 -23914
rect 394082 -23970 394138 -23914
rect 393940 -24112 393996 -24056
rect 394082 -24112 394138 -24056
rect 393940 -24254 393996 -24198
rect 394082 -24254 394138 -24198
rect 393940 -24396 393996 -24340
rect 394082 -24396 394138 -24340
rect 393940 -24538 393996 -24482
rect 394082 -24538 394138 -24482
rect 393940 -24680 393996 -24624
rect 394082 -24680 394138 -24624
rect 393940 -24822 393996 -24766
rect 394082 -24822 394138 -24766
rect 393940 -24964 393996 -24908
rect 394082 -24964 394138 -24908
rect 393940 -25106 393996 -25050
rect 394082 -25106 394138 -25050
rect 393940 -25248 393996 -25192
rect 394082 -25248 394138 -25192
rect 393940 -25390 393996 -25334
rect 394082 -25390 394138 -25334
rect 393940 -25532 393996 -25476
rect 394082 -25532 394138 -25476
rect 394337 -18006 394393 -17950
rect 394479 -18006 394535 -17950
rect 394337 -18148 394393 -18092
rect 394479 -18148 394535 -18092
rect 394337 -18290 394393 -18234
rect 394479 -18290 394535 -18234
rect 394337 -18432 394393 -18376
rect 394479 -18432 394535 -18376
rect 394337 -18574 394393 -18518
rect 394479 -18574 394535 -18518
rect 394337 -18716 394393 -18660
rect 394479 -18716 394535 -18660
rect 394337 -18858 394393 -18802
rect 394479 -18858 394535 -18802
rect 394337 -19000 394393 -18944
rect 394479 -19000 394535 -18944
rect 394337 -19142 394393 -19086
rect 394479 -19142 394535 -19086
rect 394337 -19284 394393 -19228
rect 394479 -19284 394535 -19228
rect 394337 -19426 394393 -19370
rect 394479 -19426 394535 -19370
rect 394337 -19568 394393 -19512
rect 394479 -19568 394535 -19512
rect 394337 -19710 394393 -19654
rect 394479 -19710 394535 -19654
rect 394337 -19852 394393 -19796
rect 394479 -19852 394535 -19796
rect 394337 -19994 394393 -19938
rect 394479 -19994 394535 -19938
rect 394337 -20136 394393 -20080
rect 394479 -20136 394535 -20080
rect 394337 -20278 394393 -20222
rect 394479 -20278 394535 -20222
rect 394337 -20420 394393 -20364
rect 394479 -20420 394535 -20364
rect 394337 -20562 394393 -20506
rect 394479 -20562 394535 -20506
rect 394337 -20704 394393 -20648
rect 394479 -20704 394535 -20648
rect 394337 -20846 394393 -20790
rect 394479 -20846 394535 -20790
rect 394337 -20988 394393 -20932
rect 394479 -20988 394535 -20932
rect 394337 -21130 394393 -21074
rect 394479 -21130 394535 -21074
rect 394337 -21272 394393 -21216
rect 394479 -21272 394535 -21216
rect 394337 -21414 394393 -21358
rect 394479 -21414 394535 -21358
rect 394337 -21556 394393 -21500
rect 394479 -21556 394535 -21500
rect 394337 -21698 394393 -21642
rect 394479 -21698 394535 -21642
rect 394337 -21840 394393 -21784
rect 394479 -21840 394535 -21784
rect 394337 -21982 394393 -21926
rect 394479 -21982 394535 -21926
rect 394337 -22124 394393 -22068
rect 394479 -22124 394535 -22068
rect 394337 -22266 394393 -22210
rect 394479 -22266 394535 -22210
rect 394337 -22408 394393 -22352
rect 394479 -22408 394535 -22352
rect 394337 -22550 394393 -22494
rect 394479 -22550 394535 -22494
rect 394337 -22692 394393 -22636
rect 394479 -22692 394535 -22636
rect 394337 -22834 394393 -22778
rect 394479 -22834 394535 -22778
rect 394337 -22976 394393 -22920
rect 394479 -22976 394535 -22920
rect 394337 -23118 394393 -23062
rect 394479 -23118 394535 -23062
rect 394337 -23260 394393 -23204
rect 394479 -23260 394535 -23204
rect 394337 -23402 394393 -23346
rect 394479 -23402 394535 -23346
rect 394337 -23544 394393 -23488
rect 394479 -23544 394535 -23488
rect 394337 -23686 394393 -23630
rect 394479 -23686 394535 -23630
rect 394337 -23828 394393 -23772
rect 394479 -23828 394535 -23772
rect 394337 -23970 394393 -23914
rect 394479 -23970 394535 -23914
rect 394337 -24112 394393 -24056
rect 394479 -24112 394535 -24056
rect 394337 -24254 394393 -24198
rect 394479 -24254 394535 -24198
rect 394337 -24396 394393 -24340
rect 394479 -24396 394535 -24340
rect 394337 -24538 394393 -24482
rect 394479 -24538 394535 -24482
rect 394337 -24680 394393 -24624
rect 394479 -24680 394535 -24624
rect 394337 -24822 394393 -24766
rect 394479 -24822 394535 -24766
rect 394337 -24964 394393 -24908
rect 394479 -24964 394535 -24908
rect 394337 -25106 394393 -25050
rect 394479 -25106 394535 -25050
rect 394337 -25248 394393 -25192
rect 394479 -25248 394535 -25192
rect 394337 -25390 394393 -25334
rect 394479 -25390 394535 -25334
rect 394337 -25532 394393 -25476
rect 394479 -25532 394535 -25476
rect 394740 -18006 394796 -17950
rect 394882 -18006 394938 -17950
rect 394740 -18148 394796 -18092
rect 394882 -18148 394938 -18092
rect 394740 -18290 394796 -18234
rect 394882 -18290 394938 -18234
rect 394740 -18432 394796 -18376
rect 394882 -18432 394938 -18376
rect 394740 -18574 394796 -18518
rect 394882 -18574 394938 -18518
rect 394740 -18716 394796 -18660
rect 394882 -18716 394938 -18660
rect 394740 -18858 394796 -18802
rect 394882 -18858 394938 -18802
rect 394740 -19000 394796 -18944
rect 394882 -19000 394938 -18944
rect 394740 -19142 394796 -19086
rect 394882 -19142 394938 -19086
rect 394740 -19284 394796 -19228
rect 394882 -19284 394938 -19228
rect 394740 -19426 394796 -19370
rect 394882 -19426 394938 -19370
rect 394740 -19568 394796 -19512
rect 394882 -19568 394938 -19512
rect 394740 -19710 394796 -19654
rect 394882 -19710 394938 -19654
rect 394740 -19852 394796 -19796
rect 394882 -19852 394938 -19796
rect 394740 -19994 394796 -19938
rect 394882 -19994 394938 -19938
rect 394740 -20136 394796 -20080
rect 394882 -20136 394938 -20080
rect 394740 -20278 394796 -20222
rect 394882 -20278 394938 -20222
rect 394740 -20420 394796 -20364
rect 394882 -20420 394938 -20364
rect 394740 -20562 394796 -20506
rect 394882 -20562 394938 -20506
rect 394740 -20704 394796 -20648
rect 394882 -20704 394938 -20648
rect 394740 -20846 394796 -20790
rect 394882 -20846 394938 -20790
rect 394740 -20988 394796 -20932
rect 394882 -20988 394938 -20932
rect 394740 -21130 394796 -21074
rect 394882 -21130 394938 -21074
rect 394740 -21272 394796 -21216
rect 394882 -21272 394938 -21216
rect 394740 -21414 394796 -21358
rect 394882 -21414 394938 -21358
rect 394740 -21556 394796 -21500
rect 394882 -21556 394938 -21500
rect 394740 -21698 394796 -21642
rect 394882 -21698 394938 -21642
rect 394740 -21840 394796 -21784
rect 394882 -21840 394938 -21784
rect 394740 -21982 394796 -21926
rect 394882 -21982 394938 -21926
rect 394740 -22124 394796 -22068
rect 394882 -22124 394938 -22068
rect 394740 -22266 394796 -22210
rect 394882 -22266 394938 -22210
rect 394740 -22408 394796 -22352
rect 394882 -22408 394938 -22352
rect 394740 -22550 394796 -22494
rect 394882 -22550 394938 -22494
rect 394740 -22692 394796 -22636
rect 394882 -22692 394938 -22636
rect 394740 -22834 394796 -22778
rect 394882 -22834 394938 -22778
rect 394740 -22976 394796 -22920
rect 394882 -22976 394938 -22920
rect 394740 -23118 394796 -23062
rect 394882 -23118 394938 -23062
rect 394740 -23260 394796 -23204
rect 394882 -23260 394938 -23204
rect 394740 -23402 394796 -23346
rect 394882 -23402 394938 -23346
rect 394740 -23544 394796 -23488
rect 394882 -23544 394938 -23488
rect 394740 -23686 394796 -23630
rect 394882 -23686 394938 -23630
rect 394740 -23828 394796 -23772
rect 394882 -23828 394938 -23772
rect 394740 -23970 394796 -23914
rect 394882 -23970 394938 -23914
rect 394740 -24112 394796 -24056
rect 394882 -24112 394938 -24056
rect 394740 -24254 394796 -24198
rect 394882 -24254 394938 -24198
rect 394740 -24396 394796 -24340
rect 394882 -24396 394938 -24340
rect 394740 -24538 394796 -24482
rect 394882 -24538 394938 -24482
rect 394740 -24680 394796 -24624
rect 394882 -24680 394938 -24624
rect 394740 -24822 394796 -24766
rect 394882 -24822 394938 -24766
rect 394740 -24964 394796 -24908
rect 394882 -24964 394938 -24908
rect 394740 -25106 394796 -25050
rect 394882 -25106 394938 -25050
rect 394740 -25248 394796 -25192
rect 394882 -25248 394938 -25192
rect 394740 -25390 394796 -25334
rect 394882 -25390 394938 -25334
rect 394740 -25532 394796 -25476
rect 394882 -25532 394938 -25476
rect 395142 -18006 395198 -17950
rect 395284 -18006 395340 -17950
rect 395142 -18148 395198 -18092
rect 395284 -18148 395340 -18092
rect 395142 -18290 395198 -18234
rect 395284 -18290 395340 -18234
rect 395142 -18432 395198 -18376
rect 395284 -18432 395340 -18376
rect 395142 -18574 395198 -18518
rect 395284 -18574 395340 -18518
rect 395142 -18716 395198 -18660
rect 395284 -18716 395340 -18660
rect 395142 -18858 395198 -18802
rect 395284 -18858 395340 -18802
rect 395142 -19000 395198 -18944
rect 395284 -19000 395340 -18944
rect 395142 -19142 395198 -19086
rect 395284 -19142 395340 -19086
rect 395142 -19284 395198 -19228
rect 395284 -19284 395340 -19228
rect 395142 -19426 395198 -19370
rect 395284 -19426 395340 -19370
rect 395142 -19568 395198 -19512
rect 395284 -19568 395340 -19512
rect 395142 -19710 395198 -19654
rect 395284 -19710 395340 -19654
rect 395142 -19852 395198 -19796
rect 395284 -19852 395340 -19796
rect 395142 -19994 395198 -19938
rect 395284 -19994 395340 -19938
rect 395142 -20136 395198 -20080
rect 395284 -20136 395340 -20080
rect 395142 -20278 395198 -20222
rect 395284 -20278 395340 -20222
rect 395142 -20420 395198 -20364
rect 395284 -20420 395340 -20364
rect 395142 -20562 395198 -20506
rect 395284 -20562 395340 -20506
rect 395142 -20704 395198 -20648
rect 395284 -20704 395340 -20648
rect 395142 -20846 395198 -20790
rect 395284 -20846 395340 -20790
rect 395142 -20988 395198 -20932
rect 395284 -20988 395340 -20932
rect 395142 -21130 395198 -21074
rect 395284 -21130 395340 -21074
rect 395142 -21272 395198 -21216
rect 395284 -21272 395340 -21216
rect 395142 -21414 395198 -21358
rect 395284 -21414 395340 -21358
rect 395142 -21556 395198 -21500
rect 395284 -21556 395340 -21500
rect 395142 -21698 395198 -21642
rect 395284 -21698 395340 -21642
rect 395142 -21840 395198 -21784
rect 395284 -21840 395340 -21784
rect 395142 -21982 395198 -21926
rect 395284 -21982 395340 -21926
rect 395142 -22124 395198 -22068
rect 395284 -22124 395340 -22068
rect 395142 -22266 395198 -22210
rect 395284 -22266 395340 -22210
rect 395142 -22408 395198 -22352
rect 395284 -22408 395340 -22352
rect 395142 -22550 395198 -22494
rect 395284 -22550 395340 -22494
rect 395142 -22692 395198 -22636
rect 395284 -22692 395340 -22636
rect 395142 -22834 395198 -22778
rect 395284 -22834 395340 -22778
rect 395142 -22976 395198 -22920
rect 395284 -22976 395340 -22920
rect 395142 -23118 395198 -23062
rect 395284 -23118 395340 -23062
rect 395142 -23260 395198 -23204
rect 395284 -23260 395340 -23204
rect 395142 -23402 395198 -23346
rect 395284 -23402 395340 -23346
rect 395142 -23544 395198 -23488
rect 395284 -23544 395340 -23488
rect 395142 -23686 395198 -23630
rect 395284 -23686 395340 -23630
rect 395142 -23828 395198 -23772
rect 395284 -23828 395340 -23772
rect 395142 -23970 395198 -23914
rect 395284 -23970 395340 -23914
rect 395142 -24112 395198 -24056
rect 395284 -24112 395340 -24056
rect 395142 -24254 395198 -24198
rect 395284 -24254 395340 -24198
rect 395142 -24396 395198 -24340
rect 395284 -24396 395340 -24340
rect 395142 -24538 395198 -24482
rect 395284 -24538 395340 -24482
rect 395142 -24680 395198 -24624
rect 395284 -24680 395340 -24624
rect 395142 -24822 395198 -24766
rect 395284 -24822 395340 -24766
rect 395142 -24964 395198 -24908
rect 395284 -24964 395340 -24908
rect 395142 -25106 395198 -25050
rect 395284 -25106 395340 -25050
rect 395142 -25248 395198 -25192
rect 395284 -25248 395340 -25192
rect 395142 -25390 395198 -25334
rect 395284 -25390 395340 -25334
rect 395142 -25532 395198 -25476
rect 395284 -25532 395340 -25476
rect 395545 -18006 395601 -17950
rect 395687 -18006 395743 -17950
rect 395545 -18148 395601 -18092
rect 395687 -18148 395743 -18092
rect 395545 -18290 395601 -18234
rect 395687 -18290 395743 -18234
rect 395545 -18432 395601 -18376
rect 395687 -18432 395743 -18376
rect 395545 -18574 395601 -18518
rect 395687 -18574 395743 -18518
rect 395545 -18716 395601 -18660
rect 395687 -18716 395743 -18660
rect 395545 -18858 395601 -18802
rect 395687 -18858 395743 -18802
rect 395545 -19000 395601 -18944
rect 395687 -19000 395743 -18944
rect 395545 -19142 395601 -19086
rect 395687 -19142 395743 -19086
rect 395545 -19284 395601 -19228
rect 395687 -19284 395743 -19228
rect 395545 -19426 395601 -19370
rect 395687 -19426 395743 -19370
rect 395545 -19568 395601 -19512
rect 395687 -19568 395743 -19512
rect 395545 -19710 395601 -19654
rect 395687 -19710 395743 -19654
rect 395545 -19852 395601 -19796
rect 395687 -19852 395743 -19796
rect 395545 -19994 395601 -19938
rect 395687 -19994 395743 -19938
rect 395545 -20136 395601 -20080
rect 395687 -20136 395743 -20080
rect 395545 -20278 395601 -20222
rect 395687 -20278 395743 -20222
rect 395545 -20420 395601 -20364
rect 395687 -20420 395743 -20364
rect 395545 -20562 395601 -20506
rect 395687 -20562 395743 -20506
rect 395545 -20704 395601 -20648
rect 395687 -20704 395743 -20648
rect 395545 -20846 395601 -20790
rect 395687 -20846 395743 -20790
rect 395545 -20988 395601 -20932
rect 395687 -20988 395743 -20932
rect 395545 -21130 395601 -21074
rect 395687 -21130 395743 -21074
rect 395545 -21272 395601 -21216
rect 395687 -21272 395743 -21216
rect 395545 -21414 395601 -21358
rect 395687 -21414 395743 -21358
rect 395545 -21556 395601 -21500
rect 395687 -21556 395743 -21500
rect 395545 -21698 395601 -21642
rect 395687 -21698 395743 -21642
rect 395545 -21840 395601 -21784
rect 395687 -21840 395743 -21784
rect 395545 -21982 395601 -21926
rect 395687 -21982 395743 -21926
rect 395545 -22124 395601 -22068
rect 395687 -22124 395743 -22068
rect 395545 -22266 395601 -22210
rect 395687 -22266 395743 -22210
rect 395545 -22408 395601 -22352
rect 395687 -22408 395743 -22352
rect 395545 -22550 395601 -22494
rect 395687 -22550 395743 -22494
rect 395545 -22692 395601 -22636
rect 395687 -22692 395743 -22636
rect 395545 -22834 395601 -22778
rect 395687 -22834 395743 -22778
rect 395545 -22976 395601 -22920
rect 395687 -22976 395743 -22920
rect 395545 -23118 395601 -23062
rect 395687 -23118 395743 -23062
rect 395545 -23260 395601 -23204
rect 395687 -23260 395743 -23204
rect 395545 -23402 395601 -23346
rect 395687 -23402 395743 -23346
rect 395545 -23544 395601 -23488
rect 395687 -23544 395743 -23488
rect 395545 -23686 395601 -23630
rect 395687 -23686 395743 -23630
rect 395545 -23828 395601 -23772
rect 395687 -23828 395743 -23772
rect 395545 -23970 395601 -23914
rect 395687 -23970 395743 -23914
rect 395545 -24112 395601 -24056
rect 395687 -24112 395743 -24056
rect 395545 -24254 395601 -24198
rect 395687 -24254 395743 -24198
rect 395545 -24396 395601 -24340
rect 395687 -24396 395743 -24340
rect 395545 -24538 395601 -24482
rect 395687 -24538 395743 -24482
rect 395545 -24680 395601 -24624
rect 395687 -24680 395743 -24624
rect 395545 -24822 395601 -24766
rect 395687 -24822 395743 -24766
rect 395545 -24964 395601 -24908
rect 395687 -24964 395743 -24908
rect 395545 -25106 395601 -25050
rect 395687 -25106 395743 -25050
rect 395545 -25248 395601 -25192
rect 395687 -25248 395743 -25192
rect 395545 -25390 395601 -25334
rect 395687 -25390 395743 -25334
rect 395545 -25532 395601 -25476
rect 395687 -25532 395743 -25476
rect 395941 -18006 395997 -17950
rect 396083 -18006 396139 -17950
rect 395941 -18148 395997 -18092
rect 396083 -18148 396139 -18092
rect 395941 -18290 395997 -18234
rect 396083 -18290 396139 -18234
rect 395941 -18432 395997 -18376
rect 396083 -18432 396139 -18376
rect 395941 -18574 395997 -18518
rect 396083 -18574 396139 -18518
rect 395941 -18716 395997 -18660
rect 396083 -18716 396139 -18660
rect 395941 -18858 395997 -18802
rect 396083 -18858 396139 -18802
rect 395941 -19000 395997 -18944
rect 396083 -19000 396139 -18944
rect 395941 -19142 395997 -19086
rect 396083 -19142 396139 -19086
rect 395941 -19284 395997 -19228
rect 396083 -19284 396139 -19228
rect 395941 -19426 395997 -19370
rect 396083 -19426 396139 -19370
rect 395941 -19568 395997 -19512
rect 396083 -19568 396139 -19512
rect 395941 -19710 395997 -19654
rect 396083 -19710 396139 -19654
rect 395941 -19852 395997 -19796
rect 396083 -19852 396139 -19796
rect 395941 -19994 395997 -19938
rect 396083 -19994 396139 -19938
rect 395941 -20136 395997 -20080
rect 396083 -20136 396139 -20080
rect 395941 -20278 395997 -20222
rect 396083 -20278 396139 -20222
rect 395941 -20420 395997 -20364
rect 396083 -20420 396139 -20364
rect 395941 -20562 395997 -20506
rect 396083 -20562 396139 -20506
rect 395941 -20704 395997 -20648
rect 396083 -20704 396139 -20648
rect 395941 -20846 395997 -20790
rect 396083 -20846 396139 -20790
rect 395941 -20988 395997 -20932
rect 396083 -20988 396139 -20932
rect 395941 -21130 395997 -21074
rect 396083 -21130 396139 -21074
rect 395941 -21272 395997 -21216
rect 396083 -21272 396139 -21216
rect 395941 -21414 395997 -21358
rect 396083 -21414 396139 -21358
rect 395941 -21556 395997 -21500
rect 396083 -21556 396139 -21500
rect 395941 -21698 395997 -21642
rect 396083 -21698 396139 -21642
rect 395941 -21840 395997 -21784
rect 396083 -21840 396139 -21784
rect 395941 -21982 395997 -21926
rect 396083 -21982 396139 -21926
rect 395941 -22124 395997 -22068
rect 396083 -22124 396139 -22068
rect 395941 -22266 395997 -22210
rect 396083 -22266 396139 -22210
rect 395941 -22408 395997 -22352
rect 396083 -22408 396139 -22352
rect 395941 -22550 395997 -22494
rect 396083 -22550 396139 -22494
rect 395941 -22692 395997 -22636
rect 396083 -22692 396139 -22636
rect 395941 -22834 395997 -22778
rect 396083 -22834 396139 -22778
rect 395941 -22976 395997 -22920
rect 396083 -22976 396139 -22920
rect 395941 -23118 395997 -23062
rect 396083 -23118 396139 -23062
rect 395941 -23260 395997 -23204
rect 396083 -23260 396139 -23204
rect 395941 -23402 395997 -23346
rect 396083 -23402 396139 -23346
rect 395941 -23544 395997 -23488
rect 396083 -23544 396139 -23488
rect 395941 -23686 395997 -23630
rect 396083 -23686 396139 -23630
rect 395941 -23828 395997 -23772
rect 396083 -23828 396139 -23772
rect 395941 -23970 395997 -23914
rect 396083 -23970 396139 -23914
rect 395941 -24112 395997 -24056
rect 396083 -24112 396139 -24056
rect 395941 -24254 395997 -24198
rect 396083 -24254 396139 -24198
rect 395941 -24396 395997 -24340
rect 396083 -24396 396139 -24340
rect 395941 -24538 395997 -24482
rect 396083 -24538 396139 -24482
rect 395941 -24680 395997 -24624
rect 396083 -24680 396139 -24624
rect 395941 -24822 395997 -24766
rect 396083 -24822 396139 -24766
rect 395941 -24964 395997 -24908
rect 396083 -24964 396139 -24908
rect 395941 -25106 395997 -25050
rect 396083 -25106 396139 -25050
rect 395941 -25248 395997 -25192
rect 396083 -25248 396139 -25192
rect 395941 -25390 395997 -25334
rect 396083 -25390 396139 -25334
rect 395941 -25532 395997 -25476
rect 396083 -25532 396139 -25476
rect 396526 -17914 396582 -17858
rect 396650 -17914 396706 -17858
rect 396774 -17914 396830 -17858
rect 396898 -17914 396954 -17858
rect 397022 -17914 397078 -17858
rect 396526 -18038 396582 -17982
rect 396650 -18038 396706 -17982
rect 396774 -18038 396830 -17982
rect 396898 -18038 396954 -17982
rect 397022 -18038 397078 -17982
rect 396526 -18162 396582 -18106
rect 396650 -18162 396706 -18106
rect 396774 -18162 396830 -18106
rect 396898 -18162 396954 -18106
rect 397022 -18162 397078 -18106
rect 396526 -18286 396582 -18230
rect 396650 -18286 396706 -18230
rect 396774 -18286 396830 -18230
rect 396898 -18286 396954 -18230
rect 397022 -18286 397078 -18230
rect 396526 -18410 396582 -18354
rect 396650 -18410 396706 -18354
rect 396774 -18410 396830 -18354
rect 396898 -18410 396954 -18354
rect 397022 -18410 397078 -18354
rect 396526 -18534 396582 -18478
rect 396650 -18534 396706 -18478
rect 396774 -18534 396830 -18478
rect 396898 -18534 396954 -18478
rect 397022 -18534 397078 -18478
rect 396526 -18658 396582 -18602
rect 396650 -18658 396706 -18602
rect 396774 -18658 396830 -18602
rect 396898 -18658 396954 -18602
rect 397022 -18658 397078 -18602
rect 396526 -18782 396582 -18726
rect 396650 -18782 396706 -18726
rect 396774 -18782 396830 -18726
rect 396898 -18782 396954 -18726
rect 397022 -18782 397078 -18726
rect 396526 -18906 396582 -18850
rect 396650 -18906 396706 -18850
rect 396774 -18906 396830 -18850
rect 396898 -18906 396954 -18850
rect 397022 -18906 397078 -18850
rect 396526 -19030 396582 -18974
rect 396650 -19030 396706 -18974
rect 396774 -19030 396830 -18974
rect 396898 -19030 396954 -18974
rect 397022 -19030 397078 -18974
rect 396526 -19154 396582 -19098
rect 396650 -19154 396706 -19098
rect 396774 -19154 396830 -19098
rect 396898 -19154 396954 -19098
rect 397022 -19154 397078 -19098
rect 396526 -19278 396582 -19222
rect 396650 -19278 396706 -19222
rect 396774 -19278 396830 -19222
rect 396898 -19278 396954 -19222
rect 397022 -19278 397078 -19222
rect 396526 -19402 396582 -19346
rect 396650 -19402 396706 -19346
rect 396774 -19402 396830 -19346
rect 396898 -19402 396954 -19346
rect 397022 -19402 397078 -19346
rect 396526 -19526 396582 -19470
rect 396650 -19526 396706 -19470
rect 396774 -19526 396830 -19470
rect 396898 -19526 396954 -19470
rect 397022 -19526 397078 -19470
rect 396526 -19650 396582 -19594
rect 396650 -19650 396706 -19594
rect 396774 -19650 396830 -19594
rect 396898 -19650 396954 -19594
rect 397022 -19650 397078 -19594
rect 396526 -19774 396582 -19718
rect 396650 -19774 396706 -19718
rect 396774 -19774 396830 -19718
rect 396898 -19774 396954 -19718
rect 397022 -19774 397078 -19718
rect 396526 -19898 396582 -19842
rect 396650 -19898 396706 -19842
rect 396774 -19898 396830 -19842
rect 396898 -19898 396954 -19842
rect 397022 -19898 397078 -19842
rect 396526 -20022 396582 -19966
rect 396650 -20022 396706 -19966
rect 396774 -20022 396830 -19966
rect 396898 -20022 396954 -19966
rect 397022 -20022 397078 -19966
rect 396526 -20146 396582 -20090
rect 396650 -20146 396706 -20090
rect 396774 -20146 396830 -20090
rect 396898 -20146 396954 -20090
rect 397022 -20146 397078 -20090
rect 396526 -20270 396582 -20214
rect 396650 -20270 396706 -20214
rect 396774 -20270 396830 -20214
rect 396898 -20270 396954 -20214
rect 397022 -20270 397078 -20214
rect 396526 -20394 396582 -20338
rect 396650 -20394 396706 -20338
rect 396774 -20394 396830 -20338
rect 396898 -20394 396954 -20338
rect 397022 -20394 397078 -20338
rect 396526 -20518 396582 -20462
rect 396650 -20518 396706 -20462
rect 396774 -20518 396830 -20462
rect 396898 -20518 396954 -20462
rect 397022 -20518 397078 -20462
rect 396526 -20642 396582 -20586
rect 396650 -20642 396706 -20586
rect 396774 -20642 396830 -20586
rect 396898 -20642 396954 -20586
rect 397022 -20642 397078 -20586
rect 396526 -20766 396582 -20710
rect 396650 -20766 396706 -20710
rect 396774 -20766 396830 -20710
rect 396898 -20766 396954 -20710
rect 397022 -20766 397078 -20710
rect 396526 -20890 396582 -20834
rect 396650 -20890 396706 -20834
rect 396774 -20890 396830 -20834
rect 396898 -20890 396954 -20834
rect 397022 -20890 397078 -20834
rect 396526 -21014 396582 -20958
rect 396650 -21014 396706 -20958
rect 396774 -21014 396830 -20958
rect 396898 -21014 396954 -20958
rect 397022 -21014 397078 -20958
rect 396526 -21138 396582 -21082
rect 396650 -21138 396706 -21082
rect 396774 -21138 396830 -21082
rect 396898 -21138 396954 -21082
rect 397022 -21138 397078 -21082
rect 396526 -21262 396582 -21206
rect 396650 -21262 396706 -21206
rect 396774 -21262 396830 -21206
rect 396898 -21262 396954 -21206
rect 397022 -21262 397078 -21206
rect 396526 -21386 396582 -21330
rect 396650 -21386 396706 -21330
rect 396774 -21386 396830 -21330
rect 396898 -21386 396954 -21330
rect 397022 -21386 397078 -21330
rect 396526 -21510 396582 -21454
rect 396650 -21510 396706 -21454
rect 396774 -21510 396830 -21454
rect 396898 -21510 396954 -21454
rect 397022 -21510 397078 -21454
rect 396526 -21634 396582 -21578
rect 396650 -21634 396706 -21578
rect 396774 -21634 396830 -21578
rect 396898 -21634 396954 -21578
rect 397022 -21634 397078 -21578
rect 396526 -21758 396582 -21702
rect 396650 -21758 396706 -21702
rect 396774 -21758 396830 -21702
rect 396898 -21758 396954 -21702
rect 397022 -21758 397078 -21702
rect 396526 -21882 396582 -21826
rect 396650 -21882 396706 -21826
rect 396774 -21882 396830 -21826
rect 396898 -21882 396954 -21826
rect 397022 -21882 397078 -21826
rect 396526 -22006 396582 -21950
rect 396650 -22006 396706 -21950
rect 396774 -22006 396830 -21950
rect 396898 -22006 396954 -21950
rect 397022 -22006 397078 -21950
rect 396526 -22130 396582 -22074
rect 396650 -22130 396706 -22074
rect 396774 -22130 396830 -22074
rect 396898 -22130 396954 -22074
rect 397022 -22130 397078 -22074
rect 396526 -22254 396582 -22198
rect 396650 -22254 396706 -22198
rect 396774 -22254 396830 -22198
rect 396898 -22254 396954 -22198
rect 397022 -22254 397078 -22198
rect 396526 -22378 396582 -22322
rect 396650 -22378 396706 -22322
rect 396774 -22378 396830 -22322
rect 396898 -22378 396954 -22322
rect 397022 -22378 397078 -22322
rect 396526 -22502 396582 -22446
rect 396650 -22502 396706 -22446
rect 396774 -22502 396830 -22446
rect 396898 -22502 396954 -22446
rect 397022 -22502 397078 -22446
rect 396526 -22626 396582 -22570
rect 396650 -22626 396706 -22570
rect 396774 -22626 396830 -22570
rect 396898 -22626 396954 -22570
rect 397022 -22626 397078 -22570
rect 396526 -22750 396582 -22694
rect 396650 -22750 396706 -22694
rect 396774 -22750 396830 -22694
rect 396898 -22750 396954 -22694
rect 397022 -22750 397078 -22694
rect 396526 -22874 396582 -22818
rect 396650 -22874 396706 -22818
rect 396774 -22874 396830 -22818
rect 396898 -22874 396954 -22818
rect 397022 -22874 397078 -22818
rect 396526 -22998 396582 -22942
rect 396650 -22998 396706 -22942
rect 396774 -22998 396830 -22942
rect 396898 -22998 396954 -22942
rect 397022 -22998 397078 -22942
rect 396526 -23122 396582 -23066
rect 396650 -23122 396706 -23066
rect 396774 -23122 396830 -23066
rect 396898 -23122 396954 -23066
rect 397022 -23122 397078 -23066
rect 396526 -23246 396582 -23190
rect 396650 -23246 396706 -23190
rect 396774 -23246 396830 -23190
rect 396898 -23246 396954 -23190
rect 397022 -23246 397078 -23190
rect 396526 -23370 396582 -23314
rect 396650 -23370 396706 -23314
rect 396774 -23370 396830 -23314
rect 396898 -23370 396954 -23314
rect 397022 -23370 397078 -23314
rect 396526 -23494 396582 -23438
rect 396650 -23494 396706 -23438
rect 396774 -23494 396830 -23438
rect 396898 -23494 396954 -23438
rect 397022 -23494 397078 -23438
rect 396526 -23618 396582 -23562
rect 396650 -23618 396706 -23562
rect 396774 -23618 396830 -23562
rect 396898 -23618 396954 -23562
rect 397022 -23618 397078 -23562
rect 396526 -23742 396582 -23686
rect 396650 -23742 396706 -23686
rect 396774 -23742 396830 -23686
rect 396898 -23742 396954 -23686
rect 397022 -23742 397078 -23686
rect 396526 -23866 396582 -23810
rect 396650 -23866 396706 -23810
rect 396774 -23866 396830 -23810
rect 396898 -23866 396954 -23810
rect 397022 -23866 397078 -23810
rect 396526 -23990 396582 -23934
rect 396650 -23990 396706 -23934
rect 396774 -23990 396830 -23934
rect 396898 -23990 396954 -23934
rect 397022 -23990 397078 -23934
rect 396526 -24114 396582 -24058
rect 396650 -24114 396706 -24058
rect 396774 -24114 396830 -24058
rect 396898 -24114 396954 -24058
rect 397022 -24114 397078 -24058
rect 396526 -24238 396582 -24182
rect 396650 -24238 396706 -24182
rect 396774 -24238 396830 -24182
rect 396898 -24238 396954 -24182
rect 397022 -24238 397078 -24182
rect 396526 -24362 396582 -24306
rect 396650 -24362 396706 -24306
rect 396774 -24362 396830 -24306
rect 396898 -24362 396954 -24306
rect 397022 -24362 397078 -24306
rect 396526 -24486 396582 -24430
rect 396650 -24486 396706 -24430
rect 396774 -24486 396830 -24430
rect 396898 -24486 396954 -24430
rect 397022 -24486 397078 -24430
rect 396526 -24610 396582 -24554
rect 396650 -24610 396706 -24554
rect 396774 -24610 396830 -24554
rect 396898 -24610 396954 -24554
rect 397022 -24610 397078 -24554
rect 396526 -24734 396582 -24678
rect 396650 -24734 396706 -24678
rect 396774 -24734 396830 -24678
rect 396898 -24734 396954 -24678
rect 397022 -24734 397078 -24678
rect 396526 -24858 396582 -24802
rect 396650 -24858 396706 -24802
rect 396774 -24858 396830 -24802
rect 396898 -24858 396954 -24802
rect 397022 -24858 397078 -24802
rect 396526 -24982 396582 -24926
rect 396650 -24982 396706 -24926
rect 396774 -24982 396830 -24926
rect 396898 -24982 396954 -24926
rect 397022 -24982 397078 -24926
rect 396526 -25106 396582 -25050
rect 396650 -25106 396706 -25050
rect 396774 -25106 396830 -25050
rect 396898 -25106 396954 -25050
rect 397022 -25106 397078 -25050
rect 396526 -25230 396582 -25174
rect 396650 -25230 396706 -25174
rect 396774 -25230 396830 -25174
rect 396898 -25230 396954 -25174
rect 397022 -25230 397078 -25174
rect 396526 -25354 396582 -25298
rect 396650 -25354 396706 -25298
rect 396774 -25354 396830 -25298
rect 396898 -25354 396954 -25298
rect 397022 -25354 397078 -25298
rect 396526 -25478 396582 -25422
rect 396650 -25478 396706 -25422
rect 396774 -25478 396830 -25422
rect 396898 -25478 396954 -25422
rect 397022 -25478 397078 -25422
rect 388146 -25777 388202 -25721
rect 388270 -25777 388326 -25721
rect 388394 -25777 388450 -25721
rect 388518 -25777 388574 -25721
rect 388642 -25777 388698 -25721
rect 388766 -25777 388822 -25721
rect 388890 -25777 388946 -25721
rect 389014 -25777 389070 -25721
rect 389138 -25777 389194 -25721
rect 389262 -25777 389318 -25721
rect 389386 -25777 389442 -25721
rect 389510 -25777 389566 -25721
rect 389634 -25777 389690 -25721
rect 389758 -25777 389814 -25721
rect 389882 -25777 389938 -25721
rect 390006 -25777 390062 -25721
rect 390130 -25777 390186 -25721
rect 390254 -25777 390310 -25721
rect 390378 -25777 390434 -25721
rect 390502 -25777 390558 -25721
rect 390626 -25777 390682 -25721
rect 390750 -25777 390806 -25721
rect 390874 -25777 390930 -25721
rect 390998 -25777 391054 -25721
rect 391122 -25777 391178 -25721
rect 391246 -25777 391302 -25721
rect 391370 -25777 391426 -25721
rect 391494 -25777 391550 -25721
rect 391618 -25777 391674 -25721
rect 391742 -25777 391798 -25721
rect 391866 -25777 391922 -25721
rect 391990 -25777 392046 -25721
rect 392114 -25777 392170 -25721
rect 392238 -25777 392294 -25721
rect 392362 -25777 392418 -25721
rect 392486 -25777 392542 -25721
rect 392610 -25777 392666 -25721
rect 392734 -25777 392790 -25721
rect 392858 -25777 392914 -25721
rect 392982 -25777 393038 -25721
rect 393106 -25777 393162 -25721
rect 393230 -25777 393286 -25721
rect 393354 -25777 393410 -25721
rect 393478 -25777 393534 -25721
rect 393602 -25777 393658 -25721
rect 393726 -25777 393782 -25721
rect 393850 -25777 393906 -25721
rect 393974 -25777 394030 -25721
rect 394098 -25777 394154 -25721
rect 394222 -25777 394278 -25721
rect 394346 -25777 394402 -25721
rect 394470 -25777 394526 -25721
rect 394594 -25777 394650 -25721
rect 394718 -25777 394774 -25721
rect 394842 -25777 394898 -25721
rect 394966 -25777 395022 -25721
rect 395090 -25777 395146 -25721
rect 395214 -25777 395270 -25721
rect 395338 -25777 395394 -25721
rect 395462 -25777 395518 -25721
rect 395586 -25777 395642 -25721
rect 395710 -25777 395766 -25721
rect 395898 -25777 395954 -25721
rect 396022 -25777 396078 -25721
rect 396146 -25777 396202 -25721
rect 396270 -25777 396326 -25721
rect 396394 -25777 396450 -25721
rect 396518 -25777 396574 -25721
rect 396642 -25777 396698 -25721
rect 396766 -25777 396822 -25721
rect 396890 -25777 396946 -25721
rect 397014 -25777 397070 -25721
rect 388146 -25901 388202 -25845
rect 388270 -25901 388326 -25845
rect 388394 -25901 388450 -25845
rect 388518 -25901 388574 -25845
rect 388642 -25901 388698 -25845
rect 388766 -25901 388822 -25845
rect 388890 -25901 388946 -25845
rect 389014 -25901 389070 -25845
rect 389138 -25901 389194 -25845
rect 389262 -25901 389318 -25845
rect 389386 -25901 389442 -25845
rect 389510 -25901 389566 -25845
rect 389634 -25901 389690 -25845
rect 389758 -25901 389814 -25845
rect 389882 -25901 389938 -25845
rect 390006 -25901 390062 -25845
rect 390130 -25901 390186 -25845
rect 390254 -25901 390310 -25845
rect 390378 -25901 390434 -25845
rect 390502 -25901 390558 -25845
rect 390626 -25901 390682 -25845
rect 390750 -25901 390806 -25845
rect 390874 -25901 390930 -25845
rect 390998 -25901 391054 -25845
rect 391122 -25901 391178 -25845
rect 391246 -25901 391302 -25845
rect 391370 -25901 391426 -25845
rect 391494 -25901 391550 -25845
rect 391618 -25901 391674 -25845
rect 391742 -25901 391798 -25845
rect 391866 -25901 391922 -25845
rect 391990 -25901 392046 -25845
rect 392114 -25901 392170 -25845
rect 392238 -25901 392294 -25845
rect 392362 -25901 392418 -25845
rect 392486 -25901 392542 -25845
rect 392610 -25901 392666 -25845
rect 392734 -25901 392790 -25845
rect 392858 -25901 392914 -25845
rect 392982 -25901 393038 -25845
rect 393106 -25901 393162 -25845
rect 393230 -25901 393286 -25845
rect 393354 -25901 393410 -25845
rect 393478 -25901 393534 -25845
rect 393602 -25901 393658 -25845
rect 393726 -25901 393782 -25845
rect 393850 -25901 393906 -25845
rect 393974 -25901 394030 -25845
rect 394098 -25901 394154 -25845
rect 394222 -25901 394278 -25845
rect 394346 -25901 394402 -25845
rect 394470 -25901 394526 -25845
rect 394594 -25901 394650 -25845
rect 394718 -25901 394774 -25845
rect 394842 -25901 394898 -25845
rect 394966 -25901 395022 -25845
rect 395090 -25901 395146 -25845
rect 395214 -25901 395270 -25845
rect 395338 -25901 395394 -25845
rect 395462 -25901 395518 -25845
rect 395586 -25901 395642 -25845
rect 395710 -25901 395766 -25845
rect 395898 -25901 395954 -25845
rect 396022 -25901 396078 -25845
rect 396146 -25901 396202 -25845
rect 396270 -25901 396326 -25845
rect 396394 -25901 396450 -25845
rect 396518 -25901 396574 -25845
rect 396642 -25901 396698 -25845
rect 396766 -25901 396822 -25845
rect 396890 -25901 396946 -25845
rect 397014 -25901 397070 -25845
rect 388146 -26025 388202 -25969
rect 388270 -26025 388326 -25969
rect 388394 -26025 388450 -25969
rect 388518 -26025 388574 -25969
rect 388642 -26025 388698 -25969
rect 388766 -26025 388822 -25969
rect 388890 -26025 388946 -25969
rect 389014 -26025 389070 -25969
rect 389138 -26025 389194 -25969
rect 389262 -26025 389318 -25969
rect 389386 -26025 389442 -25969
rect 389510 -26025 389566 -25969
rect 389634 -26025 389690 -25969
rect 389758 -26025 389814 -25969
rect 389882 -26025 389938 -25969
rect 390006 -26025 390062 -25969
rect 390130 -26025 390186 -25969
rect 390254 -26025 390310 -25969
rect 390378 -26025 390434 -25969
rect 390502 -26025 390558 -25969
rect 390626 -26025 390682 -25969
rect 390750 -26025 390806 -25969
rect 390874 -26025 390930 -25969
rect 390998 -26025 391054 -25969
rect 391122 -26025 391178 -25969
rect 391246 -26025 391302 -25969
rect 391370 -26025 391426 -25969
rect 391494 -26025 391550 -25969
rect 391618 -26025 391674 -25969
rect 391742 -26025 391798 -25969
rect 391866 -26025 391922 -25969
rect 391990 -26025 392046 -25969
rect 392114 -26025 392170 -25969
rect 392238 -26025 392294 -25969
rect 392362 -26025 392418 -25969
rect 392486 -26025 392542 -25969
rect 392610 -26025 392666 -25969
rect 392734 -26025 392790 -25969
rect 392858 -26025 392914 -25969
rect 392982 -26025 393038 -25969
rect 393106 -26025 393162 -25969
rect 393230 -26025 393286 -25969
rect 393354 -26025 393410 -25969
rect 393478 -26025 393534 -25969
rect 393602 -26025 393658 -25969
rect 393726 -26025 393782 -25969
rect 393850 -26025 393906 -25969
rect 393974 -26025 394030 -25969
rect 394098 -26025 394154 -25969
rect 394222 -26025 394278 -25969
rect 394346 -26025 394402 -25969
rect 394470 -26025 394526 -25969
rect 394594 -26025 394650 -25969
rect 394718 -26025 394774 -25969
rect 394842 -26025 394898 -25969
rect 394966 -26025 395022 -25969
rect 395090 -26025 395146 -25969
rect 395214 -26025 395270 -25969
rect 395338 -26025 395394 -25969
rect 395462 -26025 395518 -25969
rect 395586 -26025 395642 -25969
rect 395710 -26025 395766 -25969
rect 395898 -26025 395954 -25969
rect 396022 -26025 396078 -25969
rect 396146 -26025 396202 -25969
rect 396270 -26025 396326 -25969
rect 396394 -26025 396450 -25969
rect 396518 -26025 396574 -25969
rect 396642 -26025 396698 -25969
rect 396766 -26025 396822 -25969
rect 396890 -26025 396946 -25969
rect 397014 -26025 397070 -25969
rect 388146 -26149 388202 -26093
rect 388270 -26149 388326 -26093
rect 388394 -26149 388450 -26093
rect 388518 -26149 388574 -26093
rect 388642 -26149 388698 -26093
rect 388766 -26149 388822 -26093
rect 388890 -26149 388946 -26093
rect 389014 -26149 389070 -26093
rect 389138 -26149 389194 -26093
rect 389262 -26149 389318 -26093
rect 389386 -26149 389442 -26093
rect 389510 -26149 389566 -26093
rect 389634 -26149 389690 -26093
rect 389758 -26149 389814 -26093
rect 389882 -26149 389938 -26093
rect 390006 -26149 390062 -26093
rect 390130 -26149 390186 -26093
rect 390254 -26149 390310 -26093
rect 390378 -26149 390434 -26093
rect 390502 -26149 390558 -26093
rect 390626 -26149 390682 -26093
rect 390750 -26149 390806 -26093
rect 390874 -26149 390930 -26093
rect 390998 -26149 391054 -26093
rect 391122 -26149 391178 -26093
rect 391246 -26149 391302 -26093
rect 391370 -26149 391426 -26093
rect 391494 -26149 391550 -26093
rect 391618 -26149 391674 -26093
rect 391742 -26149 391798 -26093
rect 391866 -26149 391922 -26093
rect 391990 -26149 392046 -26093
rect 392114 -26149 392170 -26093
rect 392238 -26149 392294 -26093
rect 392362 -26149 392418 -26093
rect 392486 -26149 392542 -26093
rect 392610 -26149 392666 -26093
rect 392734 -26149 392790 -26093
rect 392858 -26149 392914 -26093
rect 392982 -26149 393038 -26093
rect 393106 -26149 393162 -26093
rect 393230 -26149 393286 -26093
rect 393354 -26149 393410 -26093
rect 393478 -26149 393534 -26093
rect 393602 -26149 393658 -26093
rect 393726 -26149 393782 -26093
rect 393850 -26149 393906 -26093
rect 393974 -26149 394030 -26093
rect 394098 -26149 394154 -26093
rect 394222 -26149 394278 -26093
rect 394346 -26149 394402 -26093
rect 394470 -26149 394526 -26093
rect 394594 -26149 394650 -26093
rect 394718 -26149 394774 -26093
rect 394842 -26149 394898 -26093
rect 394966 -26149 395022 -26093
rect 395090 -26149 395146 -26093
rect 395214 -26149 395270 -26093
rect 395338 -26149 395394 -26093
rect 395462 -26149 395518 -26093
rect 395586 -26149 395642 -26093
rect 395710 -26149 395766 -26093
rect 395898 -26149 395954 -26093
rect 396022 -26149 396078 -26093
rect 396146 -26149 396202 -26093
rect 396270 -26149 396326 -26093
rect 396394 -26149 396450 -26093
rect 396518 -26149 396574 -26093
rect 396642 -26149 396698 -26093
rect 396766 -26149 396822 -26093
rect 396890 -26149 396946 -26093
rect 397014 -26149 397070 -26093
<< metal3 >>
rect 388000 -17191 397200 -17070
rect 388000 -17247 388146 -17191
rect 388202 -17247 388270 -17191
rect 388326 -17247 388394 -17191
rect 388450 -17247 388518 -17191
rect 388574 -17247 388642 -17191
rect 388698 -17247 388766 -17191
rect 388822 -17247 388890 -17191
rect 388946 -17247 389014 -17191
rect 389070 -17247 389138 -17191
rect 389194 -17247 389262 -17191
rect 389318 -17247 389386 -17191
rect 389442 -17247 389510 -17191
rect 389566 -17247 389634 -17191
rect 389690 -17247 389758 -17191
rect 389814 -17247 389882 -17191
rect 389938 -17247 390006 -17191
rect 390062 -17247 390130 -17191
rect 390186 -17247 390254 -17191
rect 390310 -17247 390378 -17191
rect 390434 -17247 390502 -17191
rect 390558 -17247 390626 -17191
rect 390682 -17247 390750 -17191
rect 390806 -17247 390874 -17191
rect 390930 -17247 390998 -17191
rect 391054 -17247 391122 -17191
rect 391178 -17247 391246 -17191
rect 391302 -17247 391370 -17191
rect 391426 -17247 391494 -17191
rect 391550 -17247 391618 -17191
rect 391674 -17247 391742 -17191
rect 391798 -17247 391866 -17191
rect 391922 -17247 391990 -17191
rect 392046 -17247 392114 -17191
rect 392170 -17247 392238 -17191
rect 392294 -17247 392362 -17191
rect 392418 -17247 392486 -17191
rect 392542 -17247 392610 -17191
rect 392666 -17247 392734 -17191
rect 392790 -17247 392858 -17191
rect 392914 -17247 392982 -17191
rect 393038 -17247 393106 -17191
rect 393162 -17247 393230 -17191
rect 393286 -17247 393354 -17191
rect 393410 -17247 393478 -17191
rect 393534 -17247 393602 -17191
rect 393658 -17247 393726 -17191
rect 393782 -17247 393850 -17191
rect 393906 -17247 393974 -17191
rect 394030 -17247 394098 -17191
rect 394154 -17247 394222 -17191
rect 394278 -17247 394346 -17191
rect 394402 -17247 394470 -17191
rect 394526 -17247 394594 -17191
rect 394650 -17247 394718 -17191
rect 394774 -17247 394842 -17191
rect 394898 -17247 394966 -17191
rect 395022 -17247 395090 -17191
rect 395146 -17247 395214 -17191
rect 395270 -17247 395338 -17191
rect 395394 -17247 395462 -17191
rect 395518 -17247 395586 -17191
rect 395642 -17247 395710 -17191
rect 395766 -17247 395898 -17191
rect 395954 -17247 396022 -17191
rect 396078 -17247 396146 -17191
rect 396202 -17247 396270 -17191
rect 396326 -17247 396394 -17191
rect 396450 -17247 396518 -17191
rect 396574 -17247 396642 -17191
rect 396698 -17247 396766 -17191
rect 396822 -17247 396890 -17191
rect 396946 -17247 397014 -17191
rect 397070 -17247 397200 -17191
rect 388000 -17315 397200 -17247
rect 388000 -17371 388146 -17315
rect 388202 -17371 388270 -17315
rect 388326 -17371 388394 -17315
rect 388450 -17371 388518 -17315
rect 388574 -17371 388642 -17315
rect 388698 -17371 388766 -17315
rect 388822 -17371 388890 -17315
rect 388946 -17371 389014 -17315
rect 389070 -17371 389138 -17315
rect 389194 -17371 389262 -17315
rect 389318 -17371 389386 -17315
rect 389442 -17371 389510 -17315
rect 389566 -17371 389634 -17315
rect 389690 -17371 389758 -17315
rect 389814 -17371 389882 -17315
rect 389938 -17371 390006 -17315
rect 390062 -17371 390130 -17315
rect 390186 -17371 390254 -17315
rect 390310 -17371 390378 -17315
rect 390434 -17371 390502 -17315
rect 390558 -17371 390626 -17315
rect 390682 -17371 390750 -17315
rect 390806 -17371 390874 -17315
rect 390930 -17371 390998 -17315
rect 391054 -17371 391122 -17315
rect 391178 -17371 391246 -17315
rect 391302 -17371 391370 -17315
rect 391426 -17371 391494 -17315
rect 391550 -17371 391618 -17315
rect 391674 -17371 391742 -17315
rect 391798 -17371 391866 -17315
rect 391922 -17371 391990 -17315
rect 392046 -17371 392114 -17315
rect 392170 -17371 392238 -17315
rect 392294 -17371 392362 -17315
rect 392418 -17371 392486 -17315
rect 392542 -17371 392610 -17315
rect 392666 -17371 392734 -17315
rect 392790 -17371 392858 -17315
rect 392914 -17371 392982 -17315
rect 393038 -17371 393106 -17315
rect 393162 -17371 393230 -17315
rect 393286 -17371 393354 -17315
rect 393410 -17371 393478 -17315
rect 393534 -17371 393602 -17315
rect 393658 -17371 393726 -17315
rect 393782 -17371 393850 -17315
rect 393906 -17371 393974 -17315
rect 394030 -17371 394098 -17315
rect 394154 -17371 394222 -17315
rect 394278 -17371 394346 -17315
rect 394402 -17371 394470 -17315
rect 394526 -17371 394594 -17315
rect 394650 -17371 394718 -17315
rect 394774 -17371 394842 -17315
rect 394898 -17371 394966 -17315
rect 395022 -17371 395090 -17315
rect 395146 -17371 395214 -17315
rect 395270 -17371 395338 -17315
rect 395394 -17371 395462 -17315
rect 395518 -17371 395586 -17315
rect 395642 -17371 395710 -17315
rect 395766 -17371 395898 -17315
rect 395954 -17371 396022 -17315
rect 396078 -17371 396146 -17315
rect 396202 -17371 396270 -17315
rect 396326 -17371 396394 -17315
rect 396450 -17371 396518 -17315
rect 396574 -17371 396642 -17315
rect 396698 -17371 396766 -17315
rect 396822 -17371 396890 -17315
rect 396946 -17371 397014 -17315
rect 397070 -17371 397200 -17315
rect 388000 -17439 397200 -17371
rect 388000 -17495 388146 -17439
rect 388202 -17495 388270 -17439
rect 388326 -17495 388394 -17439
rect 388450 -17495 388518 -17439
rect 388574 -17495 388642 -17439
rect 388698 -17495 388766 -17439
rect 388822 -17495 388890 -17439
rect 388946 -17495 389014 -17439
rect 389070 -17495 389138 -17439
rect 389194 -17495 389262 -17439
rect 389318 -17495 389386 -17439
rect 389442 -17495 389510 -17439
rect 389566 -17495 389634 -17439
rect 389690 -17495 389758 -17439
rect 389814 -17495 389882 -17439
rect 389938 -17495 390006 -17439
rect 390062 -17495 390130 -17439
rect 390186 -17495 390254 -17439
rect 390310 -17495 390378 -17439
rect 390434 -17495 390502 -17439
rect 390558 -17495 390626 -17439
rect 390682 -17495 390750 -17439
rect 390806 -17495 390874 -17439
rect 390930 -17495 390998 -17439
rect 391054 -17495 391122 -17439
rect 391178 -17495 391246 -17439
rect 391302 -17495 391370 -17439
rect 391426 -17495 391494 -17439
rect 391550 -17495 391618 -17439
rect 391674 -17495 391742 -17439
rect 391798 -17495 391866 -17439
rect 391922 -17495 391990 -17439
rect 392046 -17495 392114 -17439
rect 392170 -17495 392238 -17439
rect 392294 -17495 392362 -17439
rect 392418 -17495 392486 -17439
rect 392542 -17495 392610 -17439
rect 392666 -17495 392734 -17439
rect 392790 -17495 392858 -17439
rect 392914 -17495 392982 -17439
rect 393038 -17495 393106 -17439
rect 393162 -17495 393230 -17439
rect 393286 -17495 393354 -17439
rect 393410 -17495 393478 -17439
rect 393534 -17495 393602 -17439
rect 393658 -17495 393726 -17439
rect 393782 -17495 393850 -17439
rect 393906 -17495 393974 -17439
rect 394030 -17495 394098 -17439
rect 394154 -17495 394222 -17439
rect 394278 -17495 394346 -17439
rect 394402 -17495 394470 -17439
rect 394526 -17495 394594 -17439
rect 394650 -17495 394718 -17439
rect 394774 -17495 394842 -17439
rect 394898 -17495 394966 -17439
rect 395022 -17495 395090 -17439
rect 395146 -17495 395214 -17439
rect 395270 -17495 395338 -17439
rect 395394 -17495 395462 -17439
rect 395518 -17495 395586 -17439
rect 395642 -17495 395710 -17439
rect 395766 -17495 395898 -17439
rect 395954 -17495 396022 -17439
rect 396078 -17495 396146 -17439
rect 396202 -17495 396270 -17439
rect 396326 -17495 396394 -17439
rect 396450 -17495 396518 -17439
rect 396574 -17495 396642 -17439
rect 396698 -17495 396766 -17439
rect 396822 -17495 396890 -17439
rect 396946 -17495 397014 -17439
rect 397070 -17495 397200 -17439
rect 388000 -17563 397200 -17495
rect 388000 -17619 388146 -17563
rect 388202 -17619 388270 -17563
rect 388326 -17619 388394 -17563
rect 388450 -17619 388518 -17563
rect 388574 -17619 388642 -17563
rect 388698 -17619 388766 -17563
rect 388822 -17619 388890 -17563
rect 388946 -17619 389014 -17563
rect 389070 -17619 389138 -17563
rect 389194 -17619 389262 -17563
rect 389318 -17619 389386 -17563
rect 389442 -17619 389510 -17563
rect 389566 -17619 389634 -17563
rect 389690 -17619 389758 -17563
rect 389814 -17619 389882 -17563
rect 389938 -17619 390006 -17563
rect 390062 -17619 390130 -17563
rect 390186 -17619 390254 -17563
rect 390310 -17619 390378 -17563
rect 390434 -17619 390502 -17563
rect 390558 -17619 390626 -17563
rect 390682 -17619 390750 -17563
rect 390806 -17619 390874 -17563
rect 390930 -17619 390998 -17563
rect 391054 -17619 391122 -17563
rect 391178 -17619 391246 -17563
rect 391302 -17619 391370 -17563
rect 391426 -17619 391494 -17563
rect 391550 -17619 391618 -17563
rect 391674 -17619 391742 -17563
rect 391798 -17619 391866 -17563
rect 391922 -17619 391990 -17563
rect 392046 -17619 392114 -17563
rect 392170 -17619 392238 -17563
rect 392294 -17619 392362 -17563
rect 392418 -17619 392486 -17563
rect 392542 -17619 392610 -17563
rect 392666 -17619 392734 -17563
rect 392790 -17619 392858 -17563
rect 392914 -17619 392982 -17563
rect 393038 -17619 393106 -17563
rect 393162 -17619 393230 -17563
rect 393286 -17619 393354 -17563
rect 393410 -17619 393478 -17563
rect 393534 -17619 393602 -17563
rect 393658 -17619 393726 -17563
rect 393782 -17619 393850 -17563
rect 393906 -17619 393974 -17563
rect 394030 -17619 394098 -17563
rect 394154 -17619 394222 -17563
rect 394278 -17619 394346 -17563
rect 394402 -17619 394470 -17563
rect 394526 -17619 394594 -17563
rect 394650 -17619 394718 -17563
rect 394774 -17619 394842 -17563
rect 394898 -17619 394966 -17563
rect 395022 -17619 395090 -17563
rect 395146 -17619 395214 -17563
rect 395270 -17619 395338 -17563
rect 395394 -17619 395462 -17563
rect 395518 -17619 395586 -17563
rect 395642 -17619 395710 -17563
rect 395766 -17619 395898 -17563
rect 395954 -17619 396022 -17563
rect 396078 -17619 396146 -17563
rect 396202 -17619 396270 -17563
rect 396326 -17619 396394 -17563
rect 396450 -17619 396518 -17563
rect 396574 -17619 396642 -17563
rect 396698 -17619 396766 -17563
rect 396822 -17619 396890 -17563
rect 396946 -17619 397014 -17563
rect 397070 -17619 397200 -17563
rect 388000 -17820 397200 -17619
rect 388000 -17858 388800 -17820
rect 388000 -17914 388114 -17858
rect 388170 -17914 388238 -17858
rect 388294 -17914 388362 -17858
rect 388418 -17914 388486 -17858
rect 388542 -17914 388610 -17858
rect 388666 -17914 388800 -17858
rect 388000 -17982 388800 -17914
rect 388000 -18038 388114 -17982
rect 388170 -18038 388238 -17982
rect 388294 -18038 388362 -17982
rect 388418 -18038 388486 -17982
rect 388542 -18038 388610 -17982
rect 388666 -18038 388800 -17982
rect 388000 -18106 388800 -18038
rect 388000 -18162 388114 -18106
rect 388170 -18162 388238 -18106
rect 388294 -18162 388362 -18106
rect 388418 -18162 388486 -18106
rect 388542 -18162 388610 -18106
rect 388666 -18162 388800 -18106
rect 388000 -18230 388800 -18162
rect 388000 -18286 388114 -18230
rect 388170 -18286 388238 -18230
rect 388294 -18286 388362 -18230
rect 388418 -18286 388486 -18230
rect 388542 -18286 388610 -18230
rect 388666 -18286 388800 -18230
rect 388000 -18354 388800 -18286
rect 388000 -18410 388114 -18354
rect 388170 -18410 388238 -18354
rect 388294 -18410 388362 -18354
rect 388418 -18410 388486 -18354
rect 388542 -18410 388610 -18354
rect 388666 -18410 388800 -18354
rect 388000 -18478 388800 -18410
rect 388000 -18534 388114 -18478
rect 388170 -18534 388238 -18478
rect 388294 -18534 388362 -18478
rect 388418 -18534 388486 -18478
rect 388542 -18534 388610 -18478
rect 388666 -18534 388800 -18478
rect 388000 -18602 388800 -18534
rect 388000 -18658 388114 -18602
rect 388170 -18658 388238 -18602
rect 388294 -18658 388362 -18602
rect 388418 -18658 388486 -18602
rect 388542 -18658 388610 -18602
rect 388666 -18658 388800 -18602
rect 388000 -18726 388800 -18658
rect 388000 -18782 388114 -18726
rect 388170 -18782 388238 -18726
rect 388294 -18782 388362 -18726
rect 388418 -18782 388486 -18726
rect 388542 -18782 388610 -18726
rect 388666 -18782 388800 -18726
rect 388000 -18850 388800 -18782
rect 388000 -18906 388114 -18850
rect 388170 -18906 388238 -18850
rect 388294 -18906 388362 -18850
rect 388418 -18906 388486 -18850
rect 388542 -18906 388610 -18850
rect 388666 -18906 388800 -18850
rect 388000 -18974 388800 -18906
rect 388000 -19030 388114 -18974
rect 388170 -19030 388238 -18974
rect 388294 -19030 388362 -18974
rect 388418 -19030 388486 -18974
rect 388542 -19030 388610 -18974
rect 388666 -19030 388800 -18974
rect 388000 -19098 388800 -19030
rect 388000 -19154 388114 -19098
rect 388170 -19154 388238 -19098
rect 388294 -19154 388362 -19098
rect 388418 -19154 388486 -19098
rect 388542 -19154 388610 -19098
rect 388666 -19154 388800 -19098
rect 388000 -19222 388800 -19154
rect 388000 -19278 388114 -19222
rect 388170 -19278 388238 -19222
rect 388294 -19278 388362 -19222
rect 388418 -19278 388486 -19222
rect 388542 -19278 388610 -19222
rect 388666 -19278 388800 -19222
rect 388000 -19346 388800 -19278
rect 388000 -19402 388114 -19346
rect 388170 -19402 388238 -19346
rect 388294 -19402 388362 -19346
rect 388418 -19402 388486 -19346
rect 388542 -19402 388610 -19346
rect 388666 -19402 388800 -19346
rect 388000 -19470 388800 -19402
rect 388000 -19526 388114 -19470
rect 388170 -19526 388238 -19470
rect 388294 -19526 388362 -19470
rect 388418 -19526 388486 -19470
rect 388542 -19526 388610 -19470
rect 388666 -19526 388800 -19470
rect 388000 -19594 388800 -19526
rect 388000 -19650 388114 -19594
rect 388170 -19650 388238 -19594
rect 388294 -19650 388362 -19594
rect 388418 -19650 388486 -19594
rect 388542 -19650 388610 -19594
rect 388666 -19650 388800 -19594
rect 388000 -19718 388800 -19650
rect 388000 -19774 388114 -19718
rect 388170 -19774 388238 -19718
rect 388294 -19774 388362 -19718
rect 388418 -19774 388486 -19718
rect 388542 -19774 388610 -19718
rect 388666 -19774 388800 -19718
rect 388000 -19842 388800 -19774
rect 388000 -19898 388114 -19842
rect 388170 -19898 388238 -19842
rect 388294 -19898 388362 -19842
rect 388418 -19898 388486 -19842
rect 388542 -19898 388610 -19842
rect 388666 -19898 388800 -19842
rect 388000 -19966 388800 -19898
rect 388000 -20022 388114 -19966
rect 388170 -20022 388238 -19966
rect 388294 -20022 388362 -19966
rect 388418 -20022 388486 -19966
rect 388542 -20022 388610 -19966
rect 388666 -20022 388800 -19966
rect 388000 -20090 388800 -20022
rect 388000 -20146 388114 -20090
rect 388170 -20146 388238 -20090
rect 388294 -20146 388362 -20090
rect 388418 -20146 388486 -20090
rect 388542 -20146 388610 -20090
rect 388666 -20146 388800 -20090
rect 388000 -20214 388800 -20146
rect 388000 -20270 388114 -20214
rect 388170 -20270 388238 -20214
rect 388294 -20270 388362 -20214
rect 388418 -20270 388486 -20214
rect 388542 -20270 388610 -20214
rect 388666 -20270 388800 -20214
rect 388000 -20338 388800 -20270
rect 388000 -20394 388114 -20338
rect 388170 -20394 388238 -20338
rect 388294 -20394 388362 -20338
rect 388418 -20394 388486 -20338
rect 388542 -20394 388610 -20338
rect 388666 -20394 388800 -20338
rect 388000 -20462 388800 -20394
rect 388000 -20518 388114 -20462
rect 388170 -20518 388238 -20462
rect 388294 -20518 388362 -20462
rect 388418 -20518 388486 -20462
rect 388542 -20518 388610 -20462
rect 388666 -20518 388800 -20462
rect 388000 -20586 388800 -20518
rect 388000 -20642 388114 -20586
rect 388170 -20642 388238 -20586
rect 388294 -20642 388362 -20586
rect 388418 -20642 388486 -20586
rect 388542 -20642 388610 -20586
rect 388666 -20642 388800 -20586
rect 388000 -20710 388800 -20642
rect 388000 -20766 388114 -20710
rect 388170 -20766 388238 -20710
rect 388294 -20766 388362 -20710
rect 388418 -20766 388486 -20710
rect 388542 -20766 388610 -20710
rect 388666 -20766 388800 -20710
rect 388000 -20834 388800 -20766
rect 388000 -20890 388114 -20834
rect 388170 -20890 388238 -20834
rect 388294 -20890 388362 -20834
rect 388418 -20890 388486 -20834
rect 388542 -20890 388610 -20834
rect 388666 -20890 388800 -20834
rect 388000 -20958 388800 -20890
rect 388000 -21014 388114 -20958
rect 388170 -21014 388238 -20958
rect 388294 -21014 388362 -20958
rect 388418 -21014 388486 -20958
rect 388542 -21014 388610 -20958
rect 388666 -21014 388800 -20958
rect 388000 -21082 388800 -21014
rect 388000 -21138 388114 -21082
rect 388170 -21138 388238 -21082
rect 388294 -21138 388362 -21082
rect 388418 -21138 388486 -21082
rect 388542 -21138 388610 -21082
rect 388666 -21138 388800 -21082
rect 388000 -21206 388800 -21138
rect 388000 -21262 388114 -21206
rect 388170 -21262 388238 -21206
rect 388294 -21262 388362 -21206
rect 388418 -21262 388486 -21206
rect 388542 -21262 388610 -21206
rect 388666 -21262 388800 -21206
rect 388000 -21330 388800 -21262
rect 388000 -21386 388114 -21330
rect 388170 -21386 388238 -21330
rect 388294 -21386 388362 -21330
rect 388418 -21386 388486 -21330
rect 388542 -21386 388610 -21330
rect 388666 -21386 388800 -21330
rect 388000 -21454 388800 -21386
rect 388000 -21510 388114 -21454
rect 388170 -21510 388238 -21454
rect 388294 -21510 388362 -21454
rect 388418 -21510 388486 -21454
rect 388542 -21510 388610 -21454
rect 388666 -21510 388800 -21454
rect 388000 -21578 388800 -21510
rect 388000 -21634 388114 -21578
rect 388170 -21634 388238 -21578
rect 388294 -21634 388362 -21578
rect 388418 -21634 388486 -21578
rect 388542 -21634 388610 -21578
rect 388666 -21634 388800 -21578
rect 388000 -21702 388800 -21634
rect 388000 -21758 388114 -21702
rect 388170 -21758 388238 -21702
rect 388294 -21758 388362 -21702
rect 388418 -21758 388486 -21702
rect 388542 -21758 388610 -21702
rect 388666 -21758 388800 -21702
rect 388000 -21826 388800 -21758
rect 388000 -21882 388114 -21826
rect 388170 -21882 388238 -21826
rect 388294 -21882 388362 -21826
rect 388418 -21882 388486 -21826
rect 388542 -21882 388610 -21826
rect 388666 -21882 388800 -21826
rect 388000 -21950 388800 -21882
rect 388000 -22006 388114 -21950
rect 388170 -22006 388238 -21950
rect 388294 -22006 388362 -21950
rect 388418 -22006 388486 -21950
rect 388542 -22006 388610 -21950
rect 388666 -22006 388800 -21950
rect 388000 -22074 388800 -22006
rect 388000 -22130 388114 -22074
rect 388170 -22130 388238 -22074
rect 388294 -22130 388362 -22074
rect 388418 -22130 388486 -22074
rect 388542 -22130 388610 -22074
rect 388666 -22130 388800 -22074
rect 388000 -22198 388800 -22130
rect 388000 -22254 388114 -22198
rect 388170 -22254 388238 -22198
rect 388294 -22254 388362 -22198
rect 388418 -22254 388486 -22198
rect 388542 -22254 388610 -22198
rect 388666 -22254 388800 -22198
rect 388000 -22322 388800 -22254
rect 388000 -22378 388114 -22322
rect 388170 -22378 388238 -22322
rect 388294 -22378 388362 -22322
rect 388418 -22378 388486 -22322
rect 388542 -22378 388610 -22322
rect 388666 -22378 388800 -22322
rect 388000 -22446 388800 -22378
rect 388000 -22502 388114 -22446
rect 388170 -22502 388238 -22446
rect 388294 -22502 388362 -22446
rect 388418 -22502 388486 -22446
rect 388542 -22502 388610 -22446
rect 388666 -22502 388800 -22446
rect 388000 -22570 388800 -22502
rect 388000 -22626 388114 -22570
rect 388170 -22626 388238 -22570
rect 388294 -22626 388362 -22570
rect 388418 -22626 388486 -22570
rect 388542 -22626 388610 -22570
rect 388666 -22626 388800 -22570
rect 388000 -22694 388800 -22626
rect 388000 -22750 388114 -22694
rect 388170 -22750 388238 -22694
rect 388294 -22750 388362 -22694
rect 388418 -22750 388486 -22694
rect 388542 -22750 388610 -22694
rect 388666 -22750 388800 -22694
rect 388000 -22818 388800 -22750
rect 388000 -22874 388114 -22818
rect 388170 -22874 388238 -22818
rect 388294 -22874 388362 -22818
rect 388418 -22874 388486 -22818
rect 388542 -22874 388610 -22818
rect 388666 -22874 388800 -22818
rect 388000 -22942 388800 -22874
rect 388000 -22998 388114 -22942
rect 388170 -22998 388238 -22942
rect 388294 -22998 388362 -22942
rect 388418 -22998 388486 -22942
rect 388542 -22998 388610 -22942
rect 388666 -22998 388800 -22942
rect 388000 -23066 388800 -22998
rect 388000 -23122 388114 -23066
rect 388170 -23122 388238 -23066
rect 388294 -23122 388362 -23066
rect 388418 -23122 388486 -23066
rect 388542 -23122 388610 -23066
rect 388666 -23122 388800 -23066
rect 388000 -23190 388800 -23122
rect 388000 -23246 388114 -23190
rect 388170 -23246 388238 -23190
rect 388294 -23246 388362 -23190
rect 388418 -23246 388486 -23190
rect 388542 -23246 388610 -23190
rect 388666 -23246 388800 -23190
rect 388000 -23314 388800 -23246
rect 388000 -23370 388114 -23314
rect 388170 -23370 388238 -23314
rect 388294 -23370 388362 -23314
rect 388418 -23370 388486 -23314
rect 388542 -23370 388610 -23314
rect 388666 -23370 388800 -23314
rect 388000 -23438 388800 -23370
rect 388000 -23494 388114 -23438
rect 388170 -23494 388238 -23438
rect 388294 -23494 388362 -23438
rect 388418 -23494 388486 -23438
rect 388542 -23494 388610 -23438
rect 388666 -23494 388800 -23438
rect 388000 -23562 388800 -23494
rect 388000 -23618 388114 -23562
rect 388170 -23618 388238 -23562
rect 388294 -23618 388362 -23562
rect 388418 -23618 388486 -23562
rect 388542 -23618 388610 -23562
rect 388666 -23618 388800 -23562
rect 388000 -23686 388800 -23618
rect 388000 -23742 388114 -23686
rect 388170 -23742 388238 -23686
rect 388294 -23742 388362 -23686
rect 388418 -23742 388486 -23686
rect 388542 -23742 388610 -23686
rect 388666 -23742 388800 -23686
rect 388000 -23810 388800 -23742
rect 388000 -23866 388114 -23810
rect 388170 -23866 388238 -23810
rect 388294 -23866 388362 -23810
rect 388418 -23866 388486 -23810
rect 388542 -23866 388610 -23810
rect 388666 -23866 388800 -23810
rect 388000 -23934 388800 -23866
rect 388000 -23990 388114 -23934
rect 388170 -23990 388238 -23934
rect 388294 -23990 388362 -23934
rect 388418 -23990 388486 -23934
rect 388542 -23990 388610 -23934
rect 388666 -23990 388800 -23934
rect 388000 -24058 388800 -23990
rect 388000 -24114 388114 -24058
rect 388170 -24114 388238 -24058
rect 388294 -24114 388362 -24058
rect 388418 -24114 388486 -24058
rect 388542 -24114 388610 -24058
rect 388666 -24114 388800 -24058
rect 388000 -24182 388800 -24114
rect 388000 -24238 388114 -24182
rect 388170 -24238 388238 -24182
rect 388294 -24238 388362 -24182
rect 388418 -24238 388486 -24182
rect 388542 -24238 388610 -24182
rect 388666 -24238 388800 -24182
rect 388000 -24306 388800 -24238
rect 388000 -24362 388114 -24306
rect 388170 -24362 388238 -24306
rect 388294 -24362 388362 -24306
rect 388418 -24362 388486 -24306
rect 388542 -24362 388610 -24306
rect 388666 -24362 388800 -24306
rect 388000 -24430 388800 -24362
rect 388000 -24486 388114 -24430
rect 388170 -24486 388238 -24430
rect 388294 -24486 388362 -24430
rect 388418 -24486 388486 -24430
rect 388542 -24486 388610 -24430
rect 388666 -24486 388800 -24430
rect 388000 -24554 388800 -24486
rect 388000 -24610 388114 -24554
rect 388170 -24610 388238 -24554
rect 388294 -24610 388362 -24554
rect 388418 -24610 388486 -24554
rect 388542 -24610 388610 -24554
rect 388666 -24610 388800 -24554
rect 388000 -24678 388800 -24610
rect 388000 -24734 388114 -24678
rect 388170 -24734 388238 -24678
rect 388294 -24734 388362 -24678
rect 388418 -24734 388486 -24678
rect 388542 -24734 388610 -24678
rect 388666 -24734 388800 -24678
rect 388000 -24802 388800 -24734
rect 388000 -24858 388114 -24802
rect 388170 -24858 388238 -24802
rect 388294 -24858 388362 -24802
rect 388418 -24858 388486 -24802
rect 388542 -24858 388610 -24802
rect 388666 -24858 388800 -24802
rect 388000 -24926 388800 -24858
rect 388000 -24982 388114 -24926
rect 388170 -24982 388238 -24926
rect 388294 -24982 388362 -24926
rect 388418 -24982 388486 -24926
rect 388542 -24982 388610 -24926
rect 388666 -24982 388800 -24926
rect 388000 -25050 388800 -24982
rect 388000 -25106 388114 -25050
rect 388170 -25106 388238 -25050
rect 388294 -25106 388362 -25050
rect 388418 -25106 388486 -25050
rect 388542 -25106 388610 -25050
rect 388666 -25106 388800 -25050
rect 388000 -25174 388800 -25106
rect 388000 -25230 388114 -25174
rect 388170 -25230 388238 -25174
rect 388294 -25230 388362 -25174
rect 388418 -25230 388486 -25174
rect 388542 -25230 388610 -25174
rect 388666 -25230 388800 -25174
rect 388000 -25298 388800 -25230
rect 388000 -25354 388114 -25298
rect 388170 -25354 388238 -25298
rect 388294 -25354 388362 -25298
rect 388418 -25354 388486 -25298
rect 388542 -25354 388610 -25298
rect 388666 -25354 388800 -25298
rect 388000 -25422 388800 -25354
rect 388000 -25478 388114 -25422
rect 388170 -25478 388238 -25422
rect 388294 -25478 388362 -25422
rect 388418 -25478 388486 -25422
rect 388542 -25478 388610 -25422
rect 388666 -25478 388800 -25422
rect 388000 -25542 388800 -25478
rect 389068 -17950 389408 -17820
rect 389068 -18006 389141 -17950
rect 389197 -18006 389283 -17950
rect 389339 -18006 389408 -17950
rect 389068 -18092 389408 -18006
rect 389068 -18148 389141 -18092
rect 389197 -18148 389283 -18092
rect 389339 -18148 389408 -18092
rect 389068 -18234 389408 -18148
rect 389068 -18290 389141 -18234
rect 389197 -18290 389283 -18234
rect 389339 -18290 389408 -18234
rect 389068 -18376 389408 -18290
rect 389068 -18432 389141 -18376
rect 389197 -18432 389283 -18376
rect 389339 -18432 389408 -18376
rect 389068 -18518 389408 -18432
rect 389068 -18574 389141 -18518
rect 389197 -18574 389283 -18518
rect 389339 -18574 389408 -18518
rect 389068 -18660 389408 -18574
rect 389068 -18716 389141 -18660
rect 389197 -18716 389283 -18660
rect 389339 -18716 389408 -18660
rect 389068 -18802 389408 -18716
rect 389068 -18858 389141 -18802
rect 389197 -18858 389283 -18802
rect 389339 -18858 389408 -18802
rect 389068 -18944 389408 -18858
rect 389068 -19000 389141 -18944
rect 389197 -19000 389283 -18944
rect 389339 -19000 389408 -18944
rect 389068 -19086 389408 -19000
rect 389068 -19142 389141 -19086
rect 389197 -19142 389283 -19086
rect 389339 -19142 389408 -19086
rect 389068 -19228 389408 -19142
rect 389068 -19284 389141 -19228
rect 389197 -19284 389283 -19228
rect 389339 -19284 389408 -19228
rect 389068 -19370 389408 -19284
rect 389068 -19426 389141 -19370
rect 389197 -19426 389283 -19370
rect 389339 -19426 389408 -19370
rect 389068 -19512 389408 -19426
rect 389068 -19568 389141 -19512
rect 389197 -19568 389283 -19512
rect 389339 -19568 389408 -19512
rect 389068 -19654 389408 -19568
rect 389068 -19710 389141 -19654
rect 389197 -19710 389283 -19654
rect 389339 -19710 389408 -19654
rect 389068 -19796 389408 -19710
rect 389068 -19852 389141 -19796
rect 389197 -19852 389283 -19796
rect 389339 -19852 389408 -19796
rect 389068 -19938 389408 -19852
rect 389068 -19994 389141 -19938
rect 389197 -19994 389283 -19938
rect 389339 -19994 389408 -19938
rect 389068 -20080 389408 -19994
rect 389068 -20136 389141 -20080
rect 389197 -20136 389283 -20080
rect 389339 -20136 389408 -20080
rect 389068 -20222 389408 -20136
rect 389068 -20278 389141 -20222
rect 389197 -20278 389283 -20222
rect 389339 -20278 389408 -20222
rect 389068 -20364 389408 -20278
rect 389068 -20420 389141 -20364
rect 389197 -20420 389283 -20364
rect 389339 -20420 389408 -20364
rect 389068 -20506 389408 -20420
rect 389068 -20562 389141 -20506
rect 389197 -20562 389283 -20506
rect 389339 -20562 389408 -20506
rect 389068 -20648 389408 -20562
rect 389068 -20704 389141 -20648
rect 389197 -20704 389283 -20648
rect 389339 -20704 389408 -20648
rect 389068 -20790 389408 -20704
rect 389068 -20846 389141 -20790
rect 389197 -20846 389283 -20790
rect 389339 -20846 389408 -20790
rect 389068 -20932 389408 -20846
rect 389068 -20988 389141 -20932
rect 389197 -20988 389283 -20932
rect 389339 -20988 389408 -20932
rect 389068 -21074 389408 -20988
rect 389068 -21130 389141 -21074
rect 389197 -21130 389283 -21074
rect 389339 -21130 389408 -21074
rect 389068 -21216 389408 -21130
rect 389068 -21272 389141 -21216
rect 389197 -21272 389283 -21216
rect 389339 -21272 389408 -21216
rect 389068 -21358 389408 -21272
rect 389068 -21414 389141 -21358
rect 389197 -21414 389283 -21358
rect 389339 -21414 389408 -21358
rect 389068 -21500 389408 -21414
rect 389068 -21556 389141 -21500
rect 389197 -21556 389283 -21500
rect 389339 -21556 389408 -21500
rect 389068 -21642 389408 -21556
rect 389068 -21698 389141 -21642
rect 389197 -21698 389283 -21642
rect 389339 -21698 389408 -21642
rect 389068 -21784 389408 -21698
rect 389068 -21840 389141 -21784
rect 389197 -21840 389283 -21784
rect 389339 -21840 389408 -21784
rect 389068 -21926 389408 -21840
rect 389068 -21982 389141 -21926
rect 389197 -21982 389283 -21926
rect 389339 -21982 389408 -21926
rect 389068 -22068 389408 -21982
rect 389068 -22124 389141 -22068
rect 389197 -22124 389283 -22068
rect 389339 -22124 389408 -22068
rect 389068 -22210 389408 -22124
rect 389068 -22266 389141 -22210
rect 389197 -22266 389283 -22210
rect 389339 -22266 389408 -22210
rect 389068 -22352 389408 -22266
rect 389068 -22408 389141 -22352
rect 389197 -22408 389283 -22352
rect 389339 -22408 389408 -22352
rect 389068 -22494 389408 -22408
rect 389068 -22550 389141 -22494
rect 389197 -22550 389283 -22494
rect 389339 -22550 389408 -22494
rect 389068 -22636 389408 -22550
rect 389068 -22692 389141 -22636
rect 389197 -22692 389283 -22636
rect 389339 -22692 389408 -22636
rect 389068 -22778 389408 -22692
rect 389068 -22834 389141 -22778
rect 389197 -22834 389283 -22778
rect 389339 -22834 389408 -22778
rect 389068 -22920 389408 -22834
rect 389068 -22976 389141 -22920
rect 389197 -22976 389283 -22920
rect 389339 -22976 389408 -22920
rect 389068 -23062 389408 -22976
rect 389068 -23118 389141 -23062
rect 389197 -23118 389283 -23062
rect 389339 -23118 389408 -23062
rect 389068 -23204 389408 -23118
rect 389068 -23260 389141 -23204
rect 389197 -23260 389283 -23204
rect 389339 -23260 389408 -23204
rect 389068 -23346 389408 -23260
rect 389068 -23402 389141 -23346
rect 389197 -23402 389283 -23346
rect 389339 -23402 389408 -23346
rect 389068 -23488 389408 -23402
rect 389068 -23544 389141 -23488
rect 389197 -23544 389283 -23488
rect 389339 -23544 389408 -23488
rect 389068 -23630 389408 -23544
rect 389068 -23686 389141 -23630
rect 389197 -23686 389283 -23630
rect 389339 -23686 389408 -23630
rect 389068 -23772 389408 -23686
rect 389068 -23828 389141 -23772
rect 389197 -23828 389283 -23772
rect 389339 -23828 389408 -23772
rect 389068 -23914 389408 -23828
rect 389068 -23970 389141 -23914
rect 389197 -23970 389283 -23914
rect 389339 -23970 389408 -23914
rect 389068 -24056 389408 -23970
rect 389068 -24112 389141 -24056
rect 389197 -24112 389283 -24056
rect 389339 -24112 389408 -24056
rect 389068 -24198 389408 -24112
rect 389068 -24254 389141 -24198
rect 389197 -24254 389283 -24198
rect 389339 -24254 389408 -24198
rect 389068 -24340 389408 -24254
rect 389068 -24396 389141 -24340
rect 389197 -24396 389283 -24340
rect 389339 -24396 389408 -24340
rect 389068 -24482 389408 -24396
rect 389068 -24538 389141 -24482
rect 389197 -24538 389283 -24482
rect 389339 -24538 389408 -24482
rect 389068 -24624 389408 -24538
rect 389068 -24680 389141 -24624
rect 389197 -24680 389283 -24624
rect 389339 -24680 389408 -24624
rect 389068 -24766 389408 -24680
rect 389068 -24822 389141 -24766
rect 389197 -24822 389283 -24766
rect 389339 -24822 389408 -24766
rect 389068 -24908 389408 -24822
rect 389068 -24964 389141 -24908
rect 389197 -24964 389283 -24908
rect 389339 -24964 389408 -24908
rect 389068 -25050 389408 -24964
rect 389068 -25106 389141 -25050
rect 389197 -25106 389283 -25050
rect 389339 -25106 389408 -25050
rect 389068 -25192 389408 -25106
rect 389068 -25248 389141 -25192
rect 389197 -25248 389283 -25192
rect 389339 -25248 389408 -25192
rect 389068 -25334 389408 -25248
rect 389068 -25390 389141 -25334
rect 389197 -25390 389283 -25334
rect 389339 -25390 389408 -25334
rect 389068 -25476 389408 -25390
rect 389068 -25532 389141 -25476
rect 389197 -25532 389283 -25476
rect 389339 -25532 389408 -25476
rect 389068 -25542 389408 -25532
rect 389468 -17950 389808 -17820
rect 389468 -18006 389542 -17950
rect 389598 -18006 389684 -17950
rect 389740 -18006 389808 -17950
rect 389468 -18092 389808 -18006
rect 389468 -18148 389542 -18092
rect 389598 -18148 389684 -18092
rect 389740 -18148 389808 -18092
rect 389468 -18234 389808 -18148
rect 389468 -18290 389542 -18234
rect 389598 -18290 389684 -18234
rect 389740 -18290 389808 -18234
rect 389468 -18376 389808 -18290
rect 389468 -18432 389542 -18376
rect 389598 -18432 389684 -18376
rect 389740 -18432 389808 -18376
rect 389468 -18518 389808 -18432
rect 389468 -18574 389542 -18518
rect 389598 -18574 389684 -18518
rect 389740 -18574 389808 -18518
rect 389468 -18660 389808 -18574
rect 389468 -18716 389542 -18660
rect 389598 -18716 389684 -18660
rect 389740 -18716 389808 -18660
rect 389468 -18802 389808 -18716
rect 389468 -18858 389542 -18802
rect 389598 -18858 389684 -18802
rect 389740 -18858 389808 -18802
rect 389468 -18944 389808 -18858
rect 389468 -19000 389542 -18944
rect 389598 -19000 389684 -18944
rect 389740 -19000 389808 -18944
rect 389468 -19086 389808 -19000
rect 389468 -19142 389542 -19086
rect 389598 -19142 389684 -19086
rect 389740 -19142 389808 -19086
rect 389468 -19228 389808 -19142
rect 389468 -19284 389542 -19228
rect 389598 -19284 389684 -19228
rect 389740 -19284 389808 -19228
rect 389468 -19370 389808 -19284
rect 389468 -19426 389542 -19370
rect 389598 -19426 389684 -19370
rect 389740 -19426 389808 -19370
rect 389468 -19512 389808 -19426
rect 389468 -19568 389542 -19512
rect 389598 -19568 389684 -19512
rect 389740 -19568 389808 -19512
rect 389468 -19654 389808 -19568
rect 389468 -19710 389542 -19654
rect 389598 -19710 389684 -19654
rect 389740 -19710 389808 -19654
rect 389468 -19796 389808 -19710
rect 389468 -19852 389542 -19796
rect 389598 -19852 389684 -19796
rect 389740 -19852 389808 -19796
rect 389468 -19938 389808 -19852
rect 389468 -19994 389542 -19938
rect 389598 -19994 389684 -19938
rect 389740 -19994 389808 -19938
rect 389468 -20080 389808 -19994
rect 389468 -20136 389542 -20080
rect 389598 -20136 389684 -20080
rect 389740 -20136 389808 -20080
rect 389468 -20222 389808 -20136
rect 389468 -20278 389542 -20222
rect 389598 -20278 389684 -20222
rect 389740 -20278 389808 -20222
rect 389468 -20364 389808 -20278
rect 389468 -20420 389542 -20364
rect 389598 -20420 389684 -20364
rect 389740 -20420 389808 -20364
rect 389468 -20506 389808 -20420
rect 389468 -20562 389542 -20506
rect 389598 -20562 389684 -20506
rect 389740 -20562 389808 -20506
rect 389468 -20648 389808 -20562
rect 389468 -20704 389542 -20648
rect 389598 -20704 389684 -20648
rect 389740 -20704 389808 -20648
rect 389468 -20790 389808 -20704
rect 389468 -20846 389542 -20790
rect 389598 -20846 389684 -20790
rect 389740 -20846 389808 -20790
rect 389468 -20932 389808 -20846
rect 389468 -20988 389542 -20932
rect 389598 -20988 389684 -20932
rect 389740 -20988 389808 -20932
rect 389468 -21074 389808 -20988
rect 389468 -21130 389542 -21074
rect 389598 -21130 389684 -21074
rect 389740 -21130 389808 -21074
rect 389468 -21216 389808 -21130
rect 389468 -21272 389542 -21216
rect 389598 -21272 389684 -21216
rect 389740 -21272 389808 -21216
rect 389468 -21358 389808 -21272
rect 389468 -21414 389542 -21358
rect 389598 -21414 389684 -21358
rect 389740 -21414 389808 -21358
rect 389468 -21500 389808 -21414
rect 389468 -21556 389542 -21500
rect 389598 -21556 389684 -21500
rect 389740 -21556 389808 -21500
rect 389468 -21642 389808 -21556
rect 389468 -21698 389542 -21642
rect 389598 -21698 389684 -21642
rect 389740 -21698 389808 -21642
rect 389468 -21784 389808 -21698
rect 389468 -21840 389542 -21784
rect 389598 -21840 389684 -21784
rect 389740 -21840 389808 -21784
rect 389468 -21926 389808 -21840
rect 389468 -21982 389542 -21926
rect 389598 -21982 389684 -21926
rect 389740 -21982 389808 -21926
rect 389468 -22068 389808 -21982
rect 389468 -22124 389542 -22068
rect 389598 -22124 389684 -22068
rect 389740 -22124 389808 -22068
rect 389468 -22210 389808 -22124
rect 389468 -22266 389542 -22210
rect 389598 -22266 389684 -22210
rect 389740 -22266 389808 -22210
rect 389468 -22352 389808 -22266
rect 389468 -22408 389542 -22352
rect 389598 -22408 389684 -22352
rect 389740 -22408 389808 -22352
rect 389468 -22494 389808 -22408
rect 389468 -22550 389542 -22494
rect 389598 -22550 389684 -22494
rect 389740 -22550 389808 -22494
rect 389468 -22636 389808 -22550
rect 389468 -22692 389542 -22636
rect 389598 -22692 389684 -22636
rect 389740 -22692 389808 -22636
rect 389468 -22778 389808 -22692
rect 389468 -22834 389542 -22778
rect 389598 -22834 389684 -22778
rect 389740 -22834 389808 -22778
rect 389468 -22920 389808 -22834
rect 389468 -22976 389542 -22920
rect 389598 -22976 389684 -22920
rect 389740 -22976 389808 -22920
rect 389468 -23062 389808 -22976
rect 389468 -23118 389542 -23062
rect 389598 -23118 389684 -23062
rect 389740 -23118 389808 -23062
rect 389468 -23204 389808 -23118
rect 389468 -23260 389542 -23204
rect 389598 -23260 389684 -23204
rect 389740 -23260 389808 -23204
rect 389468 -23346 389808 -23260
rect 389468 -23402 389542 -23346
rect 389598 -23402 389684 -23346
rect 389740 -23402 389808 -23346
rect 389468 -23488 389808 -23402
rect 389468 -23544 389542 -23488
rect 389598 -23544 389684 -23488
rect 389740 -23544 389808 -23488
rect 389468 -23630 389808 -23544
rect 389468 -23686 389542 -23630
rect 389598 -23686 389684 -23630
rect 389740 -23686 389808 -23630
rect 389468 -23772 389808 -23686
rect 389468 -23828 389542 -23772
rect 389598 -23828 389684 -23772
rect 389740 -23828 389808 -23772
rect 389468 -23914 389808 -23828
rect 389468 -23970 389542 -23914
rect 389598 -23970 389684 -23914
rect 389740 -23970 389808 -23914
rect 389468 -24056 389808 -23970
rect 389468 -24112 389542 -24056
rect 389598 -24112 389684 -24056
rect 389740 -24112 389808 -24056
rect 389468 -24198 389808 -24112
rect 389468 -24254 389542 -24198
rect 389598 -24254 389684 -24198
rect 389740 -24254 389808 -24198
rect 389468 -24340 389808 -24254
rect 389468 -24396 389542 -24340
rect 389598 -24396 389684 -24340
rect 389740 -24396 389808 -24340
rect 389468 -24482 389808 -24396
rect 389468 -24538 389542 -24482
rect 389598 -24538 389684 -24482
rect 389740 -24538 389808 -24482
rect 389468 -24624 389808 -24538
rect 389468 -24680 389542 -24624
rect 389598 -24680 389684 -24624
rect 389740 -24680 389808 -24624
rect 389468 -24766 389808 -24680
rect 389468 -24822 389542 -24766
rect 389598 -24822 389684 -24766
rect 389740 -24822 389808 -24766
rect 389468 -24908 389808 -24822
rect 389468 -24964 389542 -24908
rect 389598 -24964 389684 -24908
rect 389740 -24964 389808 -24908
rect 389468 -25050 389808 -24964
rect 389468 -25106 389542 -25050
rect 389598 -25106 389684 -25050
rect 389740 -25106 389808 -25050
rect 389468 -25192 389808 -25106
rect 389468 -25248 389542 -25192
rect 389598 -25248 389684 -25192
rect 389740 -25248 389808 -25192
rect 389468 -25334 389808 -25248
rect 389468 -25390 389542 -25334
rect 389598 -25390 389684 -25334
rect 389740 -25390 389808 -25334
rect 389468 -25476 389808 -25390
rect 389468 -25532 389542 -25476
rect 389598 -25532 389684 -25476
rect 389740 -25532 389808 -25476
rect 389468 -25542 389808 -25532
rect 389868 -17950 390208 -17820
rect 389868 -18006 389942 -17950
rect 389998 -18006 390084 -17950
rect 390140 -18006 390208 -17950
rect 389868 -18092 390208 -18006
rect 389868 -18148 389942 -18092
rect 389998 -18148 390084 -18092
rect 390140 -18148 390208 -18092
rect 389868 -18234 390208 -18148
rect 389868 -18290 389942 -18234
rect 389998 -18290 390084 -18234
rect 390140 -18290 390208 -18234
rect 389868 -18376 390208 -18290
rect 389868 -18432 389942 -18376
rect 389998 -18432 390084 -18376
rect 390140 -18432 390208 -18376
rect 389868 -18518 390208 -18432
rect 389868 -18574 389942 -18518
rect 389998 -18574 390084 -18518
rect 390140 -18574 390208 -18518
rect 389868 -18660 390208 -18574
rect 389868 -18716 389942 -18660
rect 389998 -18716 390084 -18660
rect 390140 -18716 390208 -18660
rect 389868 -18802 390208 -18716
rect 389868 -18858 389942 -18802
rect 389998 -18858 390084 -18802
rect 390140 -18858 390208 -18802
rect 389868 -18944 390208 -18858
rect 389868 -19000 389942 -18944
rect 389998 -19000 390084 -18944
rect 390140 -19000 390208 -18944
rect 389868 -19086 390208 -19000
rect 389868 -19142 389942 -19086
rect 389998 -19142 390084 -19086
rect 390140 -19142 390208 -19086
rect 389868 -19228 390208 -19142
rect 389868 -19284 389942 -19228
rect 389998 -19284 390084 -19228
rect 390140 -19284 390208 -19228
rect 389868 -19370 390208 -19284
rect 389868 -19426 389942 -19370
rect 389998 -19426 390084 -19370
rect 390140 -19426 390208 -19370
rect 389868 -19512 390208 -19426
rect 389868 -19568 389942 -19512
rect 389998 -19568 390084 -19512
rect 390140 -19568 390208 -19512
rect 389868 -19654 390208 -19568
rect 389868 -19710 389942 -19654
rect 389998 -19710 390084 -19654
rect 390140 -19710 390208 -19654
rect 389868 -19796 390208 -19710
rect 389868 -19852 389942 -19796
rect 389998 -19852 390084 -19796
rect 390140 -19852 390208 -19796
rect 389868 -19938 390208 -19852
rect 389868 -19994 389942 -19938
rect 389998 -19994 390084 -19938
rect 390140 -19994 390208 -19938
rect 389868 -20080 390208 -19994
rect 389868 -20136 389942 -20080
rect 389998 -20136 390084 -20080
rect 390140 -20136 390208 -20080
rect 389868 -20222 390208 -20136
rect 389868 -20278 389942 -20222
rect 389998 -20278 390084 -20222
rect 390140 -20278 390208 -20222
rect 389868 -20364 390208 -20278
rect 389868 -20420 389942 -20364
rect 389998 -20420 390084 -20364
rect 390140 -20420 390208 -20364
rect 389868 -20506 390208 -20420
rect 389868 -20562 389942 -20506
rect 389998 -20562 390084 -20506
rect 390140 -20562 390208 -20506
rect 389868 -20648 390208 -20562
rect 389868 -20704 389942 -20648
rect 389998 -20704 390084 -20648
rect 390140 -20704 390208 -20648
rect 389868 -20790 390208 -20704
rect 389868 -20846 389942 -20790
rect 389998 -20846 390084 -20790
rect 390140 -20846 390208 -20790
rect 389868 -20932 390208 -20846
rect 389868 -20988 389942 -20932
rect 389998 -20988 390084 -20932
rect 390140 -20988 390208 -20932
rect 389868 -21074 390208 -20988
rect 389868 -21130 389942 -21074
rect 389998 -21130 390084 -21074
rect 390140 -21130 390208 -21074
rect 389868 -21216 390208 -21130
rect 389868 -21272 389942 -21216
rect 389998 -21272 390084 -21216
rect 390140 -21272 390208 -21216
rect 389868 -21358 390208 -21272
rect 389868 -21414 389942 -21358
rect 389998 -21414 390084 -21358
rect 390140 -21414 390208 -21358
rect 389868 -21500 390208 -21414
rect 389868 -21556 389942 -21500
rect 389998 -21556 390084 -21500
rect 390140 -21556 390208 -21500
rect 389868 -21642 390208 -21556
rect 389868 -21698 389942 -21642
rect 389998 -21698 390084 -21642
rect 390140 -21698 390208 -21642
rect 389868 -21784 390208 -21698
rect 389868 -21840 389942 -21784
rect 389998 -21840 390084 -21784
rect 390140 -21840 390208 -21784
rect 389868 -21926 390208 -21840
rect 389868 -21982 389942 -21926
rect 389998 -21982 390084 -21926
rect 390140 -21982 390208 -21926
rect 389868 -22068 390208 -21982
rect 389868 -22124 389942 -22068
rect 389998 -22124 390084 -22068
rect 390140 -22124 390208 -22068
rect 389868 -22210 390208 -22124
rect 389868 -22266 389942 -22210
rect 389998 -22266 390084 -22210
rect 390140 -22266 390208 -22210
rect 389868 -22352 390208 -22266
rect 389868 -22408 389942 -22352
rect 389998 -22408 390084 -22352
rect 390140 -22408 390208 -22352
rect 389868 -22494 390208 -22408
rect 389868 -22550 389942 -22494
rect 389998 -22550 390084 -22494
rect 390140 -22550 390208 -22494
rect 389868 -22636 390208 -22550
rect 389868 -22692 389942 -22636
rect 389998 -22692 390084 -22636
rect 390140 -22692 390208 -22636
rect 389868 -22778 390208 -22692
rect 389868 -22834 389942 -22778
rect 389998 -22834 390084 -22778
rect 390140 -22834 390208 -22778
rect 389868 -22920 390208 -22834
rect 389868 -22976 389942 -22920
rect 389998 -22976 390084 -22920
rect 390140 -22976 390208 -22920
rect 389868 -23062 390208 -22976
rect 389868 -23118 389942 -23062
rect 389998 -23118 390084 -23062
rect 390140 -23118 390208 -23062
rect 389868 -23204 390208 -23118
rect 389868 -23260 389942 -23204
rect 389998 -23260 390084 -23204
rect 390140 -23260 390208 -23204
rect 389868 -23346 390208 -23260
rect 389868 -23402 389942 -23346
rect 389998 -23402 390084 -23346
rect 390140 -23402 390208 -23346
rect 389868 -23488 390208 -23402
rect 389868 -23544 389942 -23488
rect 389998 -23544 390084 -23488
rect 390140 -23544 390208 -23488
rect 389868 -23630 390208 -23544
rect 389868 -23686 389942 -23630
rect 389998 -23686 390084 -23630
rect 390140 -23686 390208 -23630
rect 389868 -23772 390208 -23686
rect 389868 -23828 389942 -23772
rect 389998 -23828 390084 -23772
rect 390140 -23828 390208 -23772
rect 389868 -23914 390208 -23828
rect 389868 -23970 389942 -23914
rect 389998 -23970 390084 -23914
rect 390140 -23970 390208 -23914
rect 389868 -24056 390208 -23970
rect 389868 -24112 389942 -24056
rect 389998 -24112 390084 -24056
rect 390140 -24112 390208 -24056
rect 389868 -24198 390208 -24112
rect 389868 -24254 389942 -24198
rect 389998 -24254 390084 -24198
rect 390140 -24254 390208 -24198
rect 389868 -24340 390208 -24254
rect 389868 -24396 389942 -24340
rect 389998 -24396 390084 -24340
rect 390140 -24396 390208 -24340
rect 389868 -24482 390208 -24396
rect 389868 -24538 389942 -24482
rect 389998 -24538 390084 -24482
rect 390140 -24538 390208 -24482
rect 389868 -24624 390208 -24538
rect 389868 -24680 389942 -24624
rect 389998 -24680 390084 -24624
rect 390140 -24680 390208 -24624
rect 389868 -24766 390208 -24680
rect 389868 -24822 389942 -24766
rect 389998 -24822 390084 -24766
rect 390140 -24822 390208 -24766
rect 389868 -24908 390208 -24822
rect 389868 -24964 389942 -24908
rect 389998 -24964 390084 -24908
rect 390140 -24964 390208 -24908
rect 389868 -25050 390208 -24964
rect 389868 -25106 389942 -25050
rect 389998 -25106 390084 -25050
rect 390140 -25106 390208 -25050
rect 389868 -25192 390208 -25106
rect 389868 -25248 389942 -25192
rect 389998 -25248 390084 -25192
rect 390140 -25248 390208 -25192
rect 389868 -25334 390208 -25248
rect 389868 -25390 389942 -25334
rect 389998 -25390 390084 -25334
rect 390140 -25390 390208 -25334
rect 389868 -25476 390208 -25390
rect 389868 -25532 389942 -25476
rect 389998 -25532 390084 -25476
rect 390140 -25532 390208 -25476
rect 389868 -25542 390208 -25532
rect 390268 -17950 390608 -17820
rect 390268 -18006 390339 -17950
rect 390395 -18006 390481 -17950
rect 390537 -18006 390608 -17950
rect 390268 -18092 390608 -18006
rect 390268 -18148 390339 -18092
rect 390395 -18148 390481 -18092
rect 390537 -18148 390608 -18092
rect 390268 -18234 390608 -18148
rect 390268 -18290 390339 -18234
rect 390395 -18290 390481 -18234
rect 390537 -18290 390608 -18234
rect 390268 -18376 390608 -18290
rect 390268 -18432 390339 -18376
rect 390395 -18432 390481 -18376
rect 390537 -18432 390608 -18376
rect 390268 -18518 390608 -18432
rect 390268 -18574 390339 -18518
rect 390395 -18574 390481 -18518
rect 390537 -18574 390608 -18518
rect 390268 -18660 390608 -18574
rect 390268 -18716 390339 -18660
rect 390395 -18716 390481 -18660
rect 390537 -18716 390608 -18660
rect 390268 -18802 390608 -18716
rect 390268 -18858 390339 -18802
rect 390395 -18858 390481 -18802
rect 390537 -18858 390608 -18802
rect 390268 -18944 390608 -18858
rect 390268 -19000 390339 -18944
rect 390395 -19000 390481 -18944
rect 390537 -19000 390608 -18944
rect 390268 -19086 390608 -19000
rect 390268 -19142 390339 -19086
rect 390395 -19142 390481 -19086
rect 390537 -19142 390608 -19086
rect 390268 -19228 390608 -19142
rect 390268 -19284 390339 -19228
rect 390395 -19284 390481 -19228
rect 390537 -19284 390608 -19228
rect 390268 -19370 390608 -19284
rect 390268 -19426 390339 -19370
rect 390395 -19426 390481 -19370
rect 390537 -19426 390608 -19370
rect 390268 -19512 390608 -19426
rect 390268 -19568 390339 -19512
rect 390395 -19568 390481 -19512
rect 390537 -19568 390608 -19512
rect 390268 -19654 390608 -19568
rect 390268 -19710 390339 -19654
rect 390395 -19710 390481 -19654
rect 390537 -19710 390608 -19654
rect 390268 -19796 390608 -19710
rect 390268 -19852 390339 -19796
rect 390395 -19852 390481 -19796
rect 390537 -19852 390608 -19796
rect 390268 -19938 390608 -19852
rect 390268 -19994 390339 -19938
rect 390395 -19994 390481 -19938
rect 390537 -19994 390608 -19938
rect 390268 -20080 390608 -19994
rect 390268 -20136 390339 -20080
rect 390395 -20136 390481 -20080
rect 390537 -20136 390608 -20080
rect 390268 -20222 390608 -20136
rect 390268 -20278 390339 -20222
rect 390395 -20278 390481 -20222
rect 390537 -20278 390608 -20222
rect 390268 -20364 390608 -20278
rect 390268 -20420 390339 -20364
rect 390395 -20420 390481 -20364
rect 390537 -20420 390608 -20364
rect 390268 -20506 390608 -20420
rect 390268 -20562 390339 -20506
rect 390395 -20562 390481 -20506
rect 390537 -20562 390608 -20506
rect 390268 -20648 390608 -20562
rect 390268 -20704 390339 -20648
rect 390395 -20704 390481 -20648
rect 390537 -20704 390608 -20648
rect 390268 -20790 390608 -20704
rect 390268 -20846 390339 -20790
rect 390395 -20846 390481 -20790
rect 390537 -20846 390608 -20790
rect 390268 -20932 390608 -20846
rect 390268 -20988 390339 -20932
rect 390395 -20988 390481 -20932
rect 390537 -20988 390608 -20932
rect 390268 -21074 390608 -20988
rect 390268 -21130 390339 -21074
rect 390395 -21130 390481 -21074
rect 390537 -21130 390608 -21074
rect 390268 -21216 390608 -21130
rect 390268 -21272 390339 -21216
rect 390395 -21272 390481 -21216
rect 390537 -21272 390608 -21216
rect 390268 -21358 390608 -21272
rect 390268 -21414 390339 -21358
rect 390395 -21414 390481 -21358
rect 390537 -21414 390608 -21358
rect 390268 -21500 390608 -21414
rect 390268 -21556 390339 -21500
rect 390395 -21556 390481 -21500
rect 390537 -21556 390608 -21500
rect 390268 -21642 390608 -21556
rect 390268 -21698 390339 -21642
rect 390395 -21698 390481 -21642
rect 390537 -21698 390608 -21642
rect 390268 -21784 390608 -21698
rect 390268 -21840 390339 -21784
rect 390395 -21840 390481 -21784
rect 390537 -21840 390608 -21784
rect 390268 -21926 390608 -21840
rect 390268 -21982 390339 -21926
rect 390395 -21982 390481 -21926
rect 390537 -21982 390608 -21926
rect 390268 -22068 390608 -21982
rect 390268 -22124 390339 -22068
rect 390395 -22124 390481 -22068
rect 390537 -22124 390608 -22068
rect 390268 -22210 390608 -22124
rect 390268 -22266 390339 -22210
rect 390395 -22266 390481 -22210
rect 390537 -22266 390608 -22210
rect 390268 -22352 390608 -22266
rect 390268 -22408 390339 -22352
rect 390395 -22408 390481 -22352
rect 390537 -22408 390608 -22352
rect 390268 -22494 390608 -22408
rect 390268 -22550 390339 -22494
rect 390395 -22550 390481 -22494
rect 390537 -22550 390608 -22494
rect 390268 -22636 390608 -22550
rect 390268 -22692 390339 -22636
rect 390395 -22692 390481 -22636
rect 390537 -22692 390608 -22636
rect 390268 -22778 390608 -22692
rect 390268 -22834 390339 -22778
rect 390395 -22834 390481 -22778
rect 390537 -22834 390608 -22778
rect 390268 -22920 390608 -22834
rect 390268 -22976 390339 -22920
rect 390395 -22976 390481 -22920
rect 390537 -22976 390608 -22920
rect 390268 -23062 390608 -22976
rect 390268 -23118 390339 -23062
rect 390395 -23118 390481 -23062
rect 390537 -23118 390608 -23062
rect 390268 -23204 390608 -23118
rect 390268 -23260 390339 -23204
rect 390395 -23260 390481 -23204
rect 390537 -23260 390608 -23204
rect 390268 -23346 390608 -23260
rect 390268 -23402 390339 -23346
rect 390395 -23402 390481 -23346
rect 390537 -23402 390608 -23346
rect 390268 -23488 390608 -23402
rect 390268 -23544 390339 -23488
rect 390395 -23544 390481 -23488
rect 390537 -23544 390608 -23488
rect 390268 -23630 390608 -23544
rect 390268 -23686 390339 -23630
rect 390395 -23686 390481 -23630
rect 390537 -23686 390608 -23630
rect 390268 -23772 390608 -23686
rect 390268 -23828 390339 -23772
rect 390395 -23828 390481 -23772
rect 390537 -23828 390608 -23772
rect 390268 -23914 390608 -23828
rect 390268 -23970 390339 -23914
rect 390395 -23970 390481 -23914
rect 390537 -23970 390608 -23914
rect 390268 -24056 390608 -23970
rect 390268 -24112 390339 -24056
rect 390395 -24112 390481 -24056
rect 390537 -24112 390608 -24056
rect 390268 -24198 390608 -24112
rect 390268 -24254 390339 -24198
rect 390395 -24254 390481 -24198
rect 390537 -24254 390608 -24198
rect 390268 -24340 390608 -24254
rect 390268 -24396 390339 -24340
rect 390395 -24396 390481 -24340
rect 390537 -24396 390608 -24340
rect 390268 -24482 390608 -24396
rect 390268 -24538 390339 -24482
rect 390395 -24538 390481 -24482
rect 390537 -24538 390608 -24482
rect 390268 -24624 390608 -24538
rect 390268 -24680 390339 -24624
rect 390395 -24680 390481 -24624
rect 390537 -24680 390608 -24624
rect 390268 -24766 390608 -24680
rect 390268 -24822 390339 -24766
rect 390395 -24822 390481 -24766
rect 390537 -24822 390608 -24766
rect 390268 -24908 390608 -24822
rect 390268 -24964 390339 -24908
rect 390395 -24964 390481 -24908
rect 390537 -24964 390608 -24908
rect 390268 -25050 390608 -24964
rect 390268 -25106 390339 -25050
rect 390395 -25106 390481 -25050
rect 390537 -25106 390608 -25050
rect 390268 -25192 390608 -25106
rect 390268 -25248 390339 -25192
rect 390395 -25248 390481 -25192
rect 390537 -25248 390608 -25192
rect 390268 -25334 390608 -25248
rect 390268 -25390 390339 -25334
rect 390395 -25390 390481 -25334
rect 390537 -25390 390608 -25334
rect 390268 -25476 390608 -25390
rect 390268 -25532 390339 -25476
rect 390395 -25532 390481 -25476
rect 390537 -25532 390608 -25476
rect 390268 -25542 390608 -25532
rect 390668 -17950 391008 -17820
rect 390668 -18006 390736 -17950
rect 390792 -18006 390878 -17950
rect 390934 -18006 391008 -17950
rect 390668 -18092 391008 -18006
rect 390668 -18148 390736 -18092
rect 390792 -18148 390878 -18092
rect 390934 -18148 391008 -18092
rect 390668 -18234 391008 -18148
rect 390668 -18290 390736 -18234
rect 390792 -18290 390878 -18234
rect 390934 -18290 391008 -18234
rect 390668 -18376 391008 -18290
rect 390668 -18432 390736 -18376
rect 390792 -18432 390878 -18376
rect 390934 -18432 391008 -18376
rect 390668 -18518 391008 -18432
rect 390668 -18574 390736 -18518
rect 390792 -18574 390878 -18518
rect 390934 -18574 391008 -18518
rect 390668 -18660 391008 -18574
rect 390668 -18716 390736 -18660
rect 390792 -18716 390878 -18660
rect 390934 -18716 391008 -18660
rect 390668 -18802 391008 -18716
rect 390668 -18858 390736 -18802
rect 390792 -18858 390878 -18802
rect 390934 -18858 391008 -18802
rect 390668 -18944 391008 -18858
rect 390668 -19000 390736 -18944
rect 390792 -19000 390878 -18944
rect 390934 -19000 391008 -18944
rect 390668 -19086 391008 -19000
rect 390668 -19142 390736 -19086
rect 390792 -19142 390878 -19086
rect 390934 -19142 391008 -19086
rect 390668 -19228 391008 -19142
rect 390668 -19284 390736 -19228
rect 390792 -19284 390878 -19228
rect 390934 -19284 391008 -19228
rect 390668 -19370 391008 -19284
rect 390668 -19426 390736 -19370
rect 390792 -19426 390878 -19370
rect 390934 -19426 391008 -19370
rect 390668 -19512 391008 -19426
rect 390668 -19568 390736 -19512
rect 390792 -19568 390878 -19512
rect 390934 -19568 391008 -19512
rect 390668 -19654 391008 -19568
rect 390668 -19710 390736 -19654
rect 390792 -19710 390878 -19654
rect 390934 -19710 391008 -19654
rect 390668 -19796 391008 -19710
rect 390668 -19852 390736 -19796
rect 390792 -19852 390878 -19796
rect 390934 -19852 391008 -19796
rect 390668 -19938 391008 -19852
rect 390668 -19994 390736 -19938
rect 390792 -19994 390878 -19938
rect 390934 -19994 391008 -19938
rect 390668 -20080 391008 -19994
rect 390668 -20136 390736 -20080
rect 390792 -20136 390878 -20080
rect 390934 -20136 391008 -20080
rect 390668 -20222 391008 -20136
rect 390668 -20278 390736 -20222
rect 390792 -20278 390878 -20222
rect 390934 -20278 391008 -20222
rect 390668 -20364 391008 -20278
rect 390668 -20420 390736 -20364
rect 390792 -20420 390878 -20364
rect 390934 -20420 391008 -20364
rect 390668 -20506 391008 -20420
rect 390668 -20562 390736 -20506
rect 390792 -20562 390878 -20506
rect 390934 -20562 391008 -20506
rect 390668 -20648 391008 -20562
rect 390668 -20704 390736 -20648
rect 390792 -20704 390878 -20648
rect 390934 -20704 391008 -20648
rect 390668 -20790 391008 -20704
rect 390668 -20846 390736 -20790
rect 390792 -20846 390878 -20790
rect 390934 -20846 391008 -20790
rect 390668 -20932 391008 -20846
rect 390668 -20988 390736 -20932
rect 390792 -20988 390878 -20932
rect 390934 -20988 391008 -20932
rect 390668 -21074 391008 -20988
rect 390668 -21130 390736 -21074
rect 390792 -21130 390878 -21074
rect 390934 -21130 391008 -21074
rect 390668 -21216 391008 -21130
rect 390668 -21272 390736 -21216
rect 390792 -21272 390878 -21216
rect 390934 -21272 391008 -21216
rect 390668 -21358 391008 -21272
rect 390668 -21414 390736 -21358
rect 390792 -21414 390878 -21358
rect 390934 -21414 391008 -21358
rect 390668 -21500 391008 -21414
rect 390668 -21556 390736 -21500
rect 390792 -21556 390878 -21500
rect 390934 -21556 391008 -21500
rect 390668 -21642 391008 -21556
rect 390668 -21698 390736 -21642
rect 390792 -21698 390878 -21642
rect 390934 -21698 391008 -21642
rect 390668 -21784 391008 -21698
rect 390668 -21840 390736 -21784
rect 390792 -21840 390878 -21784
rect 390934 -21840 391008 -21784
rect 390668 -21926 391008 -21840
rect 390668 -21982 390736 -21926
rect 390792 -21982 390878 -21926
rect 390934 -21982 391008 -21926
rect 390668 -22068 391008 -21982
rect 390668 -22124 390736 -22068
rect 390792 -22124 390878 -22068
rect 390934 -22124 391008 -22068
rect 390668 -22210 391008 -22124
rect 390668 -22266 390736 -22210
rect 390792 -22266 390878 -22210
rect 390934 -22266 391008 -22210
rect 390668 -22352 391008 -22266
rect 390668 -22408 390736 -22352
rect 390792 -22408 390878 -22352
rect 390934 -22408 391008 -22352
rect 390668 -22494 391008 -22408
rect 390668 -22550 390736 -22494
rect 390792 -22550 390878 -22494
rect 390934 -22550 391008 -22494
rect 390668 -22636 391008 -22550
rect 390668 -22692 390736 -22636
rect 390792 -22692 390878 -22636
rect 390934 -22692 391008 -22636
rect 390668 -22778 391008 -22692
rect 390668 -22834 390736 -22778
rect 390792 -22834 390878 -22778
rect 390934 -22834 391008 -22778
rect 390668 -22920 391008 -22834
rect 390668 -22976 390736 -22920
rect 390792 -22976 390878 -22920
rect 390934 -22976 391008 -22920
rect 390668 -23062 391008 -22976
rect 390668 -23118 390736 -23062
rect 390792 -23118 390878 -23062
rect 390934 -23118 391008 -23062
rect 390668 -23204 391008 -23118
rect 390668 -23260 390736 -23204
rect 390792 -23260 390878 -23204
rect 390934 -23260 391008 -23204
rect 390668 -23346 391008 -23260
rect 390668 -23402 390736 -23346
rect 390792 -23402 390878 -23346
rect 390934 -23402 391008 -23346
rect 390668 -23488 391008 -23402
rect 390668 -23544 390736 -23488
rect 390792 -23544 390878 -23488
rect 390934 -23544 391008 -23488
rect 390668 -23630 391008 -23544
rect 390668 -23686 390736 -23630
rect 390792 -23686 390878 -23630
rect 390934 -23686 391008 -23630
rect 390668 -23772 391008 -23686
rect 390668 -23828 390736 -23772
rect 390792 -23828 390878 -23772
rect 390934 -23828 391008 -23772
rect 390668 -23914 391008 -23828
rect 390668 -23970 390736 -23914
rect 390792 -23970 390878 -23914
rect 390934 -23970 391008 -23914
rect 390668 -24056 391008 -23970
rect 390668 -24112 390736 -24056
rect 390792 -24112 390878 -24056
rect 390934 -24112 391008 -24056
rect 390668 -24198 391008 -24112
rect 390668 -24254 390736 -24198
rect 390792 -24254 390878 -24198
rect 390934 -24254 391008 -24198
rect 390668 -24340 391008 -24254
rect 390668 -24396 390736 -24340
rect 390792 -24396 390878 -24340
rect 390934 -24396 391008 -24340
rect 390668 -24482 391008 -24396
rect 390668 -24538 390736 -24482
rect 390792 -24538 390878 -24482
rect 390934 -24538 391008 -24482
rect 390668 -24624 391008 -24538
rect 390668 -24680 390736 -24624
rect 390792 -24680 390878 -24624
rect 390934 -24680 391008 -24624
rect 390668 -24766 391008 -24680
rect 390668 -24822 390736 -24766
rect 390792 -24822 390878 -24766
rect 390934 -24822 391008 -24766
rect 390668 -24908 391008 -24822
rect 390668 -24964 390736 -24908
rect 390792 -24964 390878 -24908
rect 390934 -24964 391008 -24908
rect 390668 -25050 391008 -24964
rect 390668 -25106 390736 -25050
rect 390792 -25106 390878 -25050
rect 390934 -25106 391008 -25050
rect 390668 -25192 391008 -25106
rect 390668 -25248 390736 -25192
rect 390792 -25248 390878 -25192
rect 390934 -25248 391008 -25192
rect 390668 -25334 391008 -25248
rect 390668 -25390 390736 -25334
rect 390792 -25390 390878 -25334
rect 390934 -25390 391008 -25334
rect 390668 -25476 391008 -25390
rect 390668 -25532 390736 -25476
rect 390792 -25532 390878 -25476
rect 390934 -25532 391008 -25476
rect 390668 -25542 391008 -25532
rect 391068 -17950 391408 -17820
rect 391068 -18006 391140 -17950
rect 391196 -18006 391282 -17950
rect 391338 -18006 391408 -17950
rect 391068 -18092 391408 -18006
rect 391068 -18148 391140 -18092
rect 391196 -18148 391282 -18092
rect 391338 -18148 391408 -18092
rect 391068 -18234 391408 -18148
rect 391068 -18290 391140 -18234
rect 391196 -18290 391282 -18234
rect 391338 -18290 391408 -18234
rect 391068 -18376 391408 -18290
rect 391068 -18432 391140 -18376
rect 391196 -18432 391282 -18376
rect 391338 -18432 391408 -18376
rect 391068 -18518 391408 -18432
rect 391068 -18574 391140 -18518
rect 391196 -18574 391282 -18518
rect 391338 -18574 391408 -18518
rect 391068 -18660 391408 -18574
rect 391068 -18716 391140 -18660
rect 391196 -18716 391282 -18660
rect 391338 -18716 391408 -18660
rect 391068 -18802 391408 -18716
rect 391068 -18858 391140 -18802
rect 391196 -18858 391282 -18802
rect 391338 -18858 391408 -18802
rect 391068 -18944 391408 -18858
rect 391068 -19000 391140 -18944
rect 391196 -19000 391282 -18944
rect 391338 -19000 391408 -18944
rect 391068 -19086 391408 -19000
rect 391068 -19142 391140 -19086
rect 391196 -19142 391282 -19086
rect 391338 -19142 391408 -19086
rect 391068 -19228 391408 -19142
rect 391068 -19284 391140 -19228
rect 391196 -19284 391282 -19228
rect 391338 -19284 391408 -19228
rect 391068 -19370 391408 -19284
rect 391068 -19426 391140 -19370
rect 391196 -19426 391282 -19370
rect 391338 -19426 391408 -19370
rect 391068 -19512 391408 -19426
rect 391068 -19568 391140 -19512
rect 391196 -19568 391282 -19512
rect 391338 -19568 391408 -19512
rect 391068 -19654 391408 -19568
rect 391068 -19710 391140 -19654
rect 391196 -19710 391282 -19654
rect 391338 -19710 391408 -19654
rect 391068 -19796 391408 -19710
rect 391068 -19852 391140 -19796
rect 391196 -19852 391282 -19796
rect 391338 -19852 391408 -19796
rect 391068 -19938 391408 -19852
rect 391068 -19994 391140 -19938
rect 391196 -19994 391282 -19938
rect 391338 -19994 391408 -19938
rect 391068 -20080 391408 -19994
rect 391068 -20136 391140 -20080
rect 391196 -20136 391282 -20080
rect 391338 -20136 391408 -20080
rect 391068 -20222 391408 -20136
rect 391068 -20278 391140 -20222
rect 391196 -20278 391282 -20222
rect 391338 -20278 391408 -20222
rect 391068 -20364 391408 -20278
rect 391068 -20420 391140 -20364
rect 391196 -20420 391282 -20364
rect 391338 -20420 391408 -20364
rect 391068 -20506 391408 -20420
rect 391068 -20562 391140 -20506
rect 391196 -20562 391282 -20506
rect 391338 -20562 391408 -20506
rect 391068 -20648 391408 -20562
rect 391068 -20704 391140 -20648
rect 391196 -20704 391282 -20648
rect 391338 -20704 391408 -20648
rect 391068 -20790 391408 -20704
rect 391068 -20846 391140 -20790
rect 391196 -20846 391282 -20790
rect 391338 -20846 391408 -20790
rect 391068 -20932 391408 -20846
rect 391068 -20988 391140 -20932
rect 391196 -20988 391282 -20932
rect 391338 -20988 391408 -20932
rect 391068 -21074 391408 -20988
rect 391068 -21130 391140 -21074
rect 391196 -21130 391282 -21074
rect 391338 -21130 391408 -21074
rect 391068 -21216 391408 -21130
rect 391068 -21272 391140 -21216
rect 391196 -21272 391282 -21216
rect 391338 -21272 391408 -21216
rect 391068 -21358 391408 -21272
rect 391068 -21414 391140 -21358
rect 391196 -21414 391282 -21358
rect 391338 -21414 391408 -21358
rect 391068 -21500 391408 -21414
rect 391068 -21556 391140 -21500
rect 391196 -21556 391282 -21500
rect 391338 -21556 391408 -21500
rect 391068 -21642 391408 -21556
rect 391068 -21698 391140 -21642
rect 391196 -21698 391282 -21642
rect 391338 -21698 391408 -21642
rect 391068 -21784 391408 -21698
rect 391068 -21840 391140 -21784
rect 391196 -21840 391282 -21784
rect 391338 -21840 391408 -21784
rect 391068 -21926 391408 -21840
rect 391068 -21982 391140 -21926
rect 391196 -21982 391282 -21926
rect 391338 -21982 391408 -21926
rect 391068 -22068 391408 -21982
rect 391068 -22124 391140 -22068
rect 391196 -22124 391282 -22068
rect 391338 -22124 391408 -22068
rect 391068 -22210 391408 -22124
rect 391068 -22266 391140 -22210
rect 391196 -22266 391282 -22210
rect 391338 -22266 391408 -22210
rect 391068 -22352 391408 -22266
rect 391068 -22408 391140 -22352
rect 391196 -22408 391282 -22352
rect 391338 -22408 391408 -22352
rect 391068 -22494 391408 -22408
rect 391068 -22550 391140 -22494
rect 391196 -22550 391282 -22494
rect 391338 -22550 391408 -22494
rect 391068 -22636 391408 -22550
rect 391068 -22692 391140 -22636
rect 391196 -22692 391282 -22636
rect 391338 -22692 391408 -22636
rect 391068 -22778 391408 -22692
rect 391068 -22834 391140 -22778
rect 391196 -22834 391282 -22778
rect 391338 -22834 391408 -22778
rect 391068 -22920 391408 -22834
rect 391068 -22976 391140 -22920
rect 391196 -22976 391282 -22920
rect 391338 -22976 391408 -22920
rect 391068 -23062 391408 -22976
rect 391068 -23118 391140 -23062
rect 391196 -23118 391282 -23062
rect 391338 -23118 391408 -23062
rect 391068 -23204 391408 -23118
rect 391068 -23260 391140 -23204
rect 391196 -23260 391282 -23204
rect 391338 -23260 391408 -23204
rect 391068 -23346 391408 -23260
rect 391068 -23402 391140 -23346
rect 391196 -23402 391282 -23346
rect 391338 -23402 391408 -23346
rect 391068 -23488 391408 -23402
rect 391068 -23544 391140 -23488
rect 391196 -23544 391282 -23488
rect 391338 -23544 391408 -23488
rect 391068 -23630 391408 -23544
rect 391068 -23686 391140 -23630
rect 391196 -23686 391282 -23630
rect 391338 -23686 391408 -23630
rect 391068 -23772 391408 -23686
rect 391068 -23828 391140 -23772
rect 391196 -23828 391282 -23772
rect 391338 -23828 391408 -23772
rect 391068 -23914 391408 -23828
rect 391068 -23970 391140 -23914
rect 391196 -23970 391282 -23914
rect 391338 -23970 391408 -23914
rect 391068 -24056 391408 -23970
rect 391068 -24112 391140 -24056
rect 391196 -24112 391282 -24056
rect 391338 -24112 391408 -24056
rect 391068 -24198 391408 -24112
rect 391068 -24254 391140 -24198
rect 391196 -24254 391282 -24198
rect 391338 -24254 391408 -24198
rect 391068 -24340 391408 -24254
rect 391068 -24396 391140 -24340
rect 391196 -24396 391282 -24340
rect 391338 -24396 391408 -24340
rect 391068 -24482 391408 -24396
rect 391068 -24538 391140 -24482
rect 391196 -24538 391282 -24482
rect 391338 -24538 391408 -24482
rect 391068 -24624 391408 -24538
rect 391068 -24680 391140 -24624
rect 391196 -24680 391282 -24624
rect 391338 -24680 391408 -24624
rect 391068 -24766 391408 -24680
rect 391068 -24822 391140 -24766
rect 391196 -24822 391282 -24766
rect 391338 -24822 391408 -24766
rect 391068 -24908 391408 -24822
rect 391068 -24964 391140 -24908
rect 391196 -24964 391282 -24908
rect 391338 -24964 391408 -24908
rect 391068 -25050 391408 -24964
rect 391068 -25106 391140 -25050
rect 391196 -25106 391282 -25050
rect 391338 -25106 391408 -25050
rect 391068 -25192 391408 -25106
rect 391068 -25248 391140 -25192
rect 391196 -25248 391282 -25192
rect 391338 -25248 391408 -25192
rect 391068 -25334 391408 -25248
rect 391068 -25390 391140 -25334
rect 391196 -25390 391282 -25334
rect 391338 -25390 391408 -25334
rect 391068 -25476 391408 -25390
rect 391068 -25532 391140 -25476
rect 391196 -25532 391282 -25476
rect 391338 -25532 391408 -25476
rect 391068 -25542 391408 -25532
rect 391468 -17950 391808 -17820
rect 391468 -18006 391536 -17950
rect 391592 -18006 391678 -17950
rect 391734 -18006 391808 -17950
rect 391468 -18092 391808 -18006
rect 391468 -18148 391536 -18092
rect 391592 -18148 391678 -18092
rect 391734 -18148 391808 -18092
rect 391468 -18234 391808 -18148
rect 391468 -18290 391536 -18234
rect 391592 -18290 391678 -18234
rect 391734 -18290 391808 -18234
rect 391468 -18376 391808 -18290
rect 391468 -18432 391536 -18376
rect 391592 -18432 391678 -18376
rect 391734 -18432 391808 -18376
rect 391468 -18518 391808 -18432
rect 391468 -18574 391536 -18518
rect 391592 -18574 391678 -18518
rect 391734 -18574 391808 -18518
rect 391468 -18660 391808 -18574
rect 391468 -18716 391536 -18660
rect 391592 -18716 391678 -18660
rect 391734 -18716 391808 -18660
rect 391468 -18802 391808 -18716
rect 391468 -18858 391536 -18802
rect 391592 -18858 391678 -18802
rect 391734 -18858 391808 -18802
rect 391468 -18944 391808 -18858
rect 391468 -19000 391536 -18944
rect 391592 -19000 391678 -18944
rect 391734 -19000 391808 -18944
rect 391468 -19086 391808 -19000
rect 391468 -19142 391536 -19086
rect 391592 -19142 391678 -19086
rect 391734 -19142 391808 -19086
rect 391468 -19228 391808 -19142
rect 391468 -19284 391536 -19228
rect 391592 -19284 391678 -19228
rect 391734 -19284 391808 -19228
rect 391468 -19370 391808 -19284
rect 391468 -19426 391536 -19370
rect 391592 -19426 391678 -19370
rect 391734 -19426 391808 -19370
rect 391468 -19512 391808 -19426
rect 391468 -19568 391536 -19512
rect 391592 -19568 391678 -19512
rect 391734 -19568 391808 -19512
rect 391468 -19654 391808 -19568
rect 391468 -19710 391536 -19654
rect 391592 -19710 391678 -19654
rect 391734 -19710 391808 -19654
rect 391468 -19796 391808 -19710
rect 391468 -19852 391536 -19796
rect 391592 -19852 391678 -19796
rect 391734 -19852 391808 -19796
rect 391468 -19938 391808 -19852
rect 391468 -19994 391536 -19938
rect 391592 -19994 391678 -19938
rect 391734 -19994 391808 -19938
rect 391468 -20080 391808 -19994
rect 391468 -20136 391536 -20080
rect 391592 -20136 391678 -20080
rect 391734 -20136 391808 -20080
rect 391468 -20222 391808 -20136
rect 391468 -20278 391536 -20222
rect 391592 -20278 391678 -20222
rect 391734 -20278 391808 -20222
rect 391468 -20364 391808 -20278
rect 391468 -20420 391536 -20364
rect 391592 -20420 391678 -20364
rect 391734 -20420 391808 -20364
rect 391468 -20506 391808 -20420
rect 391468 -20562 391536 -20506
rect 391592 -20562 391678 -20506
rect 391734 -20562 391808 -20506
rect 391468 -20648 391808 -20562
rect 391468 -20704 391536 -20648
rect 391592 -20704 391678 -20648
rect 391734 -20704 391808 -20648
rect 391468 -20790 391808 -20704
rect 391468 -20846 391536 -20790
rect 391592 -20846 391678 -20790
rect 391734 -20846 391808 -20790
rect 391468 -20932 391808 -20846
rect 391468 -20988 391536 -20932
rect 391592 -20988 391678 -20932
rect 391734 -20988 391808 -20932
rect 391468 -21074 391808 -20988
rect 391468 -21130 391536 -21074
rect 391592 -21130 391678 -21074
rect 391734 -21130 391808 -21074
rect 391468 -21216 391808 -21130
rect 391468 -21272 391536 -21216
rect 391592 -21272 391678 -21216
rect 391734 -21272 391808 -21216
rect 391468 -21358 391808 -21272
rect 391468 -21414 391536 -21358
rect 391592 -21414 391678 -21358
rect 391734 -21414 391808 -21358
rect 391468 -21500 391808 -21414
rect 391468 -21556 391536 -21500
rect 391592 -21556 391678 -21500
rect 391734 -21556 391808 -21500
rect 391468 -21642 391808 -21556
rect 391468 -21698 391536 -21642
rect 391592 -21698 391678 -21642
rect 391734 -21698 391808 -21642
rect 391468 -21784 391808 -21698
rect 391468 -21840 391536 -21784
rect 391592 -21840 391678 -21784
rect 391734 -21840 391808 -21784
rect 391468 -21926 391808 -21840
rect 391468 -21982 391536 -21926
rect 391592 -21982 391678 -21926
rect 391734 -21982 391808 -21926
rect 391468 -22068 391808 -21982
rect 391468 -22124 391536 -22068
rect 391592 -22124 391678 -22068
rect 391734 -22124 391808 -22068
rect 391468 -22210 391808 -22124
rect 391468 -22266 391536 -22210
rect 391592 -22266 391678 -22210
rect 391734 -22266 391808 -22210
rect 391468 -22352 391808 -22266
rect 391468 -22408 391536 -22352
rect 391592 -22408 391678 -22352
rect 391734 -22408 391808 -22352
rect 391468 -22494 391808 -22408
rect 391468 -22550 391536 -22494
rect 391592 -22550 391678 -22494
rect 391734 -22550 391808 -22494
rect 391468 -22636 391808 -22550
rect 391468 -22692 391536 -22636
rect 391592 -22692 391678 -22636
rect 391734 -22692 391808 -22636
rect 391468 -22778 391808 -22692
rect 391468 -22834 391536 -22778
rect 391592 -22834 391678 -22778
rect 391734 -22834 391808 -22778
rect 391468 -22920 391808 -22834
rect 391468 -22976 391536 -22920
rect 391592 -22976 391678 -22920
rect 391734 -22976 391808 -22920
rect 391468 -23062 391808 -22976
rect 391468 -23118 391536 -23062
rect 391592 -23118 391678 -23062
rect 391734 -23118 391808 -23062
rect 391468 -23204 391808 -23118
rect 391468 -23260 391536 -23204
rect 391592 -23260 391678 -23204
rect 391734 -23260 391808 -23204
rect 391468 -23346 391808 -23260
rect 391468 -23402 391536 -23346
rect 391592 -23402 391678 -23346
rect 391734 -23402 391808 -23346
rect 391468 -23488 391808 -23402
rect 391468 -23544 391536 -23488
rect 391592 -23544 391678 -23488
rect 391734 -23544 391808 -23488
rect 391468 -23630 391808 -23544
rect 391468 -23686 391536 -23630
rect 391592 -23686 391678 -23630
rect 391734 -23686 391808 -23630
rect 391468 -23772 391808 -23686
rect 391468 -23828 391536 -23772
rect 391592 -23828 391678 -23772
rect 391734 -23828 391808 -23772
rect 391468 -23914 391808 -23828
rect 391468 -23970 391536 -23914
rect 391592 -23970 391678 -23914
rect 391734 -23970 391808 -23914
rect 391468 -24056 391808 -23970
rect 391468 -24112 391536 -24056
rect 391592 -24112 391678 -24056
rect 391734 -24112 391808 -24056
rect 391468 -24198 391808 -24112
rect 391468 -24254 391536 -24198
rect 391592 -24254 391678 -24198
rect 391734 -24254 391808 -24198
rect 391468 -24340 391808 -24254
rect 391468 -24396 391536 -24340
rect 391592 -24396 391678 -24340
rect 391734 -24396 391808 -24340
rect 391468 -24482 391808 -24396
rect 391468 -24538 391536 -24482
rect 391592 -24538 391678 -24482
rect 391734 -24538 391808 -24482
rect 391468 -24624 391808 -24538
rect 391468 -24680 391536 -24624
rect 391592 -24680 391678 -24624
rect 391734 -24680 391808 -24624
rect 391468 -24766 391808 -24680
rect 391468 -24822 391536 -24766
rect 391592 -24822 391678 -24766
rect 391734 -24822 391808 -24766
rect 391468 -24908 391808 -24822
rect 391468 -24964 391536 -24908
rect 391592 -24964 391678 -24908
rect 391734 -24964 391808 -24908
rect 391468 -25050 391808 -24964
rect 391468 -25106 391536 -25050
rect 391592 -25106 391678 -25050
rect 391734 -25106 391808 -25050
rect 391468 -25192 391808 -25106
rect 391468 -25248 391536 -25192
rect 391592 -25248 391678 -25192
rect 391734 -25248 391808 -25192
rect 391468 -25334 391808 -25248
rect 391468 -25390 391536 -25334
rect 391592 -25390 391678 -25334
rect 391734 -25390 391808 -25334
rect 391468 -25476 391808 -25390
rect 391468 -25532 391536 -25476
rect 391592 -25532 391678 -25476
rect 391734 -25532 391808 -25476
rect 391468 -25542 391808 -25532
rect 391868 -17950 392208 -17820
rect 391868 -18006 391936 -17950
rect 391992 -18006 392078 -17950
rect 392134 -18006 392208 -17950
rect 391868 -18092 392208 -18006
rect 391868 -18148 391936 -18092
rect 391992 -18148 392078 -18092
rect 392134 -18148 392208 -18092
rect 391868 -18234 392208 -18148
rect 391868 -18290 391936 -18234
rect 391992 -18290 392078 -18234
rect 392134 -18290 392208 -18234
rect 391868 -18376 392208 -18290
rect 391868 -18432 391936 -18376
rect 391992 -18432 392078 -18376
rect 392134 -18432 392208 -18376
rect 391868 -18518 392208 -18432
rect 391868 -18574 391936 -18518
rect 391992 -18574 392078 -18518
rect 392134 -18574 392208 -18518
rect 391868 -18660 392208 -18574
rect 391868 -18716 391936 -18660
rect 391992 -18716 392078 -18660
rect 392134 -18716 392208 -18660
rect 391868 -18802 392208 -18716
rect 391868 -18858 391936 -18802
rect 391992 -18858 392078 -18802
rect 392134 -18858 392208 -18802
rect 391868 -18944 392208 -18858
rect 391868 -19000 391936 -18944
rect 391992 -19000 392078 -18944
rect 392134 -19000 392208 -18944
rect 391868 -19086 392208 -19000
rect 391868 -19142 391936 -19086
rect 391992 -19142 392078 -19086
rect 392134 -19142 392208 -19086
rect 391868 -19228 392208 -19142
rect 391868 -19284 391936 -19228
rect 391992 -19284 392078 -19228
rect 392134 -19284 392208 -19228
rect 391868 -19370 392208 -19284
rect 391868 -19426 391936 -19370
rect 391992 -19426 392078 -19370
rect 392134 -19426 392208 -19370
rect 391868 -19512 392208 -19426
rect 391868 -19568 391936 -19512
rect 391992 -19568 392078 -19512
rect 392134 -19568 392208 -19512
rect 391868 -19654 392208 -19568
rect 391868 -19710 391936 -19654
rect 391992 -19710 392078 -19654
rect 392134 -19710 392208 -19654
rect 391868 -19796 392208 -19710
rect 391868 -19852 391936 -19796
rect 391992 -19852 392078 -19796
rect 392134 -19852 392208 -19796
rect 391868 -19938 392208 -19852
rect 391868 -19994 391936 -19938
rect 391992 -19994 392078 -19938
rect 392134 -19994 392208 -19938
rect 391868 -20080 392208 -19994
rect 391868 -20136 391936 -20080
rect 391992 -20136 392078 -20080
rect 392134 -20136 392208 -20080
rect 391868 -20222 392208 -20136
rect 391868 -20278 391936 -20222
rect 391992 -20278 392078 -20222
rect 392134 -20278 392208 -20222
rect 391868 -20364 392208 -20278
rect 391868 -20420 391936 -20364
rect 391992 -20420 392078 -20364
rect 392134 -20420 392208 -20364
rect 391868 -20506 392208 -20420
rect 391868 -20562 391936 -20506
rect 391992 -20562 392078 -20506
rect 392134 -20562 392208 -20506
rect 391868 -20648 392208 -20562
rect 391868 -20704 391936 -20648
rect 391992 -20704 392078 -20648
rect 392134 -20704 392208 -20648
rect 391868 -20790 392208 -20704
rect 391868 -20846 391936 -20790
rect 391992 -20846 392078 -20790
rect 392134 -20846 392208 -20790
rect 391868 -20932 392208 -20846
rect 391868 -20988 391936 -20932
rect 391992 -20988 392078 -20932
rect 392134 -20988 392208 -20932
rect 391868 -21074 392208 -20988
rect 391868 -21130 391936 -21074
rect 391992 -21130 392078 -21074
rect 392134 -21130 392208 -21074
rect 391868 -21216 392208 -21130
rect 391868 -21272 391936 -21216
rect 391992 -21272 392078 -21216
rect 392134 -21272 392208 -21216
rect 391868 -21358 392208 -21272
rect 391868 -21414 391936 -21358
rect 391992 -21414 392078 -21358
rect 392134 -21414 392208 -21358
rect 391868 -21500 392208 -21414
rect 391868 -21556 391936 -21500
rect 391992 -21556 392078 -21500
rect 392134 -21556 392208 -21500
rect 391868 -21642 392208 -21556
rect 391868 -21698 391936 -21642
rect 391992 -21698 392078 -21642
rect 392134 -21698 392208 -21642
rect 391868 -21784 392208 -21698
rect 391868 -21840 391936 -21784
rect 391992 -21840 392078 -21784
rect 392134 -21840 392208 -21784
rect 391868 -21926 392208 -21840
rect 391868 -21982 391936 -21926
rect 391992 -21982 392078 -21926
rect 392134 -21982 392208 -21926
rect 391868 -22068 392208 -21982
rect 391868 -22124 391936 -22068
rect 391992 -22124 392078 -22068
rect 392134 -22124 392208 -22068
rect 391868 -22210 392208 -22124
rect 391868 -22266 391936 -22210
rect 391992 -22266 392078 -22210
rect 392134 -22266 392208 -22210
rect 391868 -22352 392208 -22266
rect 391868 -22408 391936 -22352
rect 391992 -22408 392078 -22352
rect 392134 -22408 392208 -22352
rect 391868 -22494 392208 -22408
rect 391868 -22550 391936 -22494
rect 391992 -22550 392078 -22494
rect 392134 -22550 392208 -22494
rect 391868 -22636 392208 -22550
rect 391868 -22692 391936 -22636
rect 391992 -22692 392078 -22636
rect 392134 -22692 392208 -22636
rect 391868 -22778 392208 -22692
rect 391868 -22834 391936 -22778
rect 391992 -22834 392078 -22778
rect 392134 -22834 392208 -22778
rect 391868 -22920 392208 -22834
rect 391868 -22976 391936 -22920
rect 391992 -22976 392078 -22920
rect 392134 -22976 392208 -22920
rect 391868 -23062 392208 -22976
rect 391868 -23118 391936 -23062
rect 391992 -23118 392078 -23062
rect 392134 -23118 392208 -23062
rect 391868 -23204 392208 -23118
rect 391868 -23260 391936 -23204
rect 391992 -23260 392078 -23204
rect 392134 -23260 392208 -23204
rect 391868 -23346 392208 -23260
rect 391868 -23402 391936 -23346
rect 391992 -23402 392078 -23346
rect 392134 -23402 392208 -23346
rect 391868 -23488 392208 -23402
rect 391868 -23544 391936 -23488
rect 391992 -23544 392078 -23488
rect 392134 -23544 392208 -23488
rect 391868 -23630 392208 -23544
rect 391868 -23686 391936 -23630
rect 391992 -23686 392078 -23630
rect 392134 -23686 392208 -23630
rect 391868 -23772 392208 -23686
rect 391868 -23828 391936 -23772
rect 391992 -23828 392078 -23772
rect 392134 -23828 392208 -23772
rect 391868 -23914 392208 -23828
rect 391868 -23970 391936 -23914
rect 391992 -23970 392078 -23914
rect 392134 -23970 392208 -23914
rect 391868 -24056 392208 -23970
rect 391868 -24112 391936 -24056
rect 391992 -24112 392078 -24056
rect 392134 -24112 392208 -24056
rect 391868 -24198 392208 -24112
rect 391868 -24254 391936 -24198
rect 391992 -24254 392078 -24198
rect 392134 -24254 392208 -24198
rect 391868 -24340 392208 -24254
rect 391868 -24396 391936 -24340
rect 391992 -24396 392078 -24340
rect 392134 -24396 392208 -24340
rect 391868 -24482 392208 -24396
rect 391868 -24538 391936 -24482
rect 391992 -24538 392078 -24482
rect 392134 -24538 392208 -24482
rect 391868 -24624 392208 -24538
rect 391868 -24680 391936 -24624
rect 391992 -24680 392078 -24624
rect 392134 -24680 392208 -24624
rect 391868 -24766 392208 -24680
rect 391868 -24822 391936 -24766
rect 391992 -24822 392078 -24766
rect 392134 -24822 392208 -24766
rect 391868 -24908 392208 -24822
rect 391868 -24964 391936 -24908
rect 391992 -24964 392078 -24908
rect 392134 -24964 392208 -24908
rect 391868 -25050 392208 -24964
rect 391868 -25106 391936 -25050
rect 391992 -25106 392078 -25050
rect 392134 -25106 392208 -25050
rect 391868 -25192 392208 -25106
rect 391868 -25248 391936 -25192
rect 391992 -25248 392078 -25192
rect 392134 -25248 392208 -25192
rect 391868 -25334 392208 -25248
rect 391868 -25390 391936 -25334
rect 391992 -25390 392078 -25334
rect 392134 -25390 392208 -25334
rect 391868 -25476 392208 -25390
rect 391868 -25532 391936 -25476
rect 391992 -25532 392078 -25476
rect 392134 -25532 392208 -25476
rect 391868 -25542 392208 -25532
rect 392268 -17950 392608 -17820
rect 392268 -18006 392333 -17950
rect 392389 -18006 392475 -17950
rect 392531 -18006 392608 -17950
rect 392268 -18092 392608 -18006
rect 392268 -18148 392333 -18092
rect 392389 -18148 392475 -18092
rect 392531 -18148 392608 -18092
rect 392268 -18234 392608 -18148
rect 392268 -18290 392333 -18234
rect 392389 -18290 392475 -18234
rect 392531 -18290 392608 -18234
rect 392268 -18376 392608 -18290
rect 392268 -18432 392333 -18376
rect 392389 -18432 392475 -18376
rect 392531 -18432 392608 -18376
rect 392268 -18518 392608 -18432
rect 392268 -18574 392333 -18518
rect 392389 -18574 392475 -18518
rect 392531 -18574 392608 -18518
rect 392268 -18660 392608 -18574
rect 392268 -18716 392333 -18660
rect 392389 -18716 392475 -18660
rect 392531 -18716 392608 -18660
rect 392268 -18802 392608 -18716
rect 392268 -18858 392333 -18802
rect 392389 -18858 392475 -18802
rect 392531 -18858 392608 -18802
rect 392268 -18944 392608 -18858
rect 392268 -19000 392333 -18944
rect 392389 -19000 392475 -18944
rect 392531 -19000 392608 -18944
rect 392268 -19086 392608 -19000
rect 392268 -19142 392333 -19086
rect 392389 -19142 392475 -19086
rect 392531 -19142 392608 -19086
rect 392268 -19228 392608 -19142
rect 392268 -19284 392333 -19228
rect 392389 -19284 392475 -19228
rect 392531 -19284 392608 -19228
rect 392268 -19370 392608 -19284
rect 392268 -19426 392333 -19370
rect 392389 -19426 392475 -19370
rect 392531 -19426 392608 -19370
rect 392268 -19512 392608 -19426
rect 392268 -19568 392333 -19512
rect 392389 -19568 392475 -19512
rect 392531 -19568 392608 -19512
rect 392268 -19654 392608 -19568
rect 392268 -19710 392333 -19654
rect 392389 -19710 392475 -19654
rect 392531 -19710 392608 -19654
rect 392268 -19796 392608 -19710
rect 392268 -19852 392333 -19796
rect 392389 -19852 392475 -19796
rect 392531 -19852 392608 -19796
rect 392268 -19938 392608 -19852
rect 392268 -19994 392333 -19938
rect 392389 -19994 392475 -19938
rect 392531 -19994 392608 -19938
rect 392268 -20080 392608 -19994
rect 392268 -20136 392333 -20080
rect 392389 -20136 392475 -20080
rect 392531 -20136 392608 -20080
rect 392268 -20222 392608 -20136
rect 392268 -20278 392333 -20222
rect 392389 -20278 392475 -20222
rect 392531 -20278 392608 -20222
rect 392268 -20364 392608 -20278
rect 392268 -20420 392333 -20364
rect 392389 -20420 392475 -20364
rect 392531 -20420 392608 -20364
rect 392268 -20506 392608 -20420
rect 392268 -20562 392333 -20506
rect 392389 -20562 392475 -20506
rect 392531 -20562 392608 -20506
rect 392268 -20648 392608 -20562
rect 392268 -20704 392333 -20648
rect 392389 -20704 392475 -20648
rect 392531 -20704 392608 -20648
rect 392268 -20790 392608 -20704
rect 392268 -20846 392333 -20790
rect 392389 -20846 392475 -20790
rect 392531 -20846 392608 -20790
rect 392268 -20932 392608 -20846
rect 392268 -20988 392333 -20932
rect 392389 -20988 392475 -20932
rect 392531 -20988 392608 -20932
rect 392268 -21074 392608 -20988
rect 392268 -21130 392333 -21074
rect 392389 -21130 392475 -21074
rect 392531 -21130 392608 -21074
rect 392268 -21216 392608 -21130
rect 392268 -21272 392333 -21216
rect 392389 -21272 392475 -21216
rect 392531 -21272 392608 -21216
rect 392268 -21358 392608 -21272
rect 392268 -21414 392333 -21358
rect 392389 -21414 392475 -21358
rect 392531 -21414 392608 -21358
rect 392268 -21500 392608 -21414
rect 392268 -21556 392333 -21500
rect 392389 -21556 392475 -21500
rect 392531 -21556 392608 -21500
rect 392268 -21642 392608 -21556
rect 392268 -21698 392333 -21642
rect 392389 -21698 392475 -21642
rect 392531 -21698 392608 -21642
rect 392268 -21784 392608 -21698
rect 392268 -21840 392333 -21784
rect 392389 -21840 392475 -21784
rect 392531 -21840 392608 -21784
rect 392268 -21926 392608 -21840
rect 392268 -21982 392333 -21926
rect 392389 -21982 392475 -21926
rect 392531 -21982 392608 -21926
rect 392268 -22068 392608 -21982
rect 392268 -22124 392333 -22068
rect 392389 -22124 392475 -22068
rect 392531 -22124 392608 -22068
rect 392268 -22210 392608 -22124
rect 392268 -22266 392333 -22210
rect 392389 -22266 392475 -22210
rect 392531 -22266 392608 -22210
rect 392268 -22352 392608 -22266
rect 392268 -22408 392333 -22352
rect 392389 -22408 392475 -22352
rect 392531 -22408 392608 -22352
rect 392268 -22494 392608 -22408
rect 392268 -22550 392333 -22494
rect 392389 -22550 392475 -22494
rect 392531 -22550 392608 -22494
rect 392268 -22636 392608 -22550
rect 392268 -22692 392333 -22636
rect 392389 -22692 392475 -22636
rect 392531 -22692 392608 -22636
rect 392268 -22778 392608 -22692
rect 392268 -22834 392333 -22778
rect 392389 -22834 392475 -22778
rect 392531 -22834 392608 -22778
rect 392268 -22920 392608 -22834
rect 392268 -22976 392333 -22920
rect 392389 -22976 392475 -22920
rect 392531 -22976 392608 -22920
rect 392268 -23062 392608 -22976
rect 392268 -23118 392333 -23062
rect 392389 -23118 392475 -23062
rect 392531 -23118 392608 -23062
rect 392268 -23204 392608 -23118
rect 392268 -23260 392333 -23204
rect 392389 -23260 392475 -23204
rect 392531 -23260 392608 -23204
rect 392268 -23346 392608 -23260
rect 392268 -23402 392333 -23346
rect 392389 -23402 392475 -23346
rect 392531 -23402 392608 -23346
rect 392268 -23488 392608 -23402
rect 392268 -23544 392333 -23488
rect 392389 -23544 392475 -23488
rect 392531 -23544 392608 -23488
rect 392268 -23630 392608 -23544
rect 392268 -23686 392333 -23630
rect 392389 -23686 392475 -23630
rect 392531 -23686 392608 -23630
rect 392268 -23772 392608 -23686
rect 392268 -23828 392333 -23772
rect 392389 -23828 392475 -23772
rect 392531 -23828 392608 -23772
rect 392268 -23914 392608 -23828
rect 392268 -23970 392333 -23914
rect 392389 -23970 392475 -23914
rect 392531 -23970 392608 -23914
rect 392268 -24056 392608 -23970
rect 392268 -24112 392333 -24056
rect 392389 -24112 392475 -24056
rect 392531 -24112 392608 -24056
rect 392268 -24198 392608 -24112
rect 392268 -24254 392333 -24198
rect 392389 -24254 392475 -24198
rect 392531 -24254 392608 -24198
rect 392268 -24340 392608 -24254
rect 392268 -24396 392333 -24340
rect 392389 -24396 392475 -24340
rect 392531 -24396 392608 -24340
rect 392268 -24482 392608 -24396
rect 392268 -24538 392333 -24482
rect 392389 -24538 392475 -24482
rect 392531 -24538 392608 -24482
rect 392268 -24624 392608 -24538
rect 392268 -24680 392333 -24624
rect 392389 -24680 392475 -24624
rect 392531 -24680 392608 -24624
rect 392268 -24766 392608 -24680
rect 392268 -24822 392333 -24766
rect 392389 -24822 392475 -24766
rect 392531 -24822 392608 -24766
rect 392268 -24908 392608 -24822
rect 392268 -24964 392333 -24908
rect 392389 -24964 392475 -24908
rect 392531 -24964 392608 -24908
rect 392268 -25050 392608 -24964
rect 392268 -25106 392333 -25050
rect 392389 -25106 392475 -25050
rect 392531 -25106 392608 -25050
rect 392268 -25192 392608 -25106
rect 392268 -25248 392333 -25192
rect 392389 -25248 392475 -25192
rect 392531 -25248 392608 -25192
rect 392268 -25334 392608 -25248
rect 392268 -25390 392333 -25334
rect 392389 -25390 392475 -25334
rect 392531 -25390 392608 -25334
rect 392268 -25476 392608 -25390
rect 392268 -25532 392333 -25476
rect 392389 -25532 392475 -25476
rect 392531 -25532 392608 -25476
rect 392268 -25542 392608 -25532
rect 392668 -17950 393008 -17820
rect 392668 -18006 392738 -17950
rect 392794 -18006 392880 -17950
rect 392936 -18006 393008 -17950
rect 392668 -18092 393008 -18006
rect 392668 -18148 392738 -18092
rect 392794 -18148 392880 -18092
rect 392936 -18148 393008 -18092
rect 392668 -18234 393008 -18148
rect 392668 -18290 392738 -18234
rect 392794 -18290 392880 -18234
rect 392936 -18290 393008 -18234
rect 392668 -18376 393008 -18290
rect 392668 -18432 392738 -18376
rect 392794 -18432 392880 -18376
rect 392936 -18432 393008 -18376
rect 392668 -18518 393008 -18432
rect 392668 -18574 392738 -18518
rect 392794 -18574 392880 -18518
rect 392936 -18574 393008 -18518
rect 392668 -18660 393008 -18574
rect 392668 -18716 392738 -18660
rect 392794 -18716 392880 -18660
rect 392936 -18716 393008 -18660
rect 392668 -18802 393008 -18716
rect 392668 -18858 392738 -18802
rect 392794 -18858 392880 -18802
rect 392936 -18858 393008 -18802
rect 392668 -18944 393008 -18858
rect 392668 -19000 392738 -18944
rect 392794 -19000 392880 -18944
rect 392936 -19000 393008 -18944
rect 392668 -19086 393008 -19000
rect 392668 -19142 392738 -19086
rect 392794 -19142 392880 -19086
rect 392936 -19142 393008 -19086
rect 392668 -19228 393008 -19142
rect 392668 -19284 392738 -19228
rect 392794 -19284 392880 -19228
rect 392936 -19284 393008 -19228
rect 392668 -19370 393008 -19284
rect 392668 -19426 392738 -19370
rect 392794 -19426 392880 -19370
rect 392936 -19426 393008 -19370
rect 392668 -19512 393008 -19426
rect 392668 -19568 392738 -19512
rect 392794 -19568 392880 -19512
rect 392936 -19568 393008 -19512
rect 392668 -19654 393008 -19568
rect 392668 -19710 392738 -19654
rect 392794 -19710 392880 -19654
rect 392936 -19710 393008 -19654
rect 392668 -19796 393008 -19710
rect 392668 -19852 392738 -19796
rect 392794 -19852 392880 -19796
rect 392936 -19852 393008 -19796
rect 392668 -19938 393008 -19852
rect 392668 -19994 392738 -19938
rect 392794 -19994 392880 -19938
rect 392936 -19994 393008 -19938
rect 392668 -20080 393008 -19994
rect 392668 -20136 392738 -20080
rect 392794 -20136 392880 -20080
rect 392936 -20136 393008 -20080
rect 392668 -20222 393008 -20136
rect 392668 -20278 392738 -20222
rect 392794 -20278 392880 -20222
rect 392936 -20278 393008 -20222
rect 392668 -20364 393008 -20278
rect 392668 -20420 392738 -20364
rect 392794 -20420 392880 -20364
rect 392936 -20420 393008 -20364
rect 392668 -20506 393008 -20420
rect 392668 -20562 392738 -20506
rect 392794 -20562 392880 -20506
rect 392936 -20562 393008 -20506
rect 392668 -20648 393008 -20562
rect 392668 -20704 392738 -20648
rect 392794 -20704 392880 -20648
rect 392936 -20704 393008 -20648
rect 392668 -20790 393008 -20704
rect 392668 -20846 392738 -20790
rect 392794 -20846 392880 -20790
rect 392936 -20846 393008 -20790
rect 392668 -20932 393008 -20846
rect 392668 -20988 392738 -20932
rect 392794 -20988 392880 -20932
rect 392936 -20988 393008 -20932
rect 392668 -21074 393008 -20988
rect 392668 -21130 392738 -21074
rect 392794 -21130 392880 -21074
rect 392936 -21130 393008 -21074
rect 392668 -21216 393008 -21130
rect 392668 -21272 392738 -21216
rect 392794 -21272 392880 -21216
rect 392936 -21272 393008 -21216
rect 392668 -21358 393008 -21272
rect 392668 -21414 392738 -21358
rect 392794 -21414 392880 -21358
rect 392936 -21414 393008 -21358
rect 392668 -21500 393008 -21414
rect 392668 -21556 392738 -21500
rect 392794 -21556 392880 -21500
rect 392936 -21556 393008 -21500
rect 392668 -21642 393008 -21556
rect 392668 -21698 392738 -21642
rect 392794 -21698 392880 -21642
rect 392936 -21698 393008 -21642
rect 392668 -21784 393008 -21698
rect 392668 -21840 392738 -21784
rect 392794 -21840 392880 -21784
rect 392936 -21840 393008 -21784
rect 392668 -21926 393008 -21840
rect 392668 -21982 392738 -21926
rect 392794 -21982 392880 -21926
rect 392936 -21982 393008 -21926
rect 392668 -22068 393008 -21982
rect 392668 -22124 392738 -22068
rect 392794 -22124 392880 -22068
rect 392936 -22124 393008 -22068
rect 392668 -22210 393008 -22124
rect 392668 -22266 392738 -22210
rect 392794 -22266 392880 -22210
rect 392936 -22266 393008 -22210
rect 392668 -22352 393008 -22266
rect 392668 -22408 392738 -22352
rect 392794 -22408 392880 -22352
rect 392936 -22408 393008 -22352
rect 392668 -22494 393008 -22408
rect 392668 -22550 392738 -22494
rect 392794 -22550 392880 -22494
rect 392936 -22550 393008 -22494
rect 392668 -22636 393008 -22550
rect 392668 -22692 392738 -22636
rect 392794 -22692 392880 -22636
rect 392936 -22692 393008 -22636
rect 392668 -22778 393008 -22692
rect 392668 -22834 392738 -22778
rect 392794 -22834 392880 -22778
rect 392936 -22834 393008 -22778
rect 392668 -22920 393008 -22834
rect 392668 -22976 392738 -22920
rect 392794 -22976 392880 -22920
rect 392936 -22976 393008 -22920
rect 392668 -23062 393008 -22976
rect 392668 -23118 392738 -23062
rect 392794 -23118 392880 -23062
rect 392936 -23118 393008 -23062
rect 392668 -23204 393008 -23118
rect 392668 -23260 392738 -23204
rect 392794 -23260 392880 -23204
rect 392936 -23260 393008 -23204
rect 392668 -23346 393008 -23260
rect 392668 -23402 392738 -23346
rect 392794 -23402 392880 -23346
rect 392936 -23402 393008 -23346
rect 392668 -23488 393008 -23402
rect 392668 -23544 392738 -23488
rect 392794 -23544 392880 -23488
rect 392936 -23544 393008 -23488
rect 392668 -23630 393008 -23544
rect 392668 -23686 392738 -23630
rect 392794 -23686 392880 -23630
rect 392936 -23686 393008 -23630
rect 392668 -23772 393008 -23686
rect 392668 -23828 392738 -23772
rect 392794 -23828 392880 -23772
rect 392936 -23828 393008 -23772
rect 392668 -23914 393008 -23828
rect 392668 -23970 392738 -23914
rect 392794 -23970 392880 -23914
rect 392936 -23970 393008 -23914
rect 392668 -24056 393008 -23970
rect 392668 -24112 392738 -24056
rect 392794 -24112 392880 -24056
rect 392936 -24112 393008 -24056
rect 392668 -24198 393008 -24112
rect 392668 -24254 392738 -24198
rect 392794 -24254 392880 -24198
rect 392936 -24254 393008 -24198
rect 392668 -24340 393008 -24254
rect 392668 -24396 392738 -24340
rect 392794 -24396 392880 -24340
rect 392936 -24396 393008 -24340
rect 392668 -24482 393008 -24396
rect 392668 -24538 392738 -24482
rect 392794 -24538 392880 -24482
rect 392936 -24538 393008 -24482
rect 392668 -24624 393008 -24538
rect 392668 -24680 392738 -24624
rect 392794 -24680 392880 -24624
rect 392936 -24680 393008 -24624
rect 392668 -24766 393008 -24680
rect 392668 -24822 392738 -24766
rect 392794 -24822 392880 -24766
rect 392936 -24822 393008 -24766
rect 392668 -24908 393008 -24822
rect 392668 -24964 392738 -24908
rect 392794 -24964 392880 -24908
rect 392936 -24964 393008 -24908
rect 392668 -25050 393008 -24964
rect 392668 -25106 392738 -25050
rect 392794 -25106 392880 -25050
rect 392936 -25106 393008 -25050
rect 392668 -25192 393008 -25106
rect 392668 -25248 392738 -25192
rect 392794 -25248 392880 -25192
rect 392936 -25248 393008 -25192
rect 392668 -25334 393008 -25248
rect 392668 -25390 392738 -25334
rect 392794 -25390 392880 -25334
rect 392936 -25390 393008 -25334
rect 392668 -25476 393008 -25390
rect 392668 -25532 392738 -25476
rect 392794 -25532 392880 -25476
rect 392936 -25532 393008 -25476
rect 392668 -25542 393008 -25532
rect 393068 -17950 393408 -17820
rect 393068 -18006 393138 -17950
rect 393194 -18006 393280 -17950
rect 393336 -18006 393408 -17950
rect 393068 -18092 393408 -18006
rect 393068 -18148 393138 -18092
rect 393194 -18148 393280 -18092
rect 393336 -18148 393408 -18092
rect 393068 -18234 393408 -18148
rect 393068 -18290 393138 -18234
rect 393194 -18290 393280 -18234
rect 393336 -18290 393408 -18234
rect 393068 -18376 393408 -18290
rect 393068 -18432 393138 -18376
rect 393194 -18432 393280 -18376
rect 393336 -18432 393408 -18376
rect 393068 -18518 393408 -18432
rect 393068 -18574 393138 -18518
rect 393194 -18574 393280 -18518
rect 393336 -18574 393408 -18518
rect 393068 -18660 393408 -18574
rect 393068 -18716 393138 -18660
rect 393194 -18716 393280 -18660
rect 393336 -18716 393408 -18660
rect 393068 -18802 393408 -18716
rect 393068 -18858 393138 -18802
rect 393194 -18858 393280 -18802
rect 393336 -18858 393408 -18802
rect 393068 -18944 393408 -18858
rect 393068 -19000 393138 -18944
rect 393194 -19000 393280 -18944
rect 393336 -19000 393408 -18944
rect 393068 -19086 393408 -19000
rect 393068 -19142 393138 -19086
rect 393194 -19142 393280 -19086
rect 393336 -19142 393408 -19086
rect 393068 -19228 393408 -19142
rect 393068 -19284 393138 -19228
rect 393194 -19284 393280 -19228
rect 393336 -19284 393408 -19228
rect 393068 -19370 393408 -19284
rect 393068 -19426 393138 -19370
rect 393194 -19426 393280 -19370
rect 393336 -19426 393408 -19370
rect 393068 -19512 393408 -19426
rect 393068 -19568 393138 -19512
rect 393194 -19568 393280 -19512
rect 393336 -19568 393408 -19512
rect 393068 -19654 393408 -19568
rect 393068 -19710 393138 -19654
rect 393194 -19710 393280 -19654
rect 393336 -19710 393408 -19654
rect 393068 -19796 393408 -19710
rect 393068 -19852 393138 -19796
rect 393194 -19852 393280 -19796
rect 393336 -19852 393408 -19796
rect 393068 -19938 393408 -19852
rect 393068 -19994 393138 -19938
rect 393194 -19994 393280 -19938
rect 393336 -19994 393408 -19938
rect 393068 -20080 393408 -19994
rect 393068 -20136 393138 -20080
rect 393194 -20136 393280 -20080
rect 393336 -20136 393408 -20080
rect 393068 -20222 393408 -20136
rect 393068 -20278 393138 -20222
rect 393194 -20278 393280 -20222
rect 393336 -20278 393408 -20222
rect 393068 -20364 393408 -20278
rect 393068 -20420 393138 -20364
rect 393194 -20420 393280 -20364
rect 393336 -20420 393408 -20364
rect 393068 -20506 393408 -20420
rect 393068 -20562 393138 -20506
rect 393194 -20562 393280 -20506
rect 393336 -20562 393408 -20506
rect 393068 -20648 393408 -20562
rect 393068 -20704 393138 -20648
rect 393194 -20704 393280 -20648
rect 393336 -20704 393408 -20648
rect 393068 -20790 393408 -20704
rect 393068 -20846 393138 -20790
rect 393194 -20846 393280 -20790
rect 393336 -20846 393408 -20790
rect 393068 -20932 393408 -20846
rect 393068 -20988 393138 -20932
rect 393194 -20988 393280 -20932
rect 393336 -20988 393408 -20932
rect 393068 -21074 393408 -20988
rect 393068 -21130 393138 -21074
rect 393194 -21130 393280 -21074
rect 393336 -21130 393408 -21074
rect 393068 -21216 393408 -21130
rect 393068 -21272 393138 -21216
rect 393194 -21272 393280 -21216
rect 393336 -21272 393408 -21216
rect 393068 -21358 393408 -21272
rect 393068 -21414 393138 -21358
rect 393194 -21414 393280 -21358
rect 393336 -21414 393408 -21358
rect 393068 -21500 393408 -21414
rect 393068 -21556 393138 -21500
rect 393194 -21556 393280 -21500
rect 393336 -21556 393408 -21500
rect 393068 -21642 393408 -21556
rect 393068 -21698 393138 -21642
rect 393194 -21698 393280 -21642
rect 393336 -21698 393408 -21642
rect 393068 -21784 393408 -21698
rect 393068 -21840 393138 -21784
rect 393194 -21840 393280 -21784
rect 393336 -21840 393408 -21784
rect 393068 -21926 393408 -21840
rect 393068 -21982 393138 -21926
rect 393194 -21982 393280 -21926
rect 393336 -21982 393408 -21926
rect 393068 -22068 393408 -21982
rect 393068 -22124 393138 -22068
rect 393194 -22124 393280 -22068
rect 393336 -22124 393408 -22068
rect 393068 -22210 393408 -22124
rect 393068 -22266 393138 -22210
rect 393194 -22266 393280 -22210
rect 393336 -22266 393408 -22210
rect 393068 -22352 393408 -22266
rect 393068 -22408 393138 -22352
rect 393194 -22408 393280 -22352
rect 393336 -22408 393408 -22352
rect 393068 -22494 393408 -22408
rect 393068 -22550 393138 -22494
rect 393194 -22550 393280 -22494
rect 393336 -22550 393408 -22494
rect 393068 -22636 393408 -22550
rect 393068 -22692 393138 -22636
rect 393194 -22692 393280 -22636
rect 393336 -22692 393408 -22636
rect 393068 -22778 393408 -22692
rect 393068 -22834 393138 -22778
rect 393194 -22834 393280 -22778
rect 393336 -22834 393408 -22778
rect 393068 -22920 393408 -22834
rect 393068 -22976 393138 -22920
rect 393194 -22976 393280 -22920
rect 393336 -22976 393408 -22920
rect 393068 -23062 393408 -22976
rect 393068 -23118 393138 -23062
rect 393194 -23118 393280 -23062
rect 393336 -23118 393408 -23062
rect 393068 -23204 393408 -23118
rect 393068 -23260 393138 -23204
rect 393194 -23260 393280 -23204
rect 393336 -23260 393408 -23204
rect 393068 -23346 393408 -23260
rect 393068 -23402 393138 -23346
rect 393194 -23402 393280 -23346
rect 393336 -23402 393408 -23346
rect 393068 -23488 393408 -23402
rect 393068 -23544 393138 -23488
rect 393194 -23544 393280 -23488
rect 393336 -23544 393408 -23488
rect 393068 -23630 393408 -23544
rect 393068 -23686 393138 -23630
rect 393194 -23686 393280 -23630
rect 393336 -23686 393408 -23630
rect 393068 -23772 393408 -23686
rect 393068 -23828 393138 -23772
rect 393194 -23828 393280 -23772
rect 393336 -23828 393408 -23772
rect 393068 -23914 393408 -23828
rect 393068 -23970 393138 -23914
rect 393194 -23970 393280 -23914
rect 393336 -23970 393408 -23914
rect 393068 -24056 393408 -23970
rect 393068 -24112 393138 -24056
rect 393194 -24112 393280 -24056
rect 393336 -24112 393408 -24056
rect 393068 -24198 393408 -24112
rect 393068 -24254 393138 -24198
rect 393194 -24254 393280 -24198
rect 393336 -24254 393408 -24198
rect 393068 -24340 393408 -24254
rect 393068 -24396 393138 -24340
rect 393194 -24396 393280 -24340
rect 393336 -24396 393408 -24340
rect 393068 -24482 393408 -24396
rect 393068 -24538 393138 -24482
rect 393194 -24538 393280 -24482
rect 393336 -24538 393408 -24482
rect 393068 -24624 393408 -24538
rect 393068 -24680 393138 -24624
rect 393194 -24680 393280 -24624
rect 393336 -24680 393408 -24624
rect 393068 -24766 393408 -24680
rect 393068 -24822 393138 -24766
rect 393194 -24822 393280 -24766
rect 393336 -24822 393408 -24766
rect 393068 -24908 393408 -24822
rect 393068 -24964 393138 -24908
rect 393194 -24964 393280 -24908
rect 393336 -24964 393408 -24908
rect 393068 -25050 393408 -24964
rect 393068 -25106 393138 -25050
rect 393194 -25106 393280 -25050
rect 393336 -25106 393408 -25050
rect 393068 -25192 393408 -25106
rect 393068 -25248 393138 -25192
rect 393194 -25248 393280 -25192
rect 393336 -25248 393408 -25192
rect 393068 -25334 393408 -25248
rect 393068 -25390 393138 -25334
rect 393194 -25390 393280 -25334
rect 393336 -25390 393408 -25334
rect 393068 -25476 393408 -25390
rect 393068 -25532 393138 -25476
rect 393194 -25532 393280 -25476
rect 393336 -25532 393408 -25476
rect 393068 -25542 393408 -25532
rect 393468 -17950 393808 -17820
rect 393468 -18006 393543 -17950
rect 393599 -18006 393685 -17950
rect 393741 -18006 393808 -17950
rect 393468 -18092 393808 -18006
rect 393468 -18148 393543 -18092
rect 393599 -18148 393685 -18092
rect 393741 -18148 393808 -18092
rect 393468 -18234 393808 -18148
rect 393468 -18290 393543 -18234
rect 393599 -18290 393685 -18234
rect 393741 -18290 393808 -18234
rect 393468 -18376 393808 -18290
rect 393468 -18432 393543 -18376
rect 393599 -18432 393685 -18376
rect 393741 -18432 393808 -18376
rect 393468 -18518 393808 -18432
rect 393468 -18574 393543 -18518
rect 393599 -18574 393685 -18518
rect 393741 -18574 393808 -18518
rect 393468 -18660 393808 -18574
rect 393468 -18716 393543 -18660
rect 393599 -18716 393685 -18660
rect 393741 -18716 393808 -18660
rect 393468 -18802 393808 -18716
rect 393468 -18858 393543 -18802
rect 393599 -18858 393685 -18802
rect 393741 -18858 393808 -18802
rect 393468 -18944 393808 -18858
rect 393468 -19000 393543 -18944
rect 393599 -19000 393685 -18944
rect 393741 -19000 393808 -18944
rect 393468 -19086 393808 -19000
rect 393468 -19142 393543 -19086
rect 393599 -19142 393685 -19086
rect 393741 -19142 393808 -19086
rect 393468 -19228 393808 -19142
rect 393468 -19284 393543 -19228
rect 393599 -19284 393685 -19228
rect 393741 -19284 393808 -19228
rect 393468 -19370 393808 -19284
rect 393468 -19426 393543 -19370
rect 393599 -19426 393685 -19370
rect 393741 -19426 393808 -19370
rect 393468 -19512 393808 -19426
rect 393468 -19568 393543 -19512
rect 393599 -19568 393685 -19512
rect 393741 -19568 393808 -19512
rect 393468 -19654 393808 -19568
rect 393468 -19710 393543 -19654
rect 393599 -19710 393685 -19654
rect 393741 -19710 393808 -19654
rect 393468 -19796 393808 -19710
rect 393468 -19852 393543 -19796
rect 393599 -19852 393685 -19796
rect 393741 -19852 393808 -19796
rect 393468 -19938 393808 -19852
rect 393468 -19994 393543 -19938
rect 393599 -19994 393685 -19938
rect 393741 -19994 393808 -19938
rect 393468 -20080 393808 -19994
rect 393468 -20136 393543 -20080
rect 393599 -20136 393685 -20080
rect 393741 -20136 393808 -20080
rect 393468 -20222 393808 -20136
rect 393468 -20278 393543 -20222
rect 393599 -20278 393685 -20222
rect 393741 -20278 393808 -20222
rect 393468 -20364 393808 -20278
rect 393468 -20420 393543 -20364
rect 393599 -20420 393685 -20364
rect 393741 -20420 393808 -20364
rect 393468 -20506 393808 -20420
rect 393468 -20562 393543 -20506
rect 393599 -20562 393685 -20506
rect 393741 -20562 393808 -20506
rect 393468 -20648 393808 -20562
rect 393468 -20704 393543 -20648
rect 393599 -20704 393685 -20648
rect 393741 -20704 393808 -20648
rect 393468 -20790 393808 -20704
rect 393468 -20846 393543 -20790
rect 393599 -20846 393685 -20790
rect 393741 -20846 393808 -20790
rect 393468 -20932 393808 -20846
rect 393468 -20988 393543 -20932
rect 393599 -20988 393685 -20932
rect 393741 -20988 393808 -20932
rect 393468 -21074 393808 -20988
rect 393468 -21130 393543 -21074
rect 393599 -21130 393685 -21074
rect 393741 -21130 393808 -21074
rect 393468 -21216 393808 -21130
rect 393468 -21272 393543 -21216
rect 393599 -21272 393685 -21216
rect 393741 -21272 393808 -21216
rect 393468 -21358 393808 -21272
rect 393468 -21414 393543 -21358
rect 393599 -21414 393685 -21358
rect 393741 -21414 393808 -21358
rect 393468 -21500 393808 -21414
rect 393468 -21556 393543 -21500
rect 393599 -21556 393685 -21500
rect 393741 -21556 393808 -21500
rect 393468 -21642 393808 -21556
rect 393468 -21698 393543 -21642
rect 393599 -21698 393685 -21642
rect 393741 -21698 393808 -21642
rect 393468 -21784 393808 -21698
rect 393468 -21840 393543 -21784
rect 393599 -21840 393685 -21784
rect 393741 -21840 393808 -21784
rect 393468 -21926 393808 -21840
rect 393468 -21982 393543 -21926
rect 393599 -21982 393685 -21926
rect 393741 -21982 393808 -21926
rect 393468 -22068 393808 -21982
rect 393468 -22124 393543 -22068
rect 393599 -22124 393685 -22068
rect 393741 -22124 393808 -22068
rect 393468 -22210 393808 -22124
rect 393468 -22266 393543 -22210
rect 393599 -22266 393685 -22210
rect 393741 -22266 393808 -22210
rect 393468 -22352 393808 -22266
rect 393468 -22408 393543 -22352
rect 393599 -22408 393685 -22352
rect 393741 -22408 393808 -22352
rect 393468 -22494 393808 -22408
rect 393468 -22550 393543 -22494
rect 393599 -22550 393685 -22494
rect 393741 -22550 393808 -22494
rect 393468 -22636 393808 -22550
rect 393468 -22692 393543 -22636
rect 393599 -22692 393685 -22636
rect 393741 -22692 393808 -22636
rect 393468 -22778 393808 -22692
rect 393468 -22834 393543 -22778
rect 393599 -22834 393685 -22778
rect 393741 -22834 393808 -22778
rect 393468 -22920 393808 -22834
rect 393468 -22976 393543 -22920
rect 393599 -22976 393685 -22920
rect 393741 -22976 393808 -22920
rect 393468 -23062 393808 -22976
rect 393468 -23118 393543 -23062
rect 393599 -23118 393685 -23062
rect 393741 -23118 393808 -23062
rect 393468 -23204 393808 -23118
rect 393468 -23260 393543 -23204
rect 393599 -23260 393685 -23204
rect 393741 -23260 393808 -23204
rect 393468 -23346 393808 -23260
rect 393468 -23402 393543 -23346
rect 393599 -23402 393685 -23346
rect 393741 -23402 393808 -23346
rect 393468 -23488 393808 -23402
rect 393468 -23544 393543 -23488
rect 393599 -23544 393685 -23488
rect 393741 -23544 393808 -23488
rect 393468 -23630 393808 -23544
rect 393468 -23686 393543 -23630
rect 393599 -23686 393685 -23630
rect 393741 -23686 393808 -23630
rect 393468 -23772 393808 -23686
rect 393468 -23828 393543 -23772
rect 393599 -23828 393685 -23772
rect 393741 -23828 393808 -23772
rect 393468 -23914 393808 -23828
rect 393468 -23970 393543 -23914
rect 393599 -23970 393685 -23914
rect 393741 -23970 393808 -23914
rect 393468 -24056 393808 -23970
rect 393468 -24112 393543 -24056
rect 393599 -24112 393685 -24056
rect 393741 -24112 393808 -24056
rect 393468 -24198 393808 -24112
rect 393468 -24254 393543 -24198
rect 393599 -24254 393685 -24198
rect 393741 -24254 393808 -24198
rect 393468 -24340 393808 -24254
rect 393468 -24396 393543 -24340
rect 393599 -24396 393685 -24340
rect 393741 -24396 393808 -24340
rect 393468 -24482 393808 -24396
rect 393468 -24538 393543 -24482
rect 393599 -24538 393685 -24482
rect 393741 -24538 393808 -24482
rect 393468 -24624 393808 -24538
rect 393468 -24680 393543 -24624
rect 393599 -24680 393685 -24624
rect 393741 -24680 393808 -24624
rect 393468 -24766 393808 -24680
rect 393468 -24822 393543 -24766
rect 393599 -24822 393685 -24766
rect 393741 -24822 393808 -24766
rect 393468 -24908 393808 -24822
rect 393468 -24964 393543 -24908
rect 393599 -24964 393685 -24908
rect 393741 -24964 393808 -24908
rect 393468 -25050 393808 -24964
rect 393468 -25106 393543 -25050
rect 393599 -25106 393685 -25050
rect 393741 -25106 393808 -25050
rect 393468 -25192 393808 -25106
rect 393468 -25248 393543 -25192
rect 393599 -25248 393685 -25192
rect 393741 -25248 393808 -25192
rect 393468 -25334 393808 -25248
rect 393468 -25390 393543 -25334
rect 393599 -25390 393685 -25334
rect 393741 -25390 393808 -25334
rect 393468 -25476 393808 -25390
rect 393468 -25532 393543 -25476
rect 393599 -25532 393685 -25476
rect 393741 -25532 393808 -25476
rect 393468 -25542 393808 -25532
rect 393868 -17950 394208 -17820
rect 393868 -18006 393940 -17950
rect 393996 -18006 394082 -17950
rect 394138 -18006 394208 -17950
rect 393868 -18092 394208 -18006
rect 393868 -18148 393940 -18092
rect 393996 -18148 394082 -18092
rect 394138 -18148 394208 -18092
rect 393868 -18234 394208 -18148
rect 393868 -18290 393940 -18234
rect 393996 -18290 394082 -18234
rect 394138 -18290 394208 -18234
rect 393868 -18376 394208 -18290
rect 393868 -18432 393940 -18376
rect 393996 -18432 394082 -18376
rect 394138 -18432 394208 -18376
rect 393868 -18518 394208 -18432
rect 393868 -18574 393940 -18518
rect 393996 -18574 394082 -18518
rect 394138 -18574 394208 -18518
rect 393868 -18660 394208 -18574
rect 393868 -18716 393940 -18660
rect 393996 -18716 394082 -18660
rect 394138 -18716 394208 -18660
rect 393868 -18802 394208 -18716
rect 393868 -18858 393940 -18802
rect 393996 -18858 394082 -18802
rect 394138 -18858 394208 -18802
rect 393868 -18944 394208 -18858
rect 393868 -19000 393940 -18944
rect 393996 -19000 394082 -18944
rect 394138 -19000 394208 -18944
rect 393868 -19086 394208 -19000
rect 393868 -19142 393940 -19086
rect 393996 -19142 394082 -19086
rect 394138 -19142 394208 -19086
rect 393868 -19228 394208 -19142
rect 393868 -19284 393940 -19228
rect 393996 -19284 394082 -19228
rect 394138 -19284 394208 -19228
rect 393868 -19370 394208 -19284
rect 393868 -19426 393940 -19370
rect 393996 -19426 394082 -19370
rect 394138 -19426 394208 -19370
rect 393868 -19512 394208 -19426
rect 393868 -19568 393940 -19512
rect 393996 -19568 394082 -19512
rect 394138 -19568 394208 -19512
rect 393868 -19654 394208 -19568
rect 393868 -19710 393940 -19654
rect 393996 -19710 394082 -19654
rect 394138 -19710 394208 -19654
rect 393868 -19796 394208 -19710
rect 393868 -19852 393940 -19796
rect 393996 -19852 394082 -19796
rect 394138 -19852 394208 -19796
rect 393868 -19938 394208 -19852
rect 393868 -19994 393940 -19938
rect 393996 -19994 394082 -19938
rect 394138 -19994 394208 -19938
rect 393868 -20080 394208 -19994
rect 393868 -20136 393940 -20080
rect 393996 -20136 394082 -20080
rect 394138 -20136 394208 -20080
rect 393868 -20222 394208 -20136
rect 393868 -20278 393940 -20222
rect 393996 -20278 394082 -20222
rect 394138 -20278 394208 -20222
rect 393868 -20364 394208 -20278
rect 393868 -20420 393940 -20364
rect 393996 -20420 394082 -20364
rect 394138 -20420 394208 -20364
rect 393868 -20506 394208 -20420
rect 393868 -20562 393940 -20506
rect 393996 -20562 394082 -20506
rect 394138 -20562 394208 -20506
rect 393868 -20648 394208 -20562
rect 393868 -20704 393940 -20648
rect 393996 -20704 394082 -20648
rect 394138 -20704 394208 -20648
rect 393868 -20790 394208 -20704
rect 393868 -20846 393940 -20790
rect 393996 -20846 394082 -20790
rect 394138 -20846 394208 -20790
rect 393868 -20932 394208 -20846
rect 393868 -20988 393940 -20932
rect 393996 -20988 394082 -20932
rect 394138 -20988 394208 -20932
rect 393868 -21074 394208 -20988
rect 393868 -21130 393940 -21074
rect 393996 -21130 394082 -21074
rect 394138 -21130 394208 -21074
rect 393868 -21216 394208 -21130
rect 393868 -21272 393940 -21216
rect 393996 -21272 394082 -21216
rect 394138 -21272 394208 -21216
rect 393868 -21358 394208 -21272
rect 393868 -21414 393940 -21358
rect 393996 -21414 394082 -21358
rect 394138 -21414 394208 -21358
rect 393868 -21500 394208 -21414
rect 393868 -21556 393940 -21500
rect 393996 -21556 394082 -21500
rect 394138 -21556 394208 -21500
rect 393868 -21642 394208 -21556
rect 393868 -21698 393940 -21642
rect 393996 -21698 394082 -21642
rect 394138 -21698 394208 -21642
rect 393868 -21784 394208 -21698
rect 393868 -21840 393940 -21784
rect 393996 -21840 394082 -21784
rect 394138 -21840 394208 -21784
rect 393868 -21926 394208 -21840
rect 393868 -21982 393940 -21926
rect 393996 -21982 394082 -21926
rect 394138 -21982 394208 -21926
rect 393868 -22068 394208 -21982
rect 393868 -22124 393940 -22068
rect 393996 -22124 394082 -22068
rect 394138 -22124 394208 -22068
rect 393868 -22210 394208 -22124
rect 393868 -22266 393940 -22210
rect 393996 -22266 394082 -22210
rect 394138 -22266 394208 -22210
rect 393868 -22352 394208 -22266
rect 393868 -22408 393940 -22352
rect 393996 -22408 394082 -22352
rect 394138 -22408 394208 -22352
rect 393868 -22494 394208 -22408
rect 393868 -22550 393940 -22494
rect 393996 -22550 394082 -22494
rect 394138 -22550 394208 -22494
rect 393868 -22636 394208 -22550
rect 393868 -22692 393940 -22636
rect 393996 -22692 394082 -22636
rect 394138 -22692 394208 -22636
rect 393868 -22778 394208 -22692
rect 393868 -22834 393940 -22778
rect 393996 -22834 394082 -22778
rect 394138 -22834 394208 -22778
rect 393868 -22920 394208 -22834
rect 393868 -22976 393940 -22920
rect 393996 -22976 394082 -22920
rect 394138 -22976 394208 -22920
rect 393868 -23062 394208 -22976
rect 393868 -23118 393940 -23062
rect 393996 -23118 394082 -23062
rect 394138 -23118 394208 -23062
rect 393868 -23204 394208 -23118
rect 393868 -23260 393940 -23204
rect 393996 -23260 394082 -23204
rect 394138 -23260 394208 -23204
rect 393868 -23346 394208 -23260
rect 393868 -23402 393940 -23346
rect 393996 -23402 394082 -23346
rect 394138 -23402 394208 -23346
rect 393868 -23488 394208 -23402
rect 393868 -23544 393940 -23488
rect 393996 -23544 394082 -23488
rect 394138 -23544 394208 -23488
rect 393868 -23630 394208 -23544
rect 393868 -23686 393940 -23630
rect 393996 -23686 394082 -23630
rect 394138 -23686 394208 -23630
rect 393868 -23772 394208 -23686
rect 393868 -23828 393940 -23772
rect 393996 -23828 394082 -23772
rect 394138 -23828 394208 -23772
rect 393868 -23914 394208 -23828
rect 393868 -23970 393940 -23914
rect 393996 -23970 394082 -23914
rect 394138 -23970 394208 -23914
rect 393868 -24056 394208 -23970
rect 393868 -24112 393940 -24056
rect 393996 -24112 394082 -24056
rect 394138 -24112 394208 -24056
rect 393868 -24198 394208 -24112
rect 393868 -24254 393940 -24198
rect 393996 -24254 394082 -24198
rect 394138 -24254 394208 -24198
rect 393868 -24340 394208 -24254
rect 393868 -24396 393940 -24340
rect 393996 -24396 394082 -24340
rect 394138 -24396 394208 -24340
rect 393868 -24482 394208 -24396
rect 393868 -24538 393940 -24482
rect 393996 -24538 394082 -24482
rect 394138 -24538 394208 -24482
rect 393868 -24624 394208 -24538
rect 393868 -24680 393940 -24624
rect 393996 -24680 394082 -24624
rect 394138 -24680 394208 -24624
rect 393868 -24766 394208 -24680
rect 393868 -24822 393940 -24766
rect 393996 -24822 394082 -24766
rect 394138 -24822 394208 -24766
rect 393868 -24908 394208 -24822
rect 393868 -24964 393940 -24908
rect 393996 -24964 394082 -24908
rect 394138 -24964 394208 -24908
rect 393868 -25050 394208 -24964
rect 393868 -25106 393940 -25050
rect 393996 -25106 394082 -25050
rect 394138 -25106 394208 -25050
rect 393868 -25192 394208 -25106
rect 393868 -25248 393940 -25192
rect 393996 -25248 394082 -25192
rect 394138 -25248 394208 -25192
rect 393868 -25334 394208 -25248
rect 393868 -25390 393940 -25334
rect 393996 -25390 394082 -25334
rect 394138 -25390 394208 -25334
rect 393868 -25476 394208 -25390
rect 393868 -25532 393940 -25476
rect 393996 -25532 394082 -25476
rect 394138 -25532 394208 -25476
rect 393868 -25542 394208 -25532
rect 394268 -17950 394608 -17820
rect 394268 -18006 394337 -17950
rect 394393 -18006 394479 -17950
rect 394535 -18006 394608 -17950
rect 394268 -18092 394608 -18006
rect 394268 -18148 394337 -18092
rect 394393 -18148 394479 -18092
rect 394535 -18148 394608 -18092
rect 394268 -18234 394608 -18148
rect 394268 -18290 394337 -18234
rect 394393 -18290 394479 -18234
rect 394535 -18290 394608 -18234
rect 394268 -18376 394608 -18290
rect 394268 -18432 394337 -18376
rect 394393 -18432 394479 -18376
rect 394535 -18432 394608 -18376
rect 394268 -18518 394608 -18432
rect 394268 -18574 394337 -18518
rect 394393 -18574 394479 -18518
rect 394535 -18574 394608 -18518
rect 394268 -18660 394608 -18574
rect 394268 -18716 394337 -18660
rect 394393 -18716 394479 -18660
rect 394535 -18716 394608 -18660
rect 394268 -18802 394608 -18716
rect 394268 -18858 394337 -18802
rect 394393 -18858 394479 -18802
rect 394535 -18858 394608 -18802
rect 394268 -18944 394608 -18858
rect 394268 -19000 394337 -18944
rect 394393 -19000 394479 -18944
rect 394535 -19000 394608 -18944
rect 394268 -19086 394608 -19000
rect 394268 -19142 394337 -19086
rect 394393 -19142 394479 -19086
rect 394535 -19142 394608 -19086
rect 394268 -19228 394608 -19142
rect 394268 -19284 394337 -19228
rect 394393 -19284 394479 -19228
rect 394535 -19284 394608 -19228
rect 394268 -19370 394608 -19284
rect 394268 -19426 394337 -19370
rect 394393 -19426 394479 -19370
rect 394535 -19426 394608 -19370
rect 394268 -19512 394608 -19426
rect 394268 -19568 394337 -19512
rect 394393 -19568 394479 -19512
rect 394535 -19568 394608 -19512
rect 394268 -19654 394608 -19568
rect 394268 -19710 394337 -19654
rect 394393 -19710 394479 -19654
rect 394535 -19710 394608 -19654
rect 394268 -19796 394608 -19710
rect 394268 -19852 394337 -19796
rect 394393 -19852 394479 -19796
rect 394535 -19852 394608 -19796
rect 394268 -19938 394608 -19852
rect 394268 -19994 394337 -19938
rect 394393 -19994 394479 -19938
rect 394535 -19994 394608 -19938
rect 394268 -20080 394608 -19994
rect 394268 -20136 394337 -20080
rect 394393 -20136 394479 -20080
rect 394535 -20136 394608 -20080
rect 394268 -20222 394608 -20136
rect 394268 -20278 394337 -20222
rect 394393 -20278 394479 -20222
rect 394535 -20278 394608 -20222
rect 394268 -20364 394608 -20278
rect 394268 -20420 394337 -20364
rect 394393 -20420 394479 -20364
rect 394535 -20420 394608 -20364
rect 394268 -20506 394608 -20420
rect 394268 -20562 394337 -20506
rect 394393 -20562 394479 -20506
rect 394535 -20562 394608 -20506
rect 394268 -20648 394608 -20562
rect 394268 -20704 394337 -20648
rect 394393 -20704 394479 -20648
rect 394535 -20704 394608 -20648
rect 394268 -20790 394608 -20704
rect 394268 -20846 394337 -20790
rect 394393 -20846 394479 -20790
rect 394535 -20846 394608 -20790
rect 394268 -20932 394608 -20846
rect 394268 -20988 394337 -20932
rect 394393 -20988 394479 -20932
rect 394535 -20988 394608 -20932
rect 394268 -21074 394608 -20988
rect 394268 -21130 394337 -21074
rect 394393 -21130 394479 -21074
rect 394535 -21130 394608 -21074
rect 394268 -21216 394608 -21130
rect 394268 -21272 394337 -21216
rect 394393 -21272 394479 -21216
rect 394535 -21272 394608 -21216
rect 394268 -21358 394608 -21272
rect 394268 -21414 394337 -21358
rect 394393 -21414 394479 -21358
rect 394535 -21414 394608 -21358
rect 394268 -21500 394608 -21414
rect 394268 -21556 394337 -21500
rect 394393 -21556 394479 -21500
rect 394535 -21556 394608 -21500
rect 394268 -21642 394608 -21556
rect 394268 -21698 394337 -21642
rect 394393 -21698 394479 -21642
rect 394535 -21698 394608 -21642
rect 394268 -21784 394608 -21698
rect 394268 -21840 394337 -21784
rect 394393 -21840 394479 -21784
rect 394535 -21840 394608 -21784
rect 394268 -21926 394608 -21840
rect 394268 -21982 394337 -21926
rect 394393 -21982 394479 -21926
rect 394535 -21982 394608 -21926
rect 394268 -22068 394608 -21982
rect 394268 -22124 394337 -22068
rect 394393 -22124 394479 -22068
rect 394535 -22124 394608 -22068
rect 394268 -22210 394608 -22124
rect 394268 -22266 394337 -22210
rect 394393 -22266 394479 -22210
rect 394535 -22266 394608 -22210
rect 394268 -22352 394608 -22266
rect 394268 -22408 394337 -22352
rect 394393 -22408 394479 -22352
rect 394535 -22408 394608 -22352
rect 394268 -22494 394608 -22408
rect 394268 -22550 394337 -22494
rect 394393 -22550 394479 -22494
rect 394535 -22550 394608 -22494
rect 394268 -22636 394608 -22550
rect 394268 -22692 394337 -22636
rect 394393 -22692 394479 -22636
rect 394535 -22692 394608 -22636
rect 394268 -22778 394608 -22692
rect 394268 -22834 394337 -22778
rect 394393 -22834 394479 -22778
rect 394535 -22834 394608 -22778
rect 394268 -22920 394608 -22834
rect 394268 -22976 394337 -22920
rect 394393 -22976 394479 -22920
rect 394535 -22976 394608 -22920
rect 394268 -23062 394608 -22976
rect 394268 -23118 394337 -23062
rect 394393 -23118 394479 -23062
rect 394535 -23118 394608 -23062
rect 394268 -23204 394608 -23118
rect 394268 -23260 394337 -23204
rect 394393 -23260 394479 -23204
rect 394535 -23260 394608 -23204
rect 394268 -23346 394608 -23260
rect 394268 -23402 394337 -23346
rect 394393 -23402 394479 -23346
rect 394535 -23402 394608 -23346
rect 394268 -23488 394608 -23402
rect 394268 -23544 394337 -23488
rect 394393 -23544 394479 -23488
rect 394535 -23544 394608 -23488
rect 394268 -23630 394608 -23544
rect 394268 -23686 394337 -23630
rect 394393 -23686 394479 -23630
rect 394535 -23686 394608 -23630
rect 394268 -23772 394608 -23686
rect 394268 -23828 394337 -23772
rect 394393 -23828 394479 -23772
rect 394535 -23828 394608 -23772
rect 394268 -23914 394608 -23828
rect 394268 -23970 394337 -23914
rect 394393 -23970 394479 -23914
rect 394535 -23970 394608 -23914
rect 394268 -24056 394608 -23970
rect 394268 -24112 394337 -24056
rect 394393 -24112 394479 -24056
rect 394535 -24112 394608 -24056
rect 394268 -24198 394608 -24112
rect 394268 -24254 394337 -24198
rect 394393 -24254 394479 -24198
rect 394535 -24254 394608 -24198
rect 394268 -24340 394608 -24254
rect 394268 -24396 394337 -24340
rect 394393 -24396 394479 -24340
rect 394535 -24396 394608 -24340
rect 394268 -24482 394608 -24396
rect 394268 -24538 394337 -24482
rect 394393 -24538 394479 -24482
rect 394535 -24538 394608 -24482
rect 394268 -24624 394608 -24538
rect 394268 -24680 394337 -24624
rect 394393 -24680 394479 -24624
rect 394535 -24680 394608 -24624
rect 394268 -24766 394608 -24680
rect 394268 -24822 394337 -24766
rect 394393 -24822 394479 -24766
rect 394535 -24822 394608 -24766
rect 394268 -24908 394608 -24822
rect 394268 -24964 394337 -24908
rect 394393 -24964 394479 -24908
rect 394535 -24964 394608 -24908
rect 394268 -25050 394608 -24964
rect 394268 -25106 394337 -25050
rect 394393 -25106 394479 -25050
rect 394535 -25106 394608 -25050
rect 394268 -25192 394608 -25106
rect 394268 -25248 394337 -25192
rect 394393 -25248 394479 -25192
rect 394535 -25248 394608 -25192
rect 394268 -25334 394608 -25248
rect 394268 -25390 394337 -25334
rect 394393 -25390 394479 -25334
rect 394535 -25390 394608 -25334
rect 394268 -25476 394608 -25390
rect 394268 -25532 394337 -25476
rect 394393 -25532 394479 -25476
rect 394535 -25532 394608 -25476
rect 394268 -25542 394608 -25532
rect 394668 -17950 395008 -17820
rect 394668 -18006 394740 -17950
rect 394796 -18006 394882 -17950
rect 394938 -18006 395008 -17950
rect 394668 -18092 395008 -18006
rect 394668 -18148 394740 -18092
rect 394796 -18148 394882 -18092
rect 394938 -18148 395008 -18092
rect 394668 -18234 395008 -18148
rect 394668 -18290 394740 -18234
rect 394796 -18290 394882 -18234
rect 394938 -18290 395008 -18234
rect 394668 -18376 395008 -18290
rect 394668 -18432 394740 -18376
rect 394796 -18432 394882 -18376
rect 394938 -18432 395008 -18376
rect 394668 -18518 395008 -18432
rect 394668 -18574 394740 -18518
rect 394796 -18574 394882 -18518
rect 394938 -18574 395008 -18518
rect 394668 -18660 395008 -18574
rect 394668 -18716 394740 -18660
rect 394796 -18716 394882 -18660
rect 394938 -18716 395008 -18660
rect 394668 -18802 395008 -18716
rect 394668 -18858 394740 -18802
rect 394796 -18858 394882 -18802
rect 394938 -18858 395008 -18802
rect 394668 -18944 395008 -18858
rect 394668 -19000 394740 -18944
rect 394796 -19000 394882 -18944
rect 394938 -19000 395008 -18944
rect 394668 -19086 395008 -19000
rect 394668 -19142 394740 -19086
rect 394796 -19142 394882 -19086
rect 394938 -19142 395008 -19086
rect 394668 -19228 395008 -19142
rect 394668 -19284 394740 -19228
rect 394796 -19284 394882 -19228
rect 394938 -19284 395008 -19228
rect 394668 -19370 395008 -19284
rect 394668 -19426 394740 -19370
rect 394796 -19426 394882 -19370
rect 394938 -19426 395008 -19370
rect 394668 -19512 395008 -19426
rect 394668 -19568 394740 -19512
rect 394796 -19568 394882 -19512
rect 394938 -19568 395008 -19512
rect 394668 -19654 395008 -19568
rect 394668 -19710 394740 -19654
rect 394796 -19710 394882 -19654
rect 394938 -19710 395008 -19654
rect 394668 -19796 395008 -19710
rect 394668 -19852 394740 -19796
rect 394796 -19852 394882 -19796
rect 394938 -19852 395008 -19796
rect 394668 -19938 395008 -19852
rect 394668 -19994 394740 -19938
rect 394796 -19994 394882 -19938
rect 394938 -19994 395008 -19938
rect 394668 -20080 395008 -19994
rect 394668 -20136 394740 -20080
rect 394796 -20136 394882 -20080
rect 394938 -20136 395008 -20080
rect 394668 -20222 395008 -20136
rect 394668 -20278 394740 -20222
rect 394796 -20278 394882 -20222
rect 394938 -20278 395008 -20222
rect 394668 -20364 395008 -20278
rect 394668 -20420 394740 -20364
rect 394796 -20420 394882 -20364
rect 394938 -20420 395008 -20364
rect 394668 -20506 395008 -20420
rect 394668 -20562 394740 -20506
rect 394796 -20562 394882 -20506
rect 394938 -20562 395008 -20506
rect 394668 -20648 395008 -20562
rect 394668 -20704 394740 -20648
rect 394796 -20704 394882 -20648
rect 394938 -20704 395008 -20648
rect 394668 -20790 395008 -20704
rect 394668 -20846 394740 -20790
rect 394796 -20846 394882 -20790
rect 394938 -20846 395008 -20790
rect 394668 -20932 395008 -20846
rect 394668 -20988 394740 -20932
rect 394796 -20988 394882 -20932
rect 394938 -20988 395008 -20932
rect 394668 -21074 395008 -20988
rect 394668 -21130 394740 -21074
rect 394796 -21130 394882 -21074
rect 394938 -21130 395008 -21074
rect 394668 -21216 395008 -21130
rect 394668 -21272 394740 -21216
rect 394796 -21272 394882 -21216
rect 394938 -21272 395008 -21216
rect 394668 -21358 395008 -21272
rect 394668 -21414 394740 -21358
rect 394796 -21414 394882 -21358
rect 394938 -21414 395008 -21358
rect 394668 -21500 395008 -21414
rect 394668 -21556 394740 -21500
rect 394796 -21556 394882 -21500
rect 394938 -21556 395008 -21500
rect 394668 -21642 395008 -21556
rect 394668 -21698 394740 -21642
rect 394796 -21698 394882 -21642
rect 394938 -21698 395008 -21642
rect 394668 -21784 395008 -21698
rect 394668 -21840 394740 -21784
rect 394796 -21840 394882 -21784
rect 394938 -21840 395008 -21784
rect 394668 -21926 395008 -21840
rect 394668 -21982 394740 -21926
rect 394796 -21982 394882 -21926
rect 394938 -21982 395008 -21926
rect 394668 -22068 395008 -21982
rect 394668 -22124 394740 -22068
rect 394796 -22124 394882 -22068
rect 394938 -22124 395008 -22068
rect 394668 -22210 395008 -22124
rect 394668 -22266 394740 -22210
rect 394796 -22266 394882 -22210
rect 394938 -22266 395008 -22210
rect 394668 -22352 395008 -22266
rect 394668 -22408 394740 -22352
rect 394796 -22408 394882 -22352
rect 394938 -22408 395008 -22352
rect 394668 -22494 395008 -22408
rect 394668 -22550 394740 -22494
rect 394796 -22550 394882 -22494
rect 394938 -22550 395008 -22494
rect 394668 -22636 395008 -22550
rect 394668 -22692 394740 -22636
rect 394796 -22692 394882 -22636
rect 394938 -22692 395008 -22636
rect 394668 -22778 395008 -22692
rect 394668 -22834 394740 -22778
rect 394796 -22834 394882 -22778
rect 394938 -22834 395008 -22778
rect 394668 -22920 395008 -22834
rect 394668 -22976 394740 -22920
rect 394796 -22976 394882 -22920
rect 394938 -22976 395008 -22920
rect 394668 -23062 395008 -22976
rect 394668 -23118 394740 -23062
rect 394796 -23118 394882 -23062
rect 394938 -23118 395008 -23062
rect 394668 -23204 395008 -23118
rect 394668 -23260 394740 -23204
rect 394796 -23260 394882 -23204
rect 394938 -23260 395008 -23204
rect 394668 -23346 395008 -23260
rect 394668 -23402 394740 -23346
rect 394796 -23402 394882 -23346
rect 394938 -23402 395008 -23346
rect 394668 -23488 395008 -23402
rect 394668 -23544 394740 -23488
rect 394796 -23544 394882 -23488
rect 394938 -23544 395008 -23488
rect 394668 -23630 395008 -23544
rect 394668 -23686 394740 -23630
rect 394796 -23686 394882 -23630
rect 394938 -23686 395008 -23630
rect 394668 -23772 395008 -23686
rect 394668 -23828 394740 -23772
rect 394796 -23828 394882 -23772
rect 394938 -23828 395008 -23772
rect 394668 -23914 395008 -23828
rect 394668 -23970 394740 -23914
rect 394796 -23970 394882 -23914
rect 394938 -23970 395008 -23914
rect 394668 -24056 395008 -23970
rect 394668 -24112 394740 -24056
rect 394796 -24112 394882 -24056
rect 394938 -24112 395008 -24056
rect 394668 -24198 395008 -24112
rect 394668 -24254 394740 -24198
rect 394796 -24254 394882 -24198
rect 394938 -24254 395008 -24198
rect 394668 -24340 395008 -24254
rect 394668 -24396 394740 -24340
rect 394796 -24396 394882 -24340
rect 394938 -24396 395008 -24340
rect 394668 -24482 395008 -24396
rect 394668 -24538 394740 -24482
rect 394796 -24538 394882 -24482
rect 394938 -24538 395008 -24482
rect 394668 -24624 395008 -24538
rect 394668 -24680 394740 -24624
rect 394796 -24680 394882 -24624
rect 394938 -24680 395008 -24624
rect 394668 -24766 395008 -24680
rect 394668 -24822 394740 -24766
rect 394796 -24822 394882 -24766
rect 394938 -24822 395008 -24766
rect 394668 -24908 395008 -24822
rect 394668 -24964 394740 -24908
rect 394796 -24964 394882 -24908
rect 394938 -24964 395008 -24908
rect 394668 -25050 395008 -24964
rect 394668 -25106 394740 -25050
rect 394796 -25106 394882 -25050
rect 394938 -25106 395008 -25050
rect 394668 -25192 395008 -25106
rect 394668 -25248 394740 -25192
rect 394796 -25248 394882 -25192
rect 394938 -25248 395008 -25192
rect 394668 -25334 395008 -25248
rect 394668 -25390 394740 -25334
rect 394796 -25390 394882 -25334
rect 394938 -25390 395008 -25334
rect 394668 -25476 395008 -25390
rect 394668 -25532 394740 -25476
rect 394796 -25532 394882 -25476
rect 394938 -25532 395008 -25476
rect 394668 -25542 395008 -25532
rect 395068 -17950 395408 -17820
rect 395068 -18006 395142 -17950
rect 395198 -18006 395284 -17950
rect 395340 -18006 395408 -17950
rect 395068 -18092 395408 -18006
rect 395068 -18148 395142 -18092
rect 395198 -18148 395284 -18092
rect 395340 -18148 395408 -18092
rect 395068 -18234 395408 -18148
rect 395068 -18290 395142 -18234
rect 395198 -18290 395284 -18234
rect 395340 -18290 395408 -18234
rect 395068 -18376 395408 -18290
rect 395068 -18432 395142 -18376
rect 395198 -18432 395284 -18376
rect 395340 -18432 395408 -18376
rect 395068 -18518 395408 -18432
rect 395068 -18574 395142 -18518
rect 395198 -18574 395284 -18518
rect 395340 -18574 395408 -18518
rect 395068 -18660 395408 -18574
rect 395068 -18716 395142 -18660
rect 395198 -18716 395284 -18660
rect 395340 -18716 395408 -18660
rect 395068 -18802 395408 -18716
rect 395068 -18858 395142 -18802
rect 395198 -18858 395284 -18802
rect 395340 -18858 395408 -18802
rect 395068 -18944 395408 -18858
rect 395068 -19000 395142 -18944
rect 395198 -19000 395284 -18944
rect 395340 -19000 395408 -18944
rect 395068 -19086 395408 -19000
rect 395068 -19142 395142 -19086
rect 395198 -19142 395284 -19086
rect 395340 -19142 395408 -19086
rect 395068 -19228 395408 -19142
rect 395068 -19284 395142 -19228
rect 395198 -19284 395284 -19228
rect 395340 -19284 395408 -19228
rect 395068 -19370 395408 -19284
rect 395068 -19426 395142 -19370
rect 395198 -19426 395284 -19370
rect 395340 -19426 395408 -19370
rect 395068 -19512 395408 -19426
rect 395068 -19568 395142 -19512
rect 395198 -19568 395284 -19512
rect 395340 -19568 395408 -19512
rect 395068 -19654 395408 -19568
rect 395068 -19710 395142 -19654
rect 395198 -19710 395284 -19654
rect 395340 -19710 395408 -19654
rect 395068 -19796 395408 -19710
rect 395068 -19852 395142 -19796
rect 395198 -19852 395284 -19796
rect 395340 -19852 395408 -19796
rect 395068 -19938 395408 -19852
rect 395068 -19994 395142 -19938
rect 395198 -19994 395284 -19938
rect 395340 -19994 395408 -19938
rect 395068 -20080 395408 -19994
rect 395068 -20136 395142 -20080
rect 395198 -20136 395284 -20080
rect 395340 -20136 395408 -20080
rect 395068 -20222 395408 -20136
rect 395068 -20278 395142 -20222
rect 395198 -20278 395284 -20222
rect 395340 -20278 395408 -20222
rect 395068 -20364 395408 -20278
rect 395068 -20420 395142 -20364
rect 395198 -20420 395284 -20364
rect 395340 -20420 395408 -20364
rect 395068 -20506 395408 -20420
rect 395068 -20562 395142 -20506
rect 395198 -20562 395284 -20506
rect 395340 -20562 395408 -20506
rect 395068 -20648 395408 -20562
rect 395068 -20704 395142 -20648
rect 395198 -20704 395284 -20648
rect 395340 -20704 395408 -20648
rect 395068 -20790 395408 -20704
rect 395068 -20846 395142 -20790
rect 395198 -20846 395284 -20790
rect 395340 -20846 395408 -20790
rect 395068 -20932 395408 -20846
rect 395068 -20988 395142 -20932
rect 395198 -20988 395284 -20932
rect 395340 -20988 395408 -20932
rect 395068 -21074 395408 -20988
rect 395068 -21130 395142 -21074
rect 395198 -21130 395284 -21074
rect 395340 -21130 395408 -21074
rect 395068 -21216 395408 -21130
rect 395068 -21272 395142 -21216
rect 395198 -21272 395284 -21216
rect 395340 -21272 395408 -21216
rect 395068 -21358 395408 -21272
rect 395068 -21414 395142 -21358
rect 395198 -21414 395284 -21358
rect 395340 -21414 395408 -21358
rect 395068 -21500 395408 -21414
rect 395068 -21556 395142 -21500
rect 395198 -21556 395284 -21500
rect 395340 -21556 395408 -21500
rect 395068 -21642 395408 -21556
rect 395068 -21698 395142 -21642
rect 395198 -21698 395284 -21642
rect 395340 -21698 395408 -21642
rect 395068 -21784 395408 -21698
rect 395068 -21840 395142 -21784
rect 395198 -21840 395284 -21784
rect 395340 -21840 395408 -21784
rect 395068 -21926 395408 -21840
rect 395068 -21982 395142 -21926
rect 395198 -21982 395284 -21926
rect 395340 -21982 395408 -21926
rect 395068 -22068 395408 -21982
rect 395068 -22124 395142 -22068
rect 395198 -22124 395284 -22068
rect 395340 -22124 395408 -22068
rect 395068 -22210 395408 -22124
rect 395068 -22266 395142 -22210
rect 395198 -22266 395284 -22210
rect 395340 -22266 395408 -22210
rect 395068 -22352 395408 -22266
rect 395068 -22408 395142 -22352
rect 395198 -22408 395284 -22352
rect 395340 -22408 395408 -22352
rect 395068 -22494 395408 -22408
rect 395068 -22550 395142 -22494
rect 395198 -22550 395284 -22494
rect 395340 -22550 395408 -22494
rect 395068 -22636 395408 -22550
rect 395068 -22692 395142 -22636
rect 395198 -22692 395284 -22636
rect 395340 -22692 395408 -22636
rect 395068 -22778 395408 -22692
rect 395068 -22834 395142 -22778
rect 395198 -22834 395284 -22778
rect 395340 -22834 395408 -22778
rect 395068 -22920 395408 -22834
rect 395068 -22976 395142 -22920
rect 395198 -22976 395284 -22920
rect 395340 -22976 395408 -22920
rect 395068 -23062 395408 -22976
rect 395068 -23118 395142 -23062
rect 395198 -23118 395284 -23062
rect 395340 -23118 395408 -23062
rect 395068 -23204 395408 -23118
rect 395068 -23260 395142 -23204
rect 395198 -23260 395284 -23204
rect 395340 -23260 395408 -23204
rect 395068 -23346 395408 -23260
rect 395068 -23402 395142 -23346
rect 395198 -23402 395284 -23346
rect 395340 -23402 395408 -23346
rect 395068 -23488 395408 -23402
rect 395068 -23544 395142 -23488
rect 395198 -23544 395284 -23488
rect 395340 -23544 395408 -23488
rect 395068 -23630 395408 -23544
rect 395068 -23686 395142 -23630
rect 395198 -23686 395284 -23630
rect 395340 -23686 395408 -23630
rect 395068 -23772 395408 -23686
rect 395068 -23828 395142 -23772
rect 395198 -23828 395284 -23772
rect 395340 -23828 395408 -23772
rect 395068 -23914 395408 -23828
rect 395068 -23970 395142 -23914
rect 395198 -23970 395284 -23914
rect 395340 -23970 395408 -23914
rect 395068 -24056 395408 -23970
rect 395068 -24112 395142 -24056
rect 395198 -24112 395284 -24056
rect 395340 -24112 395408 -24056
rect 395068 -24198 395408 -24112
rect 395068 -24254 395142 -24198
rect 395198 -24254 395284 -24198
rect 395340 -24254 395408 -24198
rect 395068 -24340 395408 -24254
rect 395068 -24396 395142 -24340
rect 395198 -24396 395284 -24340
rect 395340 -24396 395408 -24340
rect 395068 -24482 395408 -24396
rect 395068 -24538 395142 -24482
rect 395198 -24538 395284 -24482
rect 395340 -24538 395408 -24482
rect 395068 -24624 395408 -24538
rect 395068 -24680 395142 -24624
rect 395198 -24680 395284 -24624
rect 395340 -24680 395408 -24624
rect 395068 -24766 395408 -24680
rect 395068 -24822 395142 -24766
rect 395198 -24822 395284 -24766
rect 395340 -24822 395408 -24766
rect 395068 -24908 395408 -24822
rect 395068 -24964 395142 -24908
rect 395198 -24964 395284 -24908
rect 395340 -24964 395408 -24908
rect 395068 -25050 395408 -24964
rect 395068 -25106 395142 -25050
rect 395198 -25106 395284 -25050
rect 395340 -25106 395408 -25050
rect 395068 -25192 395408 -25106
rect 395068 -25248 395142 -25192
rect 395198 -25248 395284 -25192
rect 395340 -25248 395408 -25192
rect 395068 -25334 395408 -25248
rect 395068 -25390 395142 -25334
rect 395198 -25390 395284 -25334
rect 395340 -25390 395408 -25334
rect 395068 -25476 395408 -25390
rect 395068 -25532 395142 -25476
rect 395198 -25532 395284 -25476
rect 395340 -25532 395408 -25476
rect 395068 -25542 395408 -25532
rect 395468 -17950 395808 -17820
rect 395468 -18006 395545 -17950
rect 395601 -18006 395687 -17950
rect 395743 -18006 395808 -17950
rect 395468 -18092 395808 -18006
rect 395468 -18148 395545 -18092
rect 395601 -18148 395687 -18092
rect 395743 -18148 395808 -18092
rect 395468 -18234 395808 -18148
rect 395468 -18290 395545 -18234
rect 395601 -18290 395687 -18234
rect 395743 -18290 395808 -18234
rect 395468 -18376 395808 -18290
rect 395468 -18432 395545 -18376
rect 395601 -18432 395687 -18376
rect 395743 -18432 395808 -18376
rect 395468 -18518 395808 -18432
rect 395468 -18574 395545 -18518
rect 395601 -18574 395687 -18518
rect 395743 -18574 395808 -18518
rect 395468 -18660 395808 -18574
rect 395468 -18716 395545 -18660
rect 395601 -18716 395687 -18660
rect 395743 -18716 395808 -18660
rect 395468 -18802 395808 -18716
rect 395468 -18858 395545 -18802
rect 395601 -18858 395687 -18802
rect 395743 -18858 395808 -18802
rect 395468 -18944 395808 -18858
rect 395468 -19000 395545 -18944
rect 395601 -19000 395687 -18944
rect 395743 -19000 395808 -18944
rect 395468 -19086 395808 -19000
rect 395468 -19142 395545 -19086
rect 395601 -19142 395687 -19086
rect 395743 -19142 395808 -19086
rect 395468 -19228 395808 -19142
rect 395468 -19284 395545 -19228
rect 395601 -19284 395687 -19228
rect 395743 -19284 395808 -19228
rect 395468 -19370 395808 -19284
rect 395468 -19426 395545 -19370
rect 395601 -19426 395687 -19370
rect 395743 -19426 395808 -19370
rect 395468 -19512 395808 -19426
rect 395468 -19568 395545 -19512
rect 395601 -19568 395687 -19512
rect 395743 -19568 395808 -19512
rect 395468 -19654 395808 -19568
rect 395468 -19710 395545 -19654
rect 395601 -19710 395687 -19654
rect 395743 -19710 395808 -19654
rect 395468 -19796 395808 -19710
rect 395468 -19852 395545 -19796
rect 395601 -19852 395687 -19796
rect 395743 -19852 395808 -19796
rect 395468 -19938 395808 -19852
rect 395468 -19994 395545 -19938
rect 395601 -19994 395687 -19938
rect 395743 -19994 395808 -19938
rect 395468 -20080 395808 -19994
rect 395468 -20136 395545 -20080
rect 395601 -20136 395687 -20080
rect 395743 -20136 395808 -20080
rect 395468 -20222 395808 -20136
rect 395468 -20278 395545 -20222
rect 395601 -20278 395687 -20222
rect 395743 -20278 395808 -20222
rect 395468 -20364 395808 -20278
rect 395468 -20420 395545 -20364
rect 395601 -20420 395687 -20364
rect 395743 -20420 395808 -20364
rect 395468 -20506 395808 -20420
rect 395468 -20562 395545 -20506
rect 395601 -20562 395687 -20506
rect 395743 -20562 395808 -20506
rect 395468 -20648 395808 -20562
rect 395468 -20704 395545 -20648
rect 395601 -20704 395687 -20648
rect 395743 -20704 395808 -20648
rect 395468 -20790 395808 -20704
rect 395468 -20846 395545 -20790
rect 395601 -20846 395687 -20790
rect 395743 -20846 395808 -20790
rect 395468 -20932 395808 -20846
rect 395468 -20988 395545 -20932
rect 395601 -20988 395687 -20932
rect 395743 -20988 395808 -20932
rect 395468 -21074 395808 -20988
rect 395468 -21130 395545 -21074
rect 395601 -21130 395687 -21074
rect 395743 -21130 395808 -21074
rect 395468 -21216 395808 -21130
rect 395468 -21272 395545 -21216
rect 395601 -21272 395687 -21216
rect 395743 -21272 395808 -21216
rect 395468 -21358 395808 -21272
rect 395468 -21414 395545 -21358
rect 395601 -21414 395687 -21358
rect 395743 -21414 395808 -21358
rect 395468 -21500 395808 -21414
rect 395468 -21556 395545 -21500
rect 395601 -21556 395687 -21500
rect 395743 -21556 395808 -21500
rect 395468 -21642 395808 -21556
rect 395468 -21698 395545 -21642
rect 395601 -21698 395687 -21642
rect 395743 -21698 395808 -21642
rect 395468 -21784 395808 -21698
rect 395468 -21840 395545 -21784
rect 395601 -21840 395687 -21784
rect 395743 -21840 395808 -21784
rect 395468 -21926 395808 -21840
rect 395468 -21982 395545 -21926
rect 395601 -21982 395687 -21926
rect 395743 -21982 395808 -21926
rect 395468 -22068 395808 -21982
rect 395468 -22124 395545 -22068
rect 395601 -22124 395687 -22068
rect 395743 -22124 395808 -22068
rect 395468 -22210 395808 -22124
rect 395468 -22266 395545 -22210
rect 395601 -22266 395687 -22210
rect 395743 -22266 395808 -22210
rect 395468 -22352 395808 -22266
rect 395468 -22408 395545 -22352
rect 395601 -22408 395687 -22352
rect 395743 -22408 395808 -22352
rect 395468 -22494 395808 -22408
rect 395468 -22550 395545 -22494
rect 395601 -22550 395687 -22494
rect 395743 -22550 395808 -22494
rect 395468 -22636 395808 -22550
rect 395468 -22692 395545 -22636
rect 395601 -22692 395687 -22636
rect 395743 -22692 395808 -22636
rect 395468 -22778 395808 -22692
rect 395468 -22834 395545 -22778
rect 395601 -22834 395687 -22778
rect 395743 -22834 395808 -22778
rect 395468 -22920 395808 -22834
rect 395468 -22976 395545 -22920
rect 395601 -22976 395687 -22920
rect 395743 -22976 395808 -22920
rect 395468 -23062 395808 -22976
rect 395468 -23118 395545 -23062
rect 395601 -23118 395687 -23062
rect 395743 -23118 395808 -23062
rect 395468 -23204 395808 -23118
rect 395468 -23260 395545 -23204
rect 395601 -23260 395687 -23204
rect 395743 -23260 395808 -23204
rect 395468 -23346 395808 -23260
rect 395468 -23402 395545 -23346
rect 395601 -23402 395687 -23346
rect 395743 -23402 395808 -23346
rect 395468 -23488 395808 -23402
rect 395468 -23544 395545 -23488
rect 395601 -23544 395687 -23488
rect 395743 -23544 395808 -23488
rect 395468 -23630 395808 -23544
rect 395468 -23686 395545 -23630
rect 395601 -23686 395687 -23630
rect 395743 -23686 395808 -23630
rect 395468 -23772 395808 -23686
rect 395468 -23828 395545 -23772
rect 395601 -23828 395687 -23772
rect 395743 -23828 395808 -23772
rect 395468 -23914 395808 -23828
rect 395468 -23970 395545 -23914
rect 395601 -23970 395687 -23914
rect 395743 -23970 395808 -23914
rect 395468 -24056 395808 -23970
rect 395468 -24112 395545 -24056
rect 395601 -24112 395687 -24056
rect 395743 -24112 395808 -24056
rect 395468 -24198 395808 -24112
rect 395468 -24254 395545 -24198
rect 395601 -24254 395687 -24198
rect 395743 -24254 395808 -24198
rect 395468 -24340 395808 -24254
rect 395468 -24396 395545 -24340
rect 395601 -24396 395687 -24340
rect 395743 -24396 395808 -24340
rect 395468 -24482 395808 -24396
rect 395468 -24538 395545 -24482
rect 395601 -24538 395687 -24482
rect 395743 -24538 395808 -24482
rect 395468 -24624 395808 -24538
rect 395468 -24680 395545 -24624
rect 395601 -24680 395687 -24624
rect 395743 -24680 395808 -24624
rect 395468 -24766 395808 -24680
rect 395468 -24822 395545 -24766
rect 395601 -24822 395687 -24766
rect 395743 -24822 395808 -24766
rect 395468 -24908 395808 -24822
rect 395468 -24964 395545 -24908
rect 395601 -24964 395687 -24908
rect 395743 -24964 395808 -24908
rect 395468 -25050 395808 -24964
rect 395468 -25106 395545 -25050
rect 395601 -25106 395687 -25050
rect 395743 -25106 395808 -25050
rect 395468 -25192 395808 -25106
rect 395468 -25248 395545 -25192
rect 395601 -25248 395687 -25192
rect 395743 -25248 395808 -25192
rect 395468 -25334 395808 -25248
rect 395468 -25390 395545 -25334
rect 395601 -25390 395687 -25334
rect 395743 -25390 395808 -25334
rect 395468 -25476 395808 -25390
rect 395468 -25532 395545 -25476
rect 395601 -25532 395687 -25476
rect 395743 -25532 395808 -25476
rect 395468 -25542 395808 -25532
rect 395868 -17950 396208 -17820
rect 395868 -18006 395941 -17950
rect 395997 -18006 396083 -17950
rect 396139 -18006 396208 -17950
rect 395868 -18092 396208 -18006
rect 395868 -18148 395941 -18092
rect 395997 -18148 396083 -18092
rect 396139 -18148 396208 -18092
rect 395868 -18234 396208 -18148
rect 395868 -18290 395941 -18234
rect 395997 -18290 396083 -18234
rect 396139 -18290 396208 -18234
rect 395868 -18376 396208 -18290
rect 395868 -18432 395941 -18376
rect 395997 -18432 396083 -18376
rect 396139 -18432 396208 -18376
rect 395868 -18518 396208 -18432
rect 395868 -18574 395941 -18518
rect 395997 -18574 396083 -18518
rect 396139 -18574 396208 -18518
rect 395868 -18660 396208 -18574
rect 395868 -18716 395941 -18660
rect 395997 -18716 396083 -18660
rect 396139 -18716 396208 -18660
rect 395868 -18802 396208 -18716
rect 395868 -18858 395941 -18802
rect 395997 -18858 396083 -18802
rect 396139 -18858 396208 -18802
rect 395868 -18944 396208 -18858
rect 395868 -19000 395941 -18944
rect 395997 -19000 396083 -18944
rect 396139 -19000 396208 -18944
rect 395868 -19086 396208 -19000
rect 395868 -19142 395941 -19086
rect 395997 -19142 396083 -19086
rect 396139 -19142 396208 -19086
rect 395868 -19228 396208 -19142
rect 395868 -19284 395941 -19228
rect 395997 -19284 396083 -19228
rect 396139 -19284 396208 -19228
rect 395868 -19370 396208 -19284
rect 395868 -19426 395941 -19370
rect 395997 -19426 396083 -19370
rect 396139 -19426 396208 -19370
rect 395868 -19512 396208 -19426
rect 395868 -19568 395941 -19512
rect 395997 -19568 396083 -19512
rect 396139 -19568 396208 -19512
rect 395868 -19654 396208 -19568
rect 395868 -19710 395941 -19654
rect 395997 -19710 396083 -19654
rect 396139 -19710 396208 -19654
rect 395868 -19796 396208 -19710
rect 395868 -19852 395941 -19796
rect 395997 -19852 396083 -19796
rect 396139 -19852 396208 -19796
rect 395868 -19938 396208 -19852
rect 395868 -19994 395941 -19938
rect 395997 -19994 396083 -19938
rect 396139 -19994 396208 -19938
rect 395868 -20080 396208 -19994
rect 395868 -20136 395941 -20080
rect 395997 -20136 396083 -20080
rect 396139 -20136 396208 -20080
rect 395868 -20222 396208 -20136
rect 395868 -20278 395941 -20222
rect 395997 -20278 396083 -20222
rect 396139 -20278 396208 -20222
rect 395868 -20364 396208 -20278
rect 395868 -20420 395941 -20364
rect 395997 -20420 396083 -20364
rect 396139 -20420 396208 -20364
rect 395868 -20506 396208 -20420
rect 395868 -20562 395941 -20506
rect 395997 -20562 396083 -20506
rect 396139 -20562 396208 -20506
rect 395868 -20648 396208 -20562
rect 395868 -20704 395941 -20648
rect 395997 -20704 396083 -20648
rect 396139 -20704 396208 -20648
rect 395868 -20790 396208 -20704
rect 395868 -20846 395941 -20790
rect 395997 -20846 396083 -20790
rect 396139 -20846 396208 -20790
rect 395868 -20932 396208 -20846
rect 395868 -20988 395941 -20932
rect 395997 -20988 396083 -20932
rect 396139 -20988 396208 -20932
rect 395868 -21074 396208 -20988
rect 395868 -21130 395941 -21074
rect 395997 -21130 396083 -21074
rect 396139 -21130 396208 -21074
rect 395868 -21216 396208 -21130
rect 395868 -21272 395941 -21216
rect 395997 -21272 396083 -21216
rect 396139 -21272 396208 -21216
rect 395868 -21358 396208 -21272
rect 395868 -21414 395941 -21358
rect 395997 -21414 396083 -21358
rect 396139 -21414 396208 -21358
rect 395868 -21500 396208 -21414
rect 395868 -21556 395941 -21500
rect 395997 -21556 396083 -21500
rect 396139 -21556 396208 -21500
rect 395868 -21642 396208 -21556
rect 395868 -21698 395941 -21642
rect 395997 -21698 396083 -21642
rect 396139 -21698 396208 -21642
rect 395868 -21784 396208 -21698
rect 395868 -21840 395941 -21784
rect 395997 -21840 396083 -21784
rect 396139 -21840 396208 -21784
rect 395868 -21926 396208 -21840
rect 395868 -21982 395941 -21926
rect 395997 -21982 396083 -21926
rect 396139 -21982 396208 -21926
rect 395868 -22068 396208 -21982
rect 395868 -22124 395941 -22068
rect 395997 -22124 396083 -22068
rect 396139 -22124 396208 -22068
rect 395868 -22210 396208 -22124
rect 395868 -22266 395941 -22210
rect 395997 -22266 396083 -22210
rect 396139 -22266 396208 -22210
rect 395868 -22352 396208 -22266
rect 395868 -22408 395941 -22352
rect 395997 -22408 396083 -22352
rect 396139 -22408 396208 -22352
rect 395868 -22494 396208 -22408
rect 395868 -22550 395941 -22494
rect 395997 -22550 396083 -22494
rect 396139 -22550 396208 -22494
rect 395868 -22636 396208 -22550
rect 395868 -22692 395941 -22636
rect 395997 -22692 396083 -22636
rect 396139 -22692 396208 -22636
rect 395868 -22778 396208 -22692
rect 395868 -22834 395941 -22778
rect 395997 -22834 396083 -22778
rect 396139 -22834 396208 -22778
rect 395868 -22920 396208 -22834
rect 395868 -22976 395941 -22920
rect 395997 -22976 396083 -22920
rect 396139 -22976 396208 -22920
rect 395868 -23062 396208 -22976
rect 395868 -23118 395941 -23062
rect 395997 -23118 396083 -23062
rect 396139 -23118 396208 -23062
rect 395868 -23204 396208 -23118
rect 395868 -23260 395941 -23204
rect 395997 -23260 396083 -23204
rect 396139 -23260 396208 -23204
rect 395868 -23346 396208 -23260
rect 395868 -23402 395941 -23346
rect 395997 -23402 396083 -23346
rect 396139 -23402 396208 -23346
rect 395868 -23488 396208 -23402
rect 395868 -23544 395941 -23488
rect 395997 -23544 396083 -23488
rect 396139 -23544 396208 -23488
rect 395868 -23630 396208 -23544
rect 395868 -23686 395941 -23630
rect 395997 -23686 396083 -23630
rect 396139 -23686 396208 -23630
rect 395868 -23772 396208 -23686
rect 395868 -23828 395941 -23772
rect 395997 -23828 396083 -23772
rect 396139 -23828 396208 -23772
rect 395868 -23914 396208 -23828
rect 395868 -23970 395941 -23914
rect 395997 -23970 396083 -23914
rect 396139 -23970 396208 -23914
rect 395868 -24056 396208 -23970
rect 395868 -24112 395941 -24056
rect 395997 -24112 396083 -24056
rect 396139 -24112 396208 -24056
rect 395868 -24198 396208 -24112
rect 395868 -24254 395941 -24198
rect 395997 -24254 396083 -24198
rect 396139 -24254 396208 -24198
rect 395868 -24340 396208 -24254
rect 395868 -24396 395941 -24340
rect 395997 -24396 396083 -24340
rect 396139 -24396 396208 -24340
rect 395868 -24482 396208 -24396
rect 395868 -24538 395941 -24482
rect 395997 -24538 396083 -24482
rect 396139 -24538 396208 -24482
rect 395868 -24624 396208 -24538
rect 395868 -24680 395941 -24624
rect 395997 -24680 396083 -24624
rect 396139 -24680 396208 -24624
rect 395868 -24766 396208 -24680
rect 395868 -24822 395941 -24766
rect 395997 -24822 396083 -24766
rect 396139 -24822 396208 -24766
rect 395868 -24908 396208 -24822
rect 395868 -24964 395941 -24908
rect 395997 -24964 396083 -24908
rect 396139 -24964 396208 -24908
rect 395868 -25050 396208 -24964
rect 395868 -25106 395941 -25050
rect 395997 -25106 396083 -25050
rect 396139 -25106 396208 -25050
rect 395868 -25192 396208 -25106
rect 395868 -25248 395941 -25192
rect 395997 -25248 396083 -25192
rect 396139 -25248 396208 -25192
rect 395868 -25334 396208 -25248
rect 395868 -25390 395941 -25334
rect 395997 -25390 396083 -25334
rect 396139 -25390 396208 -25334
rect 395868 -25476 396208 -25390
rect 395868 -25532 395941 -25476
rect 395997 -25532 396083 -25476
rect 396139 -25532 396208 -25476
rect 395868 -25542 396208 -25532
rect 396400 -17858 397200 -17820
rect 396400 -17914 396526 -17858
rect 396582 -17914 396650 -17858
rect 396706 -17914 396774 -17858
rect 396830 -17914 396898 -17858
rect 396954 -17914 397022 -17858
rect 397078 -17914 397200 -17858
rect 396400 -17982 397200 -17914
rect 396400 -18038 396526 -17982
rect 396582 -18038 396650 -17982
rect 396706 -18038 396774 -17982
rect 396830 -18038 396898 -17982
rect 396954 -18038 397022 -17982
rect 397078 -18038 397200 -17982
rect 396400 -18106 397200 -18038
rect 396400 -18162 396526 -18106
rect 396582 -18162 396650 -18106
rect 396706 -18162 396774 -18106
rect 396830 -18162 396898 -18106
rect 396954 -18162 397022 -18106
rect 397078 -18162 397200 -18106
rect 396400 -18230 397200 -18162
rect 396400 -18286 396526 -18230
rect 396582 -18286 396650 -18230
rect 396706 -18286 396774 -18230
rect 396830 -18286 396898 -18230
rect 396954 -18286 397022 -18230
rect 397078 -18286 397200 -18230
rect 396400 -18354 397200 -18286
rect 396400 -18410 396526 -18354
rect 396582 -18410 396650 -18354
rect 396706 -18410 396774 -18354
rect 396830 -18410 396898 -18354
rect 396954 -18410 397022 -18354
rect 397078 -18410 397200 -18354
rect 396400 -18478 397200 -18410
rect 396400 -18534 396526 -18478
rect 396582 -18534 396650 -18478
rect 396706 -18534 396774 -18478
rect 396830 -18534 396898 -18478
rect 396954 -18534 397022 -18478
rect 397078 -18534 397200 -18478
rect 396400 -18602 397200 -18534
rect 396400 -18658 396526 -18602
rect 396582 -18658 396650 -18602
rect 396706 -18658 396774 -18602
rect 396830 -18658 396898 -18602
rect 396954 -18658 397022 -18602
rect 397078 -18658 397200 -18602
rect 396400 -18726 397200 -18658
rect 396400 -18782 396526 -18726
rect 396582 -18782 396650 -18726
rect 396706 -18782 396774 -18726
rect 396830 -18782 396898 -18726
rect 396954 -18782 397022 -18726
rect 397078 -18782 397200 -18726
rect 396400 -18850 397200 -18782
rect 396400 -18906 396526 -18850
rect 396582 -18906 396650 -18850
rect 396706 -18906 396774 -18850
rect 396830 -18906 396898 -18850
rect 396954 -18906 397022 -18850
rect 397078 -18906 397200 -18850
rect 396400 -18974 397200 -18906
rect 396400 -19030 396526 -18974
rect 396582 -19030 396650 -18974
rect 396706 -19030 396774 -18974
rect 396830 -19030 396898 -18974
rect 396954 -19030 397022 -18974
rect 397078 -19030 397200 -18974
rect 396400 -19098 397200 -19030
rect 396400 -19154 396526 -19098
rect 396582 -19154 396650 -19098
rect 396706 -19154 396774 -19098
rect 396830 -19154 396898 -19098
rect 396954 -19154 397022 -19098
rect 397078 -19154 397200 -19098
rect 396400 -19222 397200 -19154
rect 396400 -19278 396526 -19222
rect 396582 -19278 396650 -19222
rect 396706 -19278 396774 -19222
rect 396830 -19278 396898 -19222
rect 396954 -19278 397022 -19222
rect 397078 -19278 397200 -19222
rect 396400 -19346 397200 -19278
rect 396400 -19402 396526 -19346
rect 396582 -19402 396650 -19346
rect 396706 -19402 396774 -19346
rect 396830 -19402 396898 -19346
rect 396954 -19402 397022 -19346
rect 397078 -19402 397200 -19346
rect 396400 -19470 397200 -19402
rect 396400 -19526 396526 -19470
rect 396582 -19526 396650 -19470
rect 396706 -19526 396774 -19470
rect 396830 -19526 396898 -19470
rect 396954 -19526 397022 -19470
rect 397078 -19526 397200 -19470
rect 396400 -19594 397200 -19526
rect 396400 -19650 396526 -19594
rect 396582 -19650 396650 -19594
rect 396706 -19650 396774 -19594
rect 396830 -19650 396898 -19594
rect 396954 -19650 397022 -19594
rect 397078 -19650 397200 -19594
rect 396400 -19718 397200 -19650
rect 396400 -19774 396526 -19718
rect 396582 -19774 396650 -19718
rect 396706 -19774 396774 -19718
rect 396830 -19774 396898 -19718
rect 396954 -19774 397022 -19718
rect 397078 -19774 397200 -19718
rect 396400 -19842 397200 -19774
rect 396400 -19898 396526 -19842
rect 396582 -19898 396650 -19842
rect 396706 -19898 396774 -19842
rect 396830 -19898 396898 -19842
rect 396954 -19898 397022 -19842
rect 397078 -19898 397200 -19842
rect 396400 -19966 397200 -19898
rect 396400 -20022 396526 -19966
rect 396582 -20022 396650 -19966
rect 396706 -20022 396774 -19966
rect 396830 -20022 396898 -19966
rect 396954 -20022 397022 -19966
rect 397078 -20022 397200 -19966
rect 396400 -20090 397200 -20022
rect 396400 -20146 396526 -20090
rect 396582 -20146 396650 -20090
rect 396706 -20146 396774 -20090
rect 396830 -20146 396898 -20090
rect 396954 -20146 397022 -20090
rect 397078 -20146 397200 -20090
rect 396400 -20214 397200 -20146
rect 396400 -20270 396526 -20214
rect 396582 -20270 396650 -20214
rect 396706 -20270 396774 -20214
rect 396830 -20270 396898 -20214
rect 396954 -20270 397022 -20214
rect 397078 -20270 397200 -20214
rect 396400 -20338 397200 -20270
rect 396400 -20394 396526 -20338
rect 396582 -20394 396650 -20338
rect 396706 -20394 396774 -20338
rect 396830 -20394 396898 -20338
rect 396954 -20394 397022 -20338
rect 397078 -20394 397200 -20338
rect 396400 -20462 397200 -20394
rect 396400 -20518 396526 -20462
rect 396582 -20518 396650 -20462
rect 396706 -20518 396774 -20462
rect 396830 -20518 396898 -20462
rect 396954 -20518 397022 -20462
rect 397078 -20518 397200 -20462
rect 396400 -20586 397200 -20518
rect 396400 -20642 396526 -20586
rect 396582 -20642 396650 -20586
rect 396706 -20642 396774 -20586
rect 396830 -20642 396898 -20586
rect 396954 -20642 397022 -20586
rect 397078 -20642 397200 -20586
rect 396400 -20710 397200 -20642
rect 396400 -20766 396526 -20710
rect 396582 -20766 396650 -20710
rect 396706 -20766 396774 -20710
rect 396830 -20766 396898 -20710
rect 396954 -20766 397022 -20710
rect 397078 -20766 397200 -20710
rect 396400 -20834 397200 -20766
rect 396400 -20890 396526 -20834
rect 396582 -20890 396650 -20834
rect 396706 -20890 396774 -20834
rect 396830 -20890 396898 -20834
rect 396954 -20890 397022 -20834
rect 397078 -20890 397200 -20834
rect 396400 -20958 397200 -20890
rect 396400 -21014 396526 -20958
rect 396582 -21014 396650 -20958
rect 396706 -21014 396774 -20958
rect 396830 -21014 396898 -20958
rect 396954 -21014 397022 -20958
rect 397078 -21014 397200 -20958
rect 396400 -21082 397200 -21014
rect 396400 -21138 396526 -21082
rect 396582 -21138 396650 -21082
rect 396706 -21138 396774 -21082
rect 396830 -21138 396898 -21082
rect 396954 -21138 397022 -21082
rect 397078 -21138 397200 -21082
rect 396400 -21206 397200 -21138
rect 396400 -21262 396526 -21206
rect 396582 -21262 396650 -21206
rect 396706 -21262 396774 -21206
rect 396830 -21262 396898 -21206
rect 396954 -21262 397022 -21206
rect 397078 -21262 397200 -21206
rect 396400 -21330 397200 -21262
rect 396400 -21386 396526 -21330
rect 396582 -21386 396650 -21330
rect 396706 -21386 396774 -21330
rect 396830 -21386 396898 -21330
rect 396954 -21386 397022 -21330
rect 397078 -21386 397200 -21330
rect 396400 -21454 397200 -21386
rect 396400 -21510 396526 -21454
rect 396582 -21510 396650 -21454
rect 396706 -21510 396774 -21454
rect 396830 -21510 396898 -21454
rect 396954 -21510 397022 -21454
rect 397078 -21510 397200 -21454
rect 396400 -21578 397200 -21510
rect 396400 -21634 396526 -21578
rect 396582 -21634 396650 -21578
rect 396706 -21634 396774 -21578
rect 396830 -21634 396898 -21578
rect 396954 -21634 397022 -21578
rect 397078 -21634 397200 -21578
rect 396400 -21702 397200 -21634
rect 396400 -21758 396526 -21702
rect 396582 -21758 396650 -21702
rect 396706 -21758 396774 -21702
rect 396830 -21758 396898 -21702
rect 396954 -21758 397022 -21702
rect 397078 -21758 397200 -21702
rect 396400 -21826 397200 -21758
rect 396400 -21882 396526 -21826
rect 396582 -21882 396650 -21826
rect 396706 -21882 396774 -21826
rect 396830 -21882 396898 -21826
rect 396954 -21882 397022 -21826
rect 397078 -21882 397200 -21826
rect 396400 -21950 397200 -21882
rect 396400 -22006 396526 -21950
rect 396582 -22006 396650 -21950
rect 396706 -22006 396774 -21950
rect 396830 -22006 396898 -21950
rect 396954 -22006 397022 -21950
rect 397078 -22006 397200 -21950
rect 396400 -22074 397200 -22006
rect 396400 -22130 396526 -22074
rect 396582 -22130 396650 -22074
rect 396706 -22130 396774 -22074
rect 396830 -22130 396898 -22074
rect 396954 -22130 397022 -22074
rect 397078 -22130 397200 -22074
rect 396400 -22198 397200 -22130
rect 396400 -22254 396526 -22198
rect 396582 -22254 396650 -22198
rect 396706 -22254 396774 -22198
rect 396830 -22254 396898 -22198
rect 396954 -22254 397022 -22198
rect 397078 -22254 397200 -22198
rect 396400 -22322 397200 -22254
rect 396400 -22378 396526 -22322
rect 396582 -22378 396650 -22322
rect 396706 -22378 396774 -22322
rect 396830 -22378 396898 -22322
rect 396954 -22378 397022 -22322
rect 397078 -22378 397200 -22322
rect 396400 -22446 397200 -22378
rect 396400 -22502 396526 -22446
rect 396582 -22502 396650 -22446
rect 396706 -22502 396774 -22446
rect 396830 -22502 396898 -22446
rect 396954 -22502 397022 -22446
rect 397078 -22502 397200 -22446
rect 396400 -22570 397200 -22502
rect 396400 -22626 396526 -22570
rect 396582 -22626 396650 -22570
rect 396706 -22626 396774 -22570
rect 396830 -22626 396898 -22570
rect 396954 -22626 397022 -22570
rect 397078 -22626 397200 -22570
rect 396400 -22694 397200 -22626
rect 396400 -22750 396526 -22694
rect 396582 -22750 396650 -22694
rect 396706 -22750 396774 -22694
rect 396830 -22750 396898 -22694
rect 396954 -22750 397022 -22694
rect 397078 -22750 397200 -22694
rect 396400 -22818 397200 -22750
rect 396400 -22874 396526 -22818
rect 396582 -22874 396650 -22818
rect 396706 -22874 396774 -22818
rect 396830 -22874 396898 -22818
rect 396954 -22874 397022 -22818
rect 397078 -22874 397200 -22818
rect 396400 -22942 397200 -22874
rect 396400 -22998 396526 -22942
rect 396582 -22998 396650 -22942
rect 396706 -22998 396774 -22942
rect 396830 -22998 396898 -22942
rect 396954 -22998 397022 -22942
rect 397078 -22998 397200 -22942
rect 396400 -23066 397200 -22998
rect 396400 -23122 396526 -23066
rect 396582 -23122 396650 -23066
rect 396706 -23122 396774 -23066
rect 396830 -23122 396898 -23066
rect 396954 -23122 397022 -23066
rect 397078 -23122 397200 -23066
rect 396400 -23190 397200 -23122
rect 396400 -23246 396526 -23190
rect 396582 -23246 396650 -23190
rect 396706 -23246 396774 -23190
rect 396830 -23246 396898 -23190
rect 396954 -23246 397022 -23190
rect 397078 -23246 397200 -23190
rect 396400 -23314 397200 -23246
rect 396400 -23370 396526 -23314
rect 396582 -23370 396650 -23314
rect 396706 -23370 396774 -23314
rect 396830 -23370 396898 -23314
rect 396954 -23370 397022 -23314
rect 397078 -23370 397200 -23314
rect 396400 -23438 397200 -23370
rect 396400 -23494 396526 -23438
rect 396582 -23494 396650 -23438
rect 396706 -23494 396774 -23438
rect 396830 -23494 396898 -23438
rect 396954 -23494 397022 -23438
rect 397078 -23494 397200 -23438
rect 396400 -23562 397200 -23494
rect 396400 -23618 396526 -23562
rect 396582 -23618 396650 -23562
rect 396706 -23618 396774 -23562
rect 396830 -23618 396898 -23562
rect 396954 -23618 397022 -23562
rect 397078 -23618 397200 -23562
rect 396400 -23686 397200 -23618
rect 396400 -23742 396526 -23686
rect 396582 -23742 396650 -23686
rect 396706 -23742 396774 -23686
rect 396830 -23742 396898 -23686
rect 396954 -23742 397022 -23686
rect 397078 -23742 397200 -23686
rect 396400 -23810 397200 -23742
rect 396400 -23866 396526 -23810
rect 396582 -23866 396650 -23810
rect 396706 -23866 396774 -23810
rect 396830 -23866 396898 -23810
rect 396954 -23866 397022 -23810
rect 397078 -23866 397200 -23810
rect 396400 -23934 397200 -23866
rect 396400 -23990 396526 -23934
rect 396582 -23990 396650 -23934
rect 396706 -23990 396774 -23934
rect 396830 -23990 396898 -23934
rect 396954 -23990 397022 -23934
rect 397078 -23990 397200 -23934
rect 396400 -24058 397200 -23990
rect 396400 -24114 396526 -24058
rect 396582 -24114 396650 -24058
rect 396706 -24114 396774 -24058
rect 396830 -24114 396898 -24058
rect 396954 -24114 397022 -24058
rect 397078 -24114 397200 -24058
rect 396400 -24182 397200 -24114
rect 396400 -24238 396526 -24182
rect 396582 -24238 396650 -24182
rect 396706 -24238 396774 -24182
rect 396830 -24238 396898 -24182
rect 396954 -24238 397022 -24182
rect 397078 -24238 397200 -24182
rect 396400 -24306 397200 -24238
rect 396400 -24362 396526 -24306
rect 396582 -24362 396650 -24306
rect 396706 -24362 396774 -24306
rect 396830 -24362 396898 -24306
rect 396954 -24362 397022 -24306
rect 397078 -24362 397200 -24306
rect 396400 -24430 397200 -24362
rect 396400 -24486 396526 -24430
rect 396582 -24486 396650 -24430
rect 396706 -24486 396774 -24430
rect 396830 -24486 396898 -24430
rect 396954 -24486 397022 -24430
rect 397078 -24486 397200 -24430
rect 396400 -24554 397200 -24486
rect 396400 -24610 396526 -24554
rect 396582 -24610 396650 -24554
rect 396706 -24610 396774 -24554
rect 396830 -24610 396898 -24554
rect 396954 -24610 397022 -24554
rect 397078 -24610 397200 -24554
rect 396400 -24678 397200 -24610
rect 396400 -24734 396526 -24678
rect 396582 -24734 396650 -24678
rect 396706 -24734 396774 -24678
rect 396830 -24734 396898 -24678
rect 396954 -24734 397022 -24678
rect 397078 -24734 397200 -24678
rect 396400 -24802 397200 -24734
rect 396400 -24858 396526 -24802
rect 396582 -24858 396650 -24802
rect 396706 -24858 396774 -24802
rect 396830 -24858 396898 -24802
rect 396954 -24858 397022 -24802
rect 397078 -24858 397200 -24802
rect 396400 -24926 397200 -24858
rect 396400 -24982 396526 -24926
rect 396582 -24982 396650 -24926
rect 396706 -24982 396774 -24926
rect 396830 -24982 396898 -24926
rect 396954 -24982 397022 -24926
rect 397078 -24982 397200 -24926
rect 396400 -25050 397200 -24982
rect 396400 -25106 396526 -25050
rect 396582 -25106 396650 -25050
rect 396706 -25106 396774 -25050
rect 396830 -25106 396898 -25050
rect 396954 -25106 397022 -25050
rect 397078 -25106 397200 -25050
rect 396400 -25174 397200 -25106
rect 396400 -25230 396526 -25174
rect 396582 -25230 396650 -25174
rect 396706 -25230 396774 -25174
rect 396830 -25230 396898 -25174
rect 396954 -25230 397022 -25174
rect 397078 -25230 397200 -25174
rect 396400 -25298 397200 -25230
rect 396400 -25354 396526 -25298
rect 396582 -25354 396650 -25298
rect 396706 -25354 396774 -25298
rect 396830 -25354 396898 -25298
rect 396954 -25354 397022 -25298
rect 397078 -25354 397200 -25298
rect 396400 -25422 397200 -25354
rect 396400 -25478 396526 -25422
rect 396582 -25478 396650 -25422
rect 396706 -25478 396774 -25422
rect 396830 -25478 396898 -25422
rect 396954 -25478 397022 -25422
rect 397078 -25478 397200 -25422
rect 396400 -25542 397200 -25478
rect 388000 -25721 397200 -25542
rect 388000 -25777 388146 -25721
rect 388202 -25777 388270 -25721
rect 388326 -25777 388394 -25721
rect 388450 -25777 388518 -25721
rect 388574 -25777 388642 -25721
rect 388698 -25777 388766 -25721
rect 388822 -25777 388890 -25721
rect 388946 -25777 389014 -25721
rect 389070 -25777 389138 -25721
rect 389194 -25777 389262 -25721
rect 389318 -25777 389386 -25721
rect 389442 -25777 389510 -25721
rect 389566 -25777 389634 -25721
rect 389690 -25777 389758 -25721
rect 389814 -25777 389882 -25721
rect 389938 -25777 390006 -25721
rect 390062 -25777 390130 -25721
rect 390186 -25777 390254 -25721
rect 390310 -25777 390378 -25721
rect 390434 -25777 390502 -25721
rect 390558 -25777 390626 -25721
rect 390682 -25777 390750 -25721
rect 390806 -25777 390874 -25721
rect 390930 -25777 390998 -25721
rect 391054 -25777 391122 -25721
rect 391178 -25777 391246 -25721
rect 391302 -25777 391370 -25721
rect 391426 -25777 391494 -25721
rect 391550 -25777 391618 -25721
rect 391674 -25777 391742 -25721
rect 391798 -25777 391866 -25721
rect 391922 -25777 391990 -25721
rect 392046 -25777 392114 -25721
rect 392170 -25777 392238 -25721
rect 392294 -25777 392362 -25721
rect 392418 -25777 392486 -25721
rect 392542 -25777 392610 -25721
rect 392666 -25777 392734 -25721
rect 392790 -25777 392858 -25721
rect 392914 -25777 392982 -25721
rect 393038 -25777 393106 -25721
rect 393162 -25777 393230 -25721
rect 393286 -25777 393354 -25721
rect 393410 -25777 393478 -25721
rect 393534 -25777 393602 -25721
rect 393658 -25777 393726 -25721
rect 393782 -25777 393850 -25721
rect 393906 -25777 393974 -25721
rect 394030 -25777 394098 -25721
rect 394154 -25777 394222 -25721
rect 394278 -25777 394346 -25721
rect 394402 -25777 394470 -25721
rect 394526 -25777 394594 -25721
rect 394650 -25777 394718 -25721
rect 394774 -25777 394842 -25721
rect 394898 -25777 394966 -25721
rect 395022 -25777 395090 -25721
rect 395146 -25777 395214 -25721
rect 395270 -25777 395338 -25721
rect 395394 -25777 395462 -25721
rect 395518 -25777 395586 -25721
rect 395642 -25777 395710 -25721
rect 395766 -25777 395898 -25721
rect 395954 -25777 396022 -25721
rect 396078 -25777 396146 -25721
rect 396202 -25777 396270 -25721
rect 396326 -25777 396394 -25721
rect 396450 -25777 396518 -25721
rect 396574 -25777 396642 -25721
rect 396698 -25777 396766 -25721
rect 396822 -25777 396890 -25721
rect 396946 -25777 397014 -25721
rect 397070 -25777 397200 -25721
rect 388000 -25845 397200 -25777
rect 388000 -25901 388146 -25845
rect 388202 -25901 388270 -25845
rect 388326 -25901 388394 -25845
rect 388450 -25901 388518 -25845
rect 388574 -25901 388642 -25845
rect 388698 -25901 388766 -25845
rect 388822 -25901 388890 -25845
rect 388946 -25901 389014 -25845
rect 389070 -25901 389138 -25845
rect 389194 -25901 389262 -25845
rect 389318 -25901 389386 -25845
rect 389442 -25901 389510 -25845
rect 389566 -25901 389634 -25845
rect 389690 -25901 389758 -25845
rect 389814 -25901 389882 -25845
rect 389938 -25901 390006 -25845
rect 390062 -25901 390130 -25845
rect 390186 -25901 390254 -25845
rect 390310 -25901 390378 -25845
rect 390434 -25901 390502 -25845
rect 390558 -25901 390626 -25845
rect 390682 -25901 390750 -25845
rect 390806 -25901 390874 -25845
rect 390930 -25901 390998 -25845
rect 391054 -25901 391122 -25845
rect 391178 -25901 391246 -25845
rect 391302 -25901 391370 -25845
rect 391426 -25901 391494 -25845
rect 391550 -25901 391618 -25845
rect 391674 -25901 391742 -25845
rect 391798 -25901 391866 -25845
rect 391922 -25901 391990 -25845
rect 392046 -25901 392114 -25845
rect 392170 -25901 392238 -25845
rect 392294 -25901 392362 -25845
rect 392418 -25901 392486 -25845
rect 392542 -25901 392610 -25845
rect 392666 -25901 392734 -25845
rect 392790 -25901 392858 -25845
rect 392914 -25901 392982 -25845
rect 393038 -25901 393106 -25845
rect 393162 -25901 393230 -25845
rect 393286 -25901 393354 -25845
rect 393410 -25901 393478 -25845
rect 393534 -25901 393602 -25845
rect 393658 -25901 393726 -25845
rect 393782 -25901 393850 -25845
rect 393906 -25901 393974 -25845
rect 394030 -25901 394098 -25845
rect 394154 -25901 394222 -25845
rect 394278 -25901 394346 -25845
rect 394402 -25901 394470 -25845
rect 394526 -25901 394594 -25845
rect 394650 -25901 394718 -25845
rect 394774 -25901 394842 -25845
rect 394898 -25901 394966 -25845
rect 395022 -25901 395090 -25845
rect 395146 -25901 395214 -25845
rect 395270 -25901 395338 -25845
rect 395394 -25901 395462 -25845
rect 395518 -25901 395586 -25845
rect 395642 -25901 395710 -25845
rect 395766 -25901 395898 -25845
rect 395954 -25901 396022 -25845
rect 396078 -25901 396146 -25845
rect 396202 -25901 396270 -25845
rect 396326 -25901 396394 -25845
rect 396450 -25901 396518 -25845
rect 396574 -25901 396642 -25845
rect 396698 -25901 396766 -25845
rect 396822 -25901 396890 -25845
rect 396946 -25901 397014 -25845
rect 397070 -25901 397200 -25845
rect 388000 -25969 397200 -25901
rect 388000 -26025 388146 -25969
rect 388202 -26025 388270 -25969
rect 388326 -26025 388394 -25969
rect 388450 -26025 388518 -25969
rect 388574 -26025 388642 -25969
rect 388698 -26025 388766 -25969
rect 388822 -26025 388890 -25969
rect 388946 -26025 389014 -25969
rect 389070 -26025 389138 -25969
rect 389194 -26025 389262 -25969
rect 389318 -26025 389386 -25969
rect 389442 -26025 389510 -25969
rect 389566 -26025 389634 -25969
rect 389690 -26025 389758 -25969
rect 389814 -26025 389882 -25969
rect 389938 -26025 390006 -25969
rect 390062 -26025 390130 -25969
rect 390186 -26025 390254 -25969
rect 390310 -26025 390378 -25969
rect 390434 -26025 390502 -25969
rect 390558 -26025 390626 -25969
rect 390682 -26025 390750 -25969
rect 390806 -26025 390874 -25969
rect 390930 -26025 390998 -25969
rect 391054 -26025 391122 -25969
rect 391178 -26025 391246 -25969
rect 391302 -26025 391370 -25969
rect 391426 -26025 391494 -25969
rect 391550 -26025 391618 -25969
rect 391674 -26025 391742 -25969
rect 391798 -26025 391866 -25969
rect 391922 -26025 391990 -25969
rect 392046 -26025 392114 -25969
rect 392170 -26025 392238 -25969
rect 392294 -26025 392362 -25969
rect 392418 -26025 392486 -25969
rect 392542 -26025 392610 -25969
rect 392666 -26025 392734 -25969
rect 392790 -26025 392858 -25969
rect 392914 -26025 392982 -25969
rect 393038 -26025 393106 -25969
rect 393162 -26025 393230 -25969
rect 393286 -26025 393354 -25969
rect 393410 -26025 393478 -25969
rect 393534 -26025 393602 -25969
rect 393658 -26025 393726 -25969
rect 393782 -26025 393850 -25969
rect 393906 -26025 393974 -25969
rect 394030 -26025 394098 -25969
rect 394154 -26025 394222 -25969
rect 394278 -26025 394346 -25969
rect 394402 -26025 394470 -25969
rect 394526 -26025 394594 -25969
rect 394650 -26025 394718 -25969
rect 394774 -26025 394842 -25969
rect 394898 -26025 394966 -25969
rect 395022 -26025 395090 -25969
rect 395146 -26025 395214 -25969
rect 395270 -26025 395338 -25969
rect 395394 -26025 395462 -25969
rect 395518 -26025 395586 -25969
rect 395642 -26025 395710 -25969
rect 395766 -26025 395898 -25969
rect 395954 -26025 396022 -25969
rect 396078 -26025 396146 -25969
rect 396202 -26025 396270 -25969
rect 396326 -26025 396394 -25969
rect 396450 -26025 396518 -25969
rect 396574 -26025 396642 -25969
rect 396698 -26025 396766 -25969
rect 396822 -26025 396890 -25969
rect 396946 -26025 397014 -25969
rect 397070 -26025 397200 -25969
rect 388000 -26093 397200 -26025
rect 388000 -26149 388146 -26093
rect 388202 -26149 388270 -26093
rect 388326 -26149 388394 -26093
rect 388450 -26149 388518 -26093
rect 388574 -26149 388642 -26093
rect 388698 -26149 388766 -26093
rect 388822 -26149 388890 -26093
rect 388946 -26149 389014 -26093
rect 389070 -26149 389138 -26093
rect 389194 -26149 389262 -26093
rect 389318 -26149 389386 -26093
rect 389442 -26149 389510 -26093
rect 389566 -26149 389634 -26093
rect 389690 -26149 389758 -26093
rect 389814 -26149 389882 -26093
rect 389938 -26149 390006 -26093
rect 390062 -26149 390130 -26093
rect 390186 -26149 390254 -26093
rect 390310 -26149 390378 -26093
rect 390434 -26149 390502 -26093
rect 390558 -26149 390626 -26093
rect 390682 -26149 390750 -26093
rect 390806 -26149 390874 -26093
rect 390930 -26149 390998 -26093
rect 391054 -26149 391122 -26093
rect 391178 -26149 391246 -26093
rect 391302 -26149 391370 -26093
rect 391426 -26149 391494 -26093
rect 391550 -26149 391618 -26093
rect 391674 -26149 391742 -26093
rect 391798 -26149 391866 -26093
rect 391922 -26149 391990 -26093
rect 392046 -26149 392114 -26093
rect 392170 -26149 392238 -26093
rect 392294 -26149 392362 -26093
rect 392418 -26149 392486 -26093
rect 392542 -26149 392610 -26093
rect 392666 -26149 392734 -26093
rect 392790 -26149 392858 -26093
rect 392914 -26149 392982 -26093
rect 393038 -26149 393106 -26093
rect 393162 -26149 393230 -26093
rect 393286 -26149 393354 -26093
rect 393410 -26149 393478 -26093
rect 393534 -26149 393602 -26093
rect 393658 -26149 393726 -26093
rect 393782 -26149 393850 -26093
rect 393906 -26149 393974 -26093
rect 394030 -26149 394098 -26093
rect 394154 -26149 394222 -26093
rect 394278 -26149 394346 -26093
rect 394402 -26149 394470 -26093
rect 394526 -26149 394594 -26093
rect 394650 -26149 394718 -26093
rect 394774 -26149 394842 -26093
rect 394898 -26149 394966 -26093
rect 395022 -26149 395090 -26093
rect 395146 -26149 395214 -26093
rect 395270 -26149 395338 -26093
rect 395394 -26149 395462 -26093
rect 395518 -26149 395586 -26093
rect 395642 -26149 395710 -26093
rect 395766 -26149 395898 -26093
rect 395954 -26149 396022 -26093
rect 396078 -26149 396146 -26093
rect 396202 -26149 396270 -26093
rect 396326 -26149 396394 -26093
rect 396450 -26149 396518 -26093
rect 396574 -26149 396642 -26093
rect 396698 -26149 396766 -26093
rect 396822 -26149 396890 -26093
rect 396946 -26149 397014 -26093
rect 397070 -26149 397200 -26093
rect 388000 -26270 397200 -26149
<< via3 >>
rect 388146 -17247 388202 -17191
rect 388270 -17247 388326 -17191
rect 388394 -17247 388450 -17191
rect 388518 -17247 388574 -17191
rect 388642 -17247 388698 -17191
rect 388766 -17247 388822 -17191
rect 388890 -17247 388946 -17191
rect 389014 -17247 389070 -17191
rect 389138 -17247 389194 -17191
rect 389262 -17247 389318 -17191
rect 389386 -17247 389442 -17191
rect 389510 -17247 389566 -17191
rect 389634 -17247 389690 -17191
rect 389758 -17247 389814 -17191
rect 389882 -17247 389938 -17191
rect 390006 -17247 390062 -17191
rect 390130 -17247 390186 -17191
rect 390254 -17247 390310 -17191
rect 390378 -17247 390434 -17191
rect 390502 -17247 390558 -17191
rect 390626 -17247 390682 -17191
rect 390750 -17247 390806 -17191
rect 390874 -17247 390930 -17191
rect 390998 -17247 391054 -17191
rect 391122 -17247 391178 -17191
rect 391246 -17247 391302 -17191
rect 391370 -17247 391426 -17191
rect 391494 -17247 391550 -17191
rect 391618 -17247 391674 -17191
rect 391742 -17247 391798 -17191
rect 391866 -17247 391922 -17191
rect 391990 -17247 392046 -17191
rect 392114 -17247 392170 -17191
rect 392238 -17247 392294 -17191
rect 392362 -17247 392418 -17191
rect 392486 -17247 392542 -17191
rect 392610 -17247 392666 -17191
rect 392734 -17247 392790 -17191
rect 392858 -17247 392914 -17191
rect 392982 -17247 393038 -17191
rect 393106 -17247 393162 -17191
rect 393230 -17247 393286 -17191
rect 393354 -17247 393410 -17191
rect 393478 -17247 393534 -17191
rect 393602 -17247 393658 -17191
rect 393726 -17247 393782 -17191
rect 393850 -17247 393906 -17191
rect 393974 -17247 394030 -17191
rect 394098 -17247 394154 -17191
rect 394222 -17247 394278 -17191
rect 394346 -17247 394402 -17191
rect 394470 -17247 394526 -17191
rect 394594 -17247 394650 -17191
rect 394718 -17247 394774 -17191
rect 394842 -17247 394898 -17191
rect 394966 -17247 395022 -17191
rect 395090 -17247 395146 -17191
rect 395214 -17247 395270 -17191
rect 395338 -17247 395394 -17191
rect 395462 -17247 395518 -17191
rect 395586 -17247 395642 -17191
rect 395710 -17247 395766 -17191
rect 395898 -17247 395954 -17191
rect 396022 -17247 396078 -17191
rect 396146 -17247 396202 -17191
rect 396270 -17247 396326 -17191
rect 396394 -17247 396450 -17191
rect 396518 -17247 396574 -17191
rect 396642 -17247 396698 -17191
rect 396766 -17247 396822 -17191
rect 396890 -17247 396946 -17191
rect 397014 -17247 397070 -17191
rect 388146 -17371 388202 -17315
rect 388270 -17371 388326 -17315
rect 388394 -17371 388450 -17315
rect 388518 -17371 388574 -17315
rect 388642 -17371 388698 -17315
rect 388766 -17371 388822 -17315
rect 388890 -17371 388946 -17315
rect 389014 -17371 389070 -17315
rect 389138 -17371 389194 -17315
rect 389262 -17371 389318 -17315
rect 389386 -17371 389442 -17315
rect 389510 -17371 389566 -17315
rect 389634 -17371 389690 -17315
rect 389758 -17371 389814 -17315
rect 389882 -17371 389938 -17315
rect 390006 -17371 390062 -17315
rect 390130 -17371 390186 -17315
rect 390254 -17371 390310 -17315
rect 390378 -17371 390434 -17315
rect 390502 -17371 390558 -17315
rect 390626 -17371 390682 -17315
rect 390750 -17371 390806 -17315
rect 390874 -17371 390930 -17315
rect 390998 -17371 391054 -17315
rect 391122 -17371 391178 -17315
rect 391246 -17371 391302 -17315
rect 391370 -17371 391426 -17315
rect 391494 -17371 391550 -17315
rect 391618 -17371 391674 -17315
rect 391742 -17371 391798 -17315
rect 391866 -17371 391922 -17315
rect 391990 -17371 392046 -17315
rect 392114 -17371 392170 -17315
rect 392238 -17371 392294 -17315
rect 392362 -17371 392418 -17315
rect 392486 -17371 392542 -17315
rect 392610 -17371 392666 -17315
rect 392734 -17371 392790 -17315
rect 392858 -17371 392914 -17315
rect 392982 -17371 393038 -17315
rect 393106 -17371 393162 -17315
rect 393230 -17371 393286 -17315
rect 393354 -17371 393410 -17315
rect 393478 -17371 393534 -17315
rect 393602 -17371 393658 -17315
rect 393726 -17371 393782 -17315
rect 393850 -17371 393906 -17315
rect 393974 -17371 394030 -17315
rect 394098 -17371 394154 -17315
rect 394222 -17371 394278 -17315
rect 394346 -17371 394402 -17315
rect 394470 -17371 394526 -17315
rect 394594 -17371 394650 -17315
rect 394718 -17371 394774 -17315
rect 394842 -17371 394898 -17315
rect 394966 -17371 395022 -17315
rect 395090 -17371 395146 -17315
rect 395214 -17371 395270 -17315
rect 395338 -17371 395394 -17315
rect 395462 -17371 395518 -17315
rect 395586 -17371 395642 -17315
rect 395710 -17371 395766 -17315
rect 395898 -17371 395954 -17315
rect 396022 -17371 396078 -17315
rect 396146 -17371 396202 -17315
rect 396270 -17371 396326 -17315
rect 396394 -17371 396450 -17315
rect 396518 -17371 396574 -17315
rect 396642 -17371 396698 -17315
rect 396766 -17371 396822 -17315
rect 396890 -17371 396946 -17315
rect 397014 -17371 397070 -17315
rect 388146 -17495 388202 -17439
rect 388270 -17495 388326 -17439
rect 388394 -17495 388450 -17439
rect 388518 -17495 388574 -17439
rect 388642 -17495 388698 -17439
rect 388766 -17495 388822 -17439
rect 388890 -17495 388946 -17439
rect 389014 -17495 389070 -17439
rect 389138 -17495 389194 -17439
rect 389262 -17495 389318 -17439
rect 389386 -17495 389442 -17439
rect 389510 -17495 389566 -17439
rect 389634 -17495 389690 -17439
rect 389758 -17495 389814 -17439
rect 389882 -17495 389938 -17439
rect 390006 -17495 390062 -17439
rect 390130 -17495 390186 -17439
rect 390254 -17495 390310 -17439
rect 390378 -17495 390434 -17439
rect 390502 -17495 390558 -17439
rect 390626 -17495 390682 -17439
rect 390750 -17495 390806 -17439
rect 390874 -17495 390930 -17439
rect 390998 -17495 391054 -17439
rect 391122 -17495 391178 -17439
rect 391246 -17495 391302 -17439
rect 391370 -17495 391426 -17439
rect 391494 -17495 391550 -17439
rect 391618 -17495 391674 -17439
rect 391742 -17495 391798 -17439
rect 391866 -17495 391922 -17439
rect 391990 -17495 392046 -17439
rect 392114 -17495 392170 -17439
rect 392238 -17495 392294 -17439
rect 392362 -17495 392418 -17439
rect 392486 -17495 392542 -17439
rect 392610 -17495 392666 -17439
rect 392734 -17495 392790 -17439
rect 392858 -17495 392914 -17439
rect 392982 -17495 393038 -17439
rect 393106 -17495 393162 -17439
rect 393230 -17495 393286 -17439
rect 393354 -17495 393410 -17439
rect 393478 -17495 393534 -17439
rect 393602 -17495 393658 -17439
rect 393726 -17495 393782 -17439
rect 393850 -17495 393906 -17439
rect 393974 -17495 394030 -17439
rect 394098 -17495 394154 -17439
rect 394222 -17495 394278 -17439
rect 394346 -17495 394402 -17439
rect 394470 -17495 394526 -17439
rect 394594 -17495 394650 -17439
rect 394718 -17495 394774 -17439
rect 394842 -17495 394898 -17439
rect 394966 -17495 395022 -17439
rect 395090 -17495 395146 -17439
rect 395214 -17495 395270 -17439
rect 395338 -17495 395394 -17439
rect 395462 -17495 395518 -17439
rect 395586 -17495 395642 -17439
rect 395710 -17495 395766 -17439
rect 395898 -17495 395954 -17439
rect 396022 -17495 396078 -17439
rect 396146 -17495 396202 -17439
rect 396270 -17495 396326 -17439
rect 396394 -17495 396450 -17439
rect 396518 -17495 396574 -17439
rect 396642 -17495 396698 -17439
rect 396766 -17495 396822 -17439
rect 396890 -17495 396946 -17439
rect 397014 -17495 397070 -17439
rect 388146 -17619 388202 -17563
rect 388270 -17619 388326 -17563
rect 388394 -17619 388450 -17563
rect 388518 -17619 388574 -17563
rect 388642 -17619 388698 -17563
rect 388766 -17619 388822 -17563
rect 388890 -17619 388946 -17563
rect 389014 -17619 389070 -17563
rect 389138 -17619 389194 -17563
rect 389262 -17619 389318 -17563
rect 389386 -17619 389442 -17563
rect 389510 -17619 389566 -17563
rect 389634 -17619 389690 -17563
rect 389758 -17619 389814 -17563
rect 389882 -17619 389938 -17563
rect 390006 -17619 390062 -17563
rect 390130 -17619 390186 -17563
rect 390254 -17619 390310 -17563
rect 390378 -17619 390434 -17563
rect 390502 -17619 390558 -17563
rect 390626 -17619 390682 -17563
rect 390750 -17619 390806 -17563
rect 390874 -17619 390930 -17563
rect 390998 -17619 391054 -17563
rect 391122 -17619 391178 -17563
rect 391246 -17619 391302 -17563
rect 391370 -17619 391426 -17563
rect 391494 -17619 391550 -17563
rect 391618 -17619 391674 -17563
rect 391742 -17619 391798 -17563
rect 391866 -17619 391922 -17563
rect 391990 -17619 392046 -17563
rect 392114 -17619 392170 -17563
rect 392238 -17619 392294 -17563
rect 392362 -17619 392418 -17563
rect 392486 -17619 392542 -17563
rect 392610 -17619 392666 -17563
rect 392734 -17619 392790 -17563
rect 392858 -17619 392914 -17563
rect 392982 -17619 393038 -17563
rect 393106 -17619 393162 -17563
rect 393230 -17619 393286 -17563
rect 393354 -17619 393410 -17563
rect 393478 -17619 393534 -17563
rect 393602 -17619 393658 -17563
rect 393726 -17619 393782 -17563
rect 393850 -17619 393906 -17563
rect 393974 -17619 394030 -17563
rect 394098 -17619 394154 -17563
rect 394222 -17619 394278 -17563
rect 394346 -17619 394402 -17563
rect 394470 -17619 394526 -17563
rect 394594 -17619 394650 -17563
rect 394718 -17619 394774 -17563
rect 394842 -17619 394898 -17563
rect 394966 -17619 395022 -17563
rect 395090 -17619 395146 -17563
rect 395214 -17619 395270 -17563
rect 395338 -17619 395394 -17563
rect 395462 -17619 395518 -17563
rect 395586 -17619 395642 -17563
rect 395710 -17619 395766 -17563
rect 395898 -17619 395954 -17563
rect 396022 -17619 396078 -17563
rect 396146 -17619 396202 -17563
rect 396270 -17619 396326 -17563
rect 396394 -17619 396450 -17563
rect 396518 -17619 396574 -17563
rect 396642 -17619 396698 -17563
rect 396766 -17619 396822 -17563
rect 396890 -17619 396946 -17563
rect 397014 -17619 397070 -17563
rect 388114 -17914 388170 -17858
rect 388238 -17914 388294 -17858
rect 388362 -17914 388418 -17858
rect 388486 -17914 388542 -17858
rect 388610 -17914 388666 -17858
rect 388114 -18038 388170 -17982
rect 388238 -18038 388294 -17982
rect 388362 -18038 388418 -17982
rect 388486 -18038 388542 -17982
rect 388610 -18038 388666 -17982
rect 388114 -18162 388170 -18106
rect 388238 -18162 388294 -18106
rect 388362 -18162 388418 -18106
rect 388486 -18162 388542 -18106
rect 388610 -18162 388666 -18106
rect 388114 -18286 388170 -18230
rect 388238 -18286 388294 -18230
rect 388362 -18286 388418 -18230
rect 388486 -18286 388542 -18230
rect 388610 -18286 388666 -18230
rect 388114 -18410 388170 -18354
rect 388238 -18410 388294 -18354
rect 388362 -18410 388418 -18354
rect 388486 -18410 388542 -18354
rect 388610 -18410 388666 -18354
rect 388114 -18534 388170 -18478
rect 388238 -18534 388294 -18478
rect 388362 -18534 388418 -18478
rect 388486 -18534 388542 -18478
rect 388610 -18534 388666 -18478
rect 388114 -18658 388170 -18602
rect 388238 -18658 388294 -18602
rect 388362 -18658 388418 -18602
rect 388486 -18658 388542 -18602
rect 388610 -18658 388666 -18602
rect 388114 -18782 388170 -18726
rect 388238 -18782 388294 -18726
rect 388362 -18782 388418 -18726
rect 388486 -18782 388542 -18726
rect 388610 -18782 388666 -18726
rect 388114 -18906 388170 -18850
rect 388238 -18906 388294 -18850
rect 388362 -18906 388418 -18850
rect 388486 -18906 388542 -18850
rect 388610 -18906 388666 -18850
rect 388114 -19030 388170 -18974
rect 388238 -19030 388294 -18974
rect 388362 -19030 388418 -18974
rect 388486 -19030 388542 -18974
rect 388610 -19030 388666 -18974
rect 388114 -19154 388170 -19098
rect 388238 -19154 388294 -19098
rect 388362 -19154 388418 -19098
rect 388486 -19154 388542 -19098
rect 388610 -19154 388666 -19098
rect 388114 -19278 388170 -19222
rect 388238 -19278 388294 -19222
rect 388362 -19278 388418 -19222
rect 388486 -19278 388542 -19222
rect 388610 -19278 388666 -19222
rect 388114 -19402 388170 -19346
rect 388238 -19402 388294 -19346
rect 388362 -19402 388418 -19346
rect 388486 -19402 388542 -19346
rect 388610 -19402 388666 -19346
rect 388114 -19526 388170 -19470
rect 388238 -19526 388294 -19470
rect 388362 -19526 388418 -19470
rect 388486 -19526 388542 -19470
rect 388610 -19526 388666 -19470
rect 388114 -19650 388170 -19594
rect 388238 -19650 388294 -19594
rect 388362 -19650 388418 -19594
rect 388486 -19650 388542 -19594
rect 388610 -19650 388666 -19594
rect 388114 -19774 388170 -19718
rect 388238 -19774 388294 -19718
rect 388362 -19774 388418 -19718
rect 388486 -19774 388542 -19718
rect 388610 -19774 388666 -19718
rect 388114 -19898 388170 -19842
rect 388238 -19898 388294 -19842
rect 388362 -19898 388418 -19842
rect 388486 -19898 388542 -19842
rect 388610 -19898 388666 -19842
rect 388114 -20022 388170 -19966
rect 388238 -20022 388294 -19966
rect 388362 -20022 388418 -19966
rect 388486 -20022 388542 -19966
rect 388610 -20022 388666 -19966
rect 388114 -20146 388170 -20090
rect 388238 -20146 388294 -20090
rect 388362 -20146 388418 -20090
rect 388486 -20146 388542 -20090
rect 388610 -20146 388666 -20090
rect 388114 -20270 388170 -20214
rect 388238 -20270 388294 -20214
rect 388362 -20270 388418 -20214
rect 388486 -20270 388542 -20214
rect 388610 -20270 388666 -20214
rect 388114 -20394 388170 -20338
rect 388238 -20394 388294 -20338
rect 388362 -20394 388418 -20338
rect 388486 -20394 388542 -20338
rect 388610 -20394 388666 -20338
rect 388114 -20518 388170 -20462
rect 388238 -20518 388294 -20462
rect 388362 -20518 388418 -20462
rect 388486 -20518 388542 -20462
rect 388610 -20518 388666 -20462
rect 388114 -20642 388170 -20586
rect 388238 -20642 388294 -20586
rect 388362 -20642 388418 -20586
rect 388486 -20642 388542 -20586
rect 388610 -20642 388666 -20586
rect 388114 -20766 388170 -20710
rect 388238 -20766 388294 -20710
rect 388362 -20766 388418 -20710
rect 388486 -20766 388542 -20710
rect 388610 -20766 388666 -20710
rect 388114 -20890 388170 -20834
rect 388238 -20890 388294 -20834
rect 388362 -20890 388418 -20834
rect 388486 -20890 388542 -20834
rect 388610 -20890 388666 -20834
rect 388114 -21014 388170 -20958
rect 388238 -21014 388294 -20958
rect 388362 -21014 388418 -20958
rect 388486 -21014 388542 -20958
rect 388610 -21014 388666 -20958
rect 388114 -21138 388170 -21082
rect 388238 -21138 388294 -21082
rect 388362 -21138 388418 -21082
rect 388486 -21138 388542 -21082
rect 388610 -21138 388666 -21082
rect 388114 -21262 388170 -21206
rect 388238 -21262 388294 -21206
rect 388362 -21262 388418 -21206
rect 388486 -21262 388542 -21206
rect 388610 -21262 388666 -21206
rect 388114 -21386 388170 -21330
rect 388238 -21386 388294 -21330
rect 388362 -21386 388418 -21330
rect 388486 -21386 388542 -21330
rect 388610 -21386 388666 -21330
rect 388114 -21510 388170 -21454
rect 388238 -21510 388294 -21454
rect 388362 -21510 388418 -21454
rect 388486 -21510 388542 -21454
rect 388610 -21510 388666 -21454
rect 388114 -21634 388170 -21578
rect 388238 -21634 388294 -21578
rect 388362 -21634 388418 -21578
rect 388486 -21634 388542 -21578
rect 388610 -21634 388666 -21578
rect 388114 -21758 388170 -21702
rect 388238 -21758 388294 -21702
rect 388362 -21758 388418 -21702
rect 388486 -21758 388542 -21702
rect 388610 -21758 388666 -21702
rect 388114 -21882 388170 -21826
rect 388238 -21882 388294 -21826
rect 388362 -21882 388418 -21826
rect 388486 -21882 388542 -21826
rect 388610 -21882 388666 -21826
rect 388114 -22006 388170 -21950
rect 388238 -22006 388294 -21950
rect 388362 -22006 388418 -21950
rect 388486 -22006 388542 -21950
rect 388610 -22006 388666 -21950
rect 388114 -22130 388170 -22074
rect 388238 -22130 388294 -22074
rect 388362 -22130 388418 -22074
rect 388486 -22130 388542 -22074
rect 388610 -22130 388666 -22074
rect 388114 -22254 388170 -22198
rect 388238 -22254 388294 -22198
rect 388362 -22254 388418 -22198
rect 388486 -22254 388542 -22198
rect 388610 -22254 388666 -22198
rect 388114 -22378 388170 -22322
rect 388238 -22378 388294 -22322
rect 388362 -22378 388418 -22322
rect 388486 -22378 388542 -22322
rect 388610 -22378 388666 -22322
rect 388114 -22502 388170 -22446
rect 388238 -22502 388294 -22446
rect 388362 -22502 388418 -22446
rect 388486 -22502 388542 -22446
rect 388610 -22502 388666 -22446
rect 388114 -22626 388170 -22570
rect 388238 -22626 388294 -22570
rect 388362 -22626 388418 -22570
rect 388486 -22626 388542 -22570
rect 388610 -22626 388666 -22570
rect 388114 -22750 388170 -22694
rect 388238 -22750 388294 -22694
rect 388362 -22750 388418 -22694
rect 388486 -22750 388542 -22694
rect 388610 -22750 388666 -22694
rect 388114 -22874 388170 -22818
rect 388238 -22874 388294 -22818
rect 388362 -22874 388418 -22818
rect 388486 -22874 388542 -22818
rect 388610 -22874 388666 -22818
rect 388114 -22998 388170 -22942
rect 388238 -22998 388294 -22942
rect 388362 -22998 388418 -22942
rect 388486 -22998 388542 -22942
rect 388610 -22998 388666 -22942
rect 388114 -23122 388170 -23066
rect 388238 -23122 388294 -23066
rect 388362 -23122 388418 -23066
rect 388486 -23122 388542 -23066
rect 388610 -23122 388666 -23066
rect 388114 -23246 388170 -23190
rect 388238 -23246 388294 -23190
rect 388362 -23246 388418 -23190
rect 388486 -23246 388542 -23190
rect 388610 -23246 388666 -23190
rect 388114 -23370 388170 -23314
rect 388238 -23370 388294 -23314
rect 388362 -23370 388418 -23314
rect 388486 -23370 388542 -23314
rect 388610 -23370 388666 -23314
rect 388114 -23494 388170 -23438
rect 388238 -23494 388294 -23438
rect 388362 -23494 388418 -23438
rect 388486 -23494 388542 -23438
rect 388610 -23494 388666 -23438
rect 388114 -23618 388170 -23562
rect 388238 -23618 388294 -23562
rect 388362 -23618 388418 -23562
rect 388486 -23618 388542 -23562
rect 388610 -23618 388666 -23562
rect 388114 -23742 388170 -23686
rect 388238 -23742 388294 -23686
rect 388362 -23742 388418 -23686
rect 388486 -23742 388542 -23686
rect 388610 -23742 388666 -23686
rect 388114 -23866 388170 -23810
rect 388238 -23866 388294 -23810
rect 388362 -23866 388418 -23810
rect 388486 -23866 388542 -23810
rect 388610 -23866 388666 -23810
rect 388114 -23990 388170 -23934
rect 388238 -23990 388294 -23934
rect 388362 -23990 388418 -23934
rect 388486 -23990 388542 -23934
rect 388610 -23990 388666 -23934
rect 388114 -24114 388170 -24058
rect 388238 -24114 388294 -24058
rect 388362 -24114 388418 -24058
rect 388486 -24114 388542 -24058
rect 388610 -24114 388666 -24058
rect 388114 -24238 388170 -24182
rect 388238 -24238 388294 -24182
rect 388362 -24238 388418 -24182
rect 388486 -24238 388542 -24182
rect 388610 -24238 388666 -24182
rect 388114 -24362 388170 -24306
rect 388238 -24362 388294 -24306
rect 388362 -24362 388418 -24306
rect 388486 -24362 388542 -24306
rect 388610 -24362 388666 -24306
rect 388114 -24486 388170 -24430
rect 388238 -24486 388294 -24430
rect 388362 -24486 388418 -24430
rect 388486 -24486 388542 -24430
rect 388610 -24486 388666 -24430
rect 388114 -24610 388170 -24554
rect 388238 -24610 388294 -24554
rect 388362 -24610 388418 -24554
rect 388486 -24610 388542 -24554
rect 388610 -24610 388666 -24554
rect 388114 -24734 388170 -24678
rect 388238 -24734 388294 -24678
rect 388362 -24734 388418 -24678
rect 388486 -24734 388542 -24678
rect 388610 -24734 388666 -24678
rect 388114 -24858 388170 -24802
rect 388238 -24858 388294 -24802
rect 388362 -24858 388418 -24802
rect 388486 -24858 388542 -24802
rect 388610 -24858 388666 -24802
rect 388114 -24982 388170 -24926
rect 388238 -24982 388294 -24926
rect 388362 -24982 388418 -24926
rect 388486 -24982 388542 -24926
rect 388610 -24982 388666 -24926
rect 388114 -25106 388170 -25050
rect 388238 -25106 388294 -25050
rect 388362 -25106 388418 -25050
rect 388486 -25106 388542 -25050
rect 388610 -25106 388666 -25050
rect 388114 -25230 388170 -25174
rect 388238 -25230 388294 -25174
rect 388362 -25230 388418 -25174
rect 388486 -25230 388542 -25174
rect 388610 -25230 388666 -25174
rect 388114 -25354 388170 -25298
rect 388238 -25354 388294 -25298
rect 388362 -25354 388418 -25298
rect 388486 -25354 388542 -25298
rect 388610 -25354 388666 -25298
rect 388114 -25478 388170 -25422
rect 388238 -25478 388294 -25422
rect 388362 -25478 388418 -25422
rect 388486 -25478 388542 -25422
rect 388610 -25478 388666 -25422
rect 389141 -18006 389197 -17950
rect 389283 -18006 389339 -17950
rect 389141 -18148 389197 -18092
rect 389283 -18148 389339 -18092
rect 389141 -18290 389197 -18234
rect 389283 -18290 389339 -18234
rect 389141 -18432 389197 -18376
rect 389283 -18432 389339 -18376
rect 389141 -18574 389197 -18518
rect 389283 -18574 389339 -18518
rect 389141 -18716 389197 -18660
rect 389283 -18716 389339 -18660
rect 389141 -18858 389197 -18802
rect 389283 -18858 389339 -18802
rect 389141 -19000 389197 -18944
rect 389283 -19000 389339 -18944
rect 389141 -19142 389197 -19086
rect 389283 -19142 389339 -19086
rect 389141 -19284 389197 -19228
rect 389283 -19284 389339 -19228
rect 389141 -19426 389197 -19370
rect 389283 -19426 389339 -19370
rect 389141 -19568 389197 -19512
rect 389283 -19568 389339 -19512
rect 389141 -19710 389197 -19654
rect 389283 -19710 389339 -19654
rect 389141 -19852 389197 -19796
rect 389283 -19852 389339 -19796
rect 389141 -19994 389197 -19938
rect 389283 -19994 389339 -19938
rect 389141 -20136 389197 -20080
rect 389283 -20136 389339 -20080
rect 389141 -20278 389197 -20222
rect 389283 -20278 389339 -20222
rect 389141 -20420 389197 -20364
rect 389283 -20420 389339 -20364
rect 389141 -20562 389197 -20506
rect 389283 -20562 389339 -20506
rect 389141 -20704 389197 -20648
rect 389283 -20704 389339 -20648
rect 389141 -20846 389197 -20790
rect 389283 -20846 389339 -20790
rect 389141 -20988 389197 -20932
rect 389283 -20988 389339 -20932
rect 389141 -21130 389197 -21074
rect 389283 -21130 389339 -21074
rect 389141 -21272 389197 -21216
rect 389283 -21272 389339 -21216
rect 389141 -21414 389197 -21358
rect 389283 -21414 389339 -21358
rect 389141 -21556 389197 -21500
rect 389283 -21556 389339 -21500
rect 389141 -21698 389197 -21642
rect 389283 -21698 389339 -21642
rect 389141 -21840 389197 -21784
rect 389283 -21840 389339 -21784
rect 389141 -21982 389197 -21926
rect 389283 -21982 389339 -21926
rect 389141 -22124 389197 -22068
rect 389283 -22124 389339 -22068
rect 389141 -22266 389197 -22210
rect 389283 -22266 389339 -22210
rect 389141 -22408 389197 -22352
rect 389283 -22408 389339 -22352
rect 389141 -22550 389197 -22494
rect 389283 -22550 389339 -22494
rect 389141 -22692 389197 -22636
rect 389283 -22692 389339 -22636
rect 389141 -22834 389197 -22778
rect 389283 -22834 389339 -22778
rect 389141 -22976 389197 -22920
rect 389283 -22976 389339 -22920
rect 389141 -23118 389197 -23062
rect 389283 -23118 389339 -23062
rect 389141 -23260 389197 -23204
rect 389283 -23260 389339 -23204
rect 389141 -23402 389197 -23346
rect 389283 -23402 389339 -23346
rect 389141 -23544 389197 -23488
rect 389283 -23544 389339 -23488
rect 389141 -23686 389197 -23630
rect 389283 -23686 389339 -23630
rect 389141 -23828 389197 -23772
rect 389283 -23828 389339 -23772
rect 389141 -23970 389197 -23914
rect 389283 -23970 389339 -23914
rect 389141 -24112 389197 -24056
rect 389283 -24112 389339 -24056
rect 389141 -24254 389197 -24198
rect 389283 -24254 389339 -24198
rect 389141 -24396 389197 -24340
rect 389283 -24396 389339 -24340
rect 389141 -24538 389197 -24482
rect 389283 -24538 389339 -24482
rect 389141 -24680 389197 -24624
rect 389283 -24680 389339 -24624
rect 389141 -24822 389197 -24766
rect 389283 -24822 389339 -24766
rect 389141 -24964 389197 -24908
rect 389283 -24964 389339 -24908
rect 389141 -25106 389197 -25050
rect 389283 -25106 389339 -25050
rect 389141 -25248 389197 -25192
rect 389283 -25248 389339 -25192
rect 389141 -25390 389197 -25334
rect 389283 -25390 389339 -25334
rect 389141 -25532 389197 -25476
rect 389283 -25532 389339 -25476
rect 389542 -18006 389598 -17950
rect 389684 -18006 389740 -17950
rect 389542 -18148 389598 -18092
rect 389684 -18148 389740 -18092
rect 389542 -18290 389598 -18234
rect 389684 -18290 389740 -18234
rect 389542 -18432 389598 -18376
rect 389684 -18432 389740 -18376
rect 389542 -18574 389598 -18518
rect 389684 -18574 389740 -18518
rect 389542 -18716 389598 -18660
rect 389684 -18716 389740 -18660
rect 389542 -18858 389598 -18802
rect 389684 -18858 389740 -18802
rect 389542 -19000 389598 -18944
rect 389684 -19000 389740 -18944
rect 389542 -19142 389598 -19086
rect 389684 -19142 389740 -19086
rect 389542 -19284 389598 -19228
rect 389684 -19284 389740 -19228
rect 389542 -19426 389598 -19370
rect 389684 -19426 389740 -19370
rect 389542 -19568 389598 -19512
rect 389684 -19568 389740 -19512
rect 389542 -19710 389598 -19654
rect 389684 -19710 389740 -19654
rect 389542 -19852 389598 -19796
rect 389684 -19852 389740 -19796
rect 389542 -19994 389598 -19938
rect 389684 -19994 389740 -19938
rect 389542 -20136 389598 -20080
rect 389684 -20136 389740 -20080
rect 389542 -20278 389598 -20222
rect 389684 -20278 389740 -20222
rect 389542 -20420 389598 -20364
rect 389684 -20420 389740 -20364
rect 389542 -20562 389598 -20506
rect 389684 -20562 389740 -20506
rect 389542 -20704 389598 -20648
rect 389684 -20704 389740 -20648
rect 389542 -20846 389598 -20790
rect 389684 -20846 389740 -20790
rect 389542 -20988 389598 -20932
rect 389684 -20988 389740 -20932
rect 389542 -21130 389598 -21074
rect 389684 -21130 389740 -21074
rect 389542 -21272 389598 -21216
rect 389684 -21272 389740 -21216
rect 389542 -21414 389598 -21358
rect 389684 -21414 389740 -21358
rect 389542 -21556 389598 -21500
rect 389684 -21556 389740 -21500
rect 389542 -21698 389598 -21642
rect 389684 -21698 389740 -21642
rect 389542 -21840 389598 -21784
rect 389684 -21840 389740 -21784
rect 389542 -21982 389598 -21926
rect 389684 -21982 389740 -21926
rect 389542 -22124 389598 -22068
rect 389684 -22124 389740 -22068
rect 389542 -22266 389598 -22210
rect 389684 -22266 389740 -22210
rect 389542 -22408 389598 -22352
rect 389684 -22408 389740 -22352
rect 389542 -22550 389598 -22494
rect 389684 -22550 389740 -22494
rect 389542 -22692 389598 -22636
rect 389684 -22692 389740 -22636
rect 389542 -22834 389598 -22778
rect 389684 -22834 389740 -22778
rect 389542 -22976 389598 -22920
rect 389684 -22976 389740 -22920
rect 389542 -23118 389598 -23062
rect 389684 -23118 389740 -23062
rect 389542 -23260 389598 -23204
rect 389684 -23260 389740 -23204
rect 389542 -23402 389598 -23346
rect 389684 -23402 389740 -23346
rect 389542 -23544 389598 -23488
rect 389684 -23544 389740 -23488
rect 389542 -23686 389598 -23630
rect 389684 -23686 389740 -23630
rect 389542 -23828 389598 -23772
rect 389684 -23828 389740 -23772
rect 389542 -23970 389598 -23914
rect 389684 -23970 389740 -23914
rect 389542 -24112 389598 -24056
rect 389684 -24112 389740 -24056
rect 389542 -24254 389598 -24198
rect 389684 -24254 389740 -24198
rect 389542 -24396 389598 -24340
rect 389684 -24396 389740 -24340
rect 389542 -24538 389598 -24482
rect 389684 -24538 389740 -24482
rect 389542 -24680 389598 -24624
rect 389684 -24680 389740 -24624
rect 389542 -24822 389598 -24766
rect 389684 -24822 389740 -24766
rect 389542 -24964 389598 -24908
rect 389684 -24964 389740 -24908
rect 389542 -25106 389598 -25050
rect 389684 -25106 389740 -25050
rect 389542 -25248 389598 -25192
rect 389684 -25248 389740 -25192
rect 389542 -25390 389598 -25334
rect 389684 -25390 389740 -25334
rect 389542 -25532 389598 -25476
rect 389684 -25532 389740 -25476
rect 389942 -18006 389998 -17950
rect 390084 -18006 390140 -17950
rect 389942 -18148 389998 -18092
rect 390084 -18148 390140 -18092
rect 389942 -18290 389998 -18234
rect 390084 -18290 390140 -18234
rect 389942 -18432 389998 -18376
rect 390084 -18432 390140 -18376
rect 389942 -18574 389998 -18518
rect 390084 -18574 390140 -18518
rect 389942 -18716 389998 -18660
rect 390084 -18716 390140 -18660
rect 389942 -18858 389998 -18802
rect 390084 -18858 390140 -18802
rect 389942 -19000 389998 -18944
rect 390084 -19000 390140 -18944
rect 389942 -19142 389998 -19086
rect 390084 -19142 390140 -19086
rect 389942 -19284 389998 -19228
rect 390084 -19284 390140 -19228
rect 389942 -19426 389998 -19370
rect 390084 -19426 390140 -19370
rect 389942 -19568 389998 -19512
rect 390084 -19568 390140 -19512
rect 389942 -19710 389998 -19654
rect 390084 -19710 390140 -19654
rect 389942 -19852 389998 -19796
rect 390084 -19852 390140 -19796
rect 389942 -19994 389998 -19938
rect 390084 -19994 390140 -19938
rect 389942 -20136 389998 -20080
rect 390084 -20136 390140 -20080
rect 389942 -20278 389998 -20222
rect 390084 -20278 390140 -20222
rect 389942 -20420 389998 -20364
rect 390084 -20420 390140 -20364
rect 389942 -20562 389998 -20506
rect 390084 -20562 390140 -20506
rect 389942 -20704 389998 -20648
rect 390084 -20704 390140 -20648
rect 389942 -20846 389998 -20790
rect 390084 -20846 390140 -20790
rect 389942 -20988 389998 -20932
rect 390084 -20988 390140 -20932
rect 389942 -21130 389998 -21074
rect 390084 -21130 390140 -21074
rect 389942 -21272 389998 -21216
rect 390084 -21272 390140 -21216
rect 389942 -21414 389998 -21358
rect 390084 -21414 390140 -21358
rect 389942 -21556 389998 -21500
rect 390084 -21556 390140 -21500
rect 389942 -21698 389998 -21642
rect 390084 -21698 390140 -21642
rect 389942 -21840 389998 -21784
rect 390084 -21840 390140 -21784
rect 389942 -21982 389998 -21926
rect 390084 -21982 390140 -21926
rect 389942 -22124 389998 -22068
rect 390084 -22124 390140 -22068
rect 389942 -22266 389998 -22210
rect 390084 -22266 390140 -22210
rect 389942 -22408 389998 -22352
rect 390084 -22408 390140 -22352
rect 389942 -22550 389998 -22494
rect 390084 -22550 390140 -22494
rect 389942 -22692 389998 -22636
rect 390084 -22692 390140 -22636
rect 389942 -22834 389998 -22778
rect 390084 -22834 390140 -22778
rect 389942 -22976 389998 -22920
rect 390084 -22976 390140 -22920
rect 389942 -23118 389998 -23062
rect 390084 -23118 390140 -23062
rect 389942 -23260 389998 -23204
rect 390084 -23260 390140 -23204
rect 389942 -23402 389998 -23346
rect 390084 -23402 390140 -23346
rect 389942 -23544 389998 -23488
rect 390084 -23544 390140 -23488
rect 389942 -23686 389998 -23630
rect 390084 -23686 390140 -23630
rect 389942 -23828 389998 -23772
rect 390084 -23828 390140 -23772
rect 389942 -23970 389998 -23914
rect 390084 -23970 390140 -23914
rect 389942 -24112 389998 -24056
rect 390084 -24112 390140 -24056
rect 389942 -24254 389998 -24198
rect 390084 -24254 390140 -24198
rect 389942 -24396 389998 -24340
rect 390084 -24396 390140 -24340
rect 389942 -24538 389998 -24482
rect 390084 -24538 390140 -24482
rect 389942 -24680 389998 -24624
rect 390084 -24680 390140 -24624
rect 389942 -24822 389998 -24766
rect 390084 -24822 390140 -24766
rect 389942 -24964 389998 -24908
rect 390084 -24964 390140 -24908
rect 389942 -25106 389998 -25050
rect 390084 -25106 390140 -25050
rect 389942 -25248 389998 -25192
rect 390084 -25248 390140 -25192
rect 389942 -25390 389998 -25334
rect 390084 -25390 390140 -25334
rect 389942 -25532 389998 -25476
rect 390084 -25532 390140 -25476
rect 390339 -18006 390395 -17950
rect 390481 -18006 390537 -17950
rect 390339 -18148 390395 -18092
rect 390481 -18148 390537 -18092
rect 390339 -18290 390395 -18234
rect 390481 -18290 390537 -18234
rect 390339 -18432 390395 -18376
rect 390481 -18432 390537 -18376
rect 390339 -18574 390395 -18518
rect 390481 -18574 390537 -18518
rect 390339 -18716 390395 -18660
rect 390481 -18716 390537 -18660
rect 390339 -18858 390395 -18802
rect 390481 -18858 390537 -18802
rect 390339 -19000 390395 -18944
rect 390481 -19000 390537 -18944
rect 390339 -19142 390395 -19086
rect 390481 -19142 390537 -19086
rect 390339 -19284 390395 -19228
rect 390481 -19284 390537 -19228
rect 390339 -19426 390395 -19370
rect 390481 -19426 390537 -19370
rect 390339 -19568 390395 -19512
rect 390481 -19568 390537 -19512
rect 390339 -19710 390395 -19654
rect 390481 -19710 390537 -19654
rect 390339 -19852 390395 -19796
rect 390481 -19852 390537 -19796
rect 390339 -19994 390395 -19938
rect 390481 -19994 390537 -19938
rect 390339 -20136 390395 -20080
rect 390481 -20136 390537 -20080
rect 390339 -20278 390395 -20222
rect 390481 -20278 390537 -20222
rect 390339 -20420 390395 -20364
rect 390481 -20420 390537 -20364
rect 390339 -20562 390395 -20506
rect 390481 -20562 390537 -20506
rect 390339 -20704 390395 -20648
rect 390481 -20704 390537 -20648
rect 390339 -20846 390395 -20790
rect 390481 -20846 390537 -20790
rect 390339 -20988 390395 -20932
rect 390481 -20988 390537 -20932
rect 390339 -21130 390395 -21074
rect 390481 -21130 390537 -21074
rect 390339 -21272 390395 -21216
rect 390481 -21272 390537 -21216
rect 390339 -21414 390395 -21358
rect 390481 -21414 390537 -21358
rect 390339 -21556 390395 -21500
rect 390481 -21556 390537 -21500
rect 390339 -21698 390395 -21642
rect 390481 -21698 390537 -21642
rect 390339 -21840 390395 -21784
rect 390481 -21840 390537 -21784
rect 390339 -21982 390395 -21926
rect 390481 -21982 390537 -21926
rect 390339 -22124 390395 -22068
rect 390481 -22124 390537 -22068
rect 390339 -22266 390395 -22210
rect 390481 -22266 390537 -22210
rect 390339 -22408 390395 -22352
rect 390481 -22408 390537 -22352
rect 390339 -22550 390395 -22494
rect 390481 -22550 390537 -22494
rect 390339 -22692 390395 -22636
rect 390481 -22692 390537 -22636
rect 390339 -22834 390395 -22778
rect 390481 -22834 390537 -22778
rect 390339 -22976 390395 -22920
rect 390481 -22976 390537 -22920
rect 390339 -23118 390395 -23062
rect 390481 -23118 390537 -23062
rect 390339 -23260 390395 -23204
rect 390481 -23260 390537 -23204
rect 390339 -23402 390395 -23346
rect 390481 -23402 390537 -23346
rect 390339 -23544 390395 -23488
rect 390481 -23544 390537 -23488
rect 390339 -23686 390395 -23630
rect 390481 -23686 390537 -23630
rect 390339 -23828 390395 -23772
rect 390481 -23828 390537 -23772
rect 390339 -23970 390395 -23914
rect 390481 -23970 390537 -23914
rect 390339 -24112 390395 -24056
rect 390481 -24112 390537 -24056
rect 390339 -24254 390395 -24198
rect 390481 -24254 390537 -24198
rect 390339 -24396 390395 -24340
rect 390481 -24396 390537 -24340
rect 390339 -24538 390395 -24482
rect 390481 -24538 390537 -24482
rect 390339 -24680 390395 -24624
rect 390481 -24680 390537 -24624
rect 390339 -24822 390395 -24766
rect 390481 -24822 390537 -24766
rect 390339 -24964 390395 -24908
rect 390481 -24964 390537 -24908
rect 390339 -25106 390395 -25050
rect 390481 -25106 390537 -25050
rect 390339 -25248 390395 -25192
rect 390481 -25248 390537 -25192
rect 390339 -25390 390395 -25334
rect 390481 -25390 390537 -25334
rect 390339 -25532 390395 -25476
rect 390481 -25532 390537 -25476
rect 390736 -18006 390792 -17950
rect 390878 -18006 390934 -17950
rect 390736 -18148 390792 -18092
rect 390878 -18148 390934 -18092
rect 390736 -18290 390792 -18234
rect 390878 -18290 390934 -18234
rect 390736 -18432 390792 -18376
rect 390878 -18432 390934 -18376
rect 390736 -18574 390792 -18518
rect 390878 -18574 390934 -18518
rect 390736 -18716 390792 -18660
rect 390878 -18716 390934 -18660
rect 390736 -18858 390792 -18802
rect 390878 -18858 390934 -18802
rect 390736 -19000 390792 -18944
rect 390878 -19000 390934 -18944
rect 390736 -19142 390792 -19086
rect 390878 -19142 390934 -19086
rect 390736 -19284 390792 -19228
rect 390878 -19284 390934 -19228
rect 390736 -19426 390792 -19370
rect 390878 -19426 390934 -19370
rect 390736 -19568 390792 -19512
rect 390878 -19568 390934 -19512
rect 390736 -19710 390792 -19654
rect 390878 -19710 390934 -19654
rect 390736 -19852 390792 -19796
rect 390878 -19852 390934 -19796
rect 390736 -19994 390792 -19938
rect 390878 -19994 390934 -19938
rect 390736 -20136 390792 -20080
rect 390878 -20136 390934 -20080
rect 390736 -20278 390792 -20222
rect 390878 -20278 390934 -20222
rect 390736 -20420 390792 -20364
rect 390878 -20420 390934 -20364
rect 390736 -20562 390792 -20506
rect 390878 -20562 390934 -20506
rect 390736 -20704 390792 -20648
rect 390878 -20704 390934 -20648
rect 390736 -20846 390792 -20790
rect 390878 -20846 390934 -20790
rect 390736 -20988 390792 -20932
rect 390878 -20988 390934 -20932
rect 390736 -21130 390792 -21074
rect 390878 -21130 390934 -21074
rect 390736 -21272 390792 -21216
rect 390878 -21272 390934 -21216
rect 390736 -21414 390792 -21358
rect 390878 -21414 390934 -21358
rect 390736 -21556 390792 -21500
rect 390878 -21556 390934 -21500
rect 390736 -21698 390792 -21642
rect 390878 -21698 390934 -21642
rect 390736 -21840 390792 -21784
rect 390878 -21840 390934 -21784
rect 390736 -21982 390792 -21926
rect 390878 -21982 390934 -21926
rect 390736 -22124 390792 -22068
rect 390878 -22124 390934 -22068
rect 390736 -22266 390792 -22210
rect 390878 -22266 390934 -22210
rect 390736 -22408 390792 -22352
rect 390878 -22408 390934 -22352
rect 390736 -22550 390792 -22494
rect 390878 -22550 390934 -22494
rect 390736 -22692 390792 -22636
rect 390878 -22692 390934 -22636
rect 390736 -22834 390792 -22778
rect 390878 -22834 390934 -22778
rect 390736 -22976 390792 -22920
rect 390878 -22976 390934 -22920
rect 390736 -23118 390792 -23062
rect 390878 -23118 390934 -23062
rect 390736 -23260 390792 -23204
rect 390878 -23260 390934 -23204
rect 390736 -23402 390792 -23346
rect 390878 -23402 390934 -23346
rect 390736 -23544 390792 -23488
rect 390878 -23544 390934 -23488
rect 390736 -23686 390792 -23630
rect 390878 -23686 390934 -23630
rect 390736 -23828 390792 -23772
rect 390878 -23828 390934 -23772
rect 390736 -23970 390792 -23914
rect 390878 -23970 390934 -23914
rect 390736 -24112 390792 -24056
rect 390878 -24112 390934 -24056
rect 390736 -24254 390792 -24198
rect 390878 -24254 390934 -24198
rect 390736 -24396 390792 -24340
rect 390878 -24396 390934 -24340
rect 390736 -24538 390792 -24482
rect 390878 -24538 390934 -24482
rect 390736 -24680 390792 -24624
rect 390878 -24680 390934 -24624
rect 390736 -24822 390792 -24766
rect 390878 -24822 390934 -24766
rect 390736 -24964 390792 -24908
rect 390878 -24964 390934 -24908
rect 390736 -25106 390792 -25050
rect 390878 -25106 390934 -25050
rect 390736 -25248 390792 -25192
rect 390878 -25248 390934 -25192
rect 390736 -25390 390792 -25334
rect 390878 -25390 390934 -25334
rect 390736 -25532 390792 -25476
rect 390878 -25532 390934 -25476
rect 391140 -18006 391196 -17950
rect 391282 -18006 391338 -17950
rect 391140 -18148 391196 -18092
rect 391282 -18148 391338 -18092
rect 391140 -18290 391196 -18234
rect 391282 -18290 391338 -18234
rect 391140 -18432 391196 -18376
rect 391282 -18432 391338 -18376
rect 391140 -18574 391196 -18518
rect 391282 -18574 391338 -18518
rect 391140 -18716 391196 -18660
rect 391282 -18716 391338 -18660
rect 391140 -18858 391196 -18802
rect 391282 -18858 391338 -18802
rect 391140 -19000 391196 -18944
rect 391282 -19000 391338 -18944
rect 391140 -19142 391196 -19086
rect 391282 -19142 391338 -19086
rect 391140 -19284 391196 -19228
rect 391282 -19284 391338 -19228
rect 391140 -19426 391196 -19370
rect 391282 -19426 391338 -19370
rect 391140 -19568 391196 -19512
rect 391282 -19568 391338 -19512
rect 391140 -19710 391196 -19654
rect 391282 -19710 391338 -19654
rect 391140 -19852 391196 -19796
rect 391282 -19852 391338 -19796
rect 391140 -19994 391196 -19938
rect 391282 -19994 391338 -19938
rect 391140 -20136 391196 -20080
rect 391282 -20136 391338 -20080
rect 391140 -20278 391196 -20222
rect 391282 -20278 391338 -20222
rect 391140 -20420 391196 -20364
rect 391282 -20420 391338 -20364
rect 391140 -20562 391196 -20506
rect 391282 -20562 391338 -20506
rect 391140 -20704 391196 -20648
rect 391282 -20704 391338 -20648
rect 391140 -20846 391196 -20790
rect 391282 -20846 391338 -20790
rect 391140 -20988 391196 -20932
rect 391282 -20988 391338 -20932
rect 391140 -21130 391196 -21074
rect 391282 -21130 391338 -21074
rect 391140 -21272 391196 -21216
rect 391282 -21272 391338 -21216
rect 391140 -21414 391196 -21358
rect 391282 -21414 391338 -21358
rect 391140 -21556 391196 -21500
rect 391282 -21556 391338 -21500
rect 391140 -21698 391196 -21642
rect 391282 -21698 391338 -21642
rect 391140 -21840 391196 -21784
rect 391282 -21840 391338 -21784
rect 391140 -21982 391196 -21926
rect 391282 -21982 391338 -21926
rect 391140 -22124 391196 -22068
rect 391282 -22124 391338 -22068
rect 391140 -22266 391196 -22210
rect 391282 -22266 391338 -22210
rect 391140 -22408 391196 -22352
rect 391282 -22408 391338 -22352
rect 391140 -22550 391196 -22494
rect 391282 -22550 391338 -22494
rect 391140 -22692 391196 -22636
rect 391282 -22692 391338 -22636
rect 391140 -22834 391196 -22778
rect 391282 -22834 391338 -22778
rect 391140 -22976 391196 -22920
rect 391282 -22976 391338 -22920
rect 391140 -23118 391196 -23062
rect 391282 -23118 391338 -23062
rect 391140 -23260 391196 -23204
rect 391282 -23260 391338 -23204
rect 391140 -23402 391196 -23346
rect 391282 -23402 391338 -23346
rect 391140 -23544 391196 -23488
rect 391282 -23544 391338 -23488
rect 391140 -23686 391196 -23630
rect 391282 -23686 391338 -23630
rect 391140 -23828 391196 -23772
rect 391282 -23828 391338 -23772
rect 391140 -23970 391196 -23914
rect 391282 -23970 391338 -23914
rect 391140 -24112 391196 -24056
rect 391282 -24112 391338 -24056
rect 391140 -24254 391196 -24198
rect 391282 -24254 391338 -24198
rect 391140 -24396 391196 -24340
rect 391282 -24396 391338 -24340
rect 391140 -24538 391196 -24482
rect 391282 -24538 391338 -24482
rect 391140 -24680 391196 -24624
rect 391282 -24680 391338 -24624
rect 391140 -24822 391196 -24766
rect 391282 -24822 391338 -24766
rect 391140 -24964 391196 -24908
rect 391282 -24964 391338 -24908
rect 391140 -25106 391196 -25050
rect 391282 -25106 391338 -25050
rect 391140 -25248 391196 -25192
rect 391282 -25248 391338 -25192
rect 391140 -25390 391196 -25334
rect 391282 -25390 391338 -25334
rect 391140 -25532 391196 -25476
rect 391282 -25532 391338 -25476
rect 391536 -18006 391592 -17950
rect 391678 -18006 391734 -17950
rect 391536 -18148 391592 -18092
rect 391678 -18148 391734 -18092
rect 391536 -18290 391592 -18234
rect 391678 -18290 391734 -18234
rect 391536 -18432 391592 -18376
rect 391678 -18432 391734 -18376
rect 391536 -18574 391592 -18518
rect 391678 -18574 391734 -18518
rect 391536 -18716 391592 -18660
rect 391678 -18716 391734 -18660
rect 391536 -18858 391592 -18802
rect 391678 -18858 391734 -18802
rect 391536 -19000 391592 -18944
rect 391678 -19000 391734 -18944
rect 391536 -19142 391592 -19086
rect 391678 -19142 391734 -19086
rect 391536 -19284 391592 -19228
rect 391678 -19284 391734 -19228
rect 391536 -19426 391592 -19370
rect 391678 -19426 391734 -19370
rect 391536 -19568 391592 -19512
rect 391678 -19568 391734 -19512
rect 391536 -19710 391592 -19654
rect 391678 -19710 391734 -19654
rect 391536 -19852 391592 -19796
rect 391678 -19852 391734 -19796
rect 391536 -19994 391592 -19938
rect 391678 -19994 391734 -19938
rect 391536 -20136 391592 -20080
rect 391678 -20136 391734 -20080
rect 391536 -20278 391592 -20222
rect 391678 -20278 391734 -20222
rect 391536 -20420 391592 -20364
rect 391678 -20420 391734 -20364
rect 391536 -20562 391592 -20506
rect 391678 -20562 391734 -20506
rect 391536 -20704 391592 -20648
rect 391678 -20704 391734 -20648
rect 391536 -20846 391592 -20790
rect 391678 -20846 391734 -20790
rect 391536 -20988 391592 -20932
rect 391678 -20988 391734 -20932
rect 391536 -21130 391592 -21074
rect 391678 -21130 391734 -21074
rect 391536 -21272 391592 -21216
rect 391678 -21272 391734 -21216
rect 391536 -21414 391592 -21358
rect 391678 -21414 391734 -21358
rect 391536 -21556 391592 -21500
rect 391678 -21556 391734 -21500
rect 391536 -21698 391592 -21642
rect 391678 -21698 391734 -21642
rect 391536 -21840 391592 -21784
rect 391678 -21840 391734 -21784
rect 391536 -21982 391592 -21926
rect 391678 -21982 391734 -21926
rect 391536 -22124 391592 -22068
rect 391678 -22124 391734 -22068
rect 391536 -22266 391592 -22210
rect 391678 -22266 391734 -22210
rect 391536 -22408 391592 -22352
rect 391678 -22408 391734 -22352
rect 391536 -22550 391592 -22494
rect 391678 -22550 391734 -22494
rect 391536 -22692 391592 -22636
rect 391678 -22692 391734 -22636
rect 391536 -22834 391592 -22778
rect 391678 -22834 391734 -22778
rect 391536 -22976 391592 -22920
rect 391678 -22976 391734 -22920
rect 391536 -23118 391592 -23062
rect 391678 -23118 391734 -23062
rect 391536 -23260 391592 -23204
rect 391678 -23260 391734 -23204
rect 391536 -23402 391592 -23346
rect 391678 -23402 391734 -23346
rect 391536 -23544 391592 -23488
rect 391678 -23544 391734 -23488
rect 391536 -23686 391592 -23630
rect 391678 -23686 391734 -23630
rect 391536 -23828 391592 -23772
rect 391678 -23828 391734 -23772
rect 391536 -23970 391592 -23914
rect 391678 -23970 391734 -23914
rect 391536 -24112 391592 -24056
rect 391678 -24112 391734 -24056
rect 391536 -24254 391592 -24198
rect 391678 -24254 391734 -24198
rect 391536 -24396 391592 -24340
rect 391678 -24396 391734 -24340
rect 391536 -24538 391592 -24482
rect 391678 -24538 391734 -24482
rect 391536 -24680 391592 -24624
rect 391678 -24680 391734 -24624
rect 391536 -24822 391592 -24766
rect 391678 -24822 391734 -24766
rect 391536 -24964 391592 -24908
rect 391678 -24964 391734 -24908
rect 391536 -25106 391592 -25050
rect 391678 -25106 391734 -25050
rect 391536 -25248 391592 -25192
rect 391678 -25248 391734 -25192
rect 391536 -25390 391592 -25334
rect 391678 -25390 391734 -25334
rect 391536 -25532 391592 -25476
rect 391678 -25532 391734 -25476
rect 391936 -18006 391992 -17950
rect 392078 -18006 392134 -17950
rect 391936 -18148 391992 -18092
rect 392078 -18148 392134 -18092
rect 391936 -18290 391992 -18234
rect 392078 -18290 392134 -18234
rect 391936 -18432 391992 -18376
rect 392078 -18432 392134 -18376
rect 391936 -18574 391992 -18518
rect 392078 -18574 392134 -18518
rect 391936 -18716 391992 -18660
rect 392078 -18716 392134 -18660
rect 391936 -18858 391992 -18802
rect 392078 -18858 392134 -18802
rect 391936 -19000 391992 -18944
rect 392078 -19000 392134 -18944
rect 391936 -19142 391992 -19086
rect 392078 -19142 392134 -19086
rect 391936 -19284 391992 -19228
rect 392078 -19284 392134 -19228
rect 391936 -19426 391992 -19370
rect 392078 -19426 392134 -19370
rect 391936 -19568 391992 -19512
rect 392078 -19568 392134 -19512
rect 391936 -19710 391992 -19654
rect 392078 -19710 392134 -19654
rect 391936 -19852 391992 -19796
rect 392078 -19852 392134 -19796
rect 391936 -19994 391992 -19938
rect 392078 -19994 392134 -19938
rect 391936 -20136 391992 -20080
rect 392078 -20136 392134 -20080
rect 391936 -20278 391992 -20222
rect 392078 -20278 392134 -20222
rect 391936 -20420 391992 -20364
rect 392078 -20420 392134 -20364
rect 391936 -20562 391992 -20506
rect 392078 -20562 392134 -20506
rect 391936 -20704 391992 -20648
rect 392078 -20704 392134 -20648
rect 391936 -20846 391992 -20790
rect 392078 -20846 392134 -20790
rect 391936 -20988 391992 -20932
rect 392078 -20988 392134 -20932
rect 391936 -21130 391992 -21074
rect 392078 -21130 392134 -21074
rect 391936 -21272 391992 -21216
rect 392078 -21272 392134 -21216
rect 391936 -21414 391992 -21358
rect 392078 -21414 392134 -21358
rect 391936 -21556 391992 -21500
rect 392078 -21556 392134 -21500
rect 391936 -21698 391992 -21642
rect 392078 -21698 392134 -21642
rect 391936 -21840 391992 -21784
rect 392078 -21840 392134 -21784
rect 391936 -21982 391992 -21926
rect 392078 -21982 392134 -21926
rect 391936 -22124 391992 -22068
rect 392078 -22124 392134 -22068
rect 391936 -22266 391992 -22210
rect 392078 -22266 392134 -22210
rect 391936 -22408 391992 -22352
rect 392078 -22408 392134 -22352
rect 391936 -22550 391992 -22494
rect 392078 -22550 392134 -22494
rect 391936 -22692 391992 -22636
rect 392078 -22692 392134 -22636
rect 391936 -22834 391992 -22778
rect 392078 -22834 392134 -22778
rect 391936 -22976 391992 -22920
rect 392078 -22976 392134 -22920
rect 391936 -23118 391992 -23062
rect 392078 -23118 392134 -23062
rect 391936 -23260 391992 -23204
rect 392078 -23260 392134 -23204
rect 391936 -23402 391992 -23346
rect 392078 -23402 392134 -23346
rect 391936 -23544 391992 -23488
rect 392078 -23544 392134 -23488
rect 391936 -23686 391992 -23630
rect 392078 -23686 392134 -23630
rect 391936 -23828 391992 -23772
rect 392078 -23828 392134 -23772
rect 391936 -23970 391992 -23914
rect 392078 -23970 392134 -23914
rect 391936 -24112 391992 -24056
rect 392078 -24112 392134 -24056
rect 391936 -24254 391992 -24198
rect 392078 -24254 392134 -24198
rect 391936 -24396 391992 -24340
rect 392078 -24396 392134 -24340
rect 391936 -24538 391992 -24482
rect 392078 -24538 392134 -24482
rect 391936 -24680 391992 -24624
rect 392078 -24680 392134 -24624
rect 391936 -24822 391992 -24766
rect 392078 -24822 392134 -24766
rect 391936 -24964 391992 -24908
rect 392078 -24964 392134 -24908
rect 391936 -25106 391992 -25050
rect 392078 -25106 392134 -25050
rect 391936 -25248 391992 -25192
rect 392078 -25248 392134 -25192
rect 391936 -25390 391992 -25334
rect 392078 -25390 392134 -25334
rect 391936 -25532 391992 -25476
rect 392078 -25532 392134 -25476
rect 392333 -18006 392389 -17950
rect 392475 -18006 392531 -17950
rect 392333 -18148 392389 -18092
rect 392475 -18148 392531 -18092
rect 392333 -18290 392389 -18234
rect 392475 -18290 392531 -18234
rect 392333 -18432 392389 -18376
rect 392475 -18432 392531 -18376
rect 392333 -18574 392389 -18518
rect 392475 -18574 392531 -18518
rect 392333 -18716 392389 -18660
rect 392475 -18716 392531 -18660
rect 392333 -18858 392389 -18802
rect 392475 -18858 392531 -18802
rect 392333 -19000 392389 -18944
rect 392475 -19000 392531 -18944
rect 392333 -19142 392389 -19086
rect 392475 -19142 392531 -19086
rect 392333 -19284 392389 -19228
rect 392475 -19284 392531 -19228
rect 392333 -19426 392389 -19370
rect 392475 -19426 392531 -19370
rect 392333 -19568 392389 -19512
rect 392475 -19568 392531 -19512
rect 392333 -19710 392389 -19654
rect 392475 -19710 392531 -19654
rect 392333 -19852 392389 -19796
rect 392475 -19852 392531 -19796
rect 392333 -19994 392389 -19938
rect 392475 -19994 392531 -19938
rect 392333 -20136 392389 -20080
rect 392475 -20136 392531 -20080
rect 392333 -20278 392389 -20222
rect 392475 -20278 392531 -20222
rect 392333 -20420 392389 -20364
rect 392475 -20420 392531 -20364
rect 392333 -20562 392389 -20506
rect 392475 -20562 392531 -20506
rect 392333 -20704 392389 -20648
rect 392475 -20704 392531 -20648
rect 392333 -20846 392389 -20790
rect 392475 -20846 392531 -20790
rect 392333 -20988 392389 -20932
rect 392475 -20988 392531 -20932
rect 392333 -21130 392389 -21074
rect 392475 -21130 392531 -21074
rect 392333 -21272 392389 -21216
rect 392475 -21272 392531 -21216
rect 392333 -21414 392389 -21358
rect 392475 -21414 392531 -21358
rect 392333 -21556 392389 -21500
rect 392475 -21556 392531 -21500
rect 392333 -21698 392389 -21642
rect 392475 -21698 392531 -21642
rect 392333 -21840 392389 -21784
rect 392475 -21840 392531 -21784
rect 392333 -21982 392389 -21926
rect 392475 -21982 392531 -21926
rect 392333 -22124 392389 -22068
rect 392475 -22124 392531 -22068
rect 392333 -22266 392389 -22210
rect 392475 -22266 392531 -22210
rect 392333 -22408 392389 -22352
rect 392475 -22408 392531 -22352
rect 392333 -22550 392389 -22494
rect 392475 -22550 392531 -22494
rect 392333 -22692 392389 -22636
rect 392475 -22692 392531 -22636
rect 392333 -22834 392389 -22778
rect 392475 -22834 392531 -22778
rect 392333 -22976 392389 -22920
rect 392475 -22976 392531 -22920
rect 392333 -23118 392389 -23062
rect 392475 -23118 392531 -23062
rect 392333 -23260 392389 -23204
rect 392475 -23260 392531 -23204
rect 392333 -23402 392389 -23346
rect 392475 -23402 392531 -23346
rect 392333 -23544 392389 -23488
rect 392475 -23544 392531 -23488
rect 392333 -23686 392389 -23630
rect 392475 -23686 392531 -23630
rect 392333 -23828 392389 -23772
rect 392475 -23828 392531 -23772
rect 392333 -23970 392389 -23914
rect 392475 -23970 392531 -23914
rect 392333 -24112 392389 -24056
rect 392475 -24112 392531 -24056
rect 392333 -24254 392389 -24198
rect 392475 -24254 392531 -24198
rect 392333 -24396 392389 -24340
rect 392475 -24396 392531 -24340
rect 392333 -24538 392389 -24482
rect 392475 -24538 392531 -24482
rect 392333 -24680 392389 -24624
rect 392475 -24680 392531 -24624
rect 392333 -24822 392389 -24766
rect 392475 -24822 392531 -24766
rect 392333 -24964 392389 -24908
rect 392475 -24964 392531 -24908
rect 392333 -25106 392389 -25050
rect 392475 -25106 392531 -25050
rect 392333 -25248 392389 -25192
rect 392475 -25248 392531 -25192
rect 392333 -25390 392389 -25334
rect 392475 -25390 392531 -25334
rect 392333 -25532 392389 -25476
rect 392475 -25532 392531 -25476
rect 392738 -18006 392794 -17950
rect 392880 -18006 392936 -17950
rect 392738 -18148 392794 -18092
rect 392880 -18148 392936 -18092
rect 392738 -18290 392794 -18234
rect 392880 -18290 392936 -18234
rect 392738 -18432 392794 -18376
rect 392880 -18432 392936 -18376
rect 392738 -18574 392794 -18518
rect 392880 -18574 392936 -18518
rect 392738 -18716 392794 -18660
rect 392880 -18716 392936 -18660
rect 392738 -18858 392794 -18802
rect 392880 -18858 392936 -18802
rect 392738 -19000 392794 -18944
rect 392880 -19000 392936 -18944
rect 392738 -19142 392794 -19086
rect 392880 -19142 392936 -19086
rect 392738 -19284 392794 -19228
rect 392880 -19284 392936 -19228
rect 392738 -19426 392794 -19370
rect 392880 -19426 392936 -19370
rect 392738 -19568 392794 -19512
rect 392880 -19568 392936 -19512
rect 392738 -19710 392794 -19654
rect 392880 -19710 392936 -19654
rect 392738 -19852 392794 -19796
rect 392880 -19852 392936 -19796
rect 392738 -19994 392794 -19938
rect 392880 -19994 392936 -19938
rect 392738 -20136 392794 -20080
rect 392880 -20136 392936 -20080
rect 392738 -20278 392794 -20222
rect 392880 -20278 392936 -20222
rect 392738 -20420 392794 -20364
rect 392880 -20420 392936 -20364
rect 392738 -20562 392794 -20506
rect 392880 -20562 392936 -20506
rect 392738 -20704 392794 -20648
rect 392880 -20704 392936 -20648
rect 392738 -20846 392794 -20790
rect 392880 -20846 392936 -20790
rect 392738 -20988 392794 -20932
rect 392880 -20988 392936 -20932
rect 392738 -21130 392794 -21074
rect 392880 -21130 392936 -21074
rect 392738 -21272 392794 -21216
rect 392880 -21272 392936 -21216
rect 392738 -21414 392794 -21358
rect 392880 -21414 392936 -21358
rect 392738 -21556 392794 -21500
rect 392880 -21556 392936 -21500
rect 392738 -21698 392794 -21642
rect 392880 -21698 392936 -21642
rect 392738 -21840 392794 -21784
rect 392880 -21840 392936 -21784
rect 392738 -21982 392794 -21926
rect 392880 -21982 392936 -21926
rect 392738 -22124 392794 -22068
rect 392880 -22124 392936 -22068
rect 392738 -22266 392794 -22210
rect 392880 -22266 392936 -22210
rect 392738 -22408 392794 -22352
rect 392880 -22408 392936 -22352
rect 392738 -22550 392794 -22494
rect 392880 -22550 392936 -22494
rect 392738 -22692 392794 -22636
rect 392880 -22692 392936 -22636
rect 392738 -22834 392794 -22778
rect 392880 -22834 392936 -22778
rect 392738 -22976 392794 -22920
rect 392880 -22976 392936 -22920
rect 392738 -23118 392794 -23062
rect 392880 -23118 392936 -23062
rect 392738 -23260 392794 -23204
rect 392880 -23260 392936 -23204
rect 392738 -23402 392794 -23346
rect 392880 -23402 392936 -23346
rect 392738 -23544 392794 -23488
rect 392880 -23544 392936 -23488
rect 392738 -23686 392794 -23630
rect 392880 -23686 392936 -23630
rect 392738 -23828 392794 -23772
rect 392880 -23828 392936 -23772
rect 392738 -23970 392794 -23914
rect 392880 -23970 392936 -23914
rect 392738 -24112 392794 -24056
rect 392880 -24112 392936 -24056
rect 392738 -24254 392794 -24198
rect 392880 -24254 392936 -24198
rect 392738 -24396 392794 -24340
rect 392880 -24396 392936 -24340
rect 392738 -24538 392794 -24482
rect 392880 -24538 392936 -24482
rect 392738 -24680 392794 -24624
rect 392880 -24680 392936 -24624
rect 392738 -24822 392794 -24766
rect 392880 -24822 392936 -24766
rect 392738 -24964 392794 -24908
rect 392880 -24964 392936 -24908
rect 392738 -25106 392794 -25050
rect 392880 -25106 392936 -25050
rect 392738 -25248 392794 -25192
rect 392880 -25248 392936 -25192
rect 392738 -25390 392794 -25334
rect 392880 -25390 392936 -25334
rect 392738 -25532 392794 -25476
rect 392880 -25532 392936 -25476
rect 393138 -18006 393194 -17950
rect 393280 -18006 393336 -17950
rect 393138 -18148 393194 -18092
rect 393280 -18148 393336 -18092
rect 393138 -18290 393194 -18234
rect 393280 -18290 393336 -18234
rect 393138 -18432 393194 -18376
rect 393280 -18432 393336 -18376
rect 393138 -18574 393194 -18518
rect 393280 -18574 393336 -18518
rect 393138 -18716 393194 -18660
rect 393280 -18716 393336 -18660
rect 393138 -18858 393194 -18802
rect 393280 -18858 393336 -18802
rect 393138 -19000 393194 -18944
rect 393280 -19000 393336 -18944
rect 393138 -19142 393194 -19086
rect 393280 -19142 393336 -19086
rect 393138 -19284 393194 -19228
rect 393280 -19284 393336 -19228
rect 393138 -19426 393194 -19370
rect 393280 -19426 393336 -19370
rect 393138 -19568 393194 -19512
rect 393280 -19568 393336 -19512
rect 393138 -19710 393194 -19654
rect 393280 -19710 393336 -19654
rect 393138 -19852 393194 -19796
rect 393280 -19852 393336 -19796
rect 393138 -19994 393194 -19938
rect 393280 -19994 393336 -19938
rect 393138 -20136 393194 -20080
rect 393280 -20136 393336 -20080
rect 393138 -20278 393194 -20222
rect 393280 -20278 393336 -20222
rect 393138 -20420 393194 -20364
rect 393280 -20420 393336 -20364
rect 393138 -20562 393194 -20506
rect 393280 -20562 393336 -20506
rect 393138 -20704 393194 -20648
rect 393280 -20704 393336 -20648
rect 393138 -20846 393194 -20790
rect 393280 -20846 393336 -20790
rect 393138 -20988 393194 -20932
rect 393280 -20988 393336 -20932
rect 393138 -21130 393194 -21074
rect 393280 -21130 393336 -21074
rect 393138 -21272 393194 -21216
rect 393280 -21272 393336 -21216
rect 393138 -21414 393194 -21358
rect 393280 -21414 393336 -21358
rect 393138 -21556 393194 -21500
rect 393280 -21556 393336 -21500
rect 393138 -21698 393194 -21642
rect 393280 -21698 393336 -21642
rect 393138 -21840 393194 -21784
rect 393280 -21840 393336 -21784
rect 393138 -21982 393194 -21926
rect 393280 -21982 393336 -21926
rect 393138 -22124 393194 -22068
rect 393280 -22124 393336 -22068
rect 393138 -22266 393194 -22210
rect 393280 -22266 393336 -22210
rect 393138 -22408 393194 -22352
rect 393280 -22408 393336 -22352
rect 393138 -22550 393194 -22494
rect 393280 -22550 393336 -22494
rect 393138 -22692 393194 -22636
rect 393280 -22692 393336 -22636
rect 393138 -22834 393194 -22778
rect 393280 -22834 393336 -22778
rect 393138 -22976 393194 -22920
rect 393280 -22976 393336 -22920
rect 393138 -23118 393194 -23062
rect 393280 -23118 393336 -23062
rect 393138 -23260 393194 -23204
rect 393280 -23260 393336 -23204
rect 393138 -23402 393194 -23346
rect 393280 -23402 393336 -23346
rect 393138 -23544 393194 -23488
rect 393280 -23544 393336 -23488
rect 393138 -23686 393194 -23630
rect 393280 -23686 393336 -23630
rect 393138 -23828 393194 -23772
rect 393280 -23828 393336 -23772
rect 393138 -23970 393194 -23914
rect 393280 -23970 393336 -23914
rect 393138 -24112 393194 -24056
rect 393280 -24112 393336 -24056
rect 393138 -24254 393194 -24198
rect 393280 -24254 393336 -24198
rect 393138 -24396 393194 -24340
rect 393280 -24396 393336 -24340
rect 393138 -24538 393194 -24482
rect 393280 -24538 393336 -24482
rect 393138 -24680 393194 -24624
rect 393280 -24680 393336 -24624
rect 393138 -24822 393194 -24766
rect 393280 -24822 393336 -24766
rect 393138 -24964 393194 -24908
rect 393280 -24964 393336 -24908
rect 393138 -25106 393194 -25050
rect 393280 -25106 393336 -25050
rect 393138 -25248 393194 -25192
rect 393280 -25248 393336 -25192
rect 393138 -25390 393194 -25334
rect 393280 -25390 393336 -25334
rect 393138 -25532 393194 -25476
rect 393280 -25532 393336 -25476
rect 393543 -18006 393599 -17950
rect 393685 -18006 393741 -17950
rect 393543 -18148 393599 -18092
rect 393685 -18148 393741 -18092
rect 393543 -18290 393599 -18234
rect 393685 -18290 393741 -18234
rect 393543 -18432 393599 -18376
rect 393685 -18432 393741 -18376
rect 393543 -18574 393599 -18518
rect 393685 -18574 393741 -18518
rect 393543 -18716 393599 -18660
rect 393685 -18716 393741 -18660
rect 393543 -18858 393599 -18802
rect 393685 -18858 393741 -18802
rect 393543 -19000 393599 -18944
rect 393685 -19000 393741 -18944
rect 393543 -19142 393599 -19086
rect 393685 -19142 393741 -19086
rect 393543 -19284 393599 -19228
rect 393685 -19284 393741 -19228
rect 393543 -19426 393599 -19370
rect 393685 -19426 393741 -19370
rect 393543 -19568 393599 -19512
rect 393685 -19568 393741 -19512
rect 393543 -19710 393599 -19654
rect 393685 -19710 393741 -19654
rect 393543 -19852 393599 -19796
rect 393685 -19852 393741 -19796
rect 393543 -19994 393599 -19938
rect 393685 -19994 393741 -19938
rect 393543 -20136 393599 -20080
rect 393685 -20136 393741 -20080
rect 393543 -20278 393599 -20222
rect 393685 -20278 393741 -20222
rect 393543 -20420 393599 -20364
rect 393685 -20420 393741 -20364
rect 393543 -20562 393599 -20506
rect 393685 -20562 393741 -20506
rect 393543 -20704 393599 -20648
rect 393685 -20704 393741 -20648
rect 393543 -20846 393599 -20790
rect 393685 -20846 393741 -20790
rect 393543 -20988 393599 -20932
rect 393685 -20988 393741 -20932
rect 393543 -21130 393599 -21074
rect 393685 -21130 393741 -21074
rect 393543 -21272 393599 -21216
rect 393685 -21272 393741 -21216
rect 393543 -21414 393599 -21358
rect 393685 -21414 393741 -21358
rect 393543 -21556 393599 -21500
rect 393685 -21556 393741 -21500
rect 393543 -21698 393599 -21642
rect 393685 -21698 393741 -21642
rect 393543 -21840 393599 -21784
rect 393685 -21840 393741 -21784
rect 393543 -21982 393599 -21926
rect 393685 -21982 393741 -21926
rect 393543 -22124 393599 -22068
rect 393685 -22124 393741 -22068
rect 393543 -22266 393599 -22210
rect 393685 -22266 393741 -22210
rect 393543 -22408 393599 -22352
rect 393685 -22408 393741 -22352
rect 393543 -22550 393599 -22494
rect 393685 -22550 393741 -22494
rect 393543 -22692 393599 -22636
rect 393685 -22692 393741 -22636
rect 393543 -22834 393599 -22778
rect 393685 -22834 393741 -22778
rect 393543 -22976 393599 -22920
rect 393685 -22976 393741 -22920
rect 393543 -23118 393599 -23062
rect 393685 -23118 393741 -23062
rect 393543 -23260 393599 -23204
rect 393685 -23260 393741 -23204
rect 393543 -23402 393599 -23346
rect 393685 -23402 393741 -23346
rect 393543 -23544 393599 -23488
rect 393685 -23544 393741 -23488
rect 393543 -23686 393599 -23630
rect 393685 -23686 393741 -23630
rect 393543 -23828 393599 -23772
rect 393685 -23828 393741 -23772
rect 393543 -23970 393599 -23914
rect 393685 -23970 393741 -23914
rect 393543 -24112 393599 -24056
rect 393685 -24112 393741 -24056
rect 393543 -24254 393599 -24198
rect 393685 -24254 393741 -24198
rect 393543 -24396 393599 -24340
rect 393685 -24396 393741 -24340
rect 393543 -24538 393599 -24482
rect 393685 -24538 393741 -24482
rect 393543 -24680 393599 -24624
rect 393685 -24680 393741 -24624
rect 393543 -24822 393599 -24766
rect 393685 -24822 393741 -24766
rect 393543 -24964 393599 -24908
rect 393685 -24964 393741 -24908
rect 393543 -25106 393599 -25050
rect 393685 -25106 393741 -25050
rect 393543 -25248 393599 -25192
rect 393685 -25248 393741 -25192
rect 393543 -25390 393599 -25334
rect 393685 -25390 393741 -25334
rect 393543 -25532 393599 -25476
rect 393685 -25532 393741 -25476
rect 393940 -18006 393996 -17950
rect 394082 -18006 394138 -17950
rect 393940 -18148 393996 -18092
rect 394082 -18148 394138 -18092
rect 393940 -18290 393996 -18234
rect 394082 -18290 394138 -18234
rect 393940 -18432 393996 -18376
rect 394082 -18432 394138 -18376
rect 393940 -18574 393996 -18518
rect 394082 -18574 394138 -18518
rect 393940 -18716 393996 -18660
rect 394082 -18716 394138 -18660
rect 393940 -18858 393996 -18802
rect 394082 -18858 394138 -18802
rect 393940 -19000 393996 -18944
rect 394082 -19000 394138 -18944
rect 393940 -19142 393996 -19086
rect 394082 -19142 394138 -19086
rect 393940 -19284 393996 -19228
rect 394082 -19284 394138 -19228
rect 393940 -19426 393996 -19370
rect 394082 -19426 394138 -19370
rect 393940 -19568 393996 -19512
rect 394082 -19568 394138 -19512
rect 393940 -19710 393996 -19654
rect 394082 -19710 394138 -19654
rect 393940 -19852 393996 -19796
rect 394082 -19852 394138 -19796
rect 393940 -19994 393996 -19938
rect 394082 -19994 394138 -19938
rect 393940 -20136 393996 -20080
rect 394082 -20136 394138 -20080
rect 393940 -20278 393996 -20222
rect 394082 -20278 394138 -20222
rect 393940 -20420 393996 -20364
rect 394082 -20420 394138 -20364
rect 393940 -20562 393996 -20506
rect 394082 -20562 394138 -20506
rect 393940 -20704 393996 -20648
rect 394082 -20704 394138 -20648
rect 393940 -20846 393996 -20790
rect 394082 -20846 394138 -20790
rect 393940 -20988 393996 -20932
rect 394082 -20988 394138 -20932
rect 393940 -21130 393996 -21074
rect 394082 -21130 394138 -21074
rect 393940 -21272 393996 -21216
rect 394082 -21272 394138 -21216
rect 393940 -21414 393996 -21358
rect 394082 -21414 394138 -21358
rect 393940 -21556 393996 -21500
rect 394082 -21556 394138 -21500
rect 393940 -21698 393996 -21642
rect 394082 -21698 394138 -21642
rect 393940 -21840 393996 -21784
rect 394082 -21840 394138 -21784
rect 393940 -21982 393996 -21926
rect 394082 -21982 394138 -21926
rect 393940 -22124 393996 -22068
rect 394082 -22124 394138 -22068
rect 393940 -22266 393996 -22210
rect 394082 -22266 394138 -22210
rect 393940 -22408 393996 -22352
rect 394082 -22408 394138 -22352
rect 393940 -22550 393996 -22494
rect 394082 -22550 394138 -22494
rect 393940 -22692 393996 -22636
rect 394082 -22692 394138 -22636
rect 393940 -22834 393996 -22778
rect 394082 -22834 394138 -22778
rect 393940 -22976 393996 -22920
rect 394082 -22976 394138 -22920
rect 393940 -23118 393996 -23062
rect 394082 -23118 394138 -23062
rect 393940 -23260 393996 -23204
rect 394082 -23260 394138 -23204
rect 393940 -23402 393996 -23346
rect 394082 -23402 394138 -23346
rect 393940 -23544 393996 -23488
rect 394082 -23544 394138 -23488
rect 393940 -23686 393996 -23630
rect 394082 -23686 394138 -23630
rect 393940 -23828 393996 -23772
rect 394082 -23828 394138 -23772
rect 393940 -23970 393996 -23914
rect 394082 -23970 394138 -23914
rect 393940 -24112 393996 -24056
rect 394082 -24112 394138 -24056
rect 393940 -24254 393996 -24198
rect 394082 -24254 394138 -24198
rect 393940 -24396 393996 -24340
rect 394082 -24396 394138 -24340
rect 393940 -24538 393996 -24482
rect 394082 -24538 394138 -24482
rect 393940 -24680 393996 -24624
rect 394082 -24680 394138 -24624
rect 393940 -24822 393996 -24766
rect 394082 -24822 394138 -24766
rect 393940 -24964 393996 -24908
rect 394082 -24964 394138 -24908
rect 393940 -25106 393996 -25050
rect 394082 -25106 394138 -25050
rect 393940 -25248 393996 -25192
rect 394082 -25248 394138 -25192
rect 393940 -25390 393996 -25334
rect 394082 -25390 394138 -25334
rect 393940 -25532 393996 -25476
rect 394082 -25532 394138 -25476
rect 394337 -18006 394393 -17950
rect 394479 -18006 394535 -17950
rect 394337 -18148 394393 -18092
rect 394479 -18148 394535 -18092
rect 394337 -18290 394393 -18234
rect 394479 -18290 394535 -18234
rect 394337 -18432 394393 -18376
rect 394479 -18432 394535 -18376
rect 394337 -18574 394393 -18518
rect 394479 -18574 394535 -18518
rect 394337 -18716 394393 -18660
rect 394479 -18716 394535 -18660
rect 394337 -18858 394393 -18802
rect 394479 -18858 394535 -18802
rect 394337 -19000 394393 -18944
rect 394479 -19000 394535 -18944
rect 394337 -19142 394393 -19086
rect 394479 -19142 394535 -19086
rect 394337 -19284 394393 -19228
rect 394479 -19284 394535 -19228
rect 394337 -19426 394393 -19370
rect 394479 -19426 394535 -19370
rect 394337 -19568 394393 -19512
rect 394479 -19568 394535 -19512
rect 394337 -19710 394393 -19654
rect 394479 -19710 394535 -19654
rect 394337 -19852 394393 -19796
rect 394479 -19852 394535 -19796
rect 394337 -19994 394393 -19938
rect 394479 -19994 394535 -19938
rect 394337 -20136 394393 -20080
rect 394479 -20136 394535 -20080
rect 394337 -20278 394393 -20222
rect 394479 -20278 394535 -20222
rect 394337 -20420 394393 -20364
rect 394479 -20420 394535 -20364
rect 394337 -20562 394393 -20506
rect 394479 -20562 394535 -20506
rect 394337 -20704 394393 -20648
rect 394479 -20704 394535 -20648
rect 394337 -20846 394393 -20790
rect 394479 -20846 394535 -20790
rect 394337 -20988 394393 -20932
rect 394479 -20988 394535 -20932
rect 394337 -21130 394393 -21074
rect 394479 -21130 394535 -21074
rect 394337 -21272 394393 -21216
rect 394479 -21272 394535 -21216
rect 394337 -21414 394393 -21358
rect 394479 -21414 394535 -21358
rect 394337 -21556 394393 -21500
rect 394479 -21556 394535 -21500
rect 394337 -21698 394393 -21642
rect 394479 -21698 394535 -21642
rect 394337 -21840 394393 -21784
rect 394479 -21840 394535 -21784
rect 394337 -21982 394393 -21926
rect 394479 -21982 394535 -21926
rect 394337 -22124 394393 -22068
rect 394479 -22124 394535 -22068
rect 394337 -22266 394393 -22210
rect 394479 -22266 394535 -22210
rect 394337 -22408 394393 -22352
rect 394479 -22408 394535 -22352
rect 394337 -22550 394393 -22494
rect 394479 -22550 394535 -22494
rect 394337 -22692 394393 -22636
rect 394479 -22692 394535 -22636
rect 394337 -22834 394393 -22778
rect 394479 -22834 394535 -22778
rect 394337 -22976 394393 -22920
rect 394479 -22976 394535 -22920
rect 394337 -23118 394393 -23062
rect 394479 -23118 394535 -23062
rect 394337 -23260 394393 -23204
rect 394479 -23260 394535 -23204
rect 394337 -23402 394393 -23346
rect 394479 -23402 394535 -23346
rect 394337 -23544 394393 -23488
rect 394479 -23544 394535 -23488
rect 394337 -23686 394393 -23630
rect 394479 -23686 394535 -23630
rect 394337 -23828 394393 -23772
rect 394479 -23828 394535 -23772
rect 394337 -23970 394393 -23914
rect 394479 -23970 394535 -23914
rect 394337 -24112 394393 -24056
rect 394479 -24112 394535 -24056
rect 394337 -24254 394393 -24198
rect 394479 -24254 394535 -24198
rect 394337 -24396 394393 -24340
rect 394479 -24396 394535 -24340
rect 394337 -24538 394393 -24482
rect 394479 -24538 394535 -24482
rect 394337 -24680 394393 -24624
rect 394479 -24680 394535 -24624
rect 394337 -24822 394393 -24766
rect 394479 -24822 394535 -24766
rect 394337 -24964 394393 -24908
rect 394479 -24964 394535 -24908
rect 394337 -25106 394393 -25050
rect 394479 -25106 394535 -25050
rect 394337 -25248 394393 -25192
rect 394479 -25248 394535 -25192
rect 394337 -25390 394393 -25334
rect 394479 -25390 394535 -25334
rect 394337 -25532 394393 -25476
rect 394479 -25532 394535 -25476
rect 394740 -18006 394796 -17950
rect 394882 -18006 394938 -17950
rect 394740 -18148 394796 -18092
rect 394882 -18148 394938 -18092
rect 394740 -18290 394796 -18234
rect 394882 -18290 394938 -18234
rect 394740 -18432 394796 -18376
rect 394882 -18432 394938 -18376
rect 394740 -18574 394796 -18518
rect 394882 -18574 394938 -18518
rect 394740 -18716 394796 -18660
rect 394882 -18716 394938 -18660
rect 394740 -18858 394796 -18802
rect 394882 -18858 394938 -18802
rect 394740 -19000 394796 -18944
rect 394882 -19000 394938 -18944
rect 394740 -19142 394796 -19086
rect 394882 -19142 394938 -19086
rect 394740 -19284 394796 -19228
rect 394882 -19284 394938 -19228
rect 394740 -19426 394796 -19370
rect 394882 -19426 394938 -19370
rect 394740 -19568 394796 -19512
rect 394882 -19568 394938 -19512
rect 394740 -19710 394796 -19654
rect 394882 -19710 394938 -19654
rect 394740 -19852 394796 -19796
rect 394882 -19852 394938 -19796
rect 394740 -19994 394796 -19938
rect 394882 -19994 394938 -19938
rect 394740 -20136 394796 -20080
rect 394882 -20136 394938 -20080
rect 394740 -20278 394796 -20222
rect 394882 -20278 394938 -20222
rect 394740 -20420 394796 -20364
rect 394882 -20420 394938 -20364
rect 394740 -20562 394796 -20506
rect 394882 -20562 394938 -20506
rect 394740 -20704 394796 -20648
rect 394882 -20704 394938 -20648
rect 394740 -20846 394796 -20790
rect 394882 -20846 394938 -20790
rect 394740 -20988 394796 -20932
rect 394882 -20988 394938 -20932
rect 394740 -21130 394796 -21074
rect 394882 -21130 394938 -21074
rect 394740 -21272 394796 -21216
rect 394882 -21272 394938 -21216
rect 394740 -21414 394796 -21358
rect 394882 -21414 394938 -21358
rect 394740 -21556 394796 -21500
rect 394882 -21556 394938 -21500
rect 394740 -21698 394796 -21642
rect 394882 -21698 394938 -21642
rect 394740 -21840 394796 -21784
rect 394882 -21840 394938 -21784
rect 394740 -21982 394796 -21926
rect 394882 -21982 394938 -21926
rect 394740 -22124 394796 -22068
rect 394882 -22124 394938 -22068
rect 394740 -22266 394796 -22210
rect 394882 -22266 394938 -22210
rect 394740 -22408 394796 -22352
rect 394882 -22408 394938 -22352
rect 394740 -22550 394796 -22494
rect 394882 -22550 394938 -22494
rect 394740 -22692 394796 -22636
rect 394882 -22692 394938 -22636
rect 394740 -22834 394796 -22778
rect 394882 -22834 394938 -22778
rect 394740 -22976 394796 -22920
rect 394882 -22976 394938 -22920
rect 394740 -23118 394796 -23062
rect 394882 -23118 394938 -23062
rect 394740 -23260 394796 -23204
rect 394882 -23260 394938 -23204
rect 394740 -23402 394796 -23346
rect 394882 -23402 394938 -23346
rect 394740 -23544 394796 -23488
rect 394882 -23544 394938 -23488
rect 394740 -23686 394796 -23630
rect 394882 -23686 394938 -23630
rect 394740 -23828 394796 -23772
rect 394882 -23828 394938 -23772
rect 394740 -23970 394796 -23914
rect 394882 -23970 394938 -23914
rect 394740 -24112 394796 -24056
rect 394882 -24112 394938 -24056
rect 394740 -24254 394796 -24198
rect 394882 -24254 394938 -24198
rect 394740 -24396 394796 -24340
rect 394882 -24396 394938 -24340
rect 394740 -24538 394796 -24482
rect 394882 -24538 394938 -24482
rect 394740 -24680 394796 -24624
rect 394882 -24680 394938 -24624
rect 394740 -24822 394796 -24766
rect 394882 -24822 394938 -24766
rect 394740 -24964 394796 -24908
rect 394882 -24964 394938 -24908
rect 394740 -25106 394796 -25050
rect 394882 -25106 394938 -25050
rect 394740 -25248 394796 -25192
rect 394882 -25248 394938 -25192
rect 394740 -25390 394796 -25334
rect 394882 -25390 394938 -25334
rect 394740 -25532 394796 -25476
rect 394882 -25532 394938 -25476
rect 395142 -18006 395198 -17950
rect 395284 -18006 395340 -17950
rect 395142 -18148 395198 -18092
rect 395284 -18148 395340 -18092
rect 395142 -18290 395198 -18234
rect 395284 -18290 395340 -18234
rect 395142 -18432 395198 -18376
rect 395284 -18432 395340 -18376
rect 395142 -18574 395198 -18518
rect 395284 -18574 395340 -18518
rect 395142 -18716 395198 -18660
rect 395284 -18716 395340 -18660
rect 395142 -18858 395198 -18802
rect 395284 -18858 395340 -18802
rect 395142 -19000 395198 -18944
rect 395284 -19000 395340 -18944
rect 395142 -19142 395198 -19086
rect 395284 -19142 395340 -19086
rect 395142 -19284 395198 -19228
rect 395284 -19284 395340 -19228
rect 395142 -19426 395198 -19370
rect 395284 -19426 395340 -19370
rect 395142 -19568 395198 -19512
rect 395284 -19568 395340 -19512
rect 395142 -19710 395198 -19654
rect 395284 -19710 395340 -19654
rect 395142 -19852 395198 -19796
rect 395284 -19852 395340 -19796
rect 395142 -19994 395198 -19938
rect 395284 -19994 395340 -19938
rect 395142 -20136 395198 -20080
rect 395284 -20136 395340 -20080
rect 395142 -20278 395198 -20222
rect 395284 -20278 395340 -20222
rect 395142 -20420 395198 -20364
rect 395284 -20420 395340 -20364
rect 395142 -20562 395198 -20506
rect 395284 -20562 395340 -20506
rect 395142 -20704 395198 -20648
rect 395284 -20704 395340 -20648
rect 395142 -20846 395198 -20790
rect 395284 -20846 395340 -20790
rect 395142 -20988 395198 -20932
rect 395284 -20988 395340 -20932
rect 395142 -21130 395198 -21074
rect 395284 -21130 395340 -21074
rect 395142 -21272 395198 -21216
rect 395284 -21272 395340 -21216
rect 395142 -21414 395198 -21358
rect 395284 -21414 395340 -21358
rect 395142 -21556 395198 -21500
rect 395284 -21556 395340 -21500
rect 395142 -21698 395198 -21642
rect 395284 -21698 395340 -21642
rect 395142 -21840 395198 -21784
rect 395284 -21840 395340 -21784
rect 395142 -21982 395198 -21926
rect 395284 -21982 395340 -21926
rect 395142 -22124 395198 -22068
rect 395284 -22124 395340 -22068
rect 395142 -22266 395198 -22210
rect 395284 -22266 395340 -22210
rect 395142 -22408 395198 -22352
rect 395284 -22408 395340 -22352
rect 395142 -22550 395198 -22494
rect 395284 -22550 395340 -22494
rect 395142 -22692 395198 -22636
rect 395284 -22692 395340 -22636
rect 395142 -22834 395198 -22778
rect 395284 -22834 395340 -22778
rect 395142 -22976 395198 -22920
rect 395284 -22976 395340 -22920
rect 395142 -23118 395198 -23062
rect 395284 -23118 395340 -23062
rect 395142 -23260 395198 -23204
rect 395284 -23260 395340 -23204
rect 395142 -23402 395198 -23346
rect 395284 -23402 395340 -23346
rect 395142 -23544 395198 -23488
rect 395284 -23544 395340 -23488
rect 395142 -23686 395198 -23630
rect 395284 -23686 395340 -23630
rect 395142 -23828 395198 -23772
rect 395284 -23828 395340 -23772
rect 395142 -23970 395198 -23914
rect 395284 -23970 395340 -23914
rect 395142 -24112 395198 -24056
rect 395284 -24112 395340 -24056
rect 395142 -24254 395198 -24198
rect 395284 -24254 395340 -24198
rect 395142 -24396 395198 -24340
rect 395284 -24396 395340 -24340
rect 395142 -24538 395198 -24482
rect 395284 -24538 395340 -24482
rect 395142 -24680 395198 -24624
rect 395284 -24680 395340 -24624
rect 395142 -24822 395198 -24766
rect 395284 -24822 395340 -24766
rect 395142 -24964 395198 -24908
rect 395284 -24964 395340 -24908
rect 395142 -25106 395198 -25050
rect 395284 -25106 395340 -25050
rect 395142 -25248 395198 -25192
rect 395284 -25248 395340 -25192
rect 395142 -25390 395198 -25334
rect 395284 -25390 395340 -25334
rect 395142 -25532 395198 -25476
rect 395284 -25532 395340 -25476
rect 395545 -18006 395601 -17950
rect 395687 -18006 395743 -17950
rect 395545 -18148 395601 -18092
rect 395687 -18148 395743 -18092
rect 395545 -18290 395601 -18234
rect 395687 -18290 395743 -18234
rect 395545 -18432 395601 -18376
rect 395687 -18432 395743 -18376
rect 395545 -18574 395601 -18518
rect 395687 -18574 395743 -18518
rect 395545 -18716 395601 -18660
rect 395687 -18716 395743 -18660
rect 395545 -18858 395601 -18802
rect 395687 -18858 395743 -18802
rect 395545 -19000 395601 -18944
rect 395687 -19000 395743 -18944
rect 395545 -19142 395601 -19086
rect 395687 -19142 395743 -19086
rect 395545 -19284 395601 -19228
rect 395687 -19284 395743 -19228
rect 395545 -19426 395601 -19370
rect 395687 -19426 395743 -19370
rect 395545 -19568 395601 -19512
rect 395687 -19568 395743 -19512
rect 395545 -19710 395601 -19654
rect 395687 -19710 395743 -19654
rect 395545 -19852 395601 -19796
rect 395687 -19852 395743 -19796
rect 395545 -19994 395601 -19938
rect 395687 -19994 395743 -19938
rect 395545 -20136 395601 -20080
rect 395687 -20136 395743 -20080
rect 395545 -20278 395601 -20222
rect 395687 -20278 395743 -20222
rect 395545 -20420 395601 -20364
rect 395687 -20420 395743 -20364
rect 395545 -20562 395601 -20506
rect 395687 -20562 395743 -20506
rect 395545 -20704 395601 -20648
rect 395687 -20704 395743 -20648
rect 395545 -20846 395601 -20790
rect 395687 -20846 395743 -20790
rect 395545 -20988 395601 -20932
rect 395687 -20988 395743 -20932
rect 395545 -21130 395601 -21074
rect 395687 -21130 395743 -21074
rect 395545 -21272 395601 -21216
rect 395687 -21272 395743 -21216
rect 395545 -21414 395601 -21358
rect 395687 -21414 395743 -21358
rect 395545 -21556 395601 -21500
rect 395687 -21556 395743 -21500
rect 395545 -21698 395601 -21642
rect 395687 -21698 395743 -21642
rect 395545 -21840 395601 -21784
rect 395687 -21840 395743 -21784
rect 395545 -21982 395601 -21926
rect 395687 -21982 395743 -21926
rect 395545 -22124 395601 -22068
rect 395687 -22124 395743 -22068
rect 395545 -22266 395601 -22210
rect 395687 -22266 395743 -22210
rect 395545 -22408 395601 -22352
rect 395687 -22408 395743 -22352
rect 395545 -22550 395601 -22494
rect 395687 -22550 395743 -22494
rect 395545 -22692 395601 -22636
rect 395687 -22692 395743 -22636
rect 395545 -22834 395601 -22778
rect 395687 -22834 395743 -22778
rect 395545 -22976 395601 -22920
rect 395687 -22976 395743 -22920
rect 395545 -23118 395601 -23062
rect 395687 -23118 395743 -23062
rect 395545 -23260 395601 -23204
rect 395687 -23260 395743 -23204
rect 395545 -23402 395601 -23346
rect 395687 -23402 395743 -23346
rect 395545 -23544 395601 -23488
rect 395687 -23544 395743 -23488
rect 395545 -23686 395601 -23630
rect 395687 -23686 395743 -23630
rect 395545 -23828 395601 -23772
rect 395687 -23828 395743 -23772
rect 395545 -23970 395601 -23914
rect 395687 -23970 395743 -23914
rect 395545 -24112 395601 -24056
rect 395687 -24112 395743 -24056
rect 395545 -24254 395601 -24198
rect 395687 -24254 395743 -24198
rect 395545 -24396 395601 -24340
rect 395687 -24396 395743 -24340
rect 395545 -24538 395601 -24482
rect 395687 -24538 395743 -24482
rect 395545 -24680 395601 -24624
rect 395687 -24680 395743 -24624
rect 395545 -24822 395601 -24766
rect 395687 -24822 395743 -24766
rect 395545 -24964 395601 -24908
rect 395687 -24964 395743 -24908
rect 395545 -25106 395601 -25050
rect 395687 -25106 395743 -25050
rect 395545 -25248 395601 -25192
rect 395687 -25248 395743 -25192
rect 395545 -25390 395601 -25334
rect 395687 -25390 395743 -25334
rect 395545 -25532 395601 -25476
rect 395687 -25532 395743 -25476
rect 395941 -18006 395997 -17950
rect 396083 -18006 396139 -17950
rect 395941 -18148 395997 -18092
rect 396083 -18148 396139 -18092
rect 395941 -18290 395997 -18234
rect 396083 -18290 396139 -18234
rect 395941 -18432 395997 -18376
rect 396083 -18432 396139 -18376
rect 395941 -18574 395997 -18518
rect 396083 -18574 396139 -18518
rect 395941 -18716 395997 -18660
rect 396083 -18716 396139 -18660
rect 395941 -18858 395997 -18802
rect 396083 -18858 396139 -18802
rect 395941 -19000 395997 -18944
rect 396083 -19000 396139 -18944
rect 395941 -19142 395997 -19086
rect 396083 -19142 396139 -19086
rect 395941 -19284 395997 -19228
rect 396083 -19284 396139 -19228
rect 395941 -19426 395997 -19370
rect 396083 -19426 396139 -19370
rect 395941 -19568 395997 -19512
rect 396083 -19568 396139 -19512
rect 395941 -19710 395997 -19654
rect 396083 -19710 396139 -19654
rect 395941 -19852 395997 -19796
rect 396083 -19852 396139 -19796
rect 395941 -19994 395997 -19938
rect 396083 -19994 396139 -19938
rect 395941 -20136 395997 -20080
rect 396083 -20136 396139 -20080
rect 395941 -20278 395997 -20222
rect 396083 -20278 396139 -20222
rect 395941 -20420 395997 -20364
rect 396083 -20420 396139 -20364
rect 395941 -20562 395997 -20506
rect 396083 -20562 396139 -20506
rect 395941 -20704 395997 -20648
rect 396083 -20704 396139 -20648
rect 395941 -20846 395997 -20790
rect 396083 -20846 396139 -20790
rect 395941 -20988 395997 -20932
rect 396083 -20988 396139 -20932
rect 395941 -21130 395997 -21074
rect 396083 -21130 396139 -21074
rect 395941 -21272 395997 -21216
rect 396083 -21272 396139 -21216
rect 395941 -21414 395997 -21358
rect 396083 -21414 396139 -21358
rect 395941 -21556 395997 -21500
rect 396083 -21556 396139 -21500
rect 395941 -21698 395997 -21642
rect 396083 -21698 396139 -21642
rect 395941 -21840 395997 -21784
rect 396083 -21840 396139 -21784
rect 395941 -21982 395997 -21926
rect 396083 -21982 396139 -21926
rect 395941 -22124 395997 -22068
rect 396083 -22124 396139 -22068
rect 395941 -22266 395997 -22210
rect 396083 -22266 396139 -22210
rect 395941 -22408 395997 -22352
rect 396083 -22408 396139 -22352
rect 395941 -22550 395997 -22494
rect 396083 -22550 396139 -22494
rect 395941 -22692 395997 -22636
rect 396083 -22692 396139 -22636
rect 395941 -22834 395997 -22778
rect 396083 -22834 396139 -22778
rect 395941 -22976 395997 -22920
rect 396083 -22976 396139 -22920
rect 395941 -23118 395997 -23062
rect 396083 -23118 396139 -23062
rect 395941 -23260 395997 -23204
rect 396083 -23260 396139 -23204
rect 395941 -23402 395997 -23346
rect 396083 -23402 396139 -23346
rect 395941 -23544 395997 -23488
rect 396083 -23544 396139 -23488
rect 395941 -23686 395997 -23630
rect 396083 -23686 396139 -23630
rect 395941 -23828 395997 -23772
rect 396083 -23828 396139 -23772
rect 395941 -23970 395997 -23914
rect 396083 -23970 396139 -23914
rect 395941 -24112 395997 -24056
rect 396083 -24112 396139 -24056
rect 395941 -24254 395997 -24198
rect 396083 -24254 396139 -24198
rect 395941 -24396 395997 -24340
rect 396083 -24396 396139 -24340
rect 395941 -24538 395997 -24482
rect 396083 -24538 396139 -24482
rect 395941 -24680 395997 -24624
rect 396083 -24680 396139 -24624
rect 395941 -24822 395997 -24766
rect 396083 -24822 396139 -24766
rect 395941 -24964 395997 -24908
rect 396083 -24964 396139 -24908
rect 395941 -25106 395997 -25050
rect 396083 -25106 396139 -25050
rect 395941 -25248 395997 -25192
rect 396083 -25248 396139 -25192
rect 395941 -25390 395997 -25334
rect 396083 -25390 396139 -25334
rect 395941 -25532 395997 -25476
rect 396083 -25532 396139 -25476
rect 396526 -17914 396582 -17858
rect 396650 -17914 396706 -17858
rect 396774 -17914 396830 -17858
rect 396898 -17914 396954 -17858
rect 397022 -17914 397078 -17858
rect 396526 -18038 396582 -17982
rect 396650 -18038 396706 -17982
rect 396774 -18038 396830 -17982
rect 396898 -18038 396954 -17982
rect 397022 -18038 397078 -17982
rect 396526 -18162 396582 -18106
rect 396650 -18162 396706 -18106
rect 396774 -18162 396830 -18106
rect 396898 -18162 396954 -18106
rect 397022 -18162 397078 -18106
rect 396526 -18286 396582 -18230
rect 396650 -18286 396706 -18230
rect 396774 -18286 396830 -18230
rect 396898 -18286 396954 -18230
rect 397022 -18286 397078 -18230
rect 396526 -18410 396582 -18354
rect 396650 -18410 396706 -18354
rect 396774 -18410 396830 -18354
rect 396898 -18410 396954 -18354
rect 397022 -18410 397078 -18354
rect 396526 -18534 396582 -18478
rect 396650 -18534 396706 -18478
rect 396774 -18534 396830 -18478
rect 396898 -18534 396954 -18478
rect 397022 -18534 397078 -18478
rect 396526 -18658 396582 -18602
rect 396650 -18658 396706 -18602
rect 396774 -18658 396830 -18602
rect 396898 -18658 396954 -18602
rect 397022 -18658 397078 -18602
rect 396526 -18782 396582 -18726
rect 396650 -18782 396706 -18726
rect 396774 -18782 396830 -18726
rect 396898 -18782 396954 -18726
rect 397022 -18782 397078 -18726
rect 396526 -18906 396582 -18850
rect 396650 -18906 396706 -18850
rect 396774 -18906 396830 -18850
rect 396898 -18906 396954 -18850
rect 397022 -18906 397078 -18850
rect 396526 -19030 396582 -18974
rect 396650 -19030 396706 -18974
rect 396774 -19030 396830 -18974
rect 396898 -19030 396954 -18974
rect 397022 -19030 397078 -18974
rect 396526 -19154 396582 -19098
rect 396650 -19154 396706 -19098
rect 396774 -19154 396830 -19098
rect 396898 -19154 396954 -19098
rect 397022 -19154 397078 -19098
rect 396526 -19278 396582 -19222
rect 396650 -19278 396706 -19222
rect 396774 -19278 396830 -19222
rect 396898 -19278 396954 -19222
rect 397022 -19278 397078 -19222
rect 396526 -19402 396582 -19346
rect 396650 -19402 396706 -19346
rect 396774 -19402 396830 -19346
rect 396898 -19402 396954 -19346
rect 397022 -19402 397078 -19346
rect 396526 -19526 396582 -19470
rect 396650 -19526 396706 -19470
rect 396774 -19526 396830 -19470
rect 396898 -19526 396954 -19470
rect 397022 -19526 397078 -19470
rect 396526 -19650 396582 -19594
rect 396650 -19650 396706 -19594
rect 396774 -19650 396830 -19594
rect 396898 -19650 396954 -19594
rect 397022 -19650 397078 -19594
rect 396526 -19774 396582 -19718
rect 396650 -19774 396706 -19718
rect 396774 -19774 396830 -19718
rect 396898 -19774 396954 -19718
rect 397022 -19774 397078 -19718
rect 396526 -19898 396582 -19842
rect 396650 -19898 396706 -19842
rect 396774 -19898 396830 -19842
rect 396898 -19898 396954 -19842
rect 397022 -19898 397078 -19842
rect 396526 -20022 396582 -19966
rect 396650 -20022 396706 -19966
rect 396774 -20022 396830 -19966
rect 396898 -20022 396954 -19966
rect 397022 -20022 397078 -19966
rect 396526 -20146 396582 -20090
rect 396650 -20146 396706 -20090
rect 396774 -20146 396830 -20090
rect 396898 -20146 396954 -20090
rect 397022 -20146 397078 -20090
rect 396526 -20270 396582 -20214
rect 396650 -20270 396706 -20214
rect 396774 -20270 396830 -20214
rect 396898 -20270 396954 -20214
rect 397022 -20270 397078 -20214
rect 396526 -20394 396582 -20338
rect 396650 -20394 396706 -20338
rect 396774 -20394 396830 -20338
rect 396898 -20394 396954 -20338
rect 397022 -20394 397078 -20338
rect 396526 -20518 396582 -20462
rect 396650 -20518 396706 -20462
rect 396774 -20518 396830 -20462
rect 396898 -20518 396954 -20462
rect 397022 -20518 397078 -20462
rect 396526 -20642 396582 -20586
rect 396650 -20642 396706 -20586
rect 396774 -20642 396830 -20586
rect 396898 -20642 396954 -20586
rect 397022 -20642 397078 -20586
rect 396526 -20766 396582 -20710
rect 396650 -20766 396706 -20710
rect 396774 -20766 396830 -20710
rect 396898 -20766 396954 -20710
rect 397022 -20766 397078 -20710
rect 396526 -20890 396582 -20834
rect 396650 -20890 396706 -20834
rect 396774 -20890 396830 -20834
rect 396898 -20890 396954 -20834
rect 397022 -20890 397078 -20834
rect 396526 -21014 396582 -20958
rect 396650 -21014 396706 -20958
rect 396774 -21014 396830 -20958
rect 396898 -21014 396954 -20958
rect 397022 -21014 397078 -20958
rect 396526 -21138 396582 -21082
rect 396650 -21138 396706 -21082
rect 396774 -21138 396830 -21082
rect 396898 -21138 396954 -21082
rect 397022 -21138 397078 -21082
rect 396526 -21262 396582 -21206
rect 396650 -21262 396706 -21206
rect 396774 -21262 396830 -21206
rect 396898 -21262 396954 -21206
rect 397022 -21262 397078 -21206
rect 396526 -21386 396582 -21330
rect 396650 -21386 396706 -21330
rect 396774 -21386 396830 -21330
rect 396898 -21386 396954 -21330
rect 397022 -21386 397078 -21330
rect 396526 -21510 396582 -21454
rect 396650 -21510 396706 -21454
rect 396774 -21510 396830 -21454
rect 396898 -21510 396954 -21454
rect 397022 -21510 397078 -21454
rect 396526 -21634 396582 -21578
rect 396650 -21634 396706 -21578
rect 396774 -21634 396830 -21578
rect 396898 -21634 396954 -21578
rect 397022 -21634 397078 -21578
rect 396526 -21758 396582 -21702
rect 396650 -21758 396706 -21702
rect 396774 -21758 396830 -21702
rect 396898 -21758 396954 -21702
rect 397022 -21758 397078 -21702
rect 396526 -21882 396582 -21826
rect 396650 -21882 396706 -21826
rect 396774 -21882 396830 -21826
rect 396898 -21882 396954 -21826
rect 397022 -21882 397078 -21826
rect 396526 -22006 396582 -21950
rect 396650 -22006 396706 -21950
rect 396774 -22006 396830 -21950
rect 396898 -22006 396954 -21950
rect 397022 -22006 397078 -21950
rect 396526 -22130 396582 -22074
rect 396650 -22130 396706 -22074
rect 396774 -22130 396830 -22074
rect 396898 -22130 396954 -22074
rect 397022 -22130 397078 -22074
rect 396526 -22254 396582 -22198
rect 396650 -22254 396706 -22198
rect 396774 -22254 396830 -22198
rect 396898 -22254 396954 -22198
rect 397022 -22254 397078 -22198
rect 396526 -22378 396582 -22322
rect 396650 -22378 396706 -22322
rect 396774 -22378 396830 -22322
rect 396898 -22378 396954 -22322
rect 397022 -22378 397078 -22322
rect 396526 -22502 396582 -22446
rect 396650 -22502 396706 -22446
rect 396774 -22502 396830 -22446
rect 396898 -22502 396954 -22446
rect 397022 -22502 397078 -22446
rect 396526 -22626 396582 -22570
rect 396650 -22626 396706 -22570
rect 396774 -22626 396830 -22570
rect 396898 -22626 396954 -22570
rect 397022 -22626 397078 -22570
rect 396526 -22750 396582 -22694
rect 396650 -22750 396706 -22694
rect 396774 -22750 396830 -22694
rect 396898 -22750 396954 -22694
rect 397022 -22750 397078 -22694
rect 396526 -22874 396582 -22818
rect 396650 -22874 396706 -22818
rect 396774 -22874 396830 -22818
rect 396898 -22874 396954 -22818
rect 397022 -22874 397078 -22818
rect 396526 -22998 396582 -22942
rect 396650 -22998 396706 -22942
rect 396774 -22998 396830 -22942
rect 396898 -22998 396954 -22942
rect 397022 -22998 397078 -22942
rect 396526 -23122 396582 -23066
rect 396650 -23122 396706 -23066
rect 396774 -23122 396830 -23066
rect 396898 -23122 396954 -23066
rect 397022 -23122 397078 -23066
rect 396526 -23246 396582 -23190
rect 396650 -23246 396706 -23190
rect 396774 -23246 396830 -23190
rect 396898 -23246 396954 -23190
rect 397022 -23246 397078 -23190
rect 396526 -23370 396582 -23314
rect 396650 -23370 396706 -23314
rect 396774 -23370 396830 -23314
rect 396898 -23370 396954 -23314
rect 397022 -23370 397078 -23314
rect 396526 -23494 396582 -23438
rect 396650 -23494 396706 -23438
rect 396774 -23494 396830 -23438
rect 396898 -23494 396954 -23438
rect 397022 -23494 397078 -23438
rect 396526 -23618 396582 -23562
rect 396650 -23618 396706 -23562
rect 396774 -23618 396830 -23562
rect 396898 -23618 396954 -23562
rect 397022 -23618 397078 -23562
rect 396526 -23742 396582 -23686
rect 396650 -23742 396706 -23686
rect 396774 -23742 396830 -23686
rect 396898 -23742 396954 -23686
rect 397022 -23742 397078 -23686
rect 396526 -23866 396582 -23810
rect 396650 -23866 396706 -23810
rect 396774 -23866 396830 -23810
rect 396898 -23866 396954 -23810
rect 397022 -23866 397078 -23810
rect 396526 -23990 396582 -23934
rect 396650 -23990 396706 -23934
rect 396774 -23990 396830 -23934
rect 396898 -23990 396954 -23934
rect 397022 -23990 397078 -23934
rect 396526 -24114 396582 -24058
rect 396650 -24114 396706 -24058
rect 396774 -24114 396830 -24058
rect 396898 -24114 396954 -24058
rect 397022 -24114 397078 -24058
rect 396526 -24238 396582 -24182
rect 396650 -24238 396706 -24182
rect 396774 -24238 396830 -24182
rect 396898 -24238 396954 -24182
rect 397022 -24238 397078 -24182
rect 396526 -24362 396582 -24306
rect 396650 -24362 396706 -24306
rect 396774 -24362 396830 -24306
rect 396898 -24362 396954 -24306
rect 397022 -24362 397078 -24306
rect 396526 -24486 396582 -24430
rect 396650 -24486 396706 -24430
rect 396774 -24486 396830 -24430
rect 396898 -24486 396954 -24430
rect 397022 -24486 397078 -24430
rect 396526 -24610 396582 -24554
rect 396650 -24610 396706 -24554
rect 396774 -24610 396830 -24554
rect 396898 -24610 396954 -24554
rect 397022 -24610 397078 -24554
rect 396526 -24734 396582 -24678
rect 396650 -24734 396706 -24678
rect 396774 -24734 396830 -24678
rect 396898 -24734 396954 -24678
rect 397022 -24734 397078 -24678
rect 396526 -24858 396582 -24802
rect 396650 -24858 396706 -24802
rect 396774 -24858 396830 -24802
rect 396898 -24858 396954 -24802
rect 397022 -24858 397078 -24802
rect 396526 -24982 396582 -24926
rect 396650 -24982 396706 -24926
rect 396774 -24982 396830 -24926
rect 396898 -24982 396954 -24926
rect 397022 -24982 397078 -24926
rect 396526 -25106 396582 -25050
rect 396650 -25106 396706 -25050
rect 396774 -25106 396830 -25050
rect 396898 -25106 396954 -25050
rect 397022 -25106 397078 -25050
rect 396526 -25230 396582 -25174
rect 396650 -25230 396706 -25174
rect 396774 -25230 396830 -25174
rect 396898 -25230 396954 -25174
rect 397022 -25230 397078 -25174
rect 396526 -25354 396582 -25298
rect 396650 -25354 396706 -25298
rect 396774 -25354 396830 -25298
rect 396898 -25354 396954 -25298
rect 397022 -25354 397078 -25298
rect 396526 -25478 396582 -25422
rect 396650 -25478 396706 -25422
rect 396774 -25478 396830 -25422
rect 396898 -25478 396954 -25422
rect 397022 -25478 397078 -25422
rect 388146 -25777 388202 -25721
rect 388270 -25777 388326 -25721
rect 388394 -25777 388450 -25721
rect 388518 -25777 388574 -25721
rect 388642 -25777 388698 -25721
rect 388766 -25777 388822 -25721
rect 388890 -25777 388946 -25721
rect 389014 -25777 389070 -25721
rect 389138 -25777 389194 -25721
rect 389262 -25777 389318 -25721
rect 389386 -25777 389442 -25721
rect 389510 -25777 389566 -25721
rect 389634 -25777 389690 -25721
rect 389758 -25777 389814 -25721
rect 389882 -25777 389938 -25721
rect 390006 -25777 390062 -25721
rect 390130 -25777 390186 -25721
rect 390254 -25777 390310 -25721
rect 390378 -25777 390434 -25721
rect 390502 -25777 390558 -25721
rect 390626 -25777 390682 -25721
rect 390750 -25777 390806 -25721
rect 390874 -25777 390930 -25721
rect 390998 -25777 391054 -25721
rect 391122 -25777 391178 -25721
rect 391246 -25777 391302 -25721
rect 391370 -25777 391426 -25721
rect 391494 -25777 391550 -25721
rect 391618 -25777 391674 -25721
rect 391742 -25777 391798 -25721
rect 391866 -25777 391922 -25721
rect 391990 -25777 392046 -25721
rect 392114 -25777 392170 -25721
rect 392238 -25777 392294 -25721
rect 392362 -25777 392418 -25721
rect 392486 -25777 392542 -25721
rect 392610 -25777 392666 -25721
rect 392734 -25777 392790 -25721
rect 392858 -25777 392914 -25721
rect 392982 -25777 393038 -25721
rect 393106 -25777 393162 -25721
rect 393230 -25777 393286 -25721
rect 393354 -25777 393410 -25721
rect 393478 -25777 393534 -25721
rect 393602 -25777 393658 -25721
rect 393726 -25777 393782 -25721
rect 393850 -25777 393906 -25721
rect 393974 -25777 394030 -25721
rect 394098 -25777 394154 -25721
rect 394222 -25777 394278 -25721
rect 394346 -25777 394402 -25721
rect 394470 -25777 394526 -25721
rect 394594 -25777 394650 -25721
rect 394718 -25777 394774 -25721
rect 394842 -25777 394898 -25721
rect 394966 -25777 395022 -25721
rect 395090 -25777 395146 -25721
rect 395214 -25777 395270 -25721
rect 395338 -25777 395394 -25721
rect 395462 -25777 395518 -25721
rect 395586 -25777 395642 -25721
rect 395710 -25777 395766 -25721
rect 395898 -25777 395954 -25721
rect 396022 -25777 396078 -25721
rect 396146 -25777 396202 -25721
rect 396270 -25777 396326 -25721
rect 396394 -25777 396450 -25721
rect 396518 -25777 396574 -25721
rect 396642 -25777 396698 -25721
rect 396766 -25777 396822 -25721
rect 396890 -25777 396946 -25721
rect 397014 -25777 397070 -25721
rect 388146 -25901 388202 -25845
rect 388270 -25901 388326 -25845
rect 388394 -25901 388450 -25845
rect 388518 -25901 388574 -25845
rect 388642 -25901 388698 -25845
rect 388766 -25901 388822 -25845
rect 388890 -25901 388946 -25845
rect 389014 -25901 389070 -25845
rect 389138 -25901 389194 -25845
rect 389262 -25901 389318 -25845
rect 389386 -25901 389442 -25845
rect 389510 -25901 389566 -25845
rect 389634 -25901 389690 -25845
rect 389758 -25901 389814 -25845
rect 389882 -25901 389938 -25845
rect 390006 -25901 390062 -25845
rect 390130 -25901 390186 -25845
rect 390254 -25901 390310 -25845
rect 390378 -25901 390434 -25845
rect 390502 -25901 390558 -25845
rect 390626 -25901 390682 -25845
rect 390750 -25901 390806 -25845
rect 390874 -25901 390930 -25845
rect 390998 -25901 391054 -25845
rect 391122 -25901 391178 -25845
rect 391246 -25901 391302 -25845
rect 391370 -25901 391426 -25845
rect 391494 -25901 391550 -25845
rect 391618 -25901 391674 -25845
rect 391742 -25901 391798 -25845
rect 391866 -25901 391922 -25845
rect 391990 -25901 392046 -25845
rect 392114 -25901 392170 -25845
rect 392238 -25901 392294 -25845
rect 392362 -25901 392418 -25845
rect 392486 -25901 392542 -25845
rect 392610 -25901 392666 -25845
rect 392734 -25901 392790 -25845
rect 392858 -25901 392914 -25845
rect 392982 -25901 393038 -25845
rect 393106 -25901 393162 -25845
rect 393230 -25901 393286 -25845
rect 393354 -25901 393410 -25845
rect 393478 -25901 393534 -25845
rect 393602 -25901 393658 -25845
rect 393726 -25901 393782 -25845
rect 393850 -25901 393906 -25845
rect 393974 -25901 394030 -25845
rect 394098 -25901 394154 -25845
rect 394222 -25901 394278 -25845
rect 394346 -25901 394402 -25845
rect 394470 -25901 394526 -25845
rect 394594 -25901 394650 -25845
rect 394718 -25901 394774 -25845
rect 394842 -25901 394898 -25845
rect 394966 -25901 395022 -25845
rect 395090 -25901 395146 -25845
rect 395214 -25901 395270 -25845
rect 395338 -25901 395394 -25845
rect 395462 -25901 395518 -25845
rect 395586 -25901 395642 -25845
rect 395710 -25901 395766 -25845
rect 395898 -25901 395954 -25845
rect 396022 -25901 396078 -25845
rect 396146 -25901 396202 -25845
rect 396270 -25901 396326 -25845
rect 396394 -25901 396450 -25845
rect 396518 -25901 396574 -25845
rect 396642 -25901 396698 -25845
rect 396766 -25901 396822 -25845
rect 396890 -25901 396946 -25845
rect 397014 -25901 397070 -25845
rect 388146 -26025 388202 -25969
rect 388270 -26025 388326 -25969
rect 388394 -26025 388450 -25969
rect 388518 -26025 388574 -25969
rect 388642 -26025 388698 -25969
rect 388766 -26025 388822 -25969
rect 388890 -26025 388946 -25969
rect 389014 -26025 389070 -25969
rect 389138 -26025 389194 -25969
rect 389262 -26025 389318 -25969
rect 389386 -26025 389442 -25969
rect 389510 -26025 389566 -25969
rect 389634 -26025 389690 -25969
rect 389758 -26025 389814 -25969
rect 389882 -26025 389938 -25969
rect 390006 -26025 390062 -25969
rect 390130 -26025 390186 -25969
rect 390254 -26025 390310 -25969
rect 390378 -26025 390434 -25969
rect 390502 -26025 390558 -25969
rect 390626 -26025 390682 -25969
rect 390750 -26025 390806 -25969
rect 390874 -26025 390930 -25969
rect 390998 -26025 391054 -25969
rect 391122 -26025 391178 -25969
rect 391246 -26025 391302 -25969
rect 391370 -26025 391426 -25969
rect 391494 -26025 391550 -25969
rect 391618 -26025 391674 -25969
rect 391742 -26025 391798 -25969
rect 391866 -26025 391922 -25969
rect 391990 -26025 392046 -25969
rect 392114 -26025 392170 -25969
rect 392238 -26025 392294 -25969
rect 392362 -26025 392418 -25969
rect 392486 -26025 392542 -25969
rect 392610 -26025 392666 -25969
rect 392734 -26025 392790 -25969
rect 392858 -26025 392914 -25969
rect 392982 -26025 393038 -25969
rect 393106 -26025 393162 -25969
rect 393230 -26025 393286 -25969
rect 393354 -26025 393410 -25969
rect 393478 -26025 393534 -25969
rect 393602 -26025 393658 -25969
rect 393726 -26025 393782 -25969
rect 393850 -26025 393906 -25969
rect 393974 -26025 394030 -25969
rect 394098 -26025 394154 -25969
rect 394222 -26025 394278 -25969
rect 394346 -26025 394402 -25969
rect 394470 -26025 394526 -25969
rect 394594 -26025 394650 -25969
rect 394718 -26025 394774 -25969
rect 394842 -26025 394898 -25969
rect 394966 -26025 395022 -25969
rect 395090 -26025 395146 -25969
rect 395214 -26025 395270 -25969
rect 395338 -26025 395394 -25969
rect 395462 -26025 395518 -25969
rect 395586 -26025 395642 -25969
rect 395710 -26025 395766 -25969
rect 395898 -26025 395954 -25969
rect 396022 -26025 396078 -25969
rect 396146 -26025 396202 -25969
rect 396270 -26025 396326 -25969
rect 396394 -26025 396450 -25969
rect 396518 -26025 396574 -25969
rect 396642 -26025 396698 -25969
rect 396766 -26025 396822 -25969
rect 396890 -26025 396946 -25969
rect 397014 -26025 397070 -25969
rect 388146 -26149 388202 -26093
rect 388270 -26149 388326 -26093
rect 388394 -26149 388450 -26093
rect 388518 -26149 388574 -26093
rect 388642 -26149 388698 -26093
rect 388766 -26149 388822 -26093
rect 388890 -26149 388946 -26093
rect 389014 -26149 389070 -26093
rect 389138 -26149 389194 -26093
rect 389262 -26149 389318 -26093
rect 389386 -26149 389442 -26093
rect 389510 -26149 389566 -26093
rect 389634 -26149 389690 -26093
rect 389758 -26149 389814 -26093
rect 389882 -26149 389938 -26093
rect 390006 -26149 390062 -26093
rect 390130 -26149 390186 -26093
rect 390254 -26149 390310 -26093
rect 390378 -26149 390434 -26093
rect 390502 -26149 390558 -26093
rect 390626 -26149 390682 -26093
rect 390750 -26149 390806 -26093
rect 390874 -26149 390930 -26093
rect 390998 -26149 391054 -26093
rect 391122 -26149 391178 -26093
rect 391246 -26149 391302 -26093
rect 391370 -26149 391426 -26093
rect 391494 -26149 391550 -26093
rect 391618 -26149 391674 -26093
rect 391742 -26149 391798 -26093
rect 391866 -26149 391922 -26093
rect 391990 -26149 392046 -26093
rect 392114 -26149 392170 -26093
rect 392238 -26149 392294 -26093
rect 392362 -26149 392418 -26093
rect 392486 -26149 392542 -26093
rect 392610 -26149 392666 -26093
rect 392734 -26149 392790 -26093
rect 392858 -26149 392914 -26093
rect 392982 -26149 393038 -26093
rect 393106 -26149 393162 -26093
rect 393230 -26149 393286 -26093
rect 393354 -26149 393410 -26093
rect 393478 -26149 393534 -26093
rect 393602 -26149 393658 -26093
rect 393726 -26149 393782 -26093
rect 393850 -26149 393906 -26093
rect 393974 -26149 394030 -26093
rect 394098 -26149 394154 -26093
rect 394222 -26149 394278 -26093
rect 394346 -26149 394402 -26093
rect 394470 -26149 394526 -26093
rect 394594 -26149 394650 -26093
rect 394718 -26149 394774 -26093
rect 394842 -26149 394898 -26093
rect 394966 -26149 395022 -26093
rect 395090 -26149 395146 -26093
rect 395214 -26149 395270 -26093
rect 395338 -26149 395394 -26093
rect 395462 -26149 395518 -26093
rect 395586 -26149 395642 -26093
rect 395710 -26149 395766 -26093
rect 395898 -26149 395954 -26093
rect 396022 -26149 396078 -26093
rect 396146 -26149 396202 -26093
rect 396270 -26149 396326 -26093
rect 396394 -26149 396450 -26093
rect 396518 -26149 396574 -26093
rect 396642 -26149 396698 -26093
rect 396766 -26149 396822 -26093
rect 396890 -26149 396946 -26093
rect 397014 -26149 397070 -26093
<< metal4 >>
rect 388000 -17191 397200 -17070
rect 388000 -17247 388146 -17191
rect 388202 -17247 388270 -17191
rect 388326 -17247 388394 -17191
rect 388450 -17247 388518 -17191
rect 388574 -17247 388642 -17191
rect 388698 -17247 388766 -17191
rect 388822 -17247 388890 -17191
rect 388946 -17247 389014 -17191
rect 389070 -17247 389138 -17191
rect 389194 -17247 389262 -17191
rect 389318 -17247 389386 -17191
rect 389442 -17247 389510 -17191
rect 389566 -17247 389634 -17191
rect 389690 -17247 389758 -17191
rect 389814 -17247 389882 -17191
rect 389938 -17247 390006 -17191
rect 390062 -17247 390130 -17191
rect 390186 -17247 390254 -17191
rect 390310 -17247 390378 -17191
rect 390434 -17247 390502 -17191
rect 390558 -17247 390626 -17191
rect 390682 -17247 390750 -17191
rect 390806 -17247 390874 -17191
rect 390930 -17247 390998 -17191
rect 391054 -17247 391122 -17191
rect 391178 -17247 391246 -17191
rect 391302 -17247 391370 -17191
rect 391426 -17247 391494 -17191
rect 391550 -17247 391618 -17191
rect 391674 -17247 391742 -17191
rect 391798 -17247 391866 -17191
rect 391922 -17247 391990 -17191
rect 392046 -17247 392114 -17191
rect 392170 -17247 392238 -17191
rect 392294 -17247 392362 -17191
rect 392418 -17247 392486 -17191
rect 392542 -17247 392610 -17191
rect 392666 -17247 392734 -17191
rect 392790 -17247 392858 -17191
rect 392914 -17247 392982 -17191
rect 393038 -17247 393106 -17191
rect 393162 -17247 393230 -17191
rect 393286 -17247 393354 -17191
rect 393410 -17247 393478 -17191
rect 393534 -17247 393602 -17191
rect 393658 -17247 393726 -17191
rect 393782 -17247 393850 -17191
rect 393906 -17247 393974 -17191
rect 394030 -17247 394098 -17191
rect 394154 -17247 394222 -17191
rect 394278 -17247 394346 -17191
rect 394402 -17247 394470 -17191
rect 394526 -17247 394594 -17191
rect 394650 -17247 394718 -17191
rect 394774 -17247 394842 -17191
rect 394898 -17247 394966 -17191
rect 395022 -17247 395090 -17191
rect 395146 -17247 395214 -17191
rect 395270 -17247 395338 -17191
rect 395394 -17247 395462 -17191
rect 395518 -17247 395586 -17191
rect 395642 -17247 395710 -17191
rect 395766 -17247 395898 -17191
rect 395954 -17247 396022 -17191
rect 396078 -17247 396146 -17191
rect 396202 -17247 396270 -17191
rect 396326 -17247 396394 -17191
rect 396450 -17247 396518 -17191
rect 396574 -17247 396642 -17191
rect 396698 -17247 396766 -17191
rect 396822 -17247 396890 -17191
rect 396946 -17247 397014 -17191
rect 397070 -17247 397200 -17191
rect 388000 -17315 397200 -17247
rect 388000 -17371 388146 -17315
rect 388202 -17371 388270 -17315
rect 388326 -17371 388394 -17315
rect 388450 -17371 388518 -17315
rect 388574 -17371 388642 -17315
rect 388698 -17371 388766 -17315
rect 388822 -17371 388890 -17315
rect 388946 -17371 389014 -17315
rect 389070 -17371 389138 -17315
rect 389194 -17371 389262 -17315
rect 389318 -17371 389386 -17315
rect 389442 -17371 389510 -17315
rect 389566 -17371 389634 -17315
rect 389690 -17371 389758 -17315
rect 389814 -17371 389882 -17315
rect 389938 -17371 390006 -17315
rect 390062 -17371 390130 -17315
rect 390186 -17371 390254 -17315
rect 390310 -17371 390378 -17315
rect 390434 -17371 390502 -17315
rect 390558 -17371 390626 -17315
rect 390682 -17371 390750 -17315
rect 390806 -17371 390874 -17315
rect 390930 -17371 390998 -17315
rect 391054 -17371 391122 -17315
rect 391178 -17371 391246 -17315
rect 391302 -17371 391370 -17315
rect 391426 -17371 391494 -17315
rect 391550 -17371 391618 -17315
rect 391674 -17371 391742 -17315
rect 391798 -17371 391866 -17315
rect 391922 -17371 391990 -17315
rect 392046 -17371 392114 -17315
rect 392170 -17371 392238 -17315
rect 392294 -17371 392362 -17315
rect 392418 -17371 392486 -17315
rect 392542 -17371 392610 -17315
rect 392666 -17371 392734 -17315
rect 392790 -17371 392858 -17315
rect 392914 -17371 392982 -17315
rect 393038 -17371 393106 -17315
rect 393162 -17371 393230 -17315
rect 393286 -17371 393354 -17315
rect 393410 -17371 393478 -17315
rect 393534 -17371 393602 -17315
rect 393658 -17371 393726 -17315
rect 393782 -17371 393850 -17315
rect 393906 -17371 393974 -17315
rect 394030 -17371 394098 -17315
rect 394154 -17371 394222 -17315
rect 394278 -17371 394346 -17315
rect 394402 -17371 394470 -17315
rect 394526 -17371 394594 -17315
rect 394650 -17371 394718 -17315
rect 394774 -17371 394842 -17315
rect 394898 -17371 394966 -17315
rect 395022 -17371 395090 -17315
rect 395146 -17371 395214 -17315
rect 395270 -17371 395338 -17315
rect 395394 -17371 395462 -17315
rect 395518 -17371 395586 -17315
rect 395642 -17371 395710 -17315
rect 395766 -17371 395898 -17315
rect 395954 -17371 396022 -17315
rect 396078 -17371 396146 -17315
rect 396202 -17371 396270 -17315
rect 396326 -17371 396394 -17315
rect 396450 -17371 396518 -17315
rect 396574 -17371 396642 -17315
rect 396698 -17371 396766 -17315
rect 396822 -17371 396890 -17315
rect 396946 -17371 397014 -17315
rect 397070 -17371 397200 -17315
rect 388000 -17439 397200 -17371
rect 388000 -17495 388146 -17439
rect 388202 -17495 388270 -17439
rect 388326 -17495 388394 -17439
rect 388450 -17495 388518 -17439
rect 388574 -17495 388642 -17439
rect 388698 -17495 388766 -17439
rect 388822 -17495 388890 -17439
rect 388946 -17495 389014 -17439
rect 389070 -17495 389138 -17439
rect 389194 -17495 389262 -17439
rect 389318 -17495 389386 -17439
rect 389442 -17495 389510 -17439
rect 389566 -17495 389634 -17439
rect 389690 -17495 389758 -17439
rect 389814 -17495 389882 -17439
rect 389938 -17495 390006 -17439
rect 390062 -17495 390130 -17439
rect 390186 -17495 390254 -17439
rect 390310 -17495 390378 -17439
rect 390434 -17495 390502 -17439
rect 390558 -17495 390626 -17439
rect 390682 -17495 390750 -17439
rect 390806 -17495 390874 -17439
rect 390930 -17495 390998 -17439
rect 391054 -17495 391122 -17439
rect 391178 -17495 391246 -17439
rect 391302 -17495 391370 -17439
rect 391426 -17495 391494 -17439
rect 391550 -17495 391618 -17439
rect 391674 -17495 391742 -17439
rect 391798 -17495 391866 -17439
rect 391922 -17495 391990 -17439
rect 392046 -17495 392114 -17439
rect 392170 -17495 392238 -17439
rect 392294 -17495 392362 -17439
rect 392418 -17495 392486 -17439
rect 392542 -17495 392610 -17439
rect 392666 -17495 392734 -17439
rect 392790 -17495 392858 -17439
rect 392914 -17495 392982 -17439
rect 393038 -17495 393106 -17439
rect 393162 -17495 393230 -17439
rect 393286 -17495 393354 -17439
rect 393410 -17495 393478 -17439
rect 393534 -17495 393602 -17439
rect 393658 -17495 393726 -17439
rect 393782 -17495 393850 -17439
rect 393906 -17495 393974 -17439
rect 394030 -17495 394098 -17439
rect 394154 -17495 394222 -17439
rect 394278 -17495 394346 -17439
rect 394402 -17495 394470 -17439
rect 394526 -17495 394594 -17439
rect 394650 -17495 394718 -17439
rect 394774 -17495 394842 -17439
rect 394898 -17495 394966 -17439
rect 395022 -17495 395090 -17439
rect 395146 -17495 395214 -17439
rect 395270 -17495 395338 -17439
rect 395394 -17495 395462 -17439
rect 395518 -17495 395586 -17439
rect 395642 -17495 395710 -17439
rect 395766 -17495 395898 -17439
rect 395954 -17495 396022 -17439
rect 396078 -17495 396146 -17439
rect 396202 -17495 396270 -17439
rect 396326 -17495 396394 -17439
rect 396450 -17495 396518 -17439
rect 396574 -17495 396642 -17439
rect 396698 -17495 396766 -17439
rect 396822 -17495 396890 -17439
rect 396946 -17495 397014 -17439
rect 397070 -17495 397200 -17439
rect 388000 -17563 397200 -17495
rect 388000 -17619 388146 -17563
rect 388202 -17619 388270 -17563
rect 388326 -17619 388394 -17563
rect 388450 -17619 388518 -17563
rect 388574 -17619 388642 -17563
rect 388698 -17619 388766 -17563
rect 388822 -17619 388890 -17563
rect 388946 -17619 389014 -17563
rect 389070 -17619 389138 -17563
rect 389194 -17619 389262 -17563
rect 389318 -17619 389386 -17563
rect 389442 -17619 389510 -17563
rect 389566 -17619 389634 -17563
rect 389690 -17619 389758 -17563
rect 389814 -17619 389882 -17563
rect 389938 -17619 390006 -17563
rect 390062 -17619 390130 -17563
rect 390186 -17619 390254 -17563
rect 390310 -17619 390378 -17563
rect 390434 -17619 390502 -17563
rect 390558 -17619 390626 -17563
rect 390682 -17619 390750 -17563
rect 390806 -17619 390874 -17563
rect 390930 -17619 390998 -17563
rect 391054 -17619 391122 -17563
rect 391178 -17619 391246 -17563
rect 391302 -17619 391370 -17563
rect 391426 -17619 391494 -17563
rect 391550 -17619 391618 -17563
rect 391674 -17619 391742 -17563
rect 391798 -17619 391866 -17563
rect 391922 -17619 391990 -17563
rect 392046 -17619 392114 -17563
rect 392170 -17619 392238 -17563
rect 392294 -17619 392362 -17563
rect 392418 -17619 392486 -17563
rect 392542 -17619 392610 -17563
rect 392666 -17619 392734 -17563
rect 392790 -17619 392858 -17563
rect 392914 -17619 392982 -17563
rect 393038 -17619 393106 -17563
rect 393162 -17619 393230 -17563
rect 393286 -17619 393354 -17563
rect 393410 -17619 393478 -17563
rect 393534 -17619 393602 -17563
rect 393658 -17619 393726 -17563
rect 393782 -17619 393850 -17563
rect 393906 -17619 393974 -17563
rect 394030 -17619 394098 -17563
rect 394154 -17619 394222 -17563
rect 394278 -17619 394346 -17563
rect 394402 -17619 394470 -17563
rect 394526 -17619 394594 -17563
rect 394650 -17619 394718 -17563
rect 394774 -17619 394842 -17563
rect 394898 -17619 394966 -17563
rect 395022 -17619 395090 -17563
rect 395146 -17619 395214 -17563
rect 395270 -17619 395338 -17563
rect 395394 -17619 395462 -17563
rect 395518 -17619 395586 -17563
rect 395642 -17619 395710 -17563
rect 395766 -17619 395898 -17563
rect 395954 -17619 396022 -17563
rect 396078 -17619 396146 -17563
rect 396202 -17619 396270 -17563
rect 396326 -17619 396394 -17563
rect 396450 -17619 396518 -17563
rect 396574 -17619 396642 -17563
rect 396698 -17619 396766 -17563
rect 396822 -17619 396890 -17563
rect 396946 -17619 397014 -17563
rect 397070 -17619 397200 -17563
rect 388000 -17820 397200 -17619
rect 388000 -17858 388800 -17820
rect 388000 -17914 388114 -17858
rect 388170 -17914 388238 -17858
rect 388294 -17914 388362 -17858
rect 388418 -17914 388486 -17858
rect 388542 -17914 388610 -17858
rect 388666 -17914 388800 -17858
rect 388000 -17982 388800 -17914
rect 388000 -18038 388114 -17982
rect 388170 -18038 388238 -17982
rect 388294 -18038 388362 -17982
rect 388418 -18038 388486 -17982
rect 388542 -18038 388610 -17982
rect 388666 -18038 388800 -17982
rect 388000 -18106 388800 -18038
rect 388000 -18162 388114 -18106
rect 388170 -18162 388238 -18106
rect 388294 -18162 388362 -18106
rect 388418 -18162 388486 -18106
rect 388542 -18162 388610 -18106
rect 388666 -18162 388800 -18106
rect 388000 -18230 388800 -18162
rect 388000 -18286 388114 -18230
rect 388170 -18286 388238 -18230
rect 388294 -18286 388362 -18230
rect 388418 -18286 388486 -18230
rect 388542 -18286 388610 -18230
rect 388666 -18286 388800 -18230
rect 388000 -18354 388800 -18286
rect 388000 -18410 388114 -18354
rect 388170 -18410 388238 -18354
rect 388294 -18410 388362 -18354
rect 388418 -18410 388486 -18354
rect 388542 -18410 388610 -18354
rect 388666 -18410 388800 -18354
rect 388000 -18478 388800 -18410
rect 388000 -18534 388114 -18478
rect 388170 -18534 388238 -18478
rect 388294 -18534 388362 -18478
rect 388418 -18534 388486 -18478
rect 388542 -18534 388610 -18478
rect 388666 -18534 388800 -18478
rect 388000 -18602 388800 -18534
rect 388000 -18658 388114 -18602
rect 388170 -18658 388238 -18602
rect 388294 -18658 388362 -18602
rect 388418 -18658 388486 -18602
rect 388542 -18658 388610 -18602
rect 388666 -18658 388800 -18602
rect 388000 -18726 388800 -18658
rect 388000 -18782 388114 -18726
rect 388170 -18782 388238 -18726
rect 388294 -18782 388362 -18726
rect 388418 -18782 388486 -18726
rect 388542 -18782 388610 -18726
rect 388666 -18782 388800 -18726
rect 388000 -18850 388800 -18782
rect 388000 -18906 388114 -18850
rect 388170 -18906 388238 -18850
rect 388294 -18906 388362 -18850
rect 388418 -18906 388486 -18850
rect 388542 -18906 388610 -18850
rect 388666 -18906 388800 -18850
rect 388000 -18974 388800 -18906
rect 388000 -19030 388114 -18974
rect 388170 -19030 388238 -18974
rect 388294 -19030 388362 -18974
rect 388418 -19030 388486 -18974
rect 388542 -19030 388610 -18974
rect 388666 -19030 388800 -18974
rect 388000 -19098 388800 -19030
rect 388000 -19154 388114 -19098
rect 388170 -19154 388238 -19098
rect 388294 -19154 388362 -19098
rect 388418 -19154 388486 -19098
rect 388542 -19154 388610 -19098
rect 388666 -19154 388800 -19098
rect 388000 -19222 388800 -19154
rect 388000 -19278 388114 -19222
rect 388170 -19278 388238 -19222
rect 388294 -19278 388362 -19222
rect 388418 -19278 388486 -19222
rect 388542 -19278 388610 -19222
rect 388666 -19278 388800 -19222
rect 388000 -19346 388800 -19278
rect 388000 -19402 388114 -19346
rect 388170 -19402 388238 -19346
rect 388294 -19402 388362 -19346
rect 388418 -19402 388486 -19346
rect 388542 -19402 388610 -19346
rect 388666 -19402 388800 -19346
rect 388000 -19470 388800 -19402
rect 388000 -19526 388114 -19470
rect 388170 -19526 388238 -19470
rect 388294 -19526 388362 -19470
rect 388418 -19526 388486 -19470
rect 388542 -19526 388610 -19470
rect 388666 -19526 388800 -19470
rect 388000 -19594 388800 -19526
rect 388000 -19650 388114 -19594
rect 388170 -19650 388238 -19594
rect 388294 -19650 388362 -19594
rect 388418 -19650 388486 -19594
rect 388542 -19650 388610 -19594
rect 388666 -19650 388800 -19594
rect 388000 -19718 388800 -19650
rect 388000 -19774 388114 -19718
rect 388170 -19774 388238 -19718
rect 388294 -19774 388362 -19718
rect 388418 -19774 388486 -19718
rect 388542 -19774 388610 -19718
rect 388666 -19774 388800 -19718
rect 388000 -19842 388800 -19774
rect 388000 -19898 388114 -19842
rect 388170 -19898 388238 -19842
rect 388294 -19898 388362 -19842
rect 388418 -19898 388486 -19842
rect 388542 -19898 388610 -19842
rect 388666 -19898 388800 -19842
rect 388000 -19966 388800 -19898
rect 388000 -20022 388114 -19966
rect 388170 -20022 388238 -19966
rect 388294 -20022 388362 -19966
rect 388418 -20022 388486 -19966
rect 388542 -20022 388610 -19966
rect 388666 -20022 388800 -19966
rect 388000 -20090 388800 -20022
rect 388000 -20146 388114 -20090
rect 388170 -20146 388238 -20090
rect 388294 -20146 388362 -20090
rect 388418 -20146 388486 -20090
rect 388542 -20146 388610 -20090
rect 388666 -20146 388800 -20090
rect 388000 -20214 388800 -20146
rect 388000 -20270 388114 -20214
rect 388170 -20270 388238 -20214
rect 388294 -20270 388362 -20214
rect 388418 -20270 388486 -20214
rect 388542 -20270 388610 -20214
rect 388666 -20270 388800 -20214
rect 388000 -20338 388800 -20270
rect 388000 -20394 388114 -20338
rect 388170 -20394 388238 -20338
rect 388294 -20394 388362 -20338
rect 388418 -20394 388486 -20338
rect 388542 -20394 388610 -20338
rect 388666 -20394 388800 -20338
rect 388000 -20462 388800 -20394
rect 388000 -20518 388114 -20462
rect 388170 -20518 388238 -20462
rect 388294 -20518 388362 -20462
rect 388418 -20518 388486 -20462
rect 388542 -20518 388610 -20462
rect 388666 -20518 388800 -20462
rect 388000 -20586 388800 -20518
rect 388000 -20642 388114 -20586
rect 388170 -20642 388238 -20586
rect 388294 -20642 388362 -20586
rect 388418 -20642 388486 -20586
rect 388542 -20642 388610 -20586
rect 388666 -20642 388800 -20586
rect 388000 -20710 388800 -20642
rect 388000 -20766 388114 -20710
rect 388170 -20766 388238 -20710
rect 388294 -20766 388362 -20710
rect 388418 -20766 388486 -20710
rect 388542 -20766 388610 -20710
rect 388666 -20766 388800 -20710
rect 388000 -20834 388800 -20766
rect 388000 -20890 388114 -20834
rect 388170 -20890 388238 -20834
rect 388294 -20890 388362 -20834
rect 388418 -20890 388486 -20834
rect 388542 -20890 388610 -20834
rect 388666 -20890 388800 -20834
rect 388000 -20958 388800 -20890
rect 388000 -21014 388114 -20958
rect 388170 -21014 388238 -20958
rect 388294 -21014 388362 -20958
rect 388418 -21014 388486 -20958
rect 388542 -21014 388610 -20958
rect 388666 -21014 388800 -20958
rect 388000 -21082 388800 -21014
rect 388000 -21138 388114 -21082
rect 388170 -21138 388238 -21082
rect 388294 -21138 388362 -21082
rect 388418 -21138 388486 -21082
rect 388542 -21138 388610 -21082
rect 388666 -21138 388800 -21082
rect 388000 -21206 388800 -21138
rect 388000 -21262 388114 -21206
rect 388170 -21262 388238 -21206
rect 388294 -21262 388362 -21206
rect 388418 -21262 388486 -21206
rect 388542 -21262 388610 -21206
rect 388666 -21262 388800 -21206
rect 388000 -21330 388800 -21262
rect 388000 -21386 388114 -21330
rect 388170 -21386 388238 -21330
rect 388294 -21386 388362 -21330
rect 388418 -21386 388486 -21330
rect 388542 -21386 388610 -21330
rect 388666 -21386 388800 -21330
rect 388000 -21454 388800 -21386
rect 388000 -21510 388114 -21454
rect 388170 -21510 388238 -21454
rect 388294 -21510 388362 -21454
rect 388418 -21510 388486 -21454
rect 388542 -21510 388610 -21454
rect 388666 -21510 388800 -21454
rect 388000 -21578 388800 -21510
rect 388000 -21634 388114 -21578
rect 388170 -21634 388238 -21578
rect 388294 -21634 388362 -21578
rect 388418 -21634 388486 -21578
rect 388542 -21634 388610 -21578
rect 388666 -21634 388800 -21578
rect 388000 -21702 388800 -21634
rect 388000 -21758 388114 -21702
rect 388170 -21758 388238 -21702
rect 388294 -21758 388362 -21702
rect 388418 -21758 388486 -21702
rect 388542 -21758 388610 -21702
rect 388666 -21758 388800 -21702
rect 388000 -21826 388800 -21758
rect 388000 -21882 388114 -21826
rect 388170 -21882 388238 -21826
rect 388294 -21882 388362 -21826
rect 388418 -21882 388486 -21826
rect 388542 -21882 388610 -21826
rect 388666 -21882 388800 -21826
rect 388000 -21950 388800 -21882
rect 388000 -22006 388114 -21950
rect 388170 -22006 388238 -21950
rect 388294 -22006 388362 -21950
rect 388418 -22006 388486 -21950
rect 388542 -22006 388610 -21950
rect 388666 -22006 388800 -21950
rect 388000 -22074 388800 -22006
rect 388000 -22130 388114 -22074
rect 388170 -22130 388238 -22074
rect 388294 -22130 388362 -22074
rect 388418 -22130 388486 -22074
rect 388542 -22130 388610 -22074
rect 388666 -22130 388800 -22074
rect 388000 -22198 388800 -22130
rect 388000 -22254 388114 -22198
rect 388170 -22254 388238 -22198
rect 388294 -22254 388362 -22198
rect 388418 -22254 388486 -22198
rect 388542 -22254 388610 -22198
rect 388666 -22254 388800 -22198
rect 388000 -22322 388800 -22254
rect 388000 -22378 388114 -22322
rect 388170 -22378 388238 -22322
rect 388294 -22378 388362 -22322
rect 388418 -22378 388486 -22322
rect 388542 -22378 388610 -22322
rect 388666 -22378 388800 -22322
rect 388000 -22446 388800 -22378
rect 388000 -22502 388114 -22446
rect 388170 -22502 388238 -22446
rect 388294 -22502 388362 -22446
rect 388418 -22502 388486 -22446
rect 388542 -22502 388610 -22446
rect 388666 -22502 388800 -22446
rect 388000 -22570 388800 -22502
rect 388000 -22626 388114 -22570
rect 388170 -22626 388238 -22570
rect 388294 -22626 388362 -22570
rect 388418 -22626 388486 -22570
rect 388542 -22626 388610 -22570
rect 388666 -22626 388800 -22570
rect 388000 -22694 388800 -22626
rect 388000 -22750 388114 -22694
rect 388170 -22750 388238 -22694
rect 388294 -22750 388362 -22694
rect 388418 -22750 388486 -22694
rect 388542 -22750 388610 -22694
rect 388666 -22750 388800 -22694
rect 388000 -22818 388800 -22750
rect 388000 -22874 388114 -22818
rect 388170 -22874 388238 -22818
rect 388294 -22874 388362 -22818
rect 388418 -22874 388486 -22818
rect 388542 -22874 388610 -22818
rect 388666 -22874 388800 -22818
rect 388000 -22942 388800 -22874
rect 388000 -22998 388114 -22942
rect 388170 -22998 388238 -22942
rect 388294 -22998 388362 -22942
rect 388418 -22998 388486 -22942
rect 388542 -22998 388610 -22942
rect 388666 -22998 388800 -22942
rect 388000 -23066 388800 -22998
rect 388000 -23122 388114 -23066
rect 388170 -23122 388238 -23066
rect 388294 -23122 388362 -23066
rect 388418 -23122 388486 -23066
rect 388542 -23122 388610 -23066
rect 388666 -23122 388800 -23066
rect 388000 -23190 388800 -23122
rect 388000 -23246 388114 -23190
rect 388170 -23246 388238 -23190
rect 388294 -23246 388362 -23190
rect 388418 -23246 388486 -23190
rect 388542 -23246 388610 -23190
rect 388666 -23246 388800 -23190
rect 388000 -23314 388800 -23246
rect 388000 -23370 388114 -23314
rect 388170 -23370 388238 -23314
rect 388294 -23370 388362 -23314
rect 388418 -23370 388486 -23314
rect 388542 -23370 388610 -23314
rect 388666 -23370 388800 -23314
rect 388000 -23438 388800 -23370
rect 388000 -23494 388114 -23438
rect 388170 -23494 388238 -23438
rect 388294 -23494 388362 -23438
rect 388418 -23494 388486 -23438
rect 388542 -23494 388610 -23438
rect 388666 -23494 388800 -23438
rect 388000 -23562 388800 -23494
rect 388000 -23618 388114 -23562
rect 388170 -23618 388238 -23562
rect 388294 -23618 388362 -23562
rect 388418 -23618 388486 -23562
rect 388542 -23618 388610 -23562
rect 388666 -23618 388800 -23562
rect 388000 -23686 388800 -23618
rect 388000 -23742 388114 -23686
rect 388170 -23742 388238 -23686
rect 388294 -23742 388362 -23686
rect 388418 -23742 388486 -23686
rect 388542 -23742 388610 -23686
rect 388666 -23742 388800 -23686
rect 388000 -23810 388800 -23742
rect 388000 -23866 388114 -23810
rect 388170 -23866 388238 -23810
rect 388294 -23866 388362 -23810
rect 388418 -23866 388486 -23810
rect 388542 -23866 388610 -23810
rect 388666 -23866 388800 -23810
rect 388000 -23934 388800 -23866
rect 388000 -23990 388114 -23934
rect 388170 -23990 388238 -23934
rect 388294 -23990 388362 -23934
rect 388418 -23990 388486 -23934
rect 388542 -23990 388610 -23934
rect 388666 -23990 388800 -23934
rect 388000 -24058 388800 -23990
rect 388000 -24114 388114 -24058
rect 388170 -24114 388238 -24058
rect 388294 -24114 388362 -24058
rect 388418 -24114 388486 -24058
rect 388542 -24114 388610 -24058
rect 388666 -24114 388800 -24058
rect 388000 -24182 388800 -24114
rect 388000 -24238 388114 -24182
rect 388170 -24238 388238 -24182
rect 388294 -24238 388362 -24182
rect 388418 -24238 388486 -24182
rect 388542 -24238 388610 -24182
rect 388666 -24238 388800 -24182
rect 388000 -24306 388800 -24238
rect 388000 -24362 388114 -24306
rect 388170 -24362 388238 -24306
rect 388294 -24362 388362 -24306
rect 388418 -24362 388486 -24306
rect 388542 -24362 388610 -24306
rect 388666 -24362 388800 -24306
rect 388000 -24430 388800 -24362
rect 388000 -24486 388114 -24430
rect 388170 -24486 388238 -24430
rect 388294 -24486 388362 -24430
rect 388418 -24486 388486 -24430
rect 388542 -24486 388610 -24430
rect 388666 -24486 388800 -24430
rect 388000 -24554 388800 -24486
rect 388000 -24610 388114 -24554
rect 388170 -24610 388238 -24554
rect 388294 -24610 388362 -24554
rect 388418 -24610 388486 -24554
rect 388542 -24610 388610 -24554
rect 388666 -24610 388800 -24554
rect 388000 -24678 388800 -24610
rect 388000 -24734 388114 -24678
rect 388170 -24734 388238 -24678
rect 388294 -24734 388362 -24678
rect 388418 -24734 388486 -24678
rect 388542 -24734 388610 -24678
rect 388666 -24734 388800 -24678
rect 388000 -24802 388800 -24734
rect 388000 -24858 388114 -24802
rect 388170 -24858 388238 -24802
rect 388294 -24858 388362 -24802
rect 388418 -24858 388486 -24802
rect 388542 -24858 388610 -24802
rect 388666 -24858 388800 -24802
rect 388000 -24926 388800 -24858
rect 388000 -24982 388114 -24926
rect 388170 -24982 388238 -24926
rect 388294 -24982 388362 -24926
rect 388418 -24982 388486 -24926
rect 388542 -24982 388610 -24926
rect 388666 -24982 388800 -24926
rect 388000 -25050 388800 -24982
rect 388000 -25106 388114 -25050
rect 388170 -25106 388238 -25050
rect 388294 -25106 388362 -25050
rect 388418 -25106 388486 -25050
rect 388542 -25106 388610 -25050
rect 388666 -25106 388800 -25050
rect 388000 -25174 388800 -25106
rect 388000 -25230 388114 -25174
rect 388170 -25230 388238 -25174
rect 388294 -25230 388362 -25174
rect 388418 -25230 388486 -25174
rect 388542 -25230 388610 -25174
rect 388666 -25230 388800 -25174
rect 388000 -25298 388800 -25230
rect 388000 -25354 388114 -25298
rect 388170 -25354 388238 -25298
rect 388294 -25354 388362 -25298
rect 388418 -25354 388486 -25298
rect 388542 -25354 388610 -25298
rect 388666 -25354 388800 -25298
rect 388000 -25422 388800 -25354
rect 388000 -25478 388114 -25422
rect 388170 -25478 388238 -25422
rect 388294 -25478 388362 -25422
rect 388418 -25478 388486 -25422
rect 388542 -25478 388610 -25422
rect 388666 -25478 388800 -25422
rect 388000 -25542 388800 -25478
rect 389068 -17950 389408 -17820
rect 389068 -18006 389141 -17950
rect 389197 -18006 389283 -17950
rect 389339 -18006 389408 -17950
rect 389068 -18092 389408 -18006
rect 389068 -18148 389141 -18092
rect 389197 -18148 389283 -18092
rect 389339 -18148 389408 -18092
rect 389068 -18234 389408 -18148
rect 389068 -18290 389141 -18234
rect 389197 -18290 389283 -18234
rect 389339 -18290 389408 -18234
rect 389068 -18376 389408 -18290
rect 389068 -18432 389141 -18376
rect 389197 -18432 389283 -18376
rect 389339 -18432 389408 -18376
rect 389068 -18518 389408 -18432
rect 389068 -18574 389141 -18518
rect 389197 -18574 389283 -18518
rect 389339 -18574 389408 -18518
rect 389068 -18660 389408 -18574
rect 389068 -18716 389141 -18660
rect 389197 -18716 389283 -18660
rect 389339 -18716 389408 -18660
rect 389068 -18802 389408 -18716
rect 389068 -18858 389141 -18802
rect 389197 -18858 389283 -18802
rect 389339 -18858 389408 -18802
rect 389068 -18944 389408 -18858
rect 389068 -19000 389141 -18944
rect 389197 -19000 389283 -18944
rect 389339 -19000 389408 -18944
rect 389068 -19086 389408 -19000
rect 389068 -19142 389141 -19086
rect 389197 -19142 389283 -19086
rect 389339 -19142 389408 -19086
rect 389068 -19228 389408 -19142
rect 389068 -19284 389141 -19228
rect 389197 -19284 389283 -19228
rect 389339 -19284 389408 -19228
rect 389068 -19370 389408 -19284
rect 389068 -19426 389141 -19370
rect 389197 -19426 389283 -19370
rect 389339 -19426 389408 -19370
rect 389068 -19512 389408 -19426
rect 389068 -19568 389141 -19512
rect 389197 -19568 389283 -19512
rect 389339 -19568 389408 -19512
rect 389068 -19654 389408 -19568
rect 389068 -19710 389141 -19654
rect 389197 -19710 389283 -19654
rect 389339 -19710 389408 -19654
rect 389068 -19796 389408 -19710
rect 389068 -19852 389141 -19796
rect 389197 -19852 389283 -19796
rect 389339 -19852 389408 -19796
rect 389068 -19938 389408 -19852
rect 389068 -19994 389141 -19938
rect 389197 -19994 389283 -19938
rect 389339 -19994 389408 -19938
rect 389068 -20080 389408 -19994
rect 389068 -20136 389141 -20080
rect 389197 -20136 389283 -20080
rect 389339 -20136 389408 -20080
rect 389068 -20222 389408 -20136
rect 389068 -20278 389141 -20222
rect 389197 -20278 389283 -20222
rect 389339 -20278 389408 -20222
rect 389068 -20364 389408 -20278
rect 389068 -20420 389141 -20364
rect 389197 -20420 389283 -20364
rect 389339 -20420 389408 -20364
rect 389068 -20506 389408 -20420
rect 389068 -20562 389141 -20506
rect 389197 -20562 389283 -20506
rect 389339 -20562 389408 -20506
rect 389068 -20648 389408 -20562
rect 389068 -20704 389141 -20648
rect 389197 -20704 389283 -20648
rect 389339 -20704 389408 -20648
rect 389068 -20790 389408 -20704
rect 389068 -20846 389141 -20790
rect 389197 -20846 389283 -20790
rect 389339 -20846 389408 -20790
rect 389068 -20932 389408 -20846
rect 389068 -20988 389141 -20932
rect 389197 -20988 389283 -20932
rect 389339 -20988 389408 -20932
rect 389068 -21074 389408 -20988
rect 389068 -21130 389141 -21074
rect 389197 -21130 389283 -21074
rect 389339 -21130 389408 -21074
rect 389068 -21216 389408 -21130
rect 389068 -21272 389141 -21216
rect 389197 -21272 389283 -21216
rect 389339 -21272 389408 -21216
rect 389068 -21358 389408 -21272
rect 389068 -21414 389141 -21358
rect 389197 -21414 389283 -21358
rect 389339 -21414 389408 -21358
rect 389068 -21500 389408 -21414
rect 389068 -21556 389141 -21500
rect 389197 -21556 389283 -21500
rect 389339 -21556 389408 -21500
rect 389068 -21642 389408 -21556
rect 389068 -21698 389141 -21642
rect 389197 -21698 389283 -21642
rect 389339 -21698 389408 -21642
rect 389068 -21784 389408 -21698
rect 389068 -21840 389141 -21784
rect 389197 -21840 389283 -21784
rect 389339 -21840 389408 -21784
rect 389068 -21926 389408 -21840
rect 389068 -21982 389141 -21926
rect 389197 -21982 389283 -21926
rect 389339 -21982 389408 -21926
rect 389068 -22068 389408 -21982
rect 389068 -22124 389141 -22068
rect 389197 -22124 389283 -22068
rect 389339 -22124 389408 -22068
rect 389068 -22210 389408 -22124
rect 389068 -22266 389141 -22210
rect 389197 -22266 389283 -22210
rect 389339 -22266 389408 -22210
rect 389068 -22352 389408 -22266
rect 389068 -22408 389141 -22352
rect 389197 -22408 389283 -22352
rect 389339 -22408 389408 -22352
rect 389068 -22494 389408 -22408
rect 389068 -22550 389141 -22494
rect 389197 -22550 389283 -22494
rect 389339 -22550 389408 -22494
rect 389068 -22636 389408 -22550
rect 389068 -22692 389141 -22636
rect 389197 -22692 389283 -22636
rect 389339 -22692 389408 -22636
rect 389068 -22778 389408 -22692
rect 389068 -22834 389141 -22778
rect 389197 -22834 389283 -22778
rect 389339 -22834 389408 -22778
rect 389068 -22920 389408 -22834
rect 389068 -22976 389141 -22920
rect 389197 -22976 389283 -22920
rect 389339 -22976 389408 -22920
rect 389068 -23062 389408 -22976
rect 389068 -23118 389141 -23062
rect 389197 -23118 389283 -23062
rect 389339 -23118 389408 -23062
rect 389068 -23204 389408 -23118
rect 389068 -23260 389141 -23204
rect 389197 -23260 389283 -23204
rect 389339 -23260 389408 -23204
rect 389068 -23346 389408 -23260
rect 389068 -23402 389141 -23346
rect 389197 -23402 389283 -23346
rect 389339 -23402 389408 -23346
rect 389068 -23488 389408 -23402
rect 389068 -23544 389141 -23488
rect 389197 -23544 389283 -23488
rect 389339 -23544 389408 -23488
rect 389068 -23630 389408 -23544
rect 389068 -23686 389141 -23630
rect 389197 -23686 389283 -23630
rect 389339 -23686 389408 -23630
rect 389068 -23772 389408 -23686
rect 389068 -23828 389141 -23772
rect 389197 -23828 389283 -23772
rect 389339 -23828 389408 -23772
rect 389068 -23914 389408 -23828
rect 389068 -23970 389141 -23914
rect 389197 -23970 389283 -23914
rect 389339 -23970 389408 -23914
rect 389068 -24056 389408 -23970
rect 389068 -24112 389141 -24056
rect 389197 -24112 389283 -24056
rect 389339 -24112 389408 -24056
rect 389068 -24198 389408 -24112
rect 389068 -24254 389141 -24198
rect 389197 -24254 389283 -24198
rect 389339 -24254 389408 -24198
rect 389068 -24340 389408 -24254
rect 389068 -24396 389141 -24340
rect 389197 -24396 389283 -24340
rect 389339 -24396 389408 -24340
rect 389068 -24482 389408 -24396
rect 389068 -24538 389141 -24482
rect 389197 -24538 389283 -24482
rect 389339 -24538 389408 -24482
rect 389068 -24624 389408 -24538
rect 389068 -24680 389141 -24624
rect 389197 -24680 389283 -24624
rect 389339 -24680 389408 -24624
rect 389068 -24766 389408 -24680
rect 389068 -24822 389141 -24766
rect 389197 -24822 389283 -24766
rect 389339 -24822 389408 -24766
rect 389068 -24908 389408 -24822
rect 389068 -24964 389141 -24908
rect 389197 -24964 389283 -24908
rect 389339 -24964 389408 -24908
rect 389068 -25050 389408 -24964
rect 389068 -25106 389141 -25050
rect 389197 -25106 389283 -25050
rect 389339 -25106 389408 -25050
rect 389068 -25192 389408 -25106
rect 389068 -25248 389141 -25192
rect 389197 -25248 389283 -25192
rect 389339 -25248 389408 -25192
rect 389068 -25334 389408 -25248
rect 389068 -25390 389141 -25334
rect 389197 -25390 389283 -25334
rect 389339 -25390 389408 -25334
rect 389068 -25476 389408 -25390
rect 389068 -25532 389141 -25476
rect 389197 -25532 389283 -25476
rect 389339 -25532 389408 -25476
rect 389068 -25542 389408 -25532
rect 389468 -17950 389808 -17820
rect 389468 -18006 389542 -17950
rect 389598 -18006 389684 -17950
rect 389740 -18006 389808 -17950
rect 389468 -18092 389808 -18006
rect 389468 -18148 389542 -18092
rect 389598 -18148 389684 -18092
rect 389740 -18148 389808 -18092
rect 389468 -18234 389808 -18148
rect 389468 -18290 389542 -18234
rect 389598 -18290 389684 -18234
rect 389740 -18290 389808 -18234
rect 389468 -18376 389808 -18290
rect 389468 -18432 389542 -18376
rect 389598 -18432 389684 -18376
rect 389740 -18432 389808 -18376
rect 389468 -18518 389808 -18432
rect 389468 -18574 389542 -18518
rect 389598 -18574 389684 -18518
rect 389740 -18574 389808 -18518
rect 389468 -18660 389808 -18574
rect 389468 -18716 389542 -18660
rect 389598 -18716 389684 -18660
rect 389740 -18716 389808 -18660
rect 389468 -18802 389808 -18716
rect 389468 -18858 389542 -18802
rect 389598 -18858 389684 -18802
rect 389740 -18858 389808 -18802
rect 389468 -18944 389808 -18858
rect 389468 -19000 389542 -18944
rect 389598 -19000 389684 -18944
rect 389740 -19000 389808 -18944
rect 389468 -19086 389808 -19000
rect 389468 -19142 389542 -19086
rect 389598 -19142 389684 -19086
rect 389740 -19142 389808 -19086
rect 389468 -19228 389808 -19142
rect 389468 -19284 389542 -19228
rect 389598 -19284 389684 -19228
rect 389740 -19284 389808 -19228
rect 389468 -19370 389808 -19284
rect 389468 -19426 389542 -19370
rect 389598 -19426 389684 -19370
rect 389740 -19426 389808 -19370
rect 389468 -19512 389808 -19426
rect 389468 -19568 389542 -19512
rect 389598 -19568 389684 -19512
rect 389740 -19568 389808 -19512
rect 389468 -19654 389808 -19568
rect 389468 -19710 389542 -19654
rect 389598 -19710 389684 -19654
rect 389740 -19710 389808 -19654
rect 389468 -19796 389808 -19710
rect 389468 -19852 389542 -19796
rect 389598 -19852 389684 -19796
rect 389740 -19852 389808 -19796
rect 389468 -19938 389808 -19852
rect 389468 -19994 389542 -19938
rect 389598 -19994 389684 -19938
rect 389740 -19994 389808 -19938
rect 389468 -20080 389808 -19994
rect 389468 -20136 389542 -20080
rect 389598 -20136 389684 -20080
rect 389740 -20136 389808 -20080
rect 389468 -20222 389808 -20136
rect 389468 -20278 389542 -20222
rect 389598 -20278 389684 -20222
rect 389740 -20278 389808 -20222
rect 389468 -20364 389808 -20278
rect 389468 -20420 389542 -20364
rect 389598 -20420 389684 -20364
rect 389740 -20420 389808 -20364
rect 389468 -20506 389808 -20420
rect 389468 -20562 389542 -20506
rect 389598 -20562 389684 -20506
rect 389740 -20562 389808 -20506
rect 389468 -20648 389808 -20562
rect 389468 -20704 389542 -20648
rect 389598 -20704 389684 -20648
rect 389740 -20704 389808 -20648
rect 389468 -20790 389808 -20704
rect 389468 -20846 389542 -20790
rect 389598 -20846 389684 -20790
rect 389740 -20846 389808 -20790
rect 389468 -20932 389808 -20846
rect 389468 -20988 389542 -20932
rect 389598 -20988 389684 -20932
rect 389740 -20988 389808 -20932
rect 389468 -21074 389808 -20988
rect 389468 -21130 389542 -21074
rect 389598 -21130 389684 -21074
rect 389740 -21130 389808 -21074
rect 389468 -21216 389808 -21130
rect 389468 -21272 389542 -21216
rect 389598 -21272 389684 -21216
rect 389740 -21272 389808 -21216
rect 389468 -21358 389808 -21272
rect 389468 -21414 389542 -21358
rect 389598 -21414 389684 -21358
rect 389740 -21414 389808 -21358
rect 389468 -21500 389808 -21414
rect 389468 -21556 389542 -21500
rect 389598 -21556 389684 -21500
rect 389740 -21556 389808 -21500
rect 389468 -21642 389808 -21556
rect 389468 -21698 389542 -21642
rect 389598 -21698 389684 -21642
rect 389740 -21698 389808 -21642
rect 389468 -21784 389808 -21698
rect 389468 -21840 389542 -21784
rect 389598 -21840 389684 -21784
rect 389740 -21840 389808 -21784
rect 389468 -21926 389808 -21840
rect 389468 -21982 389542 -21926
rect 389598 -21982 389684 -21926
rect 389740 -21982 389808 -21926
rect 389468 -22068 389808 -21982
rect 389468 -22124 389542 -22068
rect 389598 -22124 389684 -22068
rect 389740 -22124 389808 -22068
rect 389468 -22210 389808 -22124
rect 389468 -22266 389542 -22210
rect 389598 -22266 389684 -22210
rect 389740 -22266 389808 -22210
rect 389468 -22352 389808 -22266
rect 389468 -22408 389542 -22352
rect 389598 -22408 389684 -22352
rect 389740 -22408 389808 -22352
rect 389468 -22494 389808 -22408
rect 389468 -22550 389542 -22494
rect 389598 -22550 389684 -22494
rect 389740 -22550 389808 -22494
rect 389468 -22636 389808 -22550
rect 389468 -22692 389542 -22636
rect 389598 -22692 389684 -22636
rect 389740 -22692 389808 -22636
rect 389468 -22778 389808 -22692
rect 389468 -22834 389542 -22778
rect 389598 -22834 389684 -22778
rect 389740 -22834 389808 -22778
rect 389468 -22920 389808 -22834
rect 389468 -22976 389542 -22920
rect 389598 -22976 389684 -22920
rect 389740 -22976 389808 -22920
rect 389468 -23062 389808 -22976
rect 389468 -23118 389542 -23062
rect 389598 -23118 389684 -23062
rect 389740 -23118 389808 -23062
rect 389468 -23204 389808 -23118
rect 389468 -23260 389542 -23204
rect 389598 -23260 389684 -23204
rect 389740 -23260 389808 -23204
rect 389468 -23346 389808 -23260
rect 389468 -23402 389542 -23346
rect 389598 -23402 389684 -23346
rect 389740 -23402 389808 -23346
rect 389468 -23488 389808 -23402
rect 389468 -23544 389542 -23488
rect 389598 -23544 389684 -23488
rect 389740 -23544 389808 -23488
rect 389468 -23630 389808 -23544
rect 389468 -23686 389542 -23630
rect 389598 -23686 389684 -23630
rect 389740 -23686 389808 -23630
rect 389468 -23772 389808 -23686
rect 389468 -23828 389542 -23772
rect 389598 -23828 389684 -23772
rect 389740 -23828 389808 -23772
rect 389468 -23914 389808 -23828
rect 389468 -23970 389542 -23914
rect 389598 -23970 389684 -23914
rect 389740 -23970 389808 -23914
rect 389468 -24056 389808 -23970
rect 389468 -24112 389542 -24056
rect 389598 -24112 389684 -24056
rect 389740 -24112 389808 -24056
rect 389468 -24198 389808 -24112
rect 389468 -24254 389542 -24198
rect 389598 -24254 389684 -24198
rect 389740 -24254 389808 -24198
rect 389468 -24340 389808 -24254
rect 389468 -24396 389542 -24340
rect 389598 -24396 389684 -24340
rect 389740 -24396 389808 -24340
rect 389468 -24482 389808 -24396
rect 389468 -24538 389542 -24482
rect 389598 -24538 389684 -24482
rect 389740 -24538 389808 -24482
rect 389468 -24624 389808 -24538
rect 389468 -24680 389542 -24624
rect 389598 -24680 389684 -24624
rect 389740 -24680 389808 -24624
rect 389468 -24766 389808 -24680
rect 389468 -24822 389542 -24766
rect 389598 -24822 389684 -24766
rect 389740 -24822 389808 -24766
rect 389468 -24908 389808 -24822
rect 389468 -24964 389542 -24908
rect 389598 -24964 389684 -24908
rect 389740 -24964 389808 -24908
rect 389468 -25050 389808 -24964
rect 389468 -25106 389542 -25050
rect 389598 -25106 389684 -25050
rect 389740 -25106 389808 -25050
rect 389468 -25192 389808 -25106
rect 389468 -25248 389542 -25192
rect 389598 -25248 389684 -25192
rect 389740 -25248 389808 -25192
rect 389468 -25334 389808 -25248
rect 389468 -25390 389542 -25334
rect 389598 -25390 389684 -25334
rect 389740 -25390 389808 -25334
rect 389468 -25476 389808 -25390
rect 389468 -25532 389542 -25476
rect 389598 -25532 389684 -25476
rect 389740 -25532 389808 -25476
rect 389468 -25542 389808 -25532
rect 389868 -17950 390208 -17820
rect 389868 -18006 389942 -17950
rect 389998 -18006 390084 -17950
rect 390140 -18006 390208 -17950
rect 389868 -18092 390208 -18006
rect 389868 -18148 389942 -18092
rect 389998 -18148 390084 -18092
rect 390140 -18148 390208 -18092
rect 389868 -18234 390208 -18148
rect 389868 -18290 389942 -18234
rect 389998 -18290 390084 -18234
rect 390140 -18290 390208 -18234
rect 389868 -18376 390208 -18290
rect 389868 -18432 389942 -18376
rect 389998 -18432 390084 -18376
rect 390140 -18432 390208 -18376
rect 389868 -18518 390208 -18432
rect 389868 -18574 389942 -18518
rect 389998 -18574 390084 -18518
rect 390140 -18574 390208 -18518
rect 389868 -18660 390208 -18574
rect 389868 -18716 389942 -18660
rect 389998 -18716 390084 -18660
rect 390140 -18716 390208 -18660
rect 389868 -18802 390208 -18716
rect 389868 -18858 389942 -18802
rect 389998 -18858 390084 -18802
rect 390140 -18858 390208 -18802
rect 389868 -18944 390208 -18858
rect 389868 -19000 389942 -18944
rect 389998 -19000 390084 -18944
rect 390140 -19000 390208 -18944
rect 389868 -19086 390208 -19000
rect 389868 -19142 389942 -19086
rect 389998 -19142 390084 -19086
rect 390140 -19142 390208 -19086
rect 389868 -19228 390208 -19142
rect 389868 -19284 389942 -19228
rect 389998 -19284 390084 -19228
rect 390140 -19284 390208 -19228
rect 389868 -19370 390208 -19284
rect 389868 -19426 389942 -19370
rect 389998 -19426 390084 -19370
rect 390140 -19426 390208 -19370
rect 389868 -19512 390208 -19426
rect 389868 -19568 389942 -19512
rect 389998 -19568 390084 -19512
rect 390140 -19568 390208 -19512
rect 389868 -19654 390208 -19568
rect 389868 -19710 389942 -19654
rect 389998 -19710 390084 -19654
rect 390140 -19710 390208 -19654
rect 389868 -19796 390208 -19710
rect 389868 -19852 389942 -19796
rect 389998 -19852 390084 -19796
rect 390140 -19852 390208 -19796
rect 389868 -19938 390208 -19852
rect 389868 -19994 389942 -19938
rect 389998 -19994 390084 -19938
rect 390140 -19994 390208 -19938
rect 389868 -20080 390208 -19994
rect 389868 -20136 389942 -20080
rect 389998 -20136 390084 -20080
rect 390140 -20136 390208 -20080
rect 389868 -20222 390208 -20136
rect 389868 -20278 389942 -20222
rect 389998 -20278 390084 -20222
rect 390140 -20278 390208 -20222
rect 389868 -20364 390208 -20278
rect 389868 -20420 389942 -20364
rect 389998 -20420 390084 -20364
rect 390140 -20420 390208 -20364
rect 389868 -20506 390208 -20420
rect 389868 -20562 389942 -20506
rect 389998 -20562 390084 -20506
rect 390140 -20562 390208 -20506
rect 389868 -20648 390208 -20562
rect 389868 -20704 389942 -20648
rect 389998 -20704 390084 -20648
rect 390140 -20704 390208 -20648
rect 389868 -20790 390208 -20704
rect 389868 -20846 389942 -20790
rect 389998 -20846 390084 -20790
rect 390140 -20846 390208 -20790
rect 389868 -20932 390208 -20846
rect 389868 -20988 389942 -20932
rect 389998 -20988 390084 -20932
rect 390140 -20988 390208 -20932
rect 389868 -21074 390208 -20988
rect 389868 -21130 389942 -21074
rect 389998 -21130 390084 -21074
rect 390140 -21130 390208 -21074
rect 389868 -21216 390208 -21130
rect 389868 -21272 389942 -21216
rect 389998 -21272 390084 -21216
rect 390140 -21272 390208 -21216
rect 389868 -21358 390208 -21272
rect 389868 -21414 389942 -21358
rect 389998 -21414 390084 -21358
rect 390140 -21414 390208 -21358
rect 389868 -21500 390208 -21414
rect 389868 -21556 389942 -21500
rect 389998 -21556 390084 -21500
rect 390140 -21556 390208 -21500
rect 389868 -21642 390208 -21556
rect 389868 -21698 389942 -21642
rect 389998 -21698 390084 -21642
rect 390140 -21698 390208 -21642
rect 389868 -21784 390208 -21698
rect 389868 -21840 389942 -21784
rect 389998 -21840 390084 -21784
rect 390140 -21840 390208 -21784
rect 389868 -21926 390208 -21840
rect 389868 -21982 389942 -21926
rect 389998 -21982 390084 -21926
rect 390140 -21982 390208 -21926
rect 389868 -22068 390208 -21982
rect 389868 -22124 389942 -22068
rect 389998 -22124 390084 -22068
rect 390140 -22124 390208 -22068
rect 389868 -22210 390208 -22124
rect 389868 -22266 389942 -22210
rect 389998 -22266 390084 -22210
rect 390140 -22266 390208 -22210
rect 389868 -22352 390208 -22266
rect 389868 -22408 389942 -22352
rect 389998 -22408 390084 -22352
rect 390140 -22408 390208 -22352
rect 389868 -22494 390208 -22408
rect 389868 -22550 389942 -22494
rect 389998 -22550 390084 -22494
rect 390140 -22550 390208 -22494
rect 389868 -22636 390208 -22550
rect 389868 -22692 389942 -22636
rect 389998 -22692 390084 -22636
rect 390140 -22692 390208 -22636
rect 389868 -22778 390208 -22692
rect 389868 -22834 389942 -22778
rect 389998 -22834 390084 -22778
rect 390140 -22834 390208 -22778
rect 389868 -22920 390208 -22834
rect 389868 -22976 389942 -22920
rect 389998 -22976 390084 -22920
rect 390140 -22976 390208 -22920
rect 389868 -23062 390208 -22976
rect 389868 -23118 389942 -23062
rect 389998 -23118 390084 -23062
rect 390140 -23118 390208 -23062
rect 389868 -23204 390208 -23118
rect 389868 -23260 389942 -23204
rect 389998 -23260 390084 -23204
rect 390140 -23260 390208 -23204
rect 389868 -23346 390208 -23260
rect 389868 -23402 389942 -23346
rect 389998 -23402 390084 -23346
rect 390140 -23402 390208 -23346
rect 389868 -23488 390208 -23402
rect 389868 -23544 389942 -23488
rect 389998 -23544 390084 -23488
rect 390140 -23544 390208 -23488
rect 389868 -23630 390208 -23544
rect 389868 -23686 389942 -23630
rect 389998 -23686 390084 -23630
rect 390140 -23686 390208 -23630
rect 389868 -23772 390208 -23686
rect 389868 -23828 389942 -23772
rect 389998 -23828 390084 -23772
rect 390140 -23828 390208 -23772
rect 389868 -23914 390208 -23828
rect 389868 -23970 389942 -23914
rect 389998 -23970 390084 -23914
rect 390140 -23970 390208 -23914
rect 389868 -24056 390208 -23970
rect 389868 -24112 389942 -24056
rect 389998 -24112 390084 -24056
rect 390140 -24112 390208 -24056
rect 389868 -24198 390208 -24112
rect 389868 -24254 389942 -24198
rect 389998 -24254 390084 -24198
rect 390140 -24254 390208 -24198
rect 389868 -24340 390208 -24254
rect 389868 -24396 389942 -24340
rect 389998 -24396 390084 -24340
rect 390140 -24396 390208 -24340
rect 389868 -24482 390208 -24396
rect 389868 -24538 389942 -24482
rect 389998 -24538 390084 -24482
rect 390140 -24538 390208 -24482
rect 389868 -24624 390208 -24538
rect 389868 -24680 389942 -24624
rect 389998 -24680 390084 -24624
rect 390140 -24680 390208 -24624
rect 389868 -24766 390208 -24680
rect 389868 -24822 389942 -24766
rect 389998 -24822 390084 -24766
rect 390140 -24822 390208 -24766
rect 389868 -24908 390208 -24822
rect 389868 -24964 389942 -24908
rect 389998 -24964 390084 -24908
rect 390140 -24964 390208 -24908
rect 389868 -25050 390208 -24964
rect 389868 -25106 389942 -25050
rect 389998 -25106 390084 -25050
rect 390140 -25106 390208 -25050
rect 389868 -25192 390208 -25106
rect 389868 -25248 389942 -25192
rect 389998 -25248 390084 -25192
rect 390140 -25248 390208 -25192
rect 389868 -25334 390208 -25248
rect 389868 -25390 389942 -25334
rect 389998 -25390 390084 -25334
rect 390140 -25390 390208 -25334
rect 389868 -25476 390208 -25390
rect 389868 -25532 389942 -25476
rect 389998 -25532 390084 -25476
rect 390140 -25532 390208 -25476
rect 389868 -25542 390208 -25532
rect 390268 -17950 390608 -17820
rect 390268 -18006 390339 -17950
rect 390395 -18006 390481 -17950
rect 390537 -18006 390608 -17950
rect 390268 -18092 390608 -18006
rect 390268 -18148 390339 -18092
rect 390395 -18148 390481 -18092
rect 390537 -18148 390608 -18092
rect 390268 -18234 390608 -18148
rect 390268 -18290 390339 -18234
rect 390395 -18290 390481 -18234
rect 390537 -18290 390608 -18234
rect 390268 -18376 390608 -18290
rect 390268 -18432 390339 -18376
rect 390395 -18432 390481 -18376
rect 390537 -18432 390608 -18376
rect 390268 -18518 390608 -18432
rect 390268 -18574 390339 -18518
rect 390395 -18574 390481 -18518
rect 390537 -18574 390608 -18518
rect 390268 -18660 390608 -18574
rect 390268 -18716 390339 -18660
rect 390395 -18716 390481 -18660
rect 390537 -18716 390608 -18660
rect 390268 -18802 390608 -18716
rect 390268 -18858 390339 -18802
rect 390395 -18858 390481 -18802
rect 390537 -18858 390608 -18802
rect 390268 -18944 390608 -18858
rect 390268 -19000 390339 -18944
rect 390395 -19000 390481 -18944
rect 390537 -19000 390608 -18944
rect 390268 -19086 390608 -19000
rect 390268 -19142 390339 -19086
rect 390395 -19142 390481 -19086
rect 390537 -19142 390608 -19086
rect 390268 -19228 390608 -19142
rect 390268 -19284 390339 -19228
rect 390395 -19284 390481 -19228
rect 390537 -19284 390608 -19228
rect 390268 -19370 390608 -19284
rect 390268 -19426 390339 -19370
rect 390395 -19426 390481 -19370
rect 390537 -19426 390608 -19370
rect 390268 -19512 390608 -19426
rect 390268 -19568 390339 -19512
rect 390395 -19568 390481 -19512
rect 390537 -19568 390608 -19512
rect 390268 -19654 390608 -19568
rect 390268 -19710 390339 -19654
rect 390395 -19710 390481 -19654
rect 390537 -19710 390608 -19654
rect 390268 -19796 390608 -19710
rect 390268 -19852 390339 -19796
rect 390395 -19852 390481 -19796
rect 390537 -19852 390608 -19796
rect 390268 -19938 390608 -19852
rect 390268 -19994 390339 -19938
rect 390395 -19994 390481 -19938
rect 390537 -19994 390608 -19938
rect 390268 -20080 390608 -19994
rect 390268 -20136 390339 -20080
rect 390395 -20136 390481 -20080
rect 390537 -20136 390608 -20080
rect 390268 -20222 390608 -20136
rect 390268 -20278 390339 -20222
rect 390395 -20278 390481 -20222
rect 390537 -20278 390608 -20222
rect 390268 -20364 390608 -20278
rect 390268 -20420 390339 -20364
rect 390395 -20420 390481 -20364
rect 390537 -20420 390608 -20364
rect 390268 -20506 390608 -20420
rect 390268 -20562 390339 -20506
rect 390395 -20562 390481 -20506
rect 390537 -20562 390608 -20506
rect 390268 -20648 390608 -20562
rect 390268 -20704 390339 -20648
rect 390395 -20704 390481 -20648
rect 390537 -20704 390608 -20648
rect 390268 -20790 390608 -20704
rect 390268 -20846 390339 -20790
rect 390395 -20846 390481 -20790
rect 390537 -20846 390608 -20790
rect 390268 -20932 390608 -20846
rect 390268 -20988 390339 -20932
rect 390395 -20988 390481 -20932
rect 390537 -20988 390608 -20932
rect 390268 -21074 390608 -20988
rect 390268 -21130 390339 -21074
rect 390395 -21130 390481 -21074
rect 390537 -21130 390608 -21074
rect 390268 -21216 390608 -21130
rect 390268 -21272 390339 -21216
rect 390395 -21272 390481 -21216
rect 390537 -21272 390608 -21216
rect 390268 -21358 390608 -21272
rect 390268 -21414 390339 -21358
rect 390395 -21414 390481 -21358
rect 390537 -21414 390608 -21358
rect 390268 -21500 390608 -21414
rect 390268 -21556 390339 -21500
rect 390395 -21556 390481 -21500
rect 390537 -21556 390608 -21500
rect 390268 -21642 390608 -21556
rect 390268 -21698 390339 -21642
rect 390395 -21698 390481 -21642
rect 390537 -21698 390608 -21642
rect 390268 -21784 390608 -21698
rect 390268 -21840 390339 -21784
rect 390395 -21840 390481 -21784
rect 390537 -21840 390608 -21784
rect 390268 -21926 390608 -21840
rect 390268 -21982 390339 -21926
rect 390395 -21982 390481 -21926
rect 390537 -21982 390608 -21926
rect 390268 -22068 390608 -21982
rect 390268 -22124 390339 -22068
rect 390395 -22124 390481 -22068
rect 390537 -22124 390608 -22068
rect 390268 -22210 390608 -22124
rect 390268 -22266 390339 -22210
rect 390395 -22266 390481 -22210
rect 390537 -22266 390608 -22210
rect 390268 -22352 390608 -22266
rect 390268 -22408 390339 -22352
rect 390395 -22408 390481 -22352
rect 390537 -22408 390608 -22352
rect 390268 -22494 390608 -22408
rect 390268 -22550 390339 -22494
rect 390395 -22550 390481 -22494
rect 390537 -22550 390608 -22494
rect 390268 -22636 390608 -22550
rect 390268 -22692 390339 -22636
rect 390395 -22692 390481 -22636
rect 390537 -22692 390608 -22636
rect 390268 -22778 390608 -22692
rect 390268 -22834 390339 -22778
rect 390395 -22834 390481 -22778
rect 390537 -22834 390608 -22778
rect 390268 -22920 390608 -22834
rect 390268 -22976 390339 -22920
rect 390395 -22976 390481 -22920
rect 390537 -22976 390608 -22920
rect 390268 -23062 390608 -22976
rect 390268 -23118 390339 -23062
rect 390395 -23118 390481 -23062
rect 390537 -23118 390608 -23062
rect 390268 -23204 390608 -23118
rect 390268 -23260 390339 -23204
rect 390395 -23260 390481 -23204
rect 390537 -23260 390608 -23204
rect 390268 -23346 390608 -23260
rect 390268 -23402 390339 -23346
rect 390395 -23402 390481 -23346
rect 390537 -23402 390608 -23346
rect 390268 -23488 390608 -23402
rect 390268 -23544 390339 -23488
rect 390395 -23544 390481 -23488
rect 390537 -23544 390608 -23488
rect 390268 -23630 390608 -23544
rect 390268 -23686 390339 -23630
rect 390395 -23686 390481 -23630
rect 390537 -23686 390608 -23630
rect 390268 -23772 390608 -23686
rect 390268 -23828 390339 -23772
rect 390395 -23828 390481 -23772
rect 390537 -23828 390608 -23772
rect 390268 -23914 390608 -23828
rect 390268 -23970 390339 -23914
rect 390395 -23970 390481 -23914
rect 390537 -23970 390608 -23914
rect 390268 -24056 390608 -23970
rect 390268 -24112 390339 -24056
rect 390395 -24112 390481 -24056
rect 390537 -24112 390608 -24056
rect 390268 -24198 390608 -24112
rect 390268 -24254 390339 -24198
rect 390395 -24254 390481 -24198
rect 390537 -24254 390608 -24198
rect 390268 -24340 390608 -24254
rect 390268 -24396 390339 -24340
rect 390395 -24396 390481 -24340
rect 390537 -24396 390608 -24340
rect 390268 -24482 390608 -24396
rect 390268 -24538 390339 -24482
rect 390395 -24538 390481 -24482
rect 390537 -24538 390608 -24482
rect 390268 -24624 390608 -24538
rect 390268 -24680 390339 -24624
rect 390395 -24680 390481 -24624
rect 390537 -24680 390608 -24624
rect 390268 -24766 390608 -24680
rect 390268 -24822 390339 -24766
rect 390395 -24822 390481 -24766
rect 390537 -24822 390608 -24766
rect 390268 -24908 390608 -24822
rect 390268 -24964 390339 -24908
rect 390395 -24964 390481 -24908
rect 390537 -24964 390608 -24908
rect 390268 -25050 390608 -24964
rect 390268 -25106 390339 -25050
rect 390395 -25106 390481 -25050
rect 390537 -25106 390608 -25050
rect 390268 -25192 390608 -25106
rect 390268 -25248 390339 -25192
rect 390395 -25248 390481 -25192
rect 390537 -25248 390608 -25192
rect 390268 -25334 390608 -25248
rect 390268 -25390 390339 -25334
rect 390395 -25390 390481 -25334
rect 390537 -25390 390608 -25334
rect 390268 -25476 390608 -25390
rect 390268 -25532 390339 -25476
rect 390395 -25532 390481 -25476
rect 390537 -25532 390608 -25476
rect 390268 -25542 390608 -25532
rect 390668 -17950 391008 -17820
rect 390668 -18006 390736 -17950
rect 390792 -18006 390878 -17950
rect 390934 -18006 391008 -17950
rect 390668 -18092 391008 -18006
rect 390668 -18148 390736 -18092
rect 390792 -18148 390878 -18092
rect 390934 -18148 391008 -18092
rect 390668 -18234 391008 -18148
rect 390668 -18290 390736 -18234
rect 390792 -18290 390878 -18234
rect 390934 -18290 391008 -18234
rect 390668 -18376 391008 -18290
rect 390668 -18432 390736 -18376
rect 390792 -18432 390878 -18376
rect 390934 -18432 391008 -18376
rect 390668 -18518 391008 -18432
rect 390668 -18574 390736 -18518
rect 390792 -18574 390878 -18518
rect 390934 -18574 391008 -18518
rect 390668 -18660 391008 -18574
rect 390668 -18716 390736 -18660
rect 390792 -18716 390878 -18660
rect 390934 -18716 391008 -18660
rect 390668 -18802 391008 -18716
rect 390668 -18858 390736 -18802
rect 390792 -18858 390878 -18802
rect 390934 -18858 391008 -18802
rect 390668 -18944 391008 -18858
rect 390668 -19000 390736 -18944
rect 390792 -19000 390878 -18944
rect 390934 -19000 391008 -18944
rect 390668 -19086 391008 -19000
rect 390668 -19142 390736 -19086
rect 390792 -19142 390878 -19086
rect 390934 -19142 391008 -19086
rect 390668 -19228 391008 -19142
rect 390668 -19284 390736 -19228
rect 390792 -19284 390878 -19228
rect 390934 -19284 391008 -19228
rect 390668 -19370 391008 -19284
rect 390668 -19426 390736 -19370
rect 390792 -19426 390878 -19370
rect 390934 -19426 391008 -19370
rect 390668 -19512 391008 -19426
rect 390668 -19568 390736 -19512
rect 390792 -19568 390878 -19512
rect 390934 -19568 391008 -19512
rect 390668 -19654 391008 -19568
rect 390668 -19710 390736 -19654
rect 390792 -19710 390878 -19654
rect 390934 -19710 391008 -19654
rect 390668 -19796 391008 -19710
rect 390668 -19852 390736 -19796
rect 390792 -19852 390878 -19796
rect 390934 -19852 391008 -19796
rect 390668 -19938 391008 -19852
rect 390668 -19994 390736 -19938
rect 390792 -19994 390878 -19938
rect 390934 -19994 391008 -19938
rect 390668 -20080 391008 -19994
rect 390668 -20136 390736 -20080
rect 390792 -20136 390878 -20080
rect 390934 -20136 391008 -20080
rect 390668 -20222 391008 -20136
rect 390668 -20278 390736 -20222
rect 390792 -20278 390878 -20222
rect 390934 -20278 391008 -20222
rect 390668 -20364 391008 -20278
rect 390668 -20420 390736 -20364
rect 390792 -20420 390878 -20364
rect 390934 -20420 391008 -20364
rect 390668 -20506 391008 -20420
rect 390668 -20562 390736 -20506
rect 390792 -20562 390878 -20506
rect 390934 -20562 391008 -20506
rect 390668 -20648 391008 -20562
rect 390668 -20704 390736 -20648
rect 390792 -20704 390878 -20648
rect 390934 -20704 391008 -20648
rect 390668 -20790 391008 -20704
rect 390668 -20846 390736 -20790
rect 390792 -20846 390878 -20790
rect 390934 -20846 391008 -20790
rect 390668 -20932 391008 -20846
rect 390668 -20988 390736 -20932
rect 390792 -20988 390878 -20932
rect 390934 -20988 391008 -20932
rect 390668 -21074 391008 -20988
rect 390668 -21130 390736 -21074
rect 390792 -21130 390878 -21074
rect 390934 -21130 391008 -21074
rect 390668 -21216 391008 -21130
rect 390668 -21272 390736 -21216
rect 390792 -21272 390878 -21216
rect 390934 -21272 391008 -21216
rect 390668 -21358 391008 -21272
rect 390668 -21414 390736 -21358
rect 390792 -21414 390878 -21358
rect 390934 -21414 391008 -21358
rect 390668 -21500 391008 -21414
rect 390668 -21556 390736 -21500
rect 390792 -21556 390878 -21500
rect 390934 -21556 391008 -21500
rect 390668 -21642 391008 -21556
rect 390668 -21698 390736 -21642
rect 390792 -21698 390878 -21642
rect 390934 -21698 391008 -21642
rect 390668 -21784 391008 -21698
rect 390668 -21840 390736 -21784
rect 390792 -21840 390878 -21784
rect 390934 -21840 391008 -21784
rect 390668 -21926 391008 -21840
rect 390668 -21982 390736 -21926
rect 390792 -21982 390878 -21926
rect 390934 -21982 391008 -21926
rect 390668 -22068 391008 -21982
rect 390668 -22124 390736 -22068
rect 390792 -22124 390878 -22068
rect 390934 -22124 391008 -22068
rect 390668 -22210 391008 -22124
rect 390668 -22266 390736 -22210
rect 390792 -22266 390878 -22210
rect 390934 -22266 391008 -22210
rect 390668 -22352 391008 -22266
rect 390668 -22408 390736 -22352
rect 390792 -22408 390878 -22352
rect 390934 -22408 391008 -22352
rect 390668 -22494 391008 -22408
rect 390668 -22550 390736 -22494
rect 390792 -22550 390878 -22494
rect 390934 -22550 391008 -22494
rect 390668 -22636 391008 -22550
rect 390668 -22692 390736 -22636
rect 390792 -22692 390878 -22636
rect 390934 -22692 391008 -22636
rect 390668 -22778 391008 -22692
rect 390668 -22834 390736 -22778
rect 390792 -22834 390878 -22778
rect 390934 -22834 391008 -22778
rect 390668 -22920 391008 -22834
rect 390668 -22976 390736 -22920
rect 390792 -22976 390878 -22920
rect 390934 -22976 391008 -22920
rect 390668 -23062 391008 -22976
rect 390668 -23118 390736 -23062
rect 390792 -23118 390878 -23062
rect 390934 -23118 391008 -23062
rect 390668 -23204 391008 -23118
rect 390668 -23260 390736 -23204
rect 390792 -23260 390878 -23204
rect 390934 -23260 391008 -23204
rect 390668 -23346 391008 -23260
rect 390668 -23402 390736 -23346
rect 390792 -23402 390878 -23346
rect 390934 -23402 391008 -23346
rect 390668 -23488 391008 -23402
rect 390668 -23544 390736 -23488
rect 390792 -23544 390878 -23488
rect 390934 -23544 391008 -23488
rect 390668 -23630 391008 -23544
rect 390668 -23686 390736 -23630
rect 390792 -23686 390878 -23630
rect 390934 -23686 391008 -23630
rect 390668 -23772 391008 -23686
rect 390668 -23828 390736 -23772
rect 390792 -23828 390878 -23772
rect 390934 -23828 391008 -23772
rect 390668 -23914 391008 -23828
rect 390668 -23970 390736 -23914
rect 390792 -23970 390878 -23914
rect 390934 -23970 391008 -23914
rect 390668 -24056 391008 -23970
rect 390668 -24112 390736 -24056
rect 390792 -24112 390878 -24056
rect 390934 -24112 391008 -24056
rect 390668 -24198 391008 -24112
rect 390668 -24254 390736 -24198
rect 390792 -24254 390878 -24198
rect 390934 -24254 391008 -24198
rect 390668 -24340 391008 -24254
rect 390668 -24396 390736 -24340
rect 390792 -24396 390878 -24340
rect 390934 -24396 391008 -24340
rect 390668 -24482 391008 -24396
rect 390668 -24538 390736 -24482
rect 390792 -24538 390878 -24482
rect 390934 -24538 391008 -24482
rect 390668 -24624 391008 -24538
rect 390668 -24680 390736 -24624
rect 390792 -24680 390878 -24624
rect 390934 -24680 391008 -24624
rect 390668 -24766 391008 -24680
rect 390668 -24822 390736 -24766
rect 390792 -24822 390878 -24766
rect 390934 -24822 391008 -24766
rect 390668 -24908 391008 -24822
rect 390668 -24964 390736 -24908
rect 390792 -24964 390878 -24908
rect 390934 -24964 391008 -24908
rect 390668 -25050 391008 -24964
rect 390668 -25106 390736 -25050
rect 390792 -25106 390878 -25050
rect 390934 -25106 391008 -25050
rect 390668 -25192 391008 -25106
rect 390668 -25248 390736 -25192
rect 390792 -25248 390878 -25192
rect 390934 -25248 391008 -25192
rect 390668 -25334 391008 -25248
rect 390668 -25390 390736 -25334
rect 390792 -25390 390878 -25334
rect 390934 -25390 391008 -25334
rect 390668 -25476 391008 -25390
rect 390668 -25532 390736 -25476
rect 390792 -25532 390878 -25476
rect 390934 -25532 391008 -25476
rect 390668 -25542 391008 -25532
rect 391068 -17950 391408 -17820
rect 391068 -18006 391140 -17950
rect 391196 -18006 391282 -17950
rect 391338 -18006 391408 -17950
rect 391068 -18092 391408 -18006
rect 391068 -18148 391140 -18092
rect 391196 -18148 391282 -18092
rect 391338 -18148 391408 -18092
rect 391068 -18234 391408 -18148
rect 391068 -18290 391140 -18234
rect 391196 -18290 391282 -18234
rect 391338 -18290 391408 -18234
rect 391068 -18376 391408 -18290
rect 391068 -18432 391140 -18376
rect 391196 -18432 391282 -18376
rect 391338 -18432 391408 -18376
rect 391068 -18518 391408 -18432
rect 391068 -18574 391140 -18518
rect 391196 -18574 391282 -18518
rect 391338 -18574 391408 -18518
rect 391068 -18660 391408 -18574
rect 391068 -18716 391140 -18660
rect 391196 -18716 391282 -18660
rect 391338 -18716 391408 -18660
rect 391068 -18802 391408 -18716
rect 391068 -18858 391140 -18802
rect 391196 -18858 391282 -18802
rect 391338 -18858 391408 -18802
rect 391068 -18944 391408 -18858
rect 391068 -19000 391140 -18944
rect 391196 -19000 391282 -18944
rect 391338 -19000 391408 -18944
rect 391068 -19086 391408 -19000
rect 391068 -19142 391140 -19086
rect 391196 -19142 391282 -19086
rect 391338 -19142 391408 -19086
rect 391068 -19228 391408 -19142
rect 391068 -19284 391140 -19228
rect 391196 -19284 391282 -19228
rect 391338 -19284 391408 -19228
rect 391068 -19370 391408 -19284
rect 391068 -19426 391140 -19370
rect 391196 -19426 391282 -19370
rect 391338 -19426 391408 -19370
rect 391068 -19512 391408 -19426
rect 391068 -19568 391140 -19512
rect 391196 -19568 391282 -19512
rect 391338 -19568 391408 -19512
rect 391068 -19654 391408 -19568
rect 391068 -19710 391140 -19654
rect 391196 -19710 391282 -19654
rect 391338 -19710 391408 -19654
rect 391068 -19796 391408 -19710
rect 391068 -19852 391140 -19796
rect 391196 -19852 391282 -19796
rect 391338 -19852 391408 -19796
rect 391068 -19938 391408 -19852
rect 391068 -19994 391140 -19938
rect 391196 -19994 391282 -19938
rect 391338 -19994 391408 -19938
rect 391068 -20080 391408 -19994
rect 391068 -20136 391140 -20080
rect 391196 -20136 391282 -20080
rect 391338 -20136 391408 -20080
rect 391068 -20222 391408 -20136
rect 391068 -20278 391140 -20222
rect 391196 -20278 391282 -20222
rect 391338 -20278 391408 -20222
rect 391068 -20364 391408 -20278
rect 391068 -20420 391140 -20364
rect 391196 -20420 391282 -20364
rect 391338 -20420 391408 -20364
rect 391068 -20506 391408 -20420
rect 391068 -20562 391140 -20506
rect 391196 -20562 391282 -20506
rect 391338 -20562 391408 -20506
rect 391068 -20648 391408 -20562
rect 391068 -20704 391140 -20648
rect 391196 -20704 391282 -20648
rect 391338 -20704 391408 -20648
rect 391068 -20790 391408 -20704
rect 391068 -20846 391140 -20790
rect 391196 -20846 391282 -20790
rect 391338 -20846 391408 -20790
rect 391068 -20932 391408 -20846
rect 391068 -20988 391140 -20932
rect 391196 -20988 391282 -20932
rect 391338 -20988 391408 -20932
rect 391068 -21074 391408 -20988
rect 391068 -21130 391140 -21074
rect 391196 -21130 391282 -21074
rect 391338 -21130 391408 -21074
rect 391068 -21216 391408 -21130
rect 391068 -21272 391140 -21216
rect 391196 -21272 391282 -21216
rect 391338 -21272 391408 -21216
rect 391068 -21358 391408 -21272
rect 391068 -21414 391140 -21358
rect 391196 -21414 391282 -21358
rect 391338 -21414 391408 -21358
rect 391068 -21500 391408 -21414
rect 391068 -21556 391140 -21500
rect 391196 -21556 391282 -21500
rect 391338 -21556 391408 -21500
rect 391068 -21642 391408 -21556
rect 391068 -21698 391140 -21642
rect 391196 -21698 391282 -21642
rect 391338 -21698 391408 -21642
rect 391068 -21784 391408 -21698
rect 391068 -21840 391140 -21784
rect 391196 -21840 391282 -21784
rect 391338 -21840 391408 -21784
rect 391068 -21926 391408 -21840
rect 391068 -21982 391140 -21926
rect 391196 -21982 391282 -21926
rect 391338 -21982 391408 -21926
rect 391068 -22068 391408 -21982
rect 391068 -22124 391140 -22068
rect 391196 -22124 391282 -22068
rect 391338 -22124 391408 -22068
rect 391068 -22210 391408 -22124
rect 391068 -22266 391140 -22210
rect 391196 -22266 391282 -22210
rect 391338 -22266 391408 -22210
rect 391068 -22352 391408 -22266
rect 391068 -22408 391140 -22352
rect 391196 -22408 391282 -22352
rect 391338 -22408 391408 -22352
rect 391068 -22494 391408 -22408
rect 391068 -22550 391140 -22494
rect 391196 -22550 391282 -22494
rect 391338 -22550 391408 -22494
rect 391068 -22636 391408 -22550
rect 391068 -22692 391140 -22636
rect 391196 -22692 391282 -22636
rect 391338 -22692 391408 -22636
rect 391068 -22778 391408 -22692
rect 391068 -22834 391140 -22778
rect 391196 -22834 391282 -22778
rect 391338 -22834 391408 -22778
rect 391068 -22920 391408 -22834
rect 391068 -22976 391140 -22920
rect 391196 -22976 391282 -22920
rect 391338 -22976 391408 -22920
rect 391068 -23062 391408 -22976
rect 391068 -23118 391140 -23062
rect 391196 -23118 391282 -23062
rect 391338 -23118 391408 -23062
rect 391068 -23204 391408 -23118
rect 391068 -23260 391140 -23204
rect 391196 -23260 391282 -23204
rect 391338 -23260 391408 -23204
rect 391068 -23346 391408 -23260
rect 391068 -23402 391140 -23346
rect 391196 -23402 391282 -23346
rect 391338 -23402 391408 -23346
rect 391068 -23488 391408 -23402
rect 391068 -23544 391140 -23488
rect 391196 -23544 391282 -23488
rect 391338 -23544 391408 -23488
rect 391068 -23630 391408 -23544
rect 391068 -23686 391140 -23630
rect 391196 -23686 391282 -23630
rect 391338 -23686 391408 -23630
rect 391068 -23772 391408 -23686
rect 391068 -23828 391140 -23772
rect 391196 -23828 391282 -23772
rect 391338 -23828 391408 -23772
rect 391068 -23914 391408 -23828
rect 391068 -23970 391140 -23914
rect 391196 -23970 391282 -23914
rect 391338 -23970 391408 -23914
rect 391068 -24056 391408 -23970
rect 391068 -24112 391140 -24056
rect 391196 -24112 391282 -24056
rect 391338 -24112 391408 -24056
rect 391068 -24198 391408 -24112
rect 391068 -24254 391140 -24198
rect 391196 -24254 391282 -24198
rect 391338 -24254 391408 -24198
rect 391068 -24340 391408 -24254
rect 391068 -24396 391140 -24340
rect 391196 -24396 391282 -24340
rect 391338 -24396 391408 -24340
rect 391068 -24482 391408 -24396
rect 391068 -24538 391140 -24482
rect 391196 -24538 391282 -24482
rect 391338 -24538 391408 -24482
rect 391068 -24624 391408 -24538
rect 391068 -24680 391140 -24624
rect 391196 -24680 391282 -24624
rect 391338 -24680 391408 -24624
rect 391068 -24766 391408 -24680
rect 391068 -24822 391140 -24766
rect 391196 -24822 391282 -24766
rect 391338 -24822 391408 -24766
rect 391068 -24908 391408 -24822
rect 391068 -24964 391140 -24908
rect 391196 -24964 391282 -24908
rect 391338 -24964 391408 -24908
rect 391068 -25050 391408 -24964
rect 391068 -25106 391140 -25050
rect 391196 -25106 391282 -25050
rect 391338 -25106 391408 -25050
rect 391068 -25192 391408 -25106
rect 391068 -25248 391140 -25192
rect 391196 -25248 391282 -25192
rect 391338 -25248 391408 -25192
rect 391068 -25334 391408 -25248
rect 391068 -25390 391140 -25334
rect 391196 -25390 391282 -25334
rect 391338 -25390 391408 -25334
rect 391068 -25476 391408 -25390
rect 391068 -25532 391140 -25476
rect 391196 -25532 391282 -25476
rect 391338 -25532 391408 -25476
rect 391068 -25542 391408 -25532
rect 391468 -17950 391808 -17820
rect 391468 -18006 391536 -17950
rect 391592 -18006 391678 -17950
rect 391734 -18006 391808 -17950
rect 391468 -18092 391808 -18006
rect 391468 -18148 391536 -18092
rect 391592 -18148 391678 -18092
rect 391734 -18148 391808 -18092
rect 391468 -18234 391808 -18148
rect 391468 -18290 391536 -18234
rect 391592 -18290 391678 -18234
rect 391734 -18290 391808 -18234
rect 391468 -18376 391808 -18290
rect 391468 -18432 391536 -18376
rect 391592 -18432 391678 -18376
rect 391734 -18432 391808 -18376
rect 391468 -18518 391808 -18432
rect 391468 -18574 391536 -18518
rect 391592 -18574 391678 -18518
rect 391734 -18574 391808 -18518
rect 391468 -18660 391808 -18574
rect 391468 -18716 391536 -18660
rect 391592 -18716 391678 -18660
rect 391734 -18716 391808 -18660
rect 391468 -18802 391808 -18716
rect 391468 -18858 391536 -18802
rect 391592 -18858 391678 -18802
rect 391734 -18858 391808 -18802
rect 391468 -18944 391808 -18858
rect 391468 -19000 391536 -18944
rect 391592 -19000 391678 -18944
rect 391734 -19000 391808 -18944
rect 391468 -19086 391808 -19000
rect 391468 -19142 391536 -19086
rect 391592 -19142 391678 -19086
rect 391734 -19142 391808 -19086
rect 391468 -19228 391808 -19142
rect 391468 -19284 391536 -19228
rect 391592 -19284 391678 -19228
rect 391734 -19284 391808 -19228
rect 391468 -19370 391808 -19284
rect 391468 -19426 391536 -19370
rect 391592 -19426 391678 -19370
rect 391734 -19426 391808 -19370
rect 391468 -19512 391808 -19426
rect 391468 -19568 391536 -19512
rect 391592 -19568 391678 -19512
rect 391734 -19568 391808 -19512
rect 391468 -19654 391808 -19568
rect 391468 -19710 391536 -19654
rect 391592 -19710 391678 -19654
rect 391734 -19710 391808 -19654
rect 391468 -19796 391808 -19710
rect 391468 -19852 391536 -19796
rect 391592 -19852 391678 -19796
rect 391734 -19852 391808 -19796
rect 391468 -19938 391808 -19852
rect 391468 -19994 391536 -19938
rect 391592 -19994 391678 -19938
rect 391734 -19994 391808 -19938
rect 391468 -20080 391808 -19994
rect 391468 -20136 391536 -20080
rect 391592 -20136 391678 -20080
rect 391734 -20136 391808 -20080
rect 391468 -20222 391808 -20136
rect 391468 -20278 391536 -20222
rect 391592 -20278 391678 -20222
rect 391734 -20278 391808 -20222
rect 391468 -20364 391808 -20278
rect 391468 -20420 391536 -20364
rect 391592 -20420 391678 -20364
rect 391734 -20420 391808 -20364
rect 391468 -20506 391808 -20420
rect 391468 -20562 391536 -20506
rect 391592 -20562 391678 -20506
rect 391734 -20562 391808 -20506
rect 391468 -20648 391808 -20562
rect 391468 -20704 391536 -20648
rect 391592 -20704 391678 -20648
rect 391734 -20704 391808 -20648
rect 391468 -20790 391808 -20704
rect 391468 -20846 391536 -20790
rect 391592 -20846 391678 -20790
rect 391734 -20846 391808 -20790
rect 391468 -20932 391808 -20846
rect 391468 -20988 391536 -20932
rect 391592 -20988 391678 -20932
rect 391734 -20988 391808 -20932
rect 391468 -21074 391808 -20988
rect 391468 -21130 391536 -21074
rect 391592 -21130 391678 -21074
rect 391734 -21130 391808 -21074
rect 391468 -21216 391808 -21130
rect 391468 -21272 391536 -21216
rect 391592 -21272 391678 -21216
rect 391734 -21272 391808 -21216
rect 391468 -21358 391808 -21272
rect 391468 -21414 391536 -21358
rect 391592 -21414 391678 -21358
rect 391734 -21414 391808 -21358
rect 391468 -21500 391808 -21414
rect 391468 -21556 391536 -21500
rect 391592 -21556 391678 -21500
rect 391734 -21556 391808 -21500
rect 391468 -21642 391808 -21556
rect 391468 -21698 391536 -21642
rect 391592 -21698 391678 -21642
rect 391734 -21698 391808 -21642
rect 391468 -21784 391808 -21698
rect 391468 -21840 391536 -21784
rect 391592 -21840 391678 -21784
rect 391734 -21840 391808 -21784
rect 391468 -21926 391808 -21840
rect 391468 -21982 391536 -21926
rect 391592 -21982 391678 -21926
rect 391734 -21982 391808 -21926
rect 391468 -22068 391808 -21982
rect 391468 -22124 391536 -22068
rect 391592 -22124 391678 -22068
rect 391734 -22124 391808 -22068
rect 391468 -22210 391808 -22124
rect 391468 -22266 391536 -22210
rect 391592 -22266 391678 -22210
rect 391734 -22266 391808 -22210
rect 391468 -22352 391808 -22266
rect 391468 -22408 391536 -22352
rect 391592 -22408 391678 -22352
rect 391734 -22408 391808 -22352
rect 391468 -22494 391808 -22408
rect 391468 -22550 391536 -22494
rect 391592 -22550 391678 -22494
rect 391734 -22550 391808 -22494
rect 391468 -22636 391808 -22550
rect 391468 -22692 391536 -22636
rect 391592 -22692 391678 -22636
rect 391734 -22692 391808 -22636
rect 391468 -22778 391808 -22692
rect 391468 -22834 391536 -22778
rect 391592 -22834 391678 -22778
rect 391734 -22834 391808 -22778
rect 391468 -22920 391808 -22834
rect 391468 -22976 391536 -22920
rect 391592 -22976 391678 -22920
rect 391734 -22976 391808 -22920
rect 391468 -23062 391808 -22976
rect 391468 -23118 391536 -23062
rect 391592 -23118 391678 -23062
rect 391734 -23118 391808 -23062
rect 391468 -23204 391808 -23118
rect 391468 -23260 391536 -23204
rect 391592 -23260 391678 -23204
rect 391734 -23260 391808 -23204
rect 391468 -23346 391808 -23260
rect 391468 -23402 391536 -23346
rect 391592 -23402 391678 -23346
rect 391734 -23402 391808 -23346
rect 391468 -23488 391808 -23402
rect 391468 -23544 391536 -23488
rect 391592 -23544 391678 -23488
rect 391734 -23544 391808 -23488
rect 391468 -23630 391808 -23544
rect 391468 -23686 391536 -23630
rect 391592 -23686 391678 -23630
rect 391734 -23686 391808 -23630
rect 391468 -23772 391808 -23686
rect 391468 -23828 391536 -23772
rect 391592 -23828 391678 -23772
rect 391734 -23828 391808 -23772
rect 391468 -23914 391808 -23828
rect 391468 -23970 391536 -23914
rect 391592 -23970 391678 -23914
rect 391734 -23970 391808 -23914
rect 391468 -24056 391808 -23970
rect 391468 -24112 391536 -24056
rect 391592 -24112 391678 -24056
rect 391734 -24112 391808 -24056
rect 391468 -24198 391808 -24112
rect 391468 -24254 391536 -24198
rect 391592 -24254 391678 -24198
rect 391734 -24254 391808 -24198
rect 391468 -24340 391808 -24254
rect 391468 -24396 391536 -24340
rect 391592 -24396 391678 -24340
rect 391734 -24396 391808 -24340
rect 391468 -24482 391808 -24396
rect 391468 -24538 391536 -24482
rect 391592 -24538 391678 -24482
rect 391734 -24538 391808 -24482
rect 391468 -24624 391808 -24538
rect 391468 -24680 391536 -24624
rect 391592 -24680 391678 -24624
rect 391734 -24680 391808 -24624
rect 391468 -24766 391808 -24680
rect 391468 -24822 391536 -24766
rect 391592 -24822 391678 -24766
rect 391734 -24822 391808 -24766
rect 391468 -24908 391808 -24822
rect 391468 -24964 391536 -24908
rect 391592 -24964 391678 -24908
rect 391734 -24964 391808 -24908
rect 391468 -25050 391808 -24964
rect 391468 -25106 391536 -25050
rect 391592 -25106 391678 -25050
rect 391734 -25106 391808 -25050
rect 391468 -25192 391808 -25106
rect 391468 -25248 391536 -25192
rect 391592 -25248 391678 -25192
rect 391734 -25248 391808 -25192
rect 391468 -25334 391808 -25248
rect 391468 -25390 391536 -25334
rect 391592 -25390 391678 -25334
rect 391734 -25390 391808 -25334
rect 391468 -25476 391808 -25390
rect 391468 -25532 391536 -25476
rect 391592 -25532 391678 -25476
rect 391734 -25532 391808 -25476
rect 391468 -25542 391808 -25532
rect 391868 -17950 392208 -17820
rect 391868 -18006 391936 -17950
rect 391992 -18006 392078 -17950
rect 392134 -18006 392208 -17950
rect 391868 -18092 392208 -18006
rect 391868 -18148 391936 -18092
rect 391992 -18148 392078 -18092
rect 392134 -18148 392208 -18092
rect 391868 -18234 392208 -18148
rect 391868 -18290 391936 -18234
rect 391992 -18290 392078 -18234
rect 392134 -18290 392208 -18234
rect 391868 -18376 392208 -18290
rect 391868 -18432 391936 -18376
rect 391992 -18432 392078 -18376
rect 392134 -18432 392208 -18376
rect 391868 -18518 392208 -18432
rect 391868 -18574 391936 -18518
rect 391992 -18574 392078 -18518
rect 392134 -18574 392208 -18518
rect 391868 -18660 392208 -18574
rect 391868 -18716 391936 -18660
rect 391992 -18716 392078 -18660
rect 392134 -18716 392208 -18660
rect 391868 -18802 392208 -18716
rect 391868 -18858 391936 -18802
rect 391992 -18858 392078 -18802
rect 392134 -18858 392208 -18802
rect 391868 -18944 392208 -18858
rect 391868 -19000 391936 -18944
rect 391992 -19000 392078 -18944
rect 392134 -19000 392208 -18944
rect 391868 -19086 392208 -19000
rect 391868 -19142 391936 -19086
rect 391992 -19142 392078 -19086
rect 392134 -19142 392208 -19086
rect 391868 -19228 392208 -19142
rect 391868 -19284 391936 -19228
rect 391992 -19284 392078 -19228
rect 392134 -19284 392208 -19228
rect 391868 -19370 392208 -19284
rect 391868 -19426 391936 -19370
rect 391992 -19426 392078 -19370
rect 392134 -19426 392208 -19370
rect 391868 -19512 392208 -19426
rect 391868 -19568 391936 -19512
rect 391992 -19568 392078 -19512
rect 392134 -19568 392208 -19512
rect 391868 -19654 392208 -19568
rect 391868 -19710 391936 -19654
rect 391992 -19710 392078 -19654
rect 392134 -19710 392208 -19654
rect 391868 -19796 392208 -19710
rect 391868 -19852 391936 -19796
rect 391992 -19852 392078 -19796
rect 392134 -19852 392208 -19796
rect 391868 -19938 392208 -19852
rect 391868 -19994 391936 -19938
rect 391992 -19994 392078 -19938
rect 392134 -19994 392208 -19938
rect 391868 -20080 392208 -19994
rect 391868 -20136 391936 -20080
rect 391992 -20136 392078 -20080
rect 392134 -20136 392208 -20080
rect 391868 -20222 392208 -20136
rect 391868 -20278 391936 -20222
rect 391992 -20278 392078 -20222
rect 392134 -20278 392208 -20222
rect 391868 -20364 392208 -20278
rect 391868 -20420 391936 -20364
rect 391992 -20420 392078 -20364
rect 392134 -20420 392208 -20364
rect 391868 -20506 392208 -20420
rect 391868 -20562 391936 -20506
rect 391992 -20562 392078 -20506
rect 392134 -20562 392208 -20506
rect 391868 -20648 392208 -20562
rect 391868 -20704 391936 -20648
rect 391992 -20704 392078 -20648
rect 392134 -20704 392208 -20648
rect 391868 -20790 392208 -20704
rect 391868 -20846 391936 -20790
rect 391992 -20846 392078 -20790
rect 392134 -20846 392208 -20790
rect 391868 -20932 392208 -20846
rect 391868 -20988 391936 -20932
rect 391992 -20988 392078 -20932
rect 392134 -20988 392208 -20932
rect 391868 -21074 392208 -20988
rect 391868 -21130 391936 -21074
rect 391992 -21130 392078 -21074
rect 392134 -21130 392208 -21074
rect 391868 -21216 392208 -21130
rect 391868 -21272 391936 -21216
rect 391992 -21272 392078 -21216
rect 392134 -21272 392208 -21216
rect 391868 -21358 392208 -21272
rect 391868 -21414 391936 -21358
rect 391992 -21414 392078 -21358
rect 392134 -21414 392208 -21358
rect 391868 -21500 392208 -21414
rect 391868 -21556 391936 -21500
rect 391992 -21556 392078 -21500
rect 392134 -21556 392208 -21500
rect 391868 -21642 392208 -21556
rect 391868 -21698 391936 -21642
rect 391992 -21698 392078 -21642
rect 392134 -21698 392208 -21642
rect 391868 -21784 392208 -21698
rect 391868 -21840 391936 -21784
rect 391992 -21840 392078 -21784
rect 392134 -21840 392208 -21784
rect 391868 -21926 392208 -21840
rect 391868 -21982 391936 -21926
rect 391992 -21982 392078 -21926
rect 392134 -21982 392208 -21926
rect 391868 -22068 392208 -21982
rect 391868 -22124 391936 -22068
rect 391992 -22124 392078 -22068
rect 392134 -22124 392208 -22068
rect 391868 -22210 392208 -22124
rect 391868 -22266 391936 -22210
rect 391992 -22266 392078 -22210
rect 392134 -22266 392208 -22210
rect 391868 -22352 392208 -22266
rect 391868 -22408 391936 -22352
rect 391992 -22408 392078 -22352
rect 392134 -22408 392208 -22352
rect 391868 -22494 392208 -22408
rect 391868 -22550 391936 -22494
rect 391992 -22550 392078 -22494
rect 392134 -22550 392208 -22494
rect 391868 -22636 392208 -22550
rect 391868 -22692 391936 -22636
rect 391992 -22692 392078 -22636
rect 392134 -22692 392208 -22636
rect 391868 -22778 392208 -22692
rect 391868 -22834 391936 -22778
rect 391992 -22834 392078 -22778
rect 392134 -22834 392208 -22778
rect 391868 -22920 392208 -22834
rect 391868 -22976 391936 -22920
rect 391992 -22976 392078 -22920
rect 392134 -22976 392208 -22920
rect 391868 -23062 392208 -22976
rect 391868 -23118 391936 -23062
rect 391992 -23118 392078 -23062
rect 392134 -23118 392208 -23062
rect 391868 -23204 392208 -23118
rect 391868 -23260 391936 -23204
rect 391992 -23260 392078 -23204
rect 392134 -23260 392208 -23204
rect 391868 -23346 392208 -23260
rect 391868 -23402 391936 -23346
rect 391992 -23402 392078 -23346
rect 392134 -23402 392208 -23346
rect 391868 -23488 392208 -23402
rect 391868 -23544 391936 -23488
rect 391992 -23544 392078 -23488
rect 392134 -23544 392208 -23488
rect 391868 -23630 392208 -23544
rect 391868 -23686 391936 -23630
rect 391992 -23686 392078 -23630
rect 392134 -23686 392208 -23630
rect 391868 -23772 392208 -23686
rect 391868 -23828 391936 -23772
rect 391992 -23828 392078 -23772
rect 392134 -23828 392208 -23772
rect 391868 -23914 392208 -23828
rect 391868 -23970 391936 -23914
rect 391992 -23970 392078 -23914
rect 392134 -23970 392208 -23914
rect 391868 -24056 392208 -23970
rect 391868 -24112 391936 -24056
rect 391992 -24112 392078 -24056
rect 392134 -24112 392208 -24056
rect 391868 -24198 392208 -24112
rect 391868 -24254 391936 -24198
rect 391992 -24254 392078 -24198
rect 392134 -24254 392208 -24198
rect 391868 -24340 392208 -24254
rect 391868 -24396 391936 -24340
rect 391992 -24396 392078 -24340
rect 392134 -24396 392208 -24340
rect 391868 -24482 392208 -24396
rect 391868 -24538 391936 -24482
rect 391992 -24538 392078 -24482
rect 392134 -24538 392208 -24482
rect 391868 -24624 392208 -24538
rect 391868 -24680 391936 -24624
rect 391992 -24680 392078 -24624
rect 392134 -24680 392208 -24624
rect 391868 -24766 392208 -24680
rect 391868 -24822 391936 -24766
rect 391992 -24822 392078 -24766
rect 392134 -24822 392208 -24766
rect 391868 -24908 392208 -24822
rect 391868 -24964 391936 -24908
rect 391992 -24964 392078 -24908
rect 392134 -24964 392208 -24908
rect 391868 -25050 392208 -24964
rect 391868 -25106 391936 -25050
rect 391992 -25106 392078 -25050
rect 392134 -25106 392208 -25050
rect 391868 -25192 392208 -25106
rect 391868 -25248 391936 -25192
rect 391992 -25248 392078 -25192
rect 392134 -25248 392208 -25192
rect 391868 -25334 392208 -25248
rect 391868 -25390 391936 -25334
rect 391992 -25390 392078 -25334
rect 392134 -25390 392208 -25334
rect 391868 -25476 392208 -25390
rect 391868 -25532 391936 -25476
rect 391992 -25532 392078 -25476
rect 392134 -25532 392208 -25476
rect 391868 -25542 392208 -25532
rect 392268 -17950 392608 -17820
rect 392268 -18006 392333 -17950
rect 392389 -18006 392475 -17950
rect 392531 -18006 392608 -17950
rect 392268 -18092 392608 -18006
rect 392268 -18148 392333 -18092
rect 392389 -18148 392475 -18092
rect 392531 -18148 392608 -18092
rect 392268 -18234 392608 -18148
rect 392268 -18290 392333 -18234
rect 392389 -18290 392475 -18234
rect 392531 -18290 392608 -18234
rect 392268 -18376 392608 -18290
rect 392268 -18432 392333 -18376
rect 392389 -18432 392475 -18376
rect 392531 -18432 392608 -18376
rect 392268 -18518 392608 -18432
rect 392268 -18574 392333 -18518
rect 392389 -18574 392475 -18518
rect 392531 -18574 392608 -18518
rect 392268 -18660 392608 -18574
rect 392268 -18716 392333 -18660
rect 392389 -18716 392475 -18660
rect 392531 -18716 392608 -18660
rect 392268 -18802 392608 -18716
rect 392268 -18858 392333 -18802
rect 392389 -18858 392475 -18802
rect 392531 -18858 392608 -18802
rect 392268 -18944 392608 -18858
rect 392268 -19000 392333 -18944
rect 392389 -19000 392475 -18944
rect 392531 -19000 392608 -18944
rect 392268 -19086 392608 -19000
rect 392268 -19142 392333 -19086
rect 392389 -19142 392475 -19086
rect 392531 -19142 392608 -19086
rect 392268 -19228 392608 -19142
rect 392268 -19284 392333 -19228
rect 392389 -19284 392475 -19228
rect 392531 -19284 392608 -19228
rect 392268 -19370 392608 -19284
rect 392268 -19426 392333 -19370
rect 392389 -19426 392475 -19370
rect 392531 -19426 392608 -19370
rect 392268 -19512 392608 -19426
rect 392268 -19568 392333 -19512
rect 392389 -19568 392475 -19512
rect 392531 -19568 392608 -19512
rect 392268 -19654 392608 -19568
rect 392268 -19710 392333 -19654
rect 392389 -19710 392475 -19654
rect 392531 -19710 392608 -19654
rect 392268 -19796 392608 -19710
rect 392268 -19852 392333 -19796
rect 392389 -19852 392475 -19796
rect 392531 -19852 392608 -19796
rect 392268 -19938 392608 -19852
rect 392268 -19994 392333 -19938
rect 392389 -19994 392475 -19938
rect 392531 -19994 392608 -19938
rect 392268 -20080 392608 -19994
rect 392268 -20136 392333 -20080
rect 392389 -20136 392475 -20080
rect 392531 -20136 392608 -20080
rect 392268 -20222 392608 -20136
rect 392268 -20278 392333 -20222
rect 392389 -20278 392475 -20222
rect 392531 -20278 392608 -20222
rect 392268 -20364 392608 -20278
rect 392268 -20420 392333 -20364
rect 392389 -20420 392475 -20364
rect 392531 -20420 392608 -20364
rect 392268 -20506 392608 -20420
rect 392268 -20562 392333 -20506
rect 392389 -20562 392475 -20506
rect 392531 -20562 392608 -20506
rect 392268 -20648 392608 -20562
rect 392268 -20704 392333 -20648
rect 392389 -20704 392475 -20648
rect 392531 -20704 392608 -20648
rect 392268 -20790 392608 -20704
rect 392268 -20846 392333 -20790
rect 392389 -20846 392475 -20790
rect 392531 -20846 392608 -20790
rect 392268 -20932 392608 -20846
rect 392268 -20988 392333 -20932
rect 392389 -20988 392475 -20932
rect 392531 -20988 392608 -20932
rect 392268 -21074 392608 -20988
rect 392268 -21130 392333 -21074
rect 392389 -21130 392475 -21074
rect 392531 -21130 392608 -21074
rect 392268 -21216 392608 -21130
rect 392268 -21272 392333 -21216
rect 392389 -21272 392475 -21216
rect 392531 -21272 392608 -21216
rect 392268 -21358 392608 -21272
rect 392268 -21414 392333 -21358
rect 392389 -21414 392475 -21358
rect 392531 -21414 392608 -21358
rect 392268 -21500 392608 -21414
rect 392268 -21556 392333 -21500
rect 392389 -21556 392475 -21500
rect 392531 -21556 392608 -21500
rect 392268 -21642 392608 -21556
rect 392268 -21698 392333 -21642
rect 392389 -21698 392475 -21642
rect 392531 -21698 392608 -21642
rect 392268 -21784 392608 -21698
rect 392268 -21840 392333 -21784
rect 392389 -21840 392475 -21784
rect 392531 -21840 392608 -21784
rect 392268 -21926 392608 -21840
rect 392268 -21982 392333 -21926
rect 392389 -21982 392475 -21926
rect 392531 -21982 392608 -21926
rect 392268 -22068 392608 -21982
rect 392268 -22124 392333 -22068
rect 392389 -22124 392475 -22068
rect 392531 -22124 392608 -22068
rect 392268 -22210 392608 -22124
rect 392268 -22266 392333 -22210
rect 392389 -22266 392475 -22210
rect 392531 -22266 392608 -22210
rect 392268 -22352 392608 -22266
rect 392268 -22408 392333 -22352
rect 392389 -22408 392475 -22352
rect 392531 -22408 392608 -22352
rect 392268 -22494 392608 -22408
rect 392268 -22550 392333 -22494
rect 392389 -22550 392475 -22494
rect 392531 -22550 392608 -22494
rect 392268 -22636 392608 -22550
rect 392268 -22692 392333 -22636
rect 392389 -22692 392475 -22636
rect 392531 -22692 392608 -22636
rect 392268 -22778 392608 -22692
rect 392268 -22834 392333 -22778
rect 392389 -22834 392475 -22778
rect 392531 -22834 392608 -22778
rect 392268 -22920 392608 -22834
rect 392268 -22976 392333 -22920
rect 392389 -22976 392475 -22920
rect 392531 -22976 392608 -22920
rect 392268 -23062 392608 -22976
rect 392268 -23118 392333 -23062
rect 392389 -23118 392475 -23062
rect 392531 -23118 392608 -23062
rect 392268 -23204 392608 -23118
rect 392268 -23260 392333 -23204
rect 392389 -23260 392475 -23204
rect 392531 -23260 392608 -23204
rect 392268 -23346 392608 -23260
rect 392268 -23402 392333 -23346
rect 392389 -23402 392475 -23346
rect 392531 -23402 392608 -23346
rect 392268 -23488 392608 -23402
rect 392268 -23544 392333 -23488
rect 392389 -23544 392475 -23488
rect 392531 -23544 392608 -23488
rect 392268 -23630 392608 -23544
rect 392268 -23686 392333 -23630
rect 392389 -23686 392475 -23630
rect 392531 -23686 392608 -23630
rect 392268 -23772 392608 -23686
rect 392268 -23828 392333 -23772
rect 392389 -23828 392475 -23772
rect 392531 -23828 392608 -23772
rect 392268 -23914 392608 -23828
rect 392268 -23970 392333 -23914
rect 392389 -23970 392475 -23914
rect 392531 -23970 392608 -23914
rect 392268 -24056 392608 -23970
rect 392268 -24112 392333 -24056
rect 392389 -24112 392475 -24056
rect 392531 -24112 392608 -24056
rect 392268 -24198 392608 -24112
rect 392268 -24254 392333 -24198
rect 392389 -24254 392475 -24198
rect 392531 -24254 392608 -24198
rect 392268 -24340 392608 -24254
rect 392268 -24396 392333 -24340
rect 392389 -24396 392475 -24340
rect 392531 -24396 392608 -24340
rect 392268 -24482 392608 -24396
rect 392268 -24538 392333 -24482
rect 392389 -24538 392475 -24482
rect 392531 -24538 392608 -24482
rect 392268 -24624 392608 -24538
rect 392268 -24680 392333 -24624
rect 392389 -24680 392475 -24624
rect 392531 -24680 392608 -24624
rect 392268 -24766 392608 -24680
rect 392268 -24822 392333 -24766
rect 392389 -24822 392475 -24766
rect 392531 -24822 392608 -24766
rect 392268 -24908 392608 -24822
rect 392268 -24964 392333 -24908
rect 392389 -24964 392475 -24908
rect 392531 -24964 392608 -24908
rect 392268 -25050 392608 -24964
rect 392268 -25106 392333 -25050
rect 392389 -25106 392475 -25050
rect 392531 -25106 392608 -25050
rect 392268 -25192 392608 -25106
rect 392268 -25248 392333 -25192
rect 392389 -25248 392475 -25192
rect 392531 -25248 392608 -25192
rect 392268 -25334 392608 -25248
rect 392268 -25390 392333 -25334
rect 392389 -25390 392475 -25334
rect 392531 -25390 392608 -25334
rect 392268 -25476 392608 -25390
rect 392268 -25532 392333 -25476
rect 392389 -25532 392475 -25476
rect 392531 -25532 392608 -25476
rect 392268 -25542 392608 -25532
rect 392668 -17950 393008 -17820
rect 392668 -18006 392738 -17950
rect 392794 -18006 392880 -17950
rect 392936 -18006 393008 -17950
rect 392668 -18092 393008 -18006
rect 392668 -18148 392738 -18092
rect 392794 -18148 392880 -18092
rect 392936 -18148 393008 -18092
rect 392668 -18234 393008 -18148
rect 392668 -18290 392738 -18234
rect 392794 -18290 392880 -18234
rect 392936 -18290 393008 -18234
rect 392668 -18376 393008 -18290
rect 392668 -18432 392738 -18376
rect 392794 -18432 392880 -18376
rect 392936 -18432 393008 -18376
rect 392668 -18518 393008 -18432
rect 392668 -18574 392738 -18518
rect 392794 -18574 392880 -18518
rect 392936 -18574 393008 -18518
rect 392668 -18660 393008 -18574
rect 392668 -18716 392738 -18660
rect 392794 -18716 392880 -18660
rect 392936 -18716 393008 -18660
rect 392668 -18802 393008 -18716
rect 392668 -18858 392738 -18802
rect 392794 -18858 392880 -18802
rect 392936 -18858 393008 -18802
rect 392668 -18944 393008 -18858
rect 392668 -19000 392738 -18944
rect 392794 -19000 392880 -18944
rect 392936 -19000 393008 -18944
rect 392668 -19086 393008 -19000
rect 392668 -19142 392738 -19086
rect 392794 -19142 392880 -19086
rect 392936 -19142 393008 -19086
rect 392668 -19228 393008 -19142
rect 392668 -19284 392738 -19228
rect 392794 -19284 392880 -19228
rect 392936 -19284 393008 -19228
rect 392668 -19370 393008 -19284
rect 392668 -19426 392738 -19370
rect 392794 -19426 392880 -19370
rect 392936 -19426 393008 -19370
rect 392668 -19512 393008 -19426
rect 392668 -19568 392738 -19512
rect 392794 -19568 392880 -19512
rect 392936 -19568 393008 -19512
rect 392668 -19654 393008 -19568
rect 392668 -19710 392738 -19654
rect 392794 -19710 392880 -19654
rect 392936 -19710 393008 -19654
rect 392668 -19796 393008 -19710
rect 392668 -19852 392738 -19796
rect 392794 -19852 392880 -19796
rect 392936 -19852 393008 -19796
rect 392668 -19938 393008 -19852
rect 392668 -19994 392738 -19938
rect 392794 -19994 392880 -19938
rect 392936 -19994 393008 -19938
rect 392668 -20080 393008 -19994
rect 392668 -20136 392738 -20080
rect 392794 -20136 392880 -20080
rect 392936 -20136 393008 -20080
rect 392668 -20222 393008 -20136
rect 392668 -20278 392738 -20222
rect 392794 -20278 392880 -20222
rect 392936 -20278 393008 -20222
rect 392668 -20364 393008 -20278
rect 392668 -20420 392738 -20364
rect 392794 -20420 392880 -20364
rect 392936 -20420 393008 -20364
rect 392668 -20506 393008 -20420
rect 392668 -20562 392738 -20506
rect 392794 -20562 392880 -20506
rect 392936 -20562 393008 -20506
rect 392668 -20648 393008 -20562
rect 392668 -20704 392738 -20648
rect 392794 -20704 392880 -20648
rect 392936 -20704 393008 -20648
rect 392668 -20790 393008 -20704
rect 392668 -20846 392738 -20790
rect 392794 -20846 392880 -20790
rect 392936 -20846 393008 -20790
rect 392668 -20932 393008 -20846
rect 392668 -20988 392738 -20932
rect 392794 -20988 392880 -20932
rect 392936 -20988 393008 -20932
rect 392668 -21074 393008 -20988
rect 392668 -21130 392738 -21074
rect 392794 -21130 392880 -21074
rect 392936 -21130 393008 -21074
rect 392668 -21216 393008 -21130
rect 392668 -21272 392738 -21216
rect 392794 -21272 392880 -21216
rect 392936 -21272 393008 -21216
rect 392668 -21358 393008 -21272
rect 392668 -21414 392738 -21358
rect 392794 -21414 392880 -21358
rect 392936 -21414 393008 -21358
rect 392668 -21500 393008 -21414
rect 392668 -21556 392738 -21500
rect 392794 -21556 392880 -21500
rect 392936 -21556 393008 -21500
rect 392668 -21642 393008 -21556
rect 392668 -21698 392738 -21642
rect 392794 -21698 392880 -21642
rect 392936 -21698 393008 -21642
rect 392668 -21784 393008 -21698
rect 392668 -21840 392738 -21784
rect 392794 -21840 392880 -21784
rect 392936 -21840 393008 -21784
rect 392668 -21926 393008 -21840
rect 392668 -21982 392738 -21926
rect 392794 -21982 392880 -21926
rect 392936 -21982 393008 -21926
rect 392668 -22068 393008 -21982
rect 392668 -22124 392738 -22068
rect 392794 -22124 392880 -22068
rect 392936 -22124 393008 -22068
rect 392668 -22210 393008 -22124
rect 392668 -22266 392738 -22210
rect 392794 -22266 392880 -22210
rect 392936 -22266 393008 -22210
rect 392668 -22352 393008 -22266
rect 392668 -22408 392738 -22352
rect 392794 -22408 392880 -22352
rect 392936 -22408 393008 -22352
rect 392668 -22494 393008 -22408
rect 392668 -22550 392738 -22494
rect 392794 -22550 392880 -22494
rect 392936 -22550 393008 -22494
rect 392668 -22636 393008 -22550
rect 392668 -22692 392738 -22636
rect 392794 -22692 392880 -22636
rect 392936 -22692 393008 -22636
rect 392668 -22778 393008 -22692
rect 392668 -22834 392738 -22778
rect 392794 -22834 392880 -22778
rect 392936 -22834 393008 -22778
rect 392668 -22920 393008 -22834
rect 392668 -22976 392738 -22920
rect 392794 -22976 392880 -22920
rect 392936 -22976 393008 -22920
rect 392668 -23062 393008 -22976
rect 392668 -23118 392738 -23062
rect 392794 -23118 392880 -23062
rect 392936 -23118 393008 -23062
rect 392668 -23204 393008 -23118
rect 392668 -23260 392738 -23204
rect 392794 -23260 392880 -23204
rect 392936 -23260 393008 -23204
rect 392668 -23346 393008 -23260
rect 392668 -23402 392738 -23346
rect 392794 -23402 392880 -23346
rect 392936 -23402 393008 -23346
rect 392668 -23488 393008 -23402
rect 392668 -23544 392738 -23488
rect 392794 -23544 392880 -23488
rect 392936 -23544 393008 -23488
rect 392668 -23630 393008 -23544
rect 392668 -23686 392738 -23630
rect 392794 -23686 392880 -23630
rect 392936 -23686 393008 -23630
rect 392668 -23772 393008 -23686
rect 392668 -23828 392738 -23772
rect 392794 -23828 392880 -23772
rect 392936 -23828 393008 -23772
rect 392668 -23914 393008 -23828
rect 392668 -23970 392738 -23914
rect 392794 -23970 392880 -23914
rect 392936 -23970 393008 -23914
rect 392668 -24056 393008 -23970
rect 392668 -24112 392738 -24056
rect 392794 -24112 392880 -24056
rect 392936 -24112 393008 -24056
rect 392668 -24198 393008 -24112
rect 392668 -24254 392738 -24198
rect 392794 -24254 392880 -24198
rect 392936 -24254 393008 -24198
rect 392668 -24340 393008 -24254
rect 392668 -24396 392738 -24340
rect 392794 -24396 392880 -24340
rect 392936 -24396 393008 -24340
rect 392668 -24482 393008 -24396
rect 392668 -24538 392738 -24482
rect 392794 -24538 392880 -24482
rect 392936 -24538 393008 -24482
rect 392668 -24624 393008 -24538
rect 392668 -24680 392738 -24624
rect 392794 -24680 392880 -24624
rect 392936 -24680 393008 -24624
rect 392668 -24766 393008 -24680
rect 392668 -24822 392738 -24766
rect 392794 -24822 392880 -24766
rect 392936 -24822 393008 -24766
rect 392668 -24908 393008 -24822
rect 392668 -24964 392738 -24908
rect 392794 -24964 392880 -24908
rect 392936 -24964 393008 -24908
rect 392668 -25050 393008 -24964
rect 392668 -25106 392738 -25050
rect 392794 -25106 392880 -25050
rect 392936 -25106 393008 -25050
rect 392668 -25192 393008 -25106
rect 392668 -25248 392738 -25192
rect 392794 -25248 392880 -25192
rect 392936 -25248 393008 -25192
rect 392668 -25334 393008 -25248
rect 392668 -25390 392738 -25334
rect 392794 -25390 392880 -25334
rect 392936 -25390 393008 -25334
rect 392668 -25476 393008 -25390
rect 392668 -25532 392738 -25476
rect 392794 -25532 392880 -25476
rect 392936 -25532 393008 -25476
rect 392668 -25542 393008 -25532
rect 393068 -17950 393408 -17820
rect 393068 -18006 393138 -17950
rect 393194 -18006 393280 -17950
rect 393336 -18006 393408 -17950
rect 393068 -18092 393408 -18006
rect 393068 -18148 393138 -18092
rect 393194 -18148 393280 -18092
rect 393336 -18148 393408 -18092
rect 393068 -18234 393408 -18148
rect 393068 -18290 393138 -18234
rect 393194 -18290 393280 -18234
rect 393336 -18290 393408 -18234
rect 393068 -18376 393408 -18290
rect 393068 -18432 393138 -18376
rect 393194 -18432 393280 -18376
rect 393336 -18432 393408 -18376
rect 393068 -18518 393408 -18432
rect 393068 -18574 393138 -18518
rect 393194 -18574 393280 -18518
rect 393336 -18574 393408 -18518
rect 393068 -18660 393408 -18574
rect 393068 -18716 393138 -18660
rect 393194 -18716 393280 -18660
rect 393336 -18716 393408 -18660
rect 393068 -18802 393408 -18716
rect 393068 -18858 393138 -18802
rect 393194 -18858 393280 -18802
rect 393336 -18858 393408 -18802
rect 393068 -18944 393408 -18858
rect 393068 -19000 393138 -18944
rect 393194 -19000 393280 -18944
rect 393336 -19000 393408 -18944
rect 393068 -19086 393408 -19000
rect 393068 -19142 393138 -19086
rect 393194 -19142 393280 -19086
rect 393336 -19142 393408 -19086
rect 393068 -19228 393408 -19142
rect 393068 -19284 393138 -19228
rect 393194 -19284 393280 -19228
rect 393336 -19284 393408 -19228
rect 393068 -19370 393408 -19284
rect 393068 -19426 393138 -19370
rect 393194 -19426 393280 -19370
rect 393336 -19426 393408 -19370
rect 393068 -19512 393408 -19426
rect 393068 -19568 393138 -19512
rect 393194 -19568 393280 -19512
rect 393336 -19568 393408 -19512
rect 393068 -19654 393408 -19568
rect 393068 -19710 393138 -19654
rect 393194 -19710 393280 -19654
rect 393336 -19710 393408 -19654
rect 393068 -19796 393408 -19710
rect 393068 -19852 393138 -19796
rect 393194 -19852 393280 -19796
rect 393336 -19852 393408 -19796
rect 393068 -19938 393408 -19852
rect 393068 -19994 393138 -19938
rect 393194 -19994 393280 -19938
rect 393336 -19994 393408 -19938
rect 393068 -20080 393408 -19994
rect 393068 -20136 393138 -20080
rect 393194 -20136 393280 -20080
rect 393336 -20136 393408 -20080
rect 393068 -20222 393408 -20136
rect 393068 -20278 393138 -20222
rect 393194 -20278 393280 -20222
rect 393336 -20278 393408 -20222
rect 393068 -20364 393408 -20278
rect 393068 -20420 393138 -20364
rect 393194 -20420 393280 -20364
rect 393336 -20420 393408 -20364
rect 393068 -20506 393408 -20420
rect 393068 -20562 393138 -20506
rect 393194 -20562 393280 -20506
rect 393336 -20562 393408 -20506
rect 393068 -20648 393408 -20562
rect 393068 -20704 393138 -20648
rect 393194 -20704 393280 -20648
rect 393336 -20704 393408 -20648
rect 393068 -20790 393408 -20704
rect 393068 -20846 393138 -20790
rect 393194 -20846 393280 -20790
rect 393336 -20846 393408 -20790
rect 393068 -20932 393408 -20846
rect 393068 -20988 393138 -20932
rect 393194 -20988 393280 -20932
rect 393336 -20988 393408 -20932
rect 393068 -21074 393408 -20988
rect 393068 -21130 393138 -21074
rect 393194 -21130 393280 -21074
rect 393336 -21130 393408 -21074
rect 393068 -21216 393408 -21130
rect 393068 -21272 393138 -21216
rect 393194 -21272 393280 -21216
rect 393336 -21272 393408 -21216
rect 393068 -21358 393408 -21272
rect 393068 -21414 393138 -21358
rect 393194 -21414 393280 -21358
rect 393336 -21414 393408 -21358
rect 393068 -21500 393408 -21414
rect 393068 -21556 393138 -21500
rect 393194 -21556 393280 -21500
rect 393336 -21556 393408 -21500
rect 393068 -21642 393408 -21556
rect 393068 -21698 393138 -21642
rect 393194 -21698 393280 -21642
rect 393336 -21698 393408 -21642
rect 393068 -21784 393408 -21698
rect 393068 -21840 393138 -21784
rect 393194 -21840 393280 -21784
rect 393336 -21840 393408 -21784
rect 393068 -21926 393408 -21840
rect 393068 -21982 393138 -21926
rect 393194 -21982 393280 -21926
rect 393336 -21982 393408 -21926
rect 393068 -22068 393408 -21982
rect 393068 -22124 393138 -22068
rect 393194 -22124 393280 -22068
rect 393336 -22124 393408 -22068
rect 393068 -22210 393408 -22124
rect 393068 -22266 393138 -22210
rect 393194 -22266 393280 -22210
rect 393336 -22266 393408 -22210
rect 393068 -22352 393408 -22266
rect 393068 -22408 393138 -22352
rect 393194 -22408 393280 -22352
rect 393336 -22408 393408 -22352
rect 393068 -22494 393408 -22408
rect 393068 -22550 393138 -22494
rect 393194 -22550 393280 -22494
rect 393336 -22550 393408 -22494
rect 393068 -22636 393408 -22550
rect 393068 -22692 393138 -22636
rect 393194 -22692 393280 -22636
rect 393336 -22692 393408 -22636
rect 393068 -22778 393408 -22692
rect 393068 -22834 393138 -22778
rect 393194 -22834 393280 -22778
rect 393336 -22834 393408 -22778
rect 393068 -22920 393408 -22834
rect 393068 -22976 393138 -22920
rect 393194 -22976 393280 -22920
rect 393336 -22976 393408 -22920
rect 393068 -23062 393408 -22976
rect 393068 -23118 393138 -23062
rect 393194 -23118 393280 -23062
rect 393336 -23118 393408 -23062
rect 393068 -23204 393408 -23118
rect 393068 -23260 393138 -23204
rect 393194 -23260 393280 -23204
rect 393336 -23260 393408 -23204
rect 393068 -23346 393408 -23260
rect 393068 -23402 393138 -23346
rect 393194 -23402 393280 -23346
rect 393336 -23402 393408 -23346
rect 393068 -23488 393408 -23402
rect 393068 -23544 393138 -23488
rect 393194 -23544 393280 -23488
rect 393336 -23544 393408 -23488
rect 393068 -23630 393408 -23544
rect 393068 -23686 393138 -23630
rect 393194 -23686 393280 -23630
rect 393336 -23686 393408 -23630
rect 393068 -23772 393408 -23686
rect 393068 -23828 393138 -23772
rect 393194 -23828 393280 -23772
rect 393336 -23828 393408 -23772
rect 393068 -23914 393408 -23828
rect 393068 -23970 393138 -23914
rect 393194 -23970 393280 -23914
rect 393336 -23970 393408 -23914
rect 393068 -24056 393408 -23970
rect 393068 -24112 393138 -24056
rect 393194 -24112 393280 -24056
rect 393336 -24112 393408 -24056
rect 393068 -24198 393408 -24112
rect 393068 -24254 393138 -24198
rect 393194 -24254 393280 -24198
rect 393336 -24254 393408 -24198
rect 393068 -24340 393408 -24254
rect 393068 -24396 393138 -24340
rect 393194 -24396 393280 -24340
rect 393336 -24396 393408 -24340
rect 393068 -24482 393408 -24396
rect 393068 -24538 393138 -24482
rect 393194 -24538 393280 -24482
rect 393336 -24538 393408 -24482
rect 393068 -24624 393408 -24538
rect 393068 -24680 393138 -24624
rect 393194 -24680 393280 -24624
rect 393336 -24680 393408 -24624
rect 393068 -24766 393408 -24680
rect 393068 -24822 393138 -24766
rect 393194 -24822 393280 -24766
rect 393336 -24822 393408 -24766
rect 393068 -24908 393408 -24822
rect 393068 -24964 393138 -24908
rect 393194 -24964 393280 -24908
rect 393336 -24964 393408 -24908
rect 393068 -25050 393408 -24964
rect 393068 -25106 393138 -25050
rect 393194 -25106 393280 -25050
rect 393336 -25106 393408 -25050
rect 393068 -25192 393408 -25106
rect 393068 -25248 393138 -25192
rect 393194 -25248 393280 -25192
rect 393336 -25248 393408 -25192
rect 393068 -25334 393408 -25248
rect 393068 -25390 393138 -25334
rect 393194 -25390 393280 -25334
rect 393336 -25390 393408 -25334
rect 393068 -25476 393408 -25390
rect 393068 -25532 393138 -25476
rect 393194 -25532 393280 -25476
rect 393336 -25532 393408 -25476
rect 393068 -25542 393408 -25532
rect 393468 -17950 393808 -17820
rect 393468 -18006 393543 -17950
rect 393599 -18006 393685 -17950
rect 393741 -18006 393808 -17950
rect 393468 -18092 393808 -18006
rect 393468 -18148 393543 -18092
rect 393599 -18148 393685 -18092
rect 393741 -18148 393808 -18092
rect 393468 -18234 393808 -18148
rect 393468 -18290 393543 -18234
rect 393599 -18290 393685 -18234
rect 393741 -18290 393808 -18234
rect 393468 -18376 393808 -18290
rect 393468 -18432 393543 -18376
rect 393599 -18432 393685 -18376
rect 393741 -18432 393808 -18376
rect 393468 -18518 393808 -18432
rect 393468 -18574 393543 -18518
rect 393599 -18574 393685 -18518
rect 393741 -18574 393808 -18518
rect 393468 -18660 393808 -18574
rect 393468 -18716 393543 -18660
rect 393599 -18716 393685 -18660
rect 393741 -18716 393808 -18660
rect 393468 -18802 393808 -18716
rect 393468 -18858 393543 -18802
rect 393599 -18858 393685 -18802
rect 393741 -18858 393808 -18802
rect 393468 -18944 393808 -18858
rect 393468 -19000 393543 -18944
rect 393599 -19000 393685 -18944
rect 393741 -19000 393808 -18944
rect 393468 -19086 393808 -19000
rect 393468 -19142 393543 -19086
rect 393599 -19142 393685 -19086
rect 393741 -19142 393808 -19086
rect 393468 -19228 393808 -19142
rect 393468 -19284 393543 -19228
rect 393599 -19284 393685 -19228
rect 393741 -19284 393808 -19228
rect 393468 -19370 393808 -19284
rect 393468 -19426 393543 -19370
rect 393599 -19426 393685 -19370
rect 393741 -19426 393808 -19370
rect 393468 -19512 393808 -19426
rect 393468 -19568 393543 -19512
rect 393599 -19568 393685 -19512
rect 393741 -19568 393808 -19512
rect 393468 -19654 393808 -19568
rect 393468 -19710 393543 -19654
rect 393599 -19710 393685 -19654
rect 393741 -19710 393808 -19654
rect 393468 -19796 393808 -19710
rect 393468 -19852 393543 -19796
rect 393599 -19852 393685 -19796
rect 393741 -19852 393808 -19796
rect 393468 -19938 393808 -19852
rect 393468 -19994 393543 -19938
rect 393599 -19994 393685 -19938
rect 393741 -19994 393808 -19938
rect 393468 -20080 393808 -19994
rect 393468 -20136 393543 -20080
rect 393599 -20136 393685 -20080
rect 393741 -20136 393808 -20080
rect 393468 -20222 393808 -20136
rect 393468 -20278 393543 -20222
rect 393599 -20278 393685 -20222
rect 393741 -20278 393808 -20222
rect 393468 -20364 393808 -20278
rect 393468 -20420 393543 -20364
rect 393599 -20420 393685 -20364
rect 393741 -20420 393808 -20364
rect 393468 -20506 393808 -20420
rect 393468 -20562 393543 -20506
rect 393599 -20562 393685 -20506
rect 393741 -20562 393808 -20506
rect 393468 -20648 393808 -20562
rect 393468 -20704 393543 -20648
rect 393599 -20704 393685 -20648
rect 393741 -20704 393808 -20648
rect 393468 -20790 393808 -20704
rect 393468 -20846 393543 -20790
rect 393599 -20846 393685 -20790
rect 393741 -20846 393808 -20790
rect 393468 -20932 393808 -20846
rect 393468 -20988 393543 -20932
rect 393599 -20988 393685 -20932
rect 393741 -20988 393808 -20932
rect 393468 -21074 393808 -20988
rect 393468 -21130 393543 -21074
rect 393599 -21130 393685 -21074
rect 393741 -21130 393808 -21074
rect 393468 -21216 393808 -21130
rect 393468 -21272 393543 -21216
rect 393599 -21272 393685 -21216
rect 393741 -21272 393808 -21216
rect 393468 -21358 393808 -21272
rect 393468 -21414 393543 -21358
rect 393599 -21414 393685 -21358
rect 393741 -21414 393808 -21358
rect 393468 -21500 393808 -21414
rect 393468 -21556 393543 -21500
rect 393599 -21556 393685 -21500
rect 393741 -21556 393808 -21500
rect 393468 -21642 393808 -21556
rect 393468 -21698 393543 -21642
rect 393599 -21698 393685 -21642
rect 393741 -21698 393808 -21642
rect 393468 -21784 393808 -21698
rect 393468 -21840 393543 -21784
rect 393599 -21840 393685 -21784
rect 393741 -21840 393808 -21784
rect 393468 -21926 393808 -21840
rect 393468 -21982 393543 -21926
rect 393599 -21982 393685 -21926
rect 393741 -21982 393808 -21926
rect 393468 -22068 393808 -21982
rect 393468 -22124 393543 -22068
rect 393599 -22124 393685 -22068
rect 393741 -22124 393808 -22068
rect 393468 -22210 393808 -22124
rect 393468 -22266 393543 -22210
rect 393599 -22266 393685 -22210
rect 393741 -22266 393808 -22210
rect 393468 -22352 393808 -22266
rect 393468 -22408 393543 -22352
rect 393599 -22408 393685 -22352
rect 393741 -22408 393808 -22352
rect 393468 -22494 393808 -22408
rect 393468 -22550 393543 -22494
rect 393599 -22550 393685 -22494
rect 393741 -22550 393808 -22494
rect 393468 -22636 393808 -22550
rect 393468 -22692 393543 -22636
rect 393599 -22692 393685 -22636
rect 393741 -22692 393808 -22636
rect 393468 -22778 393808 -22692
rect 393468 -22834 393543 -22778
rect 393599 -22834 393685 -22778
rect 393741 -22834 393808 -22778
rect 393468 -22920 393808 -22834
rect 393468 -22976 393543 -22920
rect 393599 -22976 393685 -22920
rect 393741 -22976 393808 -22920
rect 393468 -23062 393808 -22976
rect 393468 -23118 393543 -23062
rect 393599 -23118 393685 -23062
rect 393741 -23118 393808 -23062
rect 393468 -23204 393808 -23118
rect 393468 -23260 393543 -23204
rect 393599 -23260 393685 -23204
rect 393741 -23260 393808 -23204
rect 393468 -23346 393808 -23260
rect 393468 -23402 393543 -23346
rect 393599 -23402 393685 -23346
rect 393741 -23402 393808 -23346
rect 393468 -23488 393808 -23402
rect 393468 -23544 393543 -23488
rect 393599 -23544 393685 -23488
rect 393741 -23544 393808 -23488
rect 393468 -23630 393808 -23544
rect 393468 -23686 393543 -23630
rect 393599 -23686 393685 -23630
rect 393741 -23686 393808 -23630
rect 393468 -23772 393808 -23686
rect 393468 -23828 393543 -23772
rect 393599 -23828 393685 -23772
rect 393741 -23828 393808 -23772
rect 393468 -23914 393808 -23828
rect 393468 -23970 393543 -23914
rect 393599 -23970 393685 -23914
rect 393741 -23970 393808 -23914
rect 393468 -24056 393808 -23970
rect 393468 -24112 393543 -24056
rect 393599 -24112 393685 -24056
rect 393741 -24112 393808 -24056
rect 393468 -24198 393808 -24112
rect 393468 -24254 393543 -24198
rect 393599 -24254 393685 -24198
rect 393741 -24254 393808 -24198
rect 393468 -24340 393808 -24254
rect 393468 -24396 393543 -24340
rect 393599 -24396 393685 -24340
rect 393741 -24396 393808 -24340
rect 393468 -24482 393808 -24396
rect 393468 -24538 393543 -24482
rect 393599 -24538 393685 -24482
rect 393741 -24538 393808 -24482
rect 393468 -24624 393808 -24538
rect 393468 -24680 393543 -24624
rect 393599 -24680 393685 -24624
rect 393741 -24680 393808 -24624
rect 393468 -24766 393808 -24680
rect 393468 -24822 393543 -24766
rect 393599 -24822 393685 -24766
rect 393741 -24822 393808 -24766
rect 393468 -24908 393808 -24822
rect 393468 -24964 393543 -24908
rect 393599 -24964 393685 -24908
rect 393741 -24964 393808 -24908
rect 393468 -25050 393808 -24964
rect 393468 -25106 393543 -25050
rect 393599 -25106 393685 -25050
rect 393741 -25106 393808 -25050
rect 393468 -25192 393808 -25106
rect 393468 -25248 393543 -25192
rect 393599 -25248 393685 -25192
rect 393741 -25248 393808 -25192
rect 393468 -25334 393808 -25248
rect 393468 -25390 393543 -25334
rect 393599 -25390 393685 -25334
rect 393741 -25390 393808 -25334
rect 393468 -25476 393808 -25390
rect 393468 -25532 393543 -25476
rect 393599 -25532 393685 -25476
rect 393741 -25532 393808 -25476
rect 393468 -25542 393808 -25532
rect 393868 -17950 394208 -17820
rect 393868 -18006 393940 -17950
rect 393996 -18006 394082 -17950
rect 394138 -18006 394208 -17950
rect 393868 -18092 394208 -18006
rect 393868 -18148 393940 -18092
rect 393996 -18148 394082 -18092
rect 394138 -18148 394208 -18092
rect 393868 -18234 394208 -18148
rect 393868 -18290 393940 -18234
rect 393996 -18290 394082 -18234
rect 394138 -18290 394208 -18234
rect 393868 -18376 394208 -18290
rect 393868 -18432 393940 -18376
rect 393996 -18432 394082 -18376
rect 394138 -18432 394208 -18376
rect 393868 -18518 394208 -18432
rect 393868 -18574 393940 -18518
rect 393996 -18574 394082 -18518
rect 394138 -18574 394208 -18518
rect 393868 -18660 394208 -18574
rect 393868 -18716 393940 -18660
rect 393996 -18716 394082 -18660
rect 394138 -18716 394208 -18660
rect 393868 -18802 394208 -18716
rect 393868 -18858 393940 -18802
rect 393996 -18858 394082 -18802
rect 394138 -18858 394208 -18802
rect 393868 -18944 394208 -18858
rect 393868 -19000 393940 -18944
rect 393996 -19000 394082 -18944
rect 394138 -19000 394208 -18944
rect 393868 -19086 394208 -19000
rect 393868 -19142 393940 -19086
rect 393996 -19142 394082 -19086
rect 394138 -19142 394208 -19086
rect 393868 -19228 394208 -19142
rect 393868 -19284 393940 -19228
rect 393996 -19284 394082 -19228
rect 394138 -19284 394208 -19228
rect 393868 -19370 394208 -19284
rect 393868 -19426 393940 -19370
rect 393996 -19426 394082 -19370
rect 394138 -19426 394208 -19370
rect 393868 -19512 394208 -19426
rect 393868 -19568 393940 -19512
rect 393996 -19568 394082 -19512
rect 394138 -19568 394208 -19512
rect 393868 -19654 394208 -19568
rect 393868 -19710 393940 -19654
rect 393996 -19710 394082 -19654
rect 394138 -19710 394208 -19654
rect 393868 -19796 394208 -19710
rect 393868 -19852 393940 -19796
rect 393996 -19852 394082 -19796
rect 394138 -19852 394208 -19796
rect 393868 -19938 394208 -19852
rect 393868 -19994 393940 -19938
rect 393996 -19994 394082 -19938
rect 394138 -19994 394208 -19938
rect 393868 -20080 394208 -19994
rect 393868 -20136 393940 -20080
rect 393996 -20136 394082 -20080
rect 394138 -20136 394208 -20080
rect 393868 -20222 394208 -20136
rect 393868 -20278 393940 -20222
rect 393996 -20278 394082 -20222
rect 394138 -20278 394208 -20222
rect 393868 -20364 394208 -20278
rect 393868 -20420 393940 -20364
rect 393996 -20420 394082 -20364
rect 394138 -20420 394208 -20364
rect 393868 -20506 394208 -20420
rect 393868 -20562 393940 -20506
rect 393996 -20562 394082 -20506
rect 394138 -20562 394208 -20506
rect 393868 -20648 394208 -20562
rect 393868 -20704 393940 -20648
rect 393996 -20704 394082 -20648
rect 394138 -20704 394208 -20648
rect 393868 -20790 394208 -20704
rect 393868 -20846 393940 -20790
rect 393996 -20846 394082 -20790
rect 394138 -20846 394208 -20790
rect 393868 -20932 394208 -20846
rect 393868 -20988 393940 -20932
rect 393996 -20988 394082 -20932
rect 394138 -20988 394208 -20932
rect 393868 -21074 394208 -20988
rect 393868 -21130 393940 -21074
rect 393996 -21130 394082 -21074
rect 394138 -21130 394208 -21074
rect 393868 -21216 394208 -21130
rect 393868 -21272 393940 -21216
rect 393996 -21272 394082 -21216
rect 394138 -21272 394208 -21216
rect 393868 -21358 394208 -21272
rect 393868 -21414 393940 -21358
rect 393996 -21414 394082 -21358
rect 394138 -21414 394208 -21358
rect 393868 -21500 394208 -21414
rect 393868 -21556 393940 -21500
rect 393996 -21556 394082 -21500
rect 394138 -21556 394208 -21500
rect 393868 -21642 394208 -21556
rect 393868 -21698 393940 -21642
rect 393996 -21698 394082 -21642
rect 394138 -21698 394208 -21642
rect 393868 -21784 394208 -21698
rect 393868 -21840 393940 -21784
rect 393996 -21840 394082 -21784
rect 394138 -21840 394208 -21784
rect 393868 -21926 394208 -21840
rect 393868 -21982 393940 -21926
rect 393996 -21982 394082 -21926
rect 394138 -21982 394208 -21926
rect 393868 -22068 394208 -21982
rect 393868 -22124 393940 -22068
rect 393996 -22124 394082 -22068
rect 394138 -22124 394208 -22068
rect 393868 -22210 394208 -22124
rect 393868 -22266 393940 -22210
rect 393996 -22266 394082 -22210
rect 394138 -22266 394208 -22210
rect 393868 -22352 394208 -22266
rect 393868 -22408 393940 -22352
rect 393996 -22408 394082 -22352
rect 394138 -22408 394208 -22352
rect 393868 -22494 394208 -22408
rect 393868 -22550 393940 -22494
rect 393996 -22550 394082 -22494
rect 394138 -22550 394208 -22494
rect 393868 -22636 394208 -22550
rect 393868 -22692 393940 -22636
rect 393996 -22692 394082 -22636
rect 394138 -22692 394208 -22636
rect 393868 -22778 394208 -22692
rect 393868 -22834 393940 -22778
rect 393996 -22834 394082 -22778
rect 394138 -22834 394208 -22778
rect 393868 -22920 394208 -22834
rect 393868 -22976 393940 -22920
rect 393996 -22976 394082 -22920
rect 394138 -22976 394208 -22920
rect 393868 -23062 394208 -22976
rect 393868 -23118 393940 -23062
rect 393996 -23118 394082 -23062
rect 394138 -23118 394208 -23062
rect 393868 -23204 394208 -23118
rect 393868 -23260 393940 -23204
rect 393996 -23260 394082 -23204
rect 394138 -23260 394208 -23204
rect 393868 -23346 394208 -23260
rect 393868 -23402 393940 -23346
rect 393996 -23402 394082 -23346
rect 394138 -23402 394208 -23346
rect 393868 -23488 394208 -23402
rect 393868 -23544 393940 -23488
rect 393996 -23544 394082 -23488
rect 394138 -23544 394208 -23488
rect 393868 -23630 394208 -23544
rect 393868 -23686 393940 -23630
rect 393996 -23686 394082 -23630
rect 394138 -23686 394208 -23630
rect 393868 -23772 394208 -23686
rect 393868 -23828 393940 -23772
rect 393996 -23828 394082 -23772
rect 394138 -23828 394208 -23772
rect 393868 -23914 394208 -23828
rect 393868 -23970 393940 -23914
rect 393996 -23970 394082 -23914
rect 394138 -23970 394208 -23914
rect 393868 -24056 394208 -23970
rect 393868 -24112 393940 -24056
rect 393996 -24112 394082 -24056
rect 394138 -24112 394208 -24056
rect 393868 -24198 394208 -24112
rect 393868 -24254 393940 -24198
rect 393996 -24254 394082 -24198
rect 394138 -24254 394208 -24198
rect 393868 -24340 394208 -24254
rect 393868 -24396 393940 -24340
rect 393996 -24396 394082 -24340
rect 394138 -24396 394208 -24340
rect 393868 -24482 394208 -24396
rect 393868 -24538 393940 -24482
rect 393996 -24538 394082 -24482
rect 394138 -24538 394208 -24482
rect 393868 -24624 394208 -24538
rect 393868 -24680 393940 -24624
rect 393996 -24680 394082 -24624
rect 394138 -24680 394208 -24624
rect 393868 -24766 394208 -24680
rect 393868 -24822 393940 -24766
rect 393996 -24822 394082 -24766
rect 394138 -24822 394208 -24766
rect 393868 -24908 394208 -24822
rect 393868 -24964 393940 -24908
rect 393996 -24964 394082 -24908
rect 394138 -24964 394208 -24908
rect 393868 -25050 394208 -24964
rect 393868 -25106 393940 -25050
rect 393996 -25106 394082 -25050
rect 394138 -25106 394208 -25050
rect 393868 -25192 394208 -25106
rect 393868 -25248 393940 -25192
rect 393996 -25248 394082 -25192
rect 394138 -25248 394208 -25192
rect 393868 -25334 394208 -25248
rect 393868 -25390 393940 -25334
rect 393996 -25390 394082 -25334
rect 394138 -25390 394208 -25334
rect 393868 -25476 394208 -25390
rect 393868 -25532 393940 -25476
rect 393996 -25532 394082 -25476
rect 394138 -25532 394208 -25476
rect 393868 -25542 394208 -25532
rect 394268 -17950 394608 -17820
rect 394268 -18006 394337 -17950
rect 394393 -18006 394479 -17950
rect 394535 -18006 394608 -17950
rect 394268 -18092 394608 -18006
rect 394268 -18148 394337 -18092
rect 394393 -18148 394479 -18092
rect 394535 -18148 394608 -18092
rect 394268 -18234 394608 -18148
rect 394268 -18290 394337 -18234
rect 394393 -18290 394479 -18234
rect 394535 -18290 394608 -18234
rect 394268 -18376 394608 -18290
rect 394268 -18432 394337 -18376
rect 394393 -18432 394479 -18376
rect 394535 -18432 394608 -18376
rect 394268 -18518 394608 -18432
rect 394268 -18574 394337 -18518
rect 394393 -18574 394479 -18518
rect 394535 -18574 394608 -18518
rect 394268 -18660 394608 -18574
rect 394268 -18716 394337 -18660
rect 394393 -18716 394479 -18660
rect 394535 -18716 394608 -18660
rect 394268 -18802 394608 -18716
rect 394268 -18858 394337 -18802
rect 394393 -18858 394479 -18802
rect 394535 -18858 394608 -18802
rect 394268 -18944 394608 -18858
rect 394268 -19000 394337 -18944
rect 394393 -19000 394479 -18944
rect 394535 -19000 394608 -18944
rect 394268 -19086 394608 -19000
rect 394268 -19142 394337 -19086
rect 394393 -19142 394479 -19086
rect 394535 -19142 394608 -19086
rect 394268 -19228 394608 -19142
rect 394268 -19284 394337 -19228
rect 394393 -19284 394479 -19228
rect 394535 -19284 394608 -19228
rect 394268 -19370 394608 -19284
rect 394268 -19426 394337 -19370
rect 394393 -19426 394479 -19370
rect 394535 -19426 394608 -19370
rect 394268 -19512 394608 -19426
rect 394268 -19568 394337 -19512
rect 394393 -19568 394479 -19512
rect 394535 -19568 394608 -19512
rect 394268 -19654 394608 -19568
rect 394268 -19710 394337 -19654
rect 394393 -19710 394479 -19654
rect 394535 -19710 394608 -19654
rect 394268 -19796 394608 -19710
rect 394268 -19852 394337 -19796
rect 394393 -19852 394479 -19796
rect 394535 -19852 394608 -19796
rect 394268 -19938 394608 -19852
rect 394268 -19994 394337 -19938
rect 394393 -19994 394479 -19938
rect 394535 -19994 394608 -19938
rect 394268 -20080 394608 -19994
rect 394268 -20136 394337 -20080
rect 394393 -20136 394479 -20080
rect 394535 -20136 394608 -20080
rect 394268 -20222 394608 -20136
rect 394268 -20278 394337 -20222
rect 394393 -20278 394479 -20222
rect 394535 -20278 394608 -20222
rect 394268 -20364 394608 -20278
rect 394268 -20420 394337 -20364
rect 394393 -20420 394479 -20364
rect 394535 -20420 394608 -20364
rect 394268 -20506 394608 -20420
rect 394268 -20562 394337 -20506
rect 394393 -20562 394479 -20506
rect 394535 -20562 394608 -20506
rect 394268 -20648 394608 -20562
rect 394268 -20704 394337 -20648
rect 394393 -20704 394479 -20648
rect 394535 -20704 394608 -20648
rect 394268 -20790 394608 -20704
rect 394268 -20846 394337 -20790
rect 394393 -20846 394479 -20790
rect 394535 -20846 394608 -20790
rect 394268 -20932 394608 -20846
rect 394268 -20988 394337 -20932
rect 394393 -20988 394479 -20932
rect 394535 -20988 394608 -20932
rect 394268 -21074 394608 -20988
rect 394268 -21130 394337 -21074
rect 394393 -21130 394479 -21074
rect 394535 -21130 394608 -21074
rect 394268 -21216 394608 -21130
rect 394268 -21272 394337 -21216
rect 394393 -21272 394479 -21216
rect 394535 -21272 394608 -21216
rect 394268 -21358 394608 -21272
rect 394268 -21414 394337 -21358
rect 394393 -21414 394479 -21358
rect 394535 -21414 394608 -21358
rect 394268 -21500 394608 -21414
rect 394268 -21556 394337 -21500
rect 394393 -21556 394479 -21500
rect 394535 -21556 394608 -21500
rect 394268 -21642 394608 -21556
rect 394268 -21698 394337 -21642
rect 394393 -21698 394479 -21642
rect 394535 -21698 394608 -21642
rect 394268 -21784 394608 -21698
rect 394268 -21840 394337 -21784
rect 394393 -21840 394479 -21784
rect 394535 -21840 394608 -21784
rect 394268 -21926 394608 -21840
rect 394268 -21982 394337 -21926
rect 394393 -21982 394479 -21926
rect 394535 -21982 394608 -21926
rect 394268 -22068 394608 -21982
rect 394268 -22124 394337 -22068
rect 394393 -22124 394479 -22068
rect 394535 -22124 394608 -22068
rect 394268 -22210 394608 -22124
rect 394268 -22266 394337 -22210
rect 394393 -22266 394479 -22210
rect 394535 -22266 394608 -22210
rect 394268 -22352 394608 -22266
rect 394268 -22408 394337 -22352
rect 394393 -22408 394479 -22352
rect 394535 -22408 394608 -22352
rect 394268 -22494 394608 -22408
rect 394268 -22550 394337 -22494
rect 394393 -22550 394479 -22494
rect 394535 -22550 394608 -22494
rect 394268 -22636 394608 -22550
rect 394268 -22692 394337 -22636
rect 394393 -22692 394479 -22636
rect 394535 -22692 394608 -22636
rect 394268 -22778 394608 -22692
rect 394268 -22834 394337 -22778
rect 394393 -22834 394479 -22778
rect 394535 -22834 394608 -22778
rect 394268 -22920 394608 -22834
rect 394268 -22976 394337 -22920
rect 394393 -22976 394479 -22920
rect 394535 -22976 394608 -22920
rect 394268 -23062 394608 -22976
rect 394268 -23118 394337 -23062
rect 394393 -23118 394479 -23062
rect 394535 -23118 394608 -23062
rect 394268 -23204 394608 -23118
rect 394268 -23260 394337 -23204
rect 394393 -23260 394479 -23204
rect 394535 -23260 394608 -23204
rect 394268 -23346 394608 -23260
rect 394268 -23402 394337 -23346
rect 394393 -23402 394479 -23346
rect 394535 -23402 394608 -23346
rect 394268 -23488 394608 -23402
rect 394268 -23544 394337 -23488
rect 394393 -23544 394479 -23488
rect 394535 -23544 394608 -23488
rect 394268 -23630 394608 -23544
rect 394268 -23686 394337 -23630
rect 394393 -23686 394479 -23630
rect 394535 -23686 394608 -23630
rect 394268 -23772 394608 -23686
rect 394268 -23828 394337 -23772
rect 394393 -23828 394479 -23772
rect 394535 -23828 394608 -23772
rect 394268 -23914 394608 -23828
rect 394268 -23970 394337 -23914
rect 394393 -23970 394479 -23914
rect 394535 -23970 394608 -23914
rect 394268 -24056 394608 -23970
rect 394268 -24112 394337 -24056
rect 394393 -24112 394479 -24056
rect 394535 -24112 394608 -24056
rect 394268 -24198 394608 -24112
rect 394268 -24254 394337 -24198
rect 394393 -24254 394479 -24198
rect 394535 -24254 394608 -24198
rect 394268 -24340 394608 -24254
rect 394268 -24396 394337 -24340
rect 394393 -24396 394479 -24340
rect 394535 -24396 394608 -24340
rect 394268 -24482 394608 -24396
rect 394268 -24538 394337 -24482
rect 394393 -24538 394479 -24482
rect 394535 -24538 394608 -24482
rect 394268 -24624 394608 -24538
rect 394268 -24680 394337 -24624
rect 394393 -24680 394479 -24624
rect 394535 -24680 394608 -24624
rect 394268 -24766 394608 -24680
rect 394268 -24822 394337 -24766
rect 394393 -24822 394479 -24766
rect 394535 -24822 394608 -24766
rect 394268 -24908 394608 -24822
rect 394268 -24964 394337 -24908
rect 394393 -24964 394479 -24908
rect 394535 -24964 394608 -24908
rect 394268 -25050 394608 -24964
rect 394268 -25106 394337 -25050
rect 394393 -25106 394479 -25050
rect 394535 -25106 394608 -25050
rect 394268 -25192 394608 -25106
rect 394268 -25248 394337 -25192
rect 394393 -25248 394479 -25192
rect 394535 -25248 394608 -25192
rect 394268 -25334 394608 -25248
rect 394268 -25390 394337 -25334
rect 394393 -25390 394479 -25334
rect 394535 -25390 394608 -25334
rect 394268 -25476 394608 -25390
rect 394268 -25532 394337 -25476
rect 394393 -25532 394479 -25476
rect 394535 -25532 394608 -25476
rect 394268 -25542 394608 -25532
rect 394668 -17950 395008 -17820
rect 394668 -18006 394740 -17950
rect 394796 -18006 394882 -17950
rect 394938 -18006 395008 -17950
rect 394668 -18092 395008 -18006
rect 394668 -18148 394740 -18092
rect 394796 -18148 394882 -18092
rect 394938 -18148 395008 -18092
rect 394668 -18234 395008 -18148
rect 394668 -18290 394740 -18234
rect 394796 -18290 394882 -18234
rect 394938 -18290 395008 -18234
rect 394668 -18376 395008 -18290
rect 394668 -18432 394740 -18376
rect 394796 -18432 394882 -18376
rect 394938 -18432 395008 -18376
rect 394668 -18518 395008 -18432
rect 394668 -18574 394740 -18518
rect 394796 -18574 394882 -18518
rect 394938 -18574 395008 -18518
rect 394668 -18660 395008 -18574
rect 394668 -18716 394740 -18660
rect 394796 -18716 394882 -18660
rect 394938 -18716 395008 -18660
rect 394668 -18802 395008 -18716
rect 394668 -18858 394740 -18802
rect 394796 -18858 394882 -18802
rect 394938 -18858 395008 -18802
rect 394668 -18944 395008 -18858
rect 394668 -19000 394740 -18944
rect 394796 -19000 394882 -18944
rect 394938 -19000 395008 -18944
rect 394668 -19086 395008 -19000
rect 394668 -19142 394740 -19086
rect 394796 -19142 394882 -19086
rect 394938 -19142 395008 -19086
rect 394668 -19228 395008 -19142
rect 394668 -19284 394740 -19228
rect 394796 -19284 394882 -19228
rect 394938 -19284 395008 -19228
rect 394668 -19370 395008 -19284
rect 394668 -19426 394740 -19370
rect 394796 -19426 394882 -19370
rect 394938 -19426 395008 -19370
rect 394668 -19512 395008 -19426
rect 394668 -19568 394740 -19512
rect 394796 -19568 394882 -19512
rect 394938 -19568 395008 -19512
rect 394668 -19654 395008 -19568
rect 394668 -19710 394740 -19654
rect 394796 -19710 394882 -19654
rect 394938 -19710 395008 -19654
rect 394668 -19796 395008 -19710
rect 394668 -19852 394740 -19796
rect 394796 -19852 394882 -19796
rect 394938 -19852 395008 -19796
rect 394668 -19938 395008 -19852
rect 394668 -19994 394740 -19938
rect 394796 -19994 394882 -19938
rect 394938 -19994 395008 -19938
rect 394668 -20080 395008 -19994
rect 394668 -20136 394740 -20080
rect 394796 -20136 394882 -20080
rect 394938 -20136 395008 -20080
rect 394668 -20222 395008 -20136
rect 394668 -20278 394740 -20222
rect 394796 -20278 394882 -20222
rect 394938 -20278 395008 -20222
rect 394668 -20364 395008 -20278
rect 394668 -20420 394740 -20364
rect 394796 -20420 394882 -20364
rect 394938 -20420 395008 -20364
rect 394668 -20506 395008 -20420
rect 394668 -20562 394740 -20506
rect 394796 -20562 394882 -20506
rect 394938 -20562 395008 -20506
rect 394668 -20648 395008 -20562
rect 394668 -20704 394740 -20648
rect 394796 -20704 394882 -20648
rect 394938 -20704 395008 -20648
rect 394668 -20790 395008 -20704
rect 394668 -20846 394740 -20790
rect 394796 -20846 394882 -20790
rect 394938 -20846 395008 -20790
rect 394668 -20932 395008 -20846
rect 394668 -20988 394740 -20932
rect 394796 -20988 394882 -20932
rect 394938 -20988 395008 -20932
rect 394668 -21074 395008 -20988
rect 394668 -21130 394740 -21074
rect 394796 -21130 394882 -21074
rect 394938 -21130 395008 -21074
rect 394668 -21216 395008 -21130
rect 394668 -21272 394740 -21216
rect 394796 -21272 394882 -21216
rect 394938 -21272 395008 -21216
rect 394668 -21358 395008 -21272
rect 394668 -21414 394740 -21358
rect 394796 -21414 394882 -21358
rect 394938 -21414 395008 -21358
rect 394668 -21500 395008 -21414
rect 394668 -21556 394740 -21500
rect 394796 -21556 394882 -21500
rect 394938 -21556 395008 -21500
rect 394668 -21642 395008 -21556
rect 394668 -21698 394740 -21642
rect 394796 -21698 394882 -21642
rect 394938 -21698 395008 -21642
rect 394668 -21784 395008 -21698
rect 394668 -21840 394740 -21784
rect 394796 -21840 394882 -21784
rect 394938 -21840 395008 -21784
rect 394668 -21926 395008 -21840
rect 394668 -21982 394740 -21926
rect 394796 -21982 394882 -21926
rect 394938 -21982 395008 -21926
rect 394668 -22068 395008 -21982
rect 394668 -22124 394740 -22068
rect 394796 -22124 394882 -22068
rect 394938 -22124 395008 -22068
rect 394668 -22210 395008 -22124
rect 394668 -22266 394740 -22210
rect 394796 -22266 394882 -22210
rect 394938 -22266 395008 -22210
rect 394668 -22352 395008 -22266
rect 394668 -22408 394740 -22352
rect 394796 -22408 394882 -22352
rect 394938 -22408 395008 -22352
rect 394668 -22494 395008 -22408
rect 394668 -22550 394740 -22494
rect 394796 -22550 394882 -22494
rect 394938 -22550 395008 -22494
rect 394668 -22636 395008 -22550
rect 394668 -22692 394740 -22636
rect 394796 -22692 394882 -22636
rect 394938 -22692 395008 -22636
rect 394668 -22778 395008 -22692
rect 394668 -22834 394740 -22778
rect 394796 -22834 394882 -22778
rect 394938 -22834 395008 -22778
rect 394668 -22920 395008 -22834
rect 394668 -22976 394740 -22920
rect 394796 -22976 394882 -22920
rect 394938 -22976 395008 -22920
rect 394668 -23062 395008 -22976
rect 394668 -23118 394740 -23062
rect 394796 -23118 394882 -23062
rect 394938 -23118 395008 -23062
rect 394668 -23204 395008 -23118
rect 394668 -23260 394740 -23204
rect 394796 -23260 394882 -23204
rect 394938 -23260 395008 -23204
rect 394668 -23346 395008 -23260
rect 394668 -23402 394740 -23346
rect 394796 -23402 394882 -23346
rect 394938 -23402 395008 -23346
rect 394668 -23488 395008 -23402
rect 394668 -23544 394740 -23488
rect 394796 -23544 394882 -23488
rect 394938 -23544 395008 -23488
rect 394668 -23630 395008 -23544
rect 394668 -23686 394740 -23630
rect 394796 -23686 394882 -23630
rect 394938 -23686 395008 -23630
rect 394668 -23772 395008 -23686
rect 394668 -23828 394740 -23772
rect 394796 -23828 394882 -23772
rect 394938 -23828 395008 -23772
rect 394668 -23914 395008 -23828
rect 394668 -23970 394740 -23914
rect 394796 -23970 394882 -23914
rect 394938 -23970 395008 -23914
rect 394668 -24056 395008 -23970
rect 394668 -24112 394740 -24056
rect 394796 -24112 394882 -24056
rect 394938 -24112 395008 -24056
rect 394668 -24198 395008 -24112
rect 394668 -24254 394740 -24198
rect 394796 -24254 394882 -24198
rect 394938 -24254 395008 -24198
rect 394668 -24340 395008 -24254
rect 394668 -24396 394740 -24340
rect 394796 -24396 394882 -24340
rect 394938 -24396 395008 -24340
rect 394668 -24482 395008 -24396
rect 394668 -24538 394740 -24482
rect 394796 -24538 394882 -24482
rect 394938 -24538 395008 -24482
rect 394668 -24624 395008 -24538
rect 394668 -24680 394740 -24624
rect 394796 -24680 394882 -24624
rect 394938 -24680 395008 -24624
rect 394668 -24766 395008 -24680
rect 394668 -24822 394740 -24766
rect 394796 -24822 394882 -24766
rect 394938 -24822 395008 -24766
rect 394668 -24908 395008 -24822
rect 394668 -24964 394740 -24908
rect 394796 -24964 394882 -24908
rect 394938 -24964 395008 -24908
rect 394668 -25050 395008 -24964
rect 394668 -25106 394740 -25050
rect 394796 -25106 394882 -25050
rect 394938 -25106 395008 -25050
rect 394668 -25192 395008 -25106
rect 394668 -25248 394740 -25192
rect 394796 -25248 394882 -25192
rect 394938 -25248 395008 -25192
rect 394668 -25334 395008 -25248
rect 394668 -25390 394740 -25334
rect 394796 -25390 394882 -25334
rect 394938 -25390 395008 -25334
rect 394668 -25476 395008 -25390
rect 394668 -25532 394740 -25476
rect 394796 -25532 394882 -25476
rect 394938 -25532 395008 -25476
rect 394668 -25542 395008 -25532
rect 395068 -17950 395408 -17820
rect 395068 -18006 395142 -17950
rect 395198 -18006 395284 -17950
rect 395340 -18006 395408 -17950
rect 395068 -18092 395408 -18006
rect 395068 -18148 395142 -18092
rect 395198 -18148 395284 -18092
rect 395340 -18148 395408 -18092
rect 395068 -18234 395408 -18148
rect 395068 -18290 395142 -18234
rect 395198 -18290 395284 -18234
rect 395340 -18290 395408 -18234
rect 395068 -18376 395408 -18290
rect 395068 -18432 395142 -18376
rect 395198 -18432 395284 -18376
rect 395340 -18432 395408 -18376
rect 395068 -18518 395408 -18432
rect 395068 -18574 395142 -18518
rect 395198 -18574 395284 -18518
rect 395340 -18574 395408 -18518
rect 395068 -18660 395408 -18574
rect 395068 -18716 395142 -18660
rect 395198 -18716 395284 -18660
rect 395340 -18716 395408 -18660
rect 395068 -18802 395408 -18716
rect 395068 -18858 395142 -18802
rect 395198 -18858 395284 -18802
rect 395340 -18858 395408 -18802
rect 395068 -18944 395408 -18858
rect 395068 -19000 395142 -18944
rect 395198 -19000 395284 -18944
rect 395340 -19000 395408 -18944
rect 395068 -19086 395408 -19000
rect 395068 -19142 395142 -19086
rect 395198 -19142 395284 -19086
rect 395340 -19142 395408 -19086
rect 395068 -19228 395408 -19142
rect 395068 -19284 395142 -19228
rect 395198 -19284 395284 -19228
rect 395340 -19284 395408 -19228
rect 395068 -19370 395408 -19284
rect 395068 -19426 395142 -19370
rect 395198 -19426 395284 -19370
rect 395340 -19426 395408 -19370
rect 395068 -19512 395408 -19426
rect 395068 -19568 395142 -19512
rect 395198 -19568 395284 -19512
rect 395340 -19568 395408 -19512
rect 395068 -19654 395408 -19568
rect 395068 -19710 395142 -19654
rect 395198 -19710 395284 -19654
rect 395340 -19710 395408 -19654
rect 395068 -19796 395408 -19710
rect 395068 -19852 395142 -19796
rect 395198 -19852 395284 -19796
rect 395340 -19852 395408 -19796
rect 395068 -19938 395408 -19852
rect 395068 -19994 395142 -19938
rect 395198 -19994 395284 -19938
rect 395340 -19994 395408 -19938
rect 395068 -20080 395408 -19994
rect 395068 -20136 395142 -20080
rect 395198 -20136 395284 -20080
rect 395340 -20136 395408 -20080
rect 395068 -20222 395408 -20136
rect 395068 -20278 395142 -20222
rect 395198 -20278 395284 -20222
rect 395340 -20278 395408 -20222
rect 395068 -20364 395408 -20278
rect 395068 -20420 395142 -20364
rect 395198 -20420 395284 -20364
rect 395340 -20420 395408 -20364
rect 395068 -20506 395408 -20420
rect 395068 -20562 395142 -20506
rect 395198 -20562 395284 -20506
rect 395340 -20562 395408 -20506
rect 395068 -20648 395408 -20562
rect 395068 -20704 395142 -20648
rect 395198 -20704 395284 -20648
rect 395340 -20704 395408 -20648
rect 395068 -20790 395408 -20704
rect 395068 -20846 395142 -20790
rect 395198 -20846 395284 -20790
rect 395340 -20846 395408 -20790
rect 395068 -20932 395408 -20846
rect 395068 -20988 395142 -20932
rect 395198 -20988 395284 -20932
rect 395340 -20988 395408 -20932
rect 395068 -21074 395408 -20988
rect 395068 -21130 395142 -21074
rect 395198 -21130 395284 -21074
rect 395340 -21130 395408 -21074
rect 395068 -21216 395408 -21130
rect 395068 -21272 395142 -21216
rect 395198 -21272 395284 -21216
rect 395340 -21272 395408 -21216
rect 395068 -21358 395408 -21272
rect 395068 -21414 395142 -21358
rect 395198 -21414 395284 -21358
rect 395340 -21414 395408 -21358
rect 395068 -21500 395408 -21414
rect 395068 -21556 395142 -21500
rect 395198 -21556 395284 -21500
rect 395340 -21556 395408 -21500
rect 395068 -21642 395408 -21556
rect 395068 -21698 395142 -21642
rect 395198 -21698 395284 -21642
rect 395340 -21698 395408 -21642
rect 395068 -21784 395408 -21698
rect 395068 -21840 395142 -21784
rect 395198 -21840 395284 -21784
rect 395340 -21840 395408 -21784
rect 395068 -21926 395408 -21840
rect 395068 -21982 395142 -21926
rect 395198 -21982 395284 -21926
rect 395340 -21982 395408 -21926
rect 395068 -22068 395408 -21982
rect 395068 -22124 395142 -22068
rect 395198 -22124 395284 -22068
rect 395340 -22124 395408 -22068
rect 395068 -22210 395408 -22124
rect 395068 -22266 395142 -22210
rect 395198 -22266 395284 -22210
rect 395340 -22266 395408 -22210
rect 395068 -22352 395408 -22266
rect 395068 -22408 395142 -22352
rect 395198 -22408 395284 -22352
rect 395340 -22408 395408 -22352
rect 395068 -22494 395408 -22408
rect 395068 -22550 395142 -22494
rect 395198 -22550 395284 -22494
rect 395340 -22550 395408 -22494
rect 395068 -22636 395408 -22550
rect 395068 -22692 395142 -22636
rect 395198 -22692 395284 -22636
rect 395340 -22692 395408 -22636
rect 395068 -22778 395408 -22692
rect 395068 -22834 395142 -22778
rect 395198 -22834 395284 -22778
rect 395340 -22834 395408 -22778
rect 395068 -22920 395408 -22834
rect 395068 -22976 395142 -22920
rect 395198 -22976 395284 -22920
rect 395340 -22976 395408 -22920
rect 395068 -23062 395408 -22976
rect 395068 -23118 395142 -23062
rect 395198 -23118 395284 -23062
rect 395340 -23118 395408 -23062
rect 395068 -23204 395408 -23118
rect 395068 -23260 395142 -23204
rect 395198 -23260 395284 -23204
rect 395340 -23260 395408 -23204
rect 395068 -23346 395408 -23260
rect 395068 -23402 395142 -23346
rect 395198 -23402 395284 -23346
rect 395340 -23402 395408 -23346
rect 395068 -23488 395408 -23402
rect 395068 -23544 395142 -23488
rect 395198 -23544 395284 -23488
rect 395340 -23544 395408 -23488
rect 395068 -23630 395408 -23544
rect 395068 -23686 395142 -23630
rect 395198 -23686 395284 -23630
rect 395340 -23686 395408 -23630
rect 395068 -23772 395408 -23686
rect 395068 -23828 395142 -23772
rect 395198 -23828 395284 -23772
rect 395340 -23828 395408 -23772
rect 395068 -23914 395408 -23828
rect 395068 -23970 395142 -23914
rect 395198 -23970 395284 -23914
rect 395340 -23970 395408 -23914
rect 395068 -24056 395408 -23970
rect 395068 -24112 395142 -24056
rect 395198 -24112 395284 -24056
rect 395340 -24112 395408 -24056
rect 395068 -24198 395408 -24112
rect 395068 -24254 395142 -24198
rect 395198 -24254 395284 -24198
rect 395340 -24254 395408 -24198
rect 395068 -24340 395408 -24254
rect 395068 -24396 395142 -24340
rect 395198 -24396 395284 -24340
rect 395340 -24396 395408 -24340
rect 395068 -24482 395408 -24396
rect 395068 -24538 395142 -24482
rect 395198 -24538 395284 -24482
rect 395340 -24538 395408 -24482
rect 395068 -24624 395408 -24538
rect 395068 -24680 395142 -24624
rect 395198 -24680 395284 -24624
rect 395340 -24680 395408 -24624
rect 395068 -24766 395408 -24680
rect 395068 -24822 395142 -24766
rect 395198 -24822 395284 -24766
rect 395340 -24822 395408 -24766
rect 395068 -24908 395408 -24822
rect 395068 -24964 395142 -24908
rect 395198 -24964 395284 -24908
rect 395340 -24964 395408 -24908
rect 395068 -25050 395408 -24964
rect 395068 -25106 395142 -25050
rect 395198 -25106 395284 -25050
rect 395340 -25106 395408 -25050
rect 395068 -25192 395408 -25106
rect 395068 -25248 395142 -25192
rect 395198 -25248 395284 -25192
rect 395340 -25248 395408 -25192
rect 395068 -25334 395408 -25248
rect 395068 -25390 395142 -25334
rect 395198 -25390 395284 -25334
rect 395340 -25390 395408 -25334
rect 395068 -25476 395408 -25390
rect 395068 -25532 395142 -25476
rect 395198 -25532 395284 -25476
rect 395340 -25532 395408 -25476
rect 395068 -25542 395408 -25532
rect 395468 -17950 395808 -17820
rect 395468 -18006 395545 -17950
rect 395601 -18006 395687 -17950
rect 395743 -18006 395808 -17950
rect 395468 -18092 395808 -18006
rect 395468 -18148 395545 -18092
rect 395601 -18148 395687 -18092
rect 395743 -18148 395808 -18092
rect 395468 -18234 395808 -18148
rect 395468 -18290 395545 -18234
rect 395601 -18290 395687 -18234
rect 395743 -18290 395808 -18234
rect 395468 -18376 395808 -18290
rect 395468 -18432 395545 -18376
rect 395601 -18432 395687 -18376
rect 395743 -18432 395808 -18376
rect 395468 -18518 395808 -18432
rect 395468 -18574 395545 -18518
rect 395601 -18574 395687 -18518
rect 395743 -18574 395808 -18518
rect 395468 -18660 395808 -18574
rect 395468 -18716 395545 -18660
rect 395601 -18716 395687 -18660
rect 395743 -18716 395808 -18660
rect 395468 -18802 395808 -18716
rect 395468 -18858 395545 -18802
rect 395601 -18858 395687 -18802
rect 395743 -18858 395808 -18802
rect 395468 -18944 395808 -18858
rect 395468 -19000 395545 -18944
rect 395601 -19000 395687 -18944
rect 395743 -19000 395808 -18944
rect 395468 -19086 395808 -19000
rect 395468 -19142 395545 -19086
rect 395601 -19142 395687 -19086
rect 395743 -19142 395808 -19086
rect 395468 -19228 395808 -19142
rect 395468 -19284 395545 -19228
rect 395601 -19284 395687 -19228
rect 395743 -19284 395808 -19228
rect 395468 -19370 395808 -19284
rect 395468 -19426 395545 -19370
rect 395601 -19426 395687 -19370
rect 395743 -19426 395808 -19370
rect 395468 -19512 395808 -19426
rect 395468 -19568 395545 -19512
rect 395601 -19568 395687 -19512
rect 395743 -19568 395808 -19512
rect 395468 -19654 395808 -19568
rect 395468 -19710 395545 -19654
rect 395601 -19710 395687 -19654
rect 395743 -19710 395808 -19654
rect 395468 -19796 395808 -19710
rect 395468 -19852 395545 -19796
rect 395601 -19852 395687 -19796
rect 395743 -19852 395808 -19796
rect 395468 -19938 395808 -19852
rect 395468 -19994 395545 -19938
rect 395601 -19994 395687 -19938
rect 395743 -19994 395808 -19938
rect 395468 -20080 395808 -19994
rect 395468 -20136 395545 -20080
rect 395601 -20136 395687 -20080
rect 395743 -20136 395808 -20080
rect 395468 -20222 395808 -20136
rect 395468 -20278 395545 -20222
rect 395601 -20278 395687 -20222
rect 395743 -20278 395808 -20222
rect 395468 -20364 395808 -20278
rect 395468 -20420 395545 -20364
rect 395601 -20420 395687 -20364
rect 395743 -20420 395808 -20364
rect 395468 -20506 395808 -20420
rect 395468 -20562 395545 -20506
rect 395601 -20562 395687 -20506
rect 395743 -20562 395808 -20506
rect 395468 -20648 395808 -20562
rect 395468 -20704 395545 -20648
rect 395601 -20704 395687 -20648
rect 395743 -20704 395808 -20648
rect 395468 -20790 395808 -20704
rect 395468 -20846 395545 -20790
rect 395601 -20846 395687 -20790
rect 395743 -20846 395808 -20790
rect 395468 -20932 395808 -20846
rect 395468 -20988 395545 -20932
rect 395601 -20988 395687 -20932
rect 395743 -20988 395808 -20932
rect 395468 -21074 395808 -20988
rect 395468 -21130 395545 -21074
rect 395601 -21130 395687 -21074
rect 395743 -21130 395808 -21074
rect 395468 -21216 395808 -21130
rect 395468 -21272 395545 -21216
rect 395601 -21272 395687 -21216
rect 395743 -21272 395808 -21216
rect 395468 -21358 395808 -21272
rect 395468 -21414 395545 -21358
rect 395601 -21414 395687 -21358
rect 395743 -21414 395808 -21358
rect 395468 -21500 395808 -21414
rect 395468 -21556 395545 -21500
rect 395601 -21556 395687 -21500
rect 395743 -21556 395808 -21500
rect 395468 -21642 395808 -21556
rect 395468 -21698 395545 -21642
rect 395601 -21698 395687 -21642
rect 395743 -21698 395808 -21642
rect 395468 -21784 395808 -21698
rect 395468 -21840 395545 -21784
rect 395601 -21840 395687 -21784
rect 395743 -21840 395808 -21784
rect 395468 -21926 395808 -21840
rect 395468 -21982 395545 -21926
rect 395601 -21982 395687 -21926
rect 395743 -21982 395808 -21926
rect 395468 -22068 395808 -21982
rect 395468 -22124 395545 -22068
rect 395601 -22124 395687 -22068
rect 395743 -22124 395808 -22068
rect 395468 -22210 395808 -22124
rect 395468 -22266 395545 -22210
rect 395601 -22266 395687 -22210
rect 395743 -22266 395808 -22210
rect 395468 -22352 395808 -22266
rect 395468 -22408 395545 -22352
rect 395601 -22408 395687 -22352
rect 395743 -22408 395808 -22352
rect 395468 -22494 395808 -22408
rect 395468 -22550 395545 -22494
rect 395601 -22550 395687 -22494
rect 395743 -22550 395808 -22494
rect 395468 -22636 395808 -22550
rect 395468 -22692 395545 -22636
rect 395601 -22692 395687 -22636
rect 395743 -22692 395808 -22636
rect 395468 -22778 395808 -22692
rect 395468 -22834 395545 -22778
rect 395601 -22834 395687 -22778
rect 395743 -22834 395808 -22778
rect 395468 -22920 395808 -22834
rect 395468 -22976 395545 -22920
rect 395601 -22976 395687 -22920
rect 395743 -22976 395808 -22920
rect 395468 -23062 395808 -22976
rect 395468 -23118 395545 -23062
rect 395601 -23118 395687 -23062
rect 395743 -23118 395808 -23062
rect 395468 -23204 395808 -23118
rect 395468 -23260 395545 -23204
rect 395601 -23260 395687 -23204
rect 395743 -23260 395808 -23204
rect 395468 -23346 395808 -23260
rect 395468 -23402 395545 -23346
rect 395601 -23402 395687 -23346
rect 395743 -23402 395808 -23346
rect 395468 -23488 395808 -23402
rect 395468 -23544 395545 -23488
rect 395601 -23544 395687 -23488
rect 395743 -23544 395808 -23488
rect 395468 -23630 395808 -23544
rect 395468 -23686 395545 -23630
rect 395601 -23686 395687 -23630
rect 395743 -23686 395808 -23630
rect 395468 -23772 395808 -23686
rect 395468 -23828 395545 -23772
rect 395601 -23828 395687 -23772
rect 395743 -23828 395808 -23772
rect 395468 -23914 395808 -23828
rect 395468 -23970 395545 -23914
rect 395601 -23970 395687 -23914
rect 395743 -23970 395808 -23914
rect 395468 -24056 395808 -23970
rect 395468 -24112 395545 -24056
rect 395601 -24112 395687 -24056
rect 395743 -24112 395808 -24056
rect 395468 -24198 395808 -24112
rect 395468 -24254 395545 -24198
rect 395601 -24254 395687 -24198
rect 395743 -24254 395808 -24198
rect 395468 -24340 395808 -24254
rect 395468 -24396 395545 -24340
rect 395601 -24396 395687 -24340
rect 395743 -24396 395808 -24340
rect 395468 -24482 395808 -24396
rect 395468 -24538 395545 -24482
rect 395601 -24538 395687 -24482
rect 395743 -24538 395808 -24482
rect 395468 -24624 395808 -24538
rect 395468 -24680 395545 -24624
rect 395601 -24680 395687 -24624
rect 395743 -24680 395808 -24624
rect 395468 -24766 395808 -24680
rect 395468 -24822 395545 -24766
rect 395601 -24822 395687 -24766
rect 395743 -24822 395808 -24766
rect 395468 -24908 395808 -24822
rect 395468 -24964 395545 -24908
rect 395601 -24964 395687 -24908
rect 395743 -24964 395808 -24908
rect 395468 -25050 395808 -24964
rect 395468 -25106 395545 -25050
rect 395601 -25106 395687 -25050
rect 395743 -25106 395808 -25050
rect 395468 -25192 395808 -25106
rect 395468 -25248 395545 -25192
rect 395601 -25248 395687 -25192
rect 395743 -25248 395808 -25192
rect 395468 -25334 395808 -25248
rect 395468 -25390 395545 -25334
rect 395601 -25390 395687 -25334
rect 395743 -25390 395808 -25334
rect 395468 -25476 395808 -25390
rect 395468 -25532 395545 -25476
rect 395601 -25532 395687 -25476
rect 395743 -25532 395808 -25476
rect 395468 -25542 395808 -25532
rect 395868 -17950 396208 -17820
rect 395868 -18006 395941 -17950
rect 395997 -18006 396083 -17950
rect 396139 -18006 396208 -17950
rect 395868 -18092 396208 -18006
rect 395868 -18148 395941 -18092
rect 395997 -18148 396083 -18092
rect 396139 -18148 396208 -18092
rect 395868 -18234 396208 -18148
rect 395868 -18290 395941 -18234
rect 395997 -18290 396083 -18234
rect 396139 -18290 396208 -18234
rect 395868 -18376 396208 -18290
rect 395868 -18432 395941 -18376
rect 395997 -18432 396083 -18376
rect 396139 -18432 396208 -18376
rect 395868 -18518 396208 -18432
rect 395868 -18574 395941 -18518
rect 395997 -18574 396083 -18518
rect 396139 -18574 396208 -18518
rect 395868 -18660 396208 -18574
rect 395868 -18716 395941 -18660
rect 395997 -18716 396083 -18660
rect 396139 -18716 396208 -18660
rect 395868 -18802 396208 -18716
rect 395868 -18858 395941 -18802
rect 395997 -18858 396083 -18802
rect 396139 -18858 396208 -18802
rect 395868 -18944 396208 -18858
rect 395868 -19000 395941 -18944
rect 395997 -19000 396083 -18944
rect 396139 -19000 396208 -18944
rect 395868 -19086 396208 -19000
rect 395868 -19142 395941 -19086
rect 395997 -19142 396083 -19086
rect 396139 -19142 396208 -19086
rect 395868 -19228 396208 -19142
rect 395868 -19284 395941 -19228
rect 395997 -19284 396083 -19228
rect 396139 -19284 396208 -19228
rect 395868 -19370 396208 -19284
rect 395868 -19426 395941 -19370
rect 395997 -19426 396083 -19370
rect 396139 -19426 396208 -19370
rect 395868 -19512 396208 -19426
rect 395868 -19568 395941 -19512
rect 395997 -19568 396083 -19512
rect 396139 -19568 396208 -19512
rect 395868 -19654 396208 -19568
rect 395868 -19710 395941 -19654
rect 395997 -19710 396083 -19654
rect 396139 -19710 396208 -19654
rect 395868 -19796 396208 -19710
rect 395868 -19852 395941 -19796
rect 395997 -19852 396083 -19796
rect 396139 -19852 396208 -19796
rect 395868 -19938 396208 -19852
rect 395868 -19994 395941 -19938
rect 395997 -19994 396083 -19938
rect 396139 -19994 396208 -19938
rect 395868 -20080 396208 -19994
rect 395868 -20136 395941 -20080
rect 395997 -20136 396083 -20080
rect 396139 -20136 396208 -20080
rect 395868 -20222 396208 -20136
rect 395868 -20278 395941 -20222
rect 395997 -20278 396083 -20222
rect 396139 -20278 396208 -20222
rect 395868 -20364 396208 -20278
rect 395868 -20420 395941 -20364
rect 395997 -20420 396083 -20364
rect 396139 -20420 396208 -20364
rect 395868 -20506 396208 -20420
rect 395868 -20562 395941 -20506
rect 395997 -20562 396083 -20506
rect 396139 -20562 396208 -20506
rect 395868 -20648 396208 -20562
rect 395868 -20704 395941 -20648
rect 395997 -20704 396083 -20648
rect 396139 -20704 396208 -20648
rect 395868 -20790 396208 -20704
rect 395868 -20846 395941 -20790
rect 395997 -20846 396083 -20790
rect 396139 -20846 396208 -20790
rect 395868 -20932 396208 -20846
rect 395868 -20988 395941 -20932
rect 395997 -20988 396083 -20932
rect 396139 -20988 396208 -20932
rect 395868 -21074 396208 -20988
rect 395868 -21130 395941 -21074
rect 395997 -21130 396083 -21074
rect 396139 -21130 396208 -21074
rect 395868 -21216 396208 -21130
rect 395868 -21272 395941 -21216
rect 395997 -21272 396083 -21216
rect 396139 -21272 396208 -21216
rect 395868 -21358 396208 -21272
rect 395868 -21414 395941 -21358
rect 395997 -21414 396083 -21358
rect 396139 -21414 396208 -21358
rect 395868 -21500 396208 -21414
rect 395868 -21556 395941 -21500
rect 395997 -21556 396083 -21500
rect 396139 -21556 396208 -21500
rect 395868 -21642 396208 -21556
rect 395868 -21698 395941 -21642
rect 395997 -21698 396083 -21642
rect 396139 -21698 396208 -21642
rect 395868 -21784 396208 -21698
rect 395868 -21840 395941 -21784
rect 395997 -21840 396083 -21784
rect 396139 -21840 396208 -21784
rect 395868 -21926 396208 -21840
rect 395868 -21982 395941 -21926
rect 395997 -21982 396083 -21926
rect 396139 -21982 396208 -21926
rect 395868 -22068 396208 -21982
rect 395868 -22124 395941 -22068
rect 395997 -22124 396083 -22068
rect 396139 -22124 396208 -22068
rect 395868 -22210 396208 -22124
rect 395868 -22266 395941 -22210
rect 395997 -22266 396083 -22210
rect 396139 -22266 396208 -22210
rect 395868 -22352 396208 -22266
rect 395868 -22408 395941 -22352
rect 395997 -22408 396083 -22352
rect 396139 -22408 396208 -22352
rect 395868 -22494 396208 -22408
rect 395868 -22550 395941 -22494
rect 395997 -22550 396083 -22494
rect 396139 -22550 396208 -22494
rect 395868 -22636 396208 -22550
rect 395868 -22692 395941 -22636
rect 395997 -22692 396083 -22636
rect 396139 -22692 396208 -22636
rect 395868 -22778 396208 -22692
rect 395868 -22834 395941 -22778
rect 395997 -22834 396083 -22778
rect 396139 -22834 396208 -22778
rect 395868 -22920 396208 -22834
rect 395868 -22976 395941 -22920
rect 395997 -22976 396083 -22920
rect 396139 -22976 396208 -22920
rect 395868 -23062 396208 -22976
rect 395868 -23118 395941 -23062
rect 395997 -23118 396083 -23062
rect 396139 -23118 396208 -23062
rect 395868 -23204 396208 -23118
rect 395868 -23260 395941 -23204
rect 395997 -23260 396083 -23204
rect 396139 -23260 396208 -23204
rect 395868 -23346 396208 -23260
rect 395868 -23402 395941 -23346
rect 395997 -23402 396083 -23346
rect 396139 -23402 396208 -23346
rect 395868 -23488 396208 -23402
rect 395868 -23544 395941 -23488
rect 395997 -23544 396083 -23488
rect 396139 -23544 396208 -23488
rect 395868 -23630 396208 -23544
rect 395868 -23686 395941 -23630
rect 395997 -23686 396083 -23630
rect 396139 -23686 396208 -23630
rect 395868 -23772 396208 -23686
rect 395868 -23828 395941 -23772
rect 395997 -23828 396083 -23772
rect 396139 -23828 396208 -23772
rect 395868 -23914 396208 -23828
rect 395868 -23970 395941 -23914
rect 395997 -23970 396083 -23914
rect 396139 -23970 396208 -23914
rect 395868 -24056 396208 -23970
rect 395868 -24112 395941 -24056
rect 395997 -24112 396083 -24056
rect 396139 -24112 396208 -24056
rect 395868 -24198 396208 -24112
rect 395868 -24254 395941 -24198
rect 395997 -24254 396083 -24198
rect 396139 -24254 396208 -24198
rect 395868 -24340 396208 -24254
rect 395868 -24396 395941 -24340
rect 395997 -24396 396083 -24340
rect 396139 -24396 396208 -24340
rect 395868 -24482 396208 -24396
rect 395868 -24538 395941 -24482
rect 395997 -24538 396083 -24482
rect 396139 -24538 396208 -24482
rect 395868 -24624 396208 -24538
rect 395868 -24680 395941 -24624
rect 395997 -24680 396083 -24624
rect 396139 -24680 396208 -24624
rect 395868 -24766 396208 -24680
rect 395868 -24822 395941 -24766
rect 395997 -24822 396083 -24766
rect 396139 -24822 396208 -24766
rect 395868 -24908 396208 -24822
rect 395868 -24964 395941 -24908
rect 395997 -24964 396083 -24908
rect 396139 -24964 396208 -24908
rect 395868 -25050 396208 -24964
rect 395868 -25106 395941 -25050
rect 395997 -25106 396083 -25050
rect 396139 -25106 396208 -25050
rect 395868 -25192 396208 -25106
rect 395868 -25248 395941 -25192
rect 395997 -25248 396083 -25192
rect 396139 -25248 396208 -25192
rect 395868 -25334 396208 -25248
rect 395868 -25390 395941 -25334
rect 395997 -25390 396083 -25334
rect 396139 -25390 396208 -25334
rect 395868 -25476 396208 -25390
rect 395868 -25532 395941 -25476
rect 395997 -25532 396083 -25476
rect 396139 -25532 396208 -25476
rect 395868 -25542 396208 -25532
rect 396400 -17858 397200 -17820
rect 396400 -17914 396526 -17858
rect 396582 -17914 396650 -17858
rect 396706 -17914 396774 -17858
rect 396830 -17914 396898 -17858
rect 396954 -17914 397022 -17858
rect 397078 -17914 397200 -17858
rect 396400 -17982 397200 -17914
rect 396400 -18038 396526 -17982
rect 396582 -18038 396650 -17982
rect 396706 -18038 396774 -17982
rect 396830 -18038 396898 -17982
rect 396954 -18038 397022 -17982
rect 397078 -18038 397200 -17982
rect 396400 -18106 397200 -18038
rect 396400 -18162 396526 -18106
rect 396582 -18162 396650 -18106
rect 396706 -18162 396774 -18106
rect 396830 -18162 396898 -18106
rect 396954 -18162 397022 -18106
rect 397078 -18162 397200 -18106
rect 396400 -18230 397200 -18162
rect 396400 -18286 396526 -18230
rect 396582 -18286 396650 -18230
rect 396706 -18286 396774 -18230
rect 396830 -18286 396898 -18230
rect 396954 -18286 397022 -18230
rect 397078 -18286 397200 -18230
rect 396400 -18354 397200 -18286
rect 396400 -18410 396526 -18354
rect 396582 -18410 396650 -18354
rect 396706 -18410 396774 -18354
rect 396830 -18410 396898 -18354
rect 396954 -18410 397022 -18354
rect 397078 -18410 397200 -18354
rect 396400 -18478 397200 -18410
rect 396400 -18534 396526 -18478
rect 396582 -18534 396650 -18478
rect 396706 -18534 396774 -18478
rect 396830 -18534 396898 -18478
rect 396954 -18534 397022 -18478
rect 397078 -18534 397200 -18478
rect 396400 -18602 397200 -18534
rect 396400 -18658 396526 -18602
rect 396582 -18658 396650 -18602
rect 396706 -18658 396774 -18602
rect 396830 -18658 396898 -18602
rect 396954 -18658 397022 -18602
rect 397078 -18658 397200 -18602
rect 396400 -18726 397200 -18658
rect 396400 -18782 396526 -18726
rect 396582 -18782 396650 -18726
rect 396706 -18782 396774 -18726
rect 396830 -18782 396898 -18726
rect 396954 -18782 397022 -18726
rect 397078 -18782 397200 -18726
rect 396400 -18850 397200 -18782
rect 396400 -18906 396526 -18850
rect 396582 -18906 396650 -18850
rect 396706 -18906 396774 -18850
rect 396830 -18906 396898 -18850
rect 396954 -18906 397022 -18850
rect 397078 -18906 397200 -18850
rect 396400 -18974 397200 -18906
rect 396400 -19030 396526 -18974
rect 396582 -19030 396650 -18974
rect 396706 -19030 396774 -18974
rect 396830 -19030 396898 -18974
rect 396954 -19030 397022 -18974
rect 397078 -19030 397200 -18974
rect 396400 -19098 397200 -19030
rect 396400 -19154 396526 -19098
rect 396582 -19154 396650 -19098
rect 396706 -19154 396774 -19098
rect 396830 -19154 396898 -19098
rect 396954 -19154 397022 -19098
rect 397078 -19154 397200 -19098
rect 396400 -19222 397200 -19154
rect 396400 -19278 396526 -19222
rect 396582 -19278 396650 -19222
rect 396706 -19278 396774 -19222
rect 396830 -19278 396898 -19222
rect 396954 -19278 397022 -19222
rect 397078 -19278 397200 -19222
rect 396400 -19346 397200 -19278
rect 396400 -19402 396526 -19346
rect 396582 -19402 396650 -19346
rect 396706 -19402 396774 -19346
rect 396830 -19402 396898 -19346
rect 396954 -19402 397022 -19346
rect 397078 -19402 397200 -19346
rect 396400 -19470 397200 -19402
rect 396400 -19526 396526 -19470
rect 396582 -19526 396650 -19470
rect 396706 -19526 396774 -19470
rect 396830 -19526 396898 -19470
rect 396954 -19526 397022 -19470
rect 397078 -19526 397200 -19470
rect 396400 -19594 397200 -19526
rect 396400 -19650 396526 -19594
rect 396582 -19650 396650 -19594
rect 396706 -19650 396774 -19594
rect 396830 -19650 396898 -19594
rect 396954 -19650 397022 -19594
rect 397078 -19650 397200 -19594
rect 396400 -19718 397200 -19650
rect 396400 -19774 396526 -19718
rect 396582 -19774 396650 -19718
rect 396706 -19774 396774 -19718
rect 396830 -19774 396898 -19718
rect 396954 -19774 397022 -19718
rect 397078 -19774 397200 -19718
rect 396400 -19842 397200 -19774
rect 396400 -19898 396526 -19842
rect 396582 -19898 396650 -19842
rect 396706 -19898 396774 -19842
rect 396830 -19898 396898 -19842
rect 396954 -19898 397022 -19842
rect 397078 -19898 397200 -19842
rect 396400 -19966 397200 -19898
rect 396400 -20022 396526 -19966
rect 396582 -20022 396650 -19966
rect 396706 -20022 396774 -19966
rect 396830 -20022 396898 -19966
rect 396954 -20022 397022 -19966
rect 397078 -20022 397200 -19966
rect 396400 -20090 397200 -20022
rect 396400 -20146 396526 -20090
rect 396582 -20146 396650 -20090
rect 396706 -20146 396774 -20090
rect 396830 -20146 396898 -20090
rect 396954 -20146 397022 -20090
rect 397078 -20146 397200 -20090
rect 396400 -20214 397200 -20146
rect 396400 -20270 396526 -20214
rect 396582 -20270 396650 -20214
rect 396706 -20270 396774 -20214
rect 396830 -20270 396898 -20214
rect 396954 -20270 397022 -20214
rect 397078 -20270 397200 -20214
rect 396400 -20338 397200 -20270
rect 396400 -20394 396526 -20338
rect 396582 -20394 396650 -20338
rect 396706 -20394 396774 -20338
rect 396830 -20394 396898 -20338
rect 396954 -20394 397022 -20338
rect 397078 -20394 397200 -20338
rect 396400 -20462 397200 -20394
rect 396400 -20518 396526 -20462
rect 396582 -20518 396650 -20462
rect 396706 -20518 396774 -20462
rect 396830 -20518 396898 -20462
rect 396954 -20518 397022 -20462
rect 397078 -20518 397200 -20462
rect 396400 -20586 397200 -20518
rect 396400 -20642 396526 -20586
rect 396582 -20642 396650 -20586
rect 396706 -20642 396774 -20586
rect 396830 -20642 396898 -20586
rect 396954 -20642 397022 -20586
rect 397078 -20642 397200 -20586
rect 396400 -20710 397200 -20642
rect 396400 -20766 396526 -20710
rect 396582 -20766 396650 -20710
rect 396706 -20766 396774 -20710
rect 396830 -20766 396898 -20710
rect 396954 -20766 397022 -20710
rect 397078 -20766 397200 -20710
rect 396400 -20834 397200 -20766
rect 396400 -20890 396526 -20834
rect 396582 -20890 396650 -20834
rect 396706 -20890 396774 -20834
rect 396830 -20890 396898 -20834
rect 396954 -20890 397022 -20834
rect 397078 -20890 397200 -20834
rect 396400 -20958 397200 -20890
rect 396400 -21014 396526 -20958
rect 396582 -21014 396650 -20958
rect 396706 -21014 396774 -20958
rect 396830 -21014 396898 -20958
rect 396954 -21014 397022 -20958
rect 397078 -21014 397200 -20958
rect 396400 -21082 397200 -21014
rect 396400 -21138 396526 -21082
rect 396582 -21138 396650 -21082
rect 396706 -21138 396774 -21082
rect 396830 -21138 396898 -21082
rect 396954 -21138 397022 -21082
rect 397078 -21138 397200 -21082
rect 396400 -21206 397200 -21138
rect 396400 -21262 396526 -21206
rect 396582 -21262 396650 -21206
rect 396706 -21262 396774 -21206
rect 396830 -21262 396898 -21206
rect 396954 -21262 397022 -21206
rect 397078 -21262 397200 -21206
rect 396400 -21330 397200 -21262
rect 396400 -21386 396526 -21330
rect 396582 -21386 396650 -21330
rect 396706 -21386 396774 -21330
rect 396830 -21386 396898 -21330
rect 396954 -21386 397022 -21330
rect 397078 -21386 397200 -21330
rect 396400 -21454 397200 -21386
rect 396400 -21510 396526 -21454
rect 396582 -21510 396650 -21454
rect 396706 -21510 396774 -21454
rect 396830 -21510 396898 -21454
rect 396954 -21510 397022 -21454
rect 397078 -21510 397200 -21454
rect 396400 -21578 397200 -21510
rect 396400 -21634 396526 -21578
rect 396582 -21634 396650 -21578
rect 396706 -21634 396774 -21578
rect 396830 -21634 396898 -21578
rect 396954 -21634 397022 -21578
rect 397078 -21634 397200 -21578
rect 396400 -21702 397200 -21634
rect 396400 -21758 396526 -21702
rect 396582 -21758 396650 -21702
rect 396706 -21758 396774 -21702
rect 396830 -21758 396898 -21702
rect 396954 -21758 397022 -21702
rect 397078 -21758 397200 -21702
rect 396400 -21826 397200 -21758
rect 396400 -21882 396526 -21826
rect 396582 -21882 396650 -21826
rect 396706 -21882 396774 -21826
rect 396830 -21882 396898 -21826
rect 396954 -21882 397022 -21826
rect 397078 -21882 397200 -21826
rect 396400 -21950 397200 -21882
rect 396400 -22006 396526 -21950
rect 396582 -22006 396650 -21950
rect 396706 -22006 396774 -21950
rect 396830 -22006 396898 -21950
rect 396954 -22006 397022 -21950
rect 397078 -22006 397200 -21950
rect 396400 -22074 397200 -22006
rect 396400 -22130 396526 -22074
rect 396582 -22130 396650 -22074
rect 396706 -22130 396774 -22074
rect 396830 -22130 396898 -22074
rect 396954 -22130 397022 -22074
rect 397078 -22130 397200 -22074
rect 396400 -22198 397200 -22130
rect 396400 -22254 396526 -22198
rect 396582 -22254 396650 -22198
rect 396706 -22254 396774 -22198
rect 396830 -22254 396898 -22198
rect 396954 -22254 397022 -22198
rect 397078 -22254 397200 -22198
rect 396400 -22322 397200 -22254
rect 396400 -22378 396526 -22322
rect 396582 -22378 396650 -22322
rect 396706 -22378 396774 -22322
rect 396830 -22378 396898 -22322
rect 396954 -22378 397022 -22322
rect 397078 -22378 397200 -22322
rect 396400 -22446 397200 -22378
rect 396400 -22502 396526 -22446
rect 396582 -22502 396650 -22446
rect 396706 -22502 396774 -22446
rect 396830 -22502 396898 -22446
rect 396954 -22502 397022 -22446
rect 397078 -22502 397200 -22446
rect 396400 -22570 397200 -22502
rect 396400 -22626 396526 -22570
rect 396582 -22626 396650 -22570
rect 396706 -22626 396774 -22570
rect 396830 -22626 396898 -22570
rect 396954 -22626 397022 -22570
rect 397078 -22626 397200 -22570
rect 396400 -22694 397200 -22626
rect 396400 -22750 396526 -22694
rect 396582 -22750 396650 -22694
rect 396706 -22750 396774 -22694
rect 396830 -22750 396898 -22694
rect 396954 -22750 397022 -22694
rect 397078 -22750 397200 -22694
rect 396400 -22818 397200 -22750
rect 396400 -22874 396526 -22818
rect 396582 -22874 396650 -22818
rect 396706 -22874 396774 -22818
rect 396830 -22874 396898 -22818
rect 396954 -22874 397022 -22818
rect 397078 -22874 397200 -22818
rect 396400 -22942 397200 -22874
rect 396400 -22998 396526 -22942
rect 396582 -22998 396650 -22942
rect 396706 -22998 396774 -22942
rect 396830 -22998 396898 -22942
rect 396954 -22998 397022 -22942
rect 397078 -22998 397200 -22942
rect 396400 -23066 397200 -22998
rect 396400 -23122 396526 -23066
rect 396582 -23122 396650 -23066
rect 396706 -23122 396774 -23066
rect 396830 -23122 396898 -23066
rect 396954 -23122 397022 -23066
rect 397078 -23122 397200 -23066
rect 396400 -23190 397200 -23122
rect 396400 -23246 396526 -23190
rect 396582 -23246 396650 -23190
rect 396706 -23246 396774 -23190
rect 396830 -23246 396898 -23190
rect 396954 -23246 397022 -23190
rect 397078 -23246 397200 -23190
rect 396400 -23314 397200 -23246
rect 396400 -23370 396526 -23314
rect 396582 -23370 396650 -23314
rect 396706 -23370 396774 -23314
rect 396830 -23370 396898 -23314
rect 396954 -23370 397022 -23314
rect 397078 -23370 397200 -23314
rect 396400 -23438 397200 -23370
rect 396400 -23494 396526 -23438
rect 396582 -23494 396650 -23438
rect 396706 -23494 396774 -23438
rect 396830 -23494 396898 -23438
rect 396954 -23494 397022 -23438
rect 397078 -23494 397200 -23438
rect 396400 -23562 397200 -23494
rect 396400 -23618 396526 -23562
rect 396582 -23618 396650 -23562
rect 396706 -23618 396774 -23562
rect 396830 -23618 396898 -23562
rect 396954 -23618 397022 -23562
rect 397078 -23618 397200 -23562
rect 396400 -23686 397200 -23618
rect 396400 -23742 396526 -23686
rect 396582 -23742 396650 -23686
rect 396706 -23742 396774 -23686
rect 396830 -23742 396898 -23686
rect 396954 -23742 397022 -23686
rect 397078 -23742 397200 -23686
rect 396400 -23810 397200 -23742
rect 396400 -23866 396526 -23810
rect 396582 -23866 396650 -23810
rect 396706 -23866 396774 -23810
rect 396830 -23866 396898 -23810
rect 396954 -23866 397022 -23810
rect 397078 -23866 397200 -23810
rect 396400 -23934 397200 -23866
rect 396400 -23990 396526 -23934
rect 396582 -23990 396650 -23934
rect 396706 -23990 396774 -23934
rect 396830 -23990 396898 -23934
rect 396954 -23990 397022 -23934
rect 397078 -23990 397200 -23934
rect 396400 -24058 397200 -23990
rect 396400 -24114 396526 -24058
rect 396582 -24114 396650 -24058
rect 396706 -24114 396774 -24058
rect 396830 -24114 396898 -24058
rect 396954 -24114 397022 -24058
rect 397078 -24114 397200 -24058
rect 396400 -24182 397200 -24114
rect 396400 -24238 396526 -24182
rect 396582 -24238 396650 -24182
rect 396706 -24238 396774 -24182
rect 396830 -24238 396898 -24182
rect 396954 -24238 397022 -24182
rect 397078 -24238 397200 -24182
rect 396400 -24306 397200 -24238
rect 396400 -24362 396526 -24306
rect 396582 -24362 396650 -24306
rect 396706 -24362 396774 -24306
rect 396830 -24362 396898 -24306
rect 396954 -24362 397022 -24306
rect 397078 -24362 397200 -24306
rect 396400 -24430 397200 -24362
rect 396400 -24486 396526 -24430
rect 396582 -24486 396650 -24430
rect 396706 -24486 396774 -24430
rect 396830 -24486 396898 -24430
rect 396954 -24486 397022 -24430
rect 397078 -24486 397200 -24430
rect 396400 -24554 397200 -24486
rect 396400 -24610 396526 -24554
rect 396582 -24610 396650 -24554
rect 396706 -24610 396774 -24554
rect 396830 -24610 396898 -24554
rect 396954 -24610 397022 -24554
rect 397078 -24610 397200 -24554
rect 396400 -24678 397200 -24610
rect 396400 -24734 396526 -24678
rect 396582 -24734 396650 -24678
rect 396706 -24734 396774 -24678
rect 396830 -24734 396898 -24678
rect 396954 -24734 397022 -24678
rect 397078 -24734 397200 -24678
rect 396400 -24802 397200 -24734
rect 396400 -24858 396526 -24802
rect 396582 -24858 396650 -24802
rect 396706 -24858 396774 -24802
rect 396830 -24858 396898 -24802
rect 396954 -24858 397022 -24802
rect 397078 -24858 397200 -24802
rect 396400 -24926 397200 -24858
rect 396400 -24982 396526 -24926
rect 396582 -24982 396650 -24926
rect 396706 -24982 396774 -24926
rect 396830 -24982 396898 -24926
rect 396954 -24982 397022 -24926
rect 397078 -24982 397200 -24926
rect 396400 -25050 397200 -24982
rect 396400 -25106 396526 -25050
rect 396582 -25106 396650 -25050
rect 396706 -25106 396774 -25050
rect 396830 -25106 396898 -25050
rect 396954 -25106 397022 -25050
rect 397078 -25106 397200 -25050
rect 396400 -25174 397200 -25106
rect 396400 -25230 396526 -25174
rect 396582 -25230 396650 -25174
rect 396706 -25230 396774 -25174
rect 396830 -25230 396898 -25174
rect 396954 -25230 397022 -25174
rect 397078 -25230 397200 -25174
rect 396400 -25298 397200 -25230
rect 396400 -25354 396526 -25298
rect 396582 -25354 396650 -25298
rect 396706 -25354 396774 -25298
rect 396830 -25354 396898 -25298
rect 396954 -25354 397022 -25298
rect 397078 -25354 397200 -25298
rect 396400 -25422 397200 -25354
rect 396400 -25478 396526 -25422
rect 396582 -25478 396650 -25422
rect 396706 -25478 396774 -25422
rect 396830 -25478 396898 -25422
rect 396954 -25478 397022 -25422
rect 397078 -25478 397200 -25422
rect 396400 -25542 397200 -25478
rect 388000 -25721 397200 -25542
rect 388000 -25777 388146 -25721
rect 388202 -25777 388270 -25721
rect 388326 -25777 388394 -25721
rect 388450 -25777 388518 -25721
rect 388574 -25777 388642 -25721
rect 388698 -25777 388766 -25721
rect 388822 -25777 388890 -25721
rect 388946 -25777 389014 -25721
rect 389070 -25777 389138 -25721
rect 389194 -25777 389262 -25721
rect 389318 -25777 389386 -25721
rect 389442 -25777 389510 -25721
rect 389566 -25777 389634 -25721
rect 389690 -25777 389758 -25721
rect 389814 -25777 389882 -25721
rect 389938 -25777 390006 -25721
rect 390062 -25777 390130 -25721
rect 390186 -25777 390254 -25721
rect 390310 -25777 390378 -25721
rect 390434 -25777 390502 -25721
rect 390558 -25777 390626 -25721
rect 390682 -25777 390750 -25721
rect 390806 -25777 390874 -25721
rect 390930 -25777 390998 -25721
rect 391054 -25777 391122 -25721
rect 391178 -25777 391246 -25721
rect 391302 -25777 391370 -25721
rect 391426 -25777 391494 -25721
rect 391550 -25777 391618 -25721
rect 391674 -25777 391742 -25721
rect 391798 -25777 391866 -25721
rect 391922 -25777 391990 -25721
rect 392046 -25777 392114 -25721
rect 392170 -25777 392238 -25721
rect 392294 -25777 392362 -25721
rect 392418 -25777 392486 -25721
rect 392542 -25777 392610 -25721
rect 392666 -25777 392734 -25721
rect 392790 -25777 392858 -25721
rect 392914 -25777 392982 -25721
rect 393038 -25777 393106 -25721
rect 393162 -25777 393230 -25721
rect 393286 -25777 393354 -25721
rect 393410 -25777 393478 -25721
rect 393534 -25777 393602 -25721
rect 393658 -25777 393726 -25721
rect 393782 -25777 393850 -25721
rect 393906 -25777 393974 -25721
rect 394030 -25777 394098 -25721
rect 394154 -25777 394222 -25721
rect 394278 -25777 394346 -25721
rect 394402 -25777 394470 -25721
rect 394526 -25777 394594 -25721
rect 394650 -25777 394718 -25721
rect 394774 -25777 394842 -25721
rect 394898 -25777 394966 -25721
rect 395022 -25777 395090 -25721
rect 395146 -25777 395214 -25721
rect 395270 -25777 395338 -25721
rect 395394 -25777 395462 -25721
rect 395518 -25777 395586 -25721
rect 395642 -25777 395710 -25721
rect 395766 -25777 395898 -25721
rect 395954 -25777 396022 -25721
rect 396078 -25777 396146 -25721
rect 396202 -25777 396270 -25721
rect 396326 -25777 396394 -25721
rect 396450 -25777 396518 -25721
rect 396574 -25777 396642 -25721
rect 396698 -25777 396766 -25721
rect 396822 -25777 396890 -25721
rect 396946 -25777 397014 -25721
rect 397070 -25777 397200 -25721
rect 388000 -25845 397200 -25777
rect 388000 -25901 388146 -25845
rect 388202 -25901 388270 -25845
rect 388326 -25901 388394 -25845
rect 388450 -25901 388518 -25845
rect 388574 -25901 388642 -25845
rect 388698 -25901 388766 -25845
rect 388822 -25901 388890 -25845
rect 388946 -25901 389014 -25845
rect 389070 -25901 389138 -25845
rect 389194 -25901 389262 -25845
rect 389318 -25901 389386 -25845
rect 389442 -25901 389510 -25845
rect 389566 -25901 389634 -25845
rect 389690 -25901 389758 -25845
rect 389814 -25901 389882 -25845
rect 389938 -25901 390006 -25845
rect 390062 -25901 390130 -25845
rect 390186 -25901 390254 -25845
rect 390310 -25901 390378 -25845
rect 390434 -25901 390502 -25845
rect 390558 -25901 390626 -25845
rect 390682 -25901 390750 -25845
rect 390806 -25901 390874 -25845
rect 390930 -25901 390998 -25845
rect 391054 -25901 391122 -25845
rect 391178 -25901 391246 -25845
rect 391302 -25901 391370 -25845
rect 391426 -25901 391494 -25845
rect 391550 -25901 391618 -25845
rect 391674 -25901 391742 -25845
rect 391798 -25901 391866 -25845
rect 391922 -25901 391990 -25845
rect 392046 -25901 392114 -25845
rect 392170 -25901 392238 -25845
rect 392294 -25901 392362 -25845
rect 392418 -25901 392486 -25845
rect 392542 -25901 392610 -25845
rect 392666 -25901 392734 -25845
rect 392790 -25901 392858 -25845
rect 392914 -25901 392982 -25845
rect 393038 -25901 393106 -25845
rect 393162 -25901 393230 -25845
rect 393286 -25901 393354 -25845
rect 393410 -25901 393478 -25845
rect 393534 -25901 393602 -25845
rect 393658 -25901 393726 -25845
rect 393782 -25901 393850 -25845
rect 393906 -25901 393974 -25845
rect 394030 -25901 394098 -25845
rect 394154 -25901 394222 -25845
rect 394278 -25901 394346 -25845
rect 394402 -25901 394470 -25845
rect 394526 -25901 394594 -25845
rect 394650 -25901 394718 -25845
rect 394774 -25901 394842 -25845
rect 394898 -25901 394966 -25845
rect 395022 -25901 395090 -25845
rect 395146 -25901 395214 -25845
rect 395270 -25901 395338 -25845
rect 395394 -25901 395462 -25845
rect 395518 -25901 395586 -25845
rect 395642 -25901 395710 -25845
rect 395766 -25901 395898 -25845
rect 395954 -25901 396022 -25845
rect 396078 -25901 396146 -25845
rect 396202 -25901 396270 -25845
rect 396326 -25901 396394 -25845
rect 396450 -25901 396518 -25845
rect 396574 -25901 396642 -25845
rect 396698 -25901 396766 -25845
rect 396822 -25901 396890 -25845
rect 396946 -25901 397014 -25845
rect 397070 -25901 397200 -25845
rect 388000 -25969 397200 -25901
rect 388000 -26025 388146 -25969
rect 388202 -26025 388270 -25969
rect 388326 -26025 388394 -25969
rect 388450 -26025 388518 -25969
rect 388574 -26025 388642 -25969
rect 388698 -26025 388766 -25969
rect 388822 -26025 388890 -25969
rect 388946 -26025 389014 -25969
rect 389070 -26025 389138 -25969
rect 389194 -26025 389262 -25969
rect 389318 -26025 389386 -25969
rect 389442 -26025 389510 -25969
rect 389566 -26025 389634 -25969
rect 389690 -26025 389758 -25969
rect 389814 -26025 389882 -25969
rect 389938 -26025 390006 -25969
rect 390062 -26025 390130 -25969
rect 390186 -26025 390254 -25969
rect 390310 -26025 390378 -25969
rect 390434 -26025 390502 -25969
rect 390558 -26025 390626 -25969
rect 390682 -26025 390750 -25969
rect 390806 -26025 390874 -25969
rect 390930 -26025 390998 -25969
rect 391054 -26025 391122 -25969
rect 391178 -26025 391246 -25969
rect 391302 -26025 391370 -25969
rect 391426 -26025 391494 -25969
rect 391550 -26025 391618 -25969
rect 391674 -26025 391742 -25969
rect 391798 -26025 391866 -25969
rect 391922 -26025 391990 -25969
rect 392046 -26025 392114 -25969
rect 392170 -26025 392238 -25969
rect 392294 -26025 392362 -25969
rect 392418 -26025 392486 -25969
rect 392542 -26025 392610 -25969
rect 392666 -26025 392734 -25969
rect 392790 -26025 392858 -25969
rect 392914 -26025 392982 -25969
rect 393038 -26025 393106 -25969
rect 393162 -26025 393230 -25969
rect 393286 -26025 393354 -25969
rect 393410 -26025 393478 -25969
rect 393534 -26025 393602 -25969
rect 393658 -26025 393726 -25969
rect 393782 -26025 393850 -25969
rect 393906 -26025 393974 -25969
rect 394030 -26025 394098 -25969
rect 394154 -26025 394222 -25969
rect 394278 -26025 394346 -25969
rect 394402 -26025 394470 -25969
rect 394526 -26025 394594 -25969
rect 394650 -26025 394718 -25969
rect 394774 -26025 394842 -25969
rect 394898 -26025 394966 -25969
rect 395022 -26025 395090 -25969
rect 395146 -26025 395214 -25969
rect 395270 -26025 395338 -25969
rect 395394 -26025 395462 -25969
rect 395518 -26025 395586 -25969
rect 395642 -26025 395710 -25969
rect 395766 -26025 395898 -25969
rect 395954 -26025 396022 -25969
rect 396078 -26025 396146 -25969
rect 396202 -26025 396270 -25969
rect 396326 -26025 396394 -25969
rect 396450 -26025 396518 -25969
rect 396574 -26025 396642 -25969
rect 396698 -26025 396766 -25969
rect 396822 -26025 396890 -25969
rect 396946 -26025 397014 -25969
rect 397070 -26025 397200 -25969
rect 388000 -26093 397200 -26025
rect 388000 -26149 388146 -26093
rect 388202 -26149 388270 -26093
rect 388326 -26149 388394 -26093
rect 388450 -26149 388518 -26093
rect 388574 -26149 388642 -26093
rect 388698 -26149 388766 -26093
rect 388822 -26149 388890 -26093
rect 388946 -26149 389014 -26093
rect 389070 -26149 389138 -26093
rect 389194 -26149 389262 -26093
rect 389318 -26149 389386 -26093
rect 389442 -26149 389510 -26093
rect 389566 -26149 389634 -26093
rect 389690 -26149 389758 -26093
rect 389814 -26149 389882 -26093
rect 389938 -26149 390006 -26093
rect 390062 -26149 390130 -26093
rect 390186 -26149 390254 -26093
rect 390310 -26149 390378 -26093
rect 390434 -26149 390502 -26093
rect 390558 -26149 390626 -26093
rect 390682 -26149 390750 -26093
rect 390806 -26149 390874 -26093
rect 390930 -26149 390998 -26093
rect 391054 -26149 391122 -26093
rect 391178 -26149 391246 -26093
rect 391302 -26149 391370 -26093
rect 391426 -26149 391494 -26093
rect 391550 -26149 391618 -26093
rect 391674 -26149 391742 -26093
rect 391798 -26149 391866 -26093
rect 391922 -26149 391990 -26093
rect 392046 -26149 392114 -26093
rect 392170 -26149 392238 -26093
rect 392294 -26149 392362 -26093
rect 392418 -26149 392486 -26093
rect 392542 -26149 392610 -26093
rect 392666 -26149 392734 -26093
rect 392790 -26149 392858 -26093
rect 392914 -26149 392982 -26093
rect 393038 -26149 393106 -26093
rect 393162 -26149 393230 -26093
rect 393286 -26149 393354 -26093
rect 393410 -26149 393478 -26093
rect 393534 -26149 393602 -26093
rect 393658 -26149 393726 -26093
rect 393782 -26149 393850 -26093
rect 393906 -26149 393974 -26093
rect 394030 -26149 394098 -26093
rect 394154 -26149 394222 -26093
rect 394278 -26149 394346 -26093
rect 394402 -26149 394470 -26093
rect 394526 -26149 394594 -26093
rect 394650 -26149 394718 -26093
rect 394774 -26149 394842 -26093
rect 394898 -26149 394966 -26093
rect 395022 -26149 395090 -26093
rect 395146 -26149 395214 -26093
rect 395270 -26149 395338 -26093
rect 395394 -26149 395462 -26093
rect 395518 -26149 395586 -26093
rect 395642 -26149 395710 -26093
rect 395766 -26149 395898 -26093
rect 395954 -26149 396022 -26093
rect 396078 -26149 396146 -26093
rect 396202 -26149 396270 -26093
rect 396326 -26149 396394 -26093
rect 396450 -26149 396518 -26093
rect 396574 -26149 396642 -26093
rect 396698 -26149 396766 -26093
rect 396822 -26149 396890 -26093
rect 396946 -26149 397014 -26093
rect 397070 -26149 397200 -26093
rect 388000 -26270 397200 -26149
<< via4 >>
rect 388146 -17247 388202 -17191
rect 388270 -17247 388326 -17191
rect 388394 -17247 388450 -17191
rect 388518 -17247 388574 -17191
rect 388642 -17247 388698 -17191
rect 388766 -17247 388822 -17191
rect 388890 -17247 388946 -17191
rect 389014 -17247 389070 -17191
rect 389138 -17247 389194 -17191
rect 389262 -17247 389318 -17191
rect 389386 -17247 389442 -17191
rect 389510 -17247 389566 -17191
rect 389634 -17247 389690 -17191
rect 389758 -17247 389814 -17191
rect 389882 -17247 389938 -17191
rect 390006 -17247 390062 -17191
rect 390130 -17247 390186 -17191
rect 390254 -17247 390310 -17191
rect 390378 -17247 390434 -17191
rect 390502 -17247 390558 -17191
rect 390626 -17247 390682 -17191
rect 390750 -17247 390806 -17191
rect 390874 -17247 390930 -17191
rect 390998 -17247 391054 -17191
rect 391122 -17247 391178 -17191
rect 391246 -17247 391302 -17191
rect 391370 -17247 391426 -17191
rect 391494 -17247 391550 -17191
rect 391618 -17247 391674 -17191
rect 391742 -17247 391798 -17191
rect 391866 -17247 391922 -17191
rect 391990 -17247 392046 -17191
rect 392114 -17247 392170 -17191
rect 392238 -17247 392294 -17191
rect 392362 -17247 392418 -17191
rect 392486 -17247 392542 -17191
rect 392610 -17247 392666 -17191
rect 392734 -17247 392790 -17191
rect 392858 -17247 392914 -17191
rect 392982 -17247 393038 -17191
rect 393106 -17247 393162 -17191
rect 393230 -17247 393286 -17191
rect 393354 -17247 393410 -17191
rect 393478 -17247 393534 -17191
rect 393602 -17247 393658 -17191
rect 393726 -17247 393782 -17191
rect 393850 -17247 393906 -17191
rect 393974 -17247 394030 -17191
rect 394098 -17247 394154 -17191
rect 394222 -17247 394278 -17191
rect 394346 -17247 394402 -17191
rect 394470 -17247 394526 -17191
rect 394594 -17247 394650 -17191
rect 394718 -17247 394774 -17191
rect 394842 -17247 394898 -17191
rect 394966 -17247 395022 -17191
rect 395090 -17247 395146 -17191
rect 395214 -17247 395270 -17191
rect 395338 -17247 395394 -17191
rect 395462 -17247 395518 -17191
rect 395586 -17247 395642 -17191
rect 395710 -17247 395766 -17191
rect 395898 -17247 395954 -17191
rect 396022 -17247 396078 -17191
rect 396146 -17247 396202 -17191
rect 396270 -17247 396326 -17191
rect 396394 -17247 396450 -17191
rect 396518 -17247 396574 -17191
rect 396642 -17247 396698 -17191
rect 396766 -17247 396822 -17191
rect 396890 -17247 396946 -17191
rect 397014 -17247 397070 -17191
rect 388146 -17371 388202 -17315
rect 388270 -17371 388326 -17315
rect 388394 -17371 388450 -17315
rect 388518 -17371 388574 -17315
rect 388642 -17371 388698 -17315
rect 388766 -17371 388822 -17315
rect 388890 -17371 388946 -17315
rect 389014 -17371 389070 -17315
rect 389138 -17371 389194 -17315
rect 389262 -17371 389318 -17315
rect 389386 -17371 389442 -17315
rect 389510 -17371 389566 -17315
rect 389634 -17371 389690 -17315
rect 389758 -17371 389814 -17315
rect 389882 -17371 389938 -17315
rect 390006 -17371 390062 -17315
rect 390130 -17371 390186 -17315
rect 390254 -17371 390310 -17315
rect 390378 -17371 390434 -17315
rect 390502 -17371 390558 -17315
rect 390626 -17371 390682 -17315
rect 390750 -17371 390806 -17315
rect 390874 -17371 390930 -17315
rect 390998 -17371 391054 -17315
rect 391122 -17371 391178 -17315
rect 391246 -17371 391302 -17315
rect 391370 -17371 391426 -17315
rect 391494 -17371 391550 -17315
rect 391618 -17371 391674 -17315
rect 391742 -17371 391798 -17315
rect 391866 -17371 391922 -17315
rect 391990 -17371 392046 -17315
rect 392114 -17371 392170 -17315
rect 392238 -17371 392294 -17315
rect 392362 -17371 392418 -17315
rect 392486 -17371 392542 -17315
rect 392610 -17371 392666 -17315
rect 392734 -17371 392790 -17315
rect 392858 -17371 392914 -17315
rect 392982 -17371 393038 -17315
rect 393106 -17371 393162 -17315
rect 393230 -17371 393286 -17315
rect 393354 -17371 393410 -17315
rect 393478 -17371 393534 -17315
rect 393602 -17371 393658 -17315
rect 393726 -17371 393782 -17315
rect 393850 -17371 393906 -17315
rect 393974 -17371 394030 -17315
rect 394098 -17371 394154 -17315
rect 394222 -17371 394278 -17315
rect 394346 -17371 394402 -17315
rect 394470 -17371 394526 -17315
rect 394594 -17371 394650 -17315
rect 394718 -17371 394774 -17315
rect 394842 -17371 394898 -17315
rect 394966 -17371 395022 -17315
rect 395090 -17371 395146 -17315
rect 395214 -17371 395270 -17315
rect 395338 -17371 395394 -17315
rect 395462 -17371 395518 -17315
rect 395586 -17371 395642 -17315
rect 395710 -17371 395766 -17315
rect 395898 -17371 395954 -17315
rect 396022 -17371 396078 -17315
rect 396146 -17371 396202 -17315
rect 396270 -17371 396326 -17315
rect 396394 -17371 396450 -17315
rect 396518 -17371 396574 -17315
rect 396642 -17371 396698 -17315
rect 396766 -17371 396822 -17315
rect 396890 -17371 396946 -17315
rect 397014 -17371 397070 -17315
rect 388146 -17495 388202 -17439
rect 388270 -17495 388326 -17439
rect 388394 -17495 388450 -17439
rect 388518 -17495 388574 -17439
rect 388642 -17495 388698 -17439
rect 388766 -17495 388822 -17439
rect 388890 -17495 388946 -17439
rect 389014 -17495 389070 -17439
rect 389138 -17495 389194 -17439
rect 389262 -17495 389318 -17439
rect 389386 -17495 389442 -17439
rect 389510 -17495 389566 -17439
rect 389634 -17495 389690 -17439
rect 389758 -17495 389814 -17439
rect 389882 -17495 389938 -17439
rect 390006 -17495 390062 -17439
rect 390130 -17495 390186 -17439
rect 390254 -17495 390310 -17439
rect 390378 -17495 390434 -17439
rect 390502 -17495 390558 -17439
rect 390626 -17495 390682 -17439
rect 390750 -17495 390806 -17439
rect 390874 -17495 390930 -17439
rect 390998 -17495 391054 -17439
rect 391122 -17495 391178 -17439
rect 391246 -17495 391302 -17439
rect 391370 -17495 391426 -17439
rect 391494 -17495 391550 -17439
rect 391618 -17495 391674 -17439
rect 391742 -17495 391798 -17439
rect 391866 -17495 391922 -17439
rect 391990 -17495 392046 -17439
rect 392114 -17495 392170 -17439
rect 392238 -17495 392294 -17439
rect 392362 -17495 392418 -17439
rect 392486 -17495 392542 -17439
rect 392610 -17495 392666 -17439
rect 392734 -17495 392790 -17439
rect 392858 -17495 392914 -17439
rect 392982 -17495 393038 -17439
rect 393106 -17495 393162 -17439
rect 393230 -17495 393286 -17439
rect 393354 -17495 393410 -17439
rect 393478 -17495 393534 -17439
rect 393602 -17495 393658 -17439
rect 393726 -17495 393782 -17439
rect 393850 -17495 393906 -17439
rect 393974 -17495 394030 -17439
rect 394098 -17495 394154 -17439
rect 394222 -17495 394278 -17439
rect 394346 -17495 394402 -17439
rect 394470 -17495 394526 -17439
rect 394594 -17495 394650 -17439
rect 394718 -17495 394774 -17439
rect 394842 -17495 394898 -17439
rect 394966 -17495 395022 -17439
rect 395090 -17495 395146 -17439
rect 395214 -17495 395270 -17439
rect 395338 -17495 395394 -17439
rect 395462 -17495 395518 -17439
rect 395586 -17495 395642 -17439
rect 395710 -17495 395766 -17439
rect 395898 -17495 395954 -17439
rect 396022 -17495 396078 -17439
rect 396146 -17495 396202 -17439
rect 396270 -17495 396326 -17439
rect 396394 -17495 396450 -17439
rect 396518 -17495 396574 -17439
rect 396642 -17495 396698 -17439
rect 396766 -17495 396822 -17439
rect 396890 -17495 396946 -17439
rect 397014 -17495 397070 -17439
rect 388146 -17619 388202 -17563
rect 388270 -17619 388326 -17563
rect 388394 -17619 388450 -17563
rect 388518 -17619 388574 -17563
rect 388642 -17619 388698 -17563
rect 388766 -17619 388822 -17563
rect 388890 -17619 388946 -17563
rect 389014 -17619 389070 -17563
rect 389138 -17619 389194 -17563
rect 389262 -17619 389318 -17563
rect 389386 -17619 389442 -17563
rect 389510 -17619 389566 -17563
rect 389634 -17619 389690 -17563
rect 389758 -17619 389814 -17563
rect 389882 -17619 389938 -17563
rect 390006 -17619 390062 -17563
rect 390130 -17619 390186 -17563
rect 390254 -17619 390310 -17563
rect 390378 -17619 390434 -17563
rect 390502 -17619 390558 -17563
rect 390626 -17619 390682 -17563
rect 390750 -17619 390806 -17563
rect 390874 -17619 390930 -17563
rect 390998 -17619 391054 -17563
rect 391122 -17619 391178 -17563
rect 391246 -17619 391302 -17563
rect 391370 -17619 391426 -17563
rect 391494 -17619 391550 -17563
rect 391618 -17619 391674 -17563
rect 391742 -17619 391798 -17563
rect 391866 -17619 391922 -17563
rect 391990 -17619 392046 -17563
rect 392114 -17619 392170 -17563
rect 392238 -17619 392294 -17563
rect 392362 -17619 392418 -17563
rect 392486 -17619 392542 -17563
rect 392610 -17619 392666 -17563
rect 392734 -17619 392790 -17563
rect 392858 -17619 392914 -17563
rect 392982 -17619 393038 -17563
rect 393106 -17619 393162 -17563
rect 393230 -17619 393286 -17563
rect 393354 -17619 393410 -17563
rect 393478 -17619 393534 -17563
rect 393602 -17619 393658 -17563
rect 393726 -17619 393782 -17563
rect 393850 -17619 393906 -17563
rect 393974 -17619 394030 -17563
rect 394098 -17619 394154 -17563
rect 394222 -17619 394278 -17563
rect 394346 -17619 394402 -17563
rect 394470 -17619 394526 -17563
rect 394594 -17619 394650 -17563
rect 394718 -17619 394774 -17563
rect 394842 -17619 394898 -17563
rect 394966 -17619 395022 -17563
rect 395090 -17619 395146 -17563
rect 395214 -17619 395270 -17563
rect 395338 -17619 395394 -17563
rect 395462 -17619 395518 -17563
rect 395586 -17619 395642 -17563
rect 395710 -17619 395766 -17563
rect 395898 -17619 395954 -17563
rect 396022 -17619 396078 -17563
rect 396146 -17619 396202 -17563
rect 396270 -17619 396326 -17563
rect 396394 -17619 396450 -17563
rect 396518 -17619 396574 -17563
rect 396642 -17619 396698 -17563
rect 396766 -17619 396822 -17563
rect 396890 -17619 396946 -17563
rect 397014 -17619 397070 -17563
rect 388114 -17914 388170 -17858
rect 388238 -17914 388294 -17858
rect 388362 -17914 388418 -17858
rect 388486 -17914 388542 -17858
rect 388610 -17914 388666 -17858
rect 388114 -18038 388170 -17982
rect 388238 -18038 388294 -17982
rect 388362 -18038 388418 -17982
rect 388486 -18038 388542 -17982
rect 388610 -18038 388666 -17982
rect 388114 -18162 388170 -18106
rect 388238 -18162 388294 -18106
rect 388362 -18162 388418 -18106
rect 388486 -18162 388542 -18106
rect 388610 -18162 388666 -18106
rect 388114 -18286 388170 -18230
rect 388238 -18286 388294 -18230
rect 388362 -18286 388418 -18230
rect 388486 -18286 388542 -18230
rect 388610 -18286 388666 -18230
rect 388114 -18410 388170 -18354
rect 388238 -18410 388294 -18354
rect 388362 -18410 388418 -18354
rect 388486 -18410 388542 -18354
rect 388610 -18410 388666 -18354
rect 388114 -18534 388170 -18478
rect 388238 -18534 388294 -18478
rect 388362 -18534 388418 -18478
rect 388486 -18534 388542 -18478
rect 388610 -18534 388666 -18478
rect 388114 -18658 388170 -18602
rect 388238 -18658 388294 -18602
rect 388362 -18658 388418 -18602
rect 388486 -18658 388542 -18602
rect 388610 -18658 388666 -18602
rect 388114 -18782 388170 -18726
rect 388238 -18782 388294 -18726
rect 388362 -18782 388418 -18726
rect 388486 -18782 388542 -18726
rect 388610 -18782 388666 -18726
rect 388114 -18906 388170 -18850
rect 388238 -18906 388294 -18850
rect 388362 -18906 388418 -18850
rect 388486 -18906 388542 -18850
rect 388610 -18906 388666 -18850
rect 388114 -19030 388170 -18974
rect 388238 -19030 388294 -18974
rect 388362 -19030 388418 -18974
rect 388486 -19030 388542 -18974
rect 388610 -19030 388666 -18974
rect 388114 -19154 388170 -19098
rect 388238 -19154 388294 -19098
rect 388362 -19154 388418 -19098
rect 388486 -19154 388542 -19098
rect 388610 -19154 388666 -19098
rect 388114 -19278 388170 -19222
rect 388238 -19278 388294 -19222
rect 388362 -19278 388418 -19222
rect 388486 -19278 388542 -19222
rect 388610 -19278 388666 -19222
rect 388114 -19402 388170 -19346
rect 388238 -19402 388294 -19346
rect 388362 -19402 388418 -19346
rect 388486 -19402 388542 -19346
rect 388610 -19402 388666 -19346
rect 388114 -19526 388170 -19470
rect 388238 -19526 388294 -19470
rect 388362 -19526 388418 -19470
rect 388486 -19526 388542 -19470
rect 388610 -19526 388666 -19470
rect 388114 -19650 388170 -19594
rect 388238 -19650 388294 -19594
rect 388362 -19650 388418 -19594
rect 388486 -19650 388542 -19594
rect 388610 -19650 388666 -19594
rect 388114 -19774 388170 -19718
rect 388238 -19774 388294 -19718
rect 388362 -19774 388418 -19718
rect 388486 -19774 388542 -19718
rect 388610 -19774 388666 -19718
rect 388114 -19898 388170 -19842
rect 388238 -19898 388294 -19842
rect 388362 -19898 388418 -19842
rect 388486 -19898 388542 -19842
rect 388610 -19898 388666 -19842
rect 388114 -20022 388170 -19966
rect 388238 -20022 388294 -19966
rect 388362 -20022 388418 -19966
rect 388486 -20022 388542 -19966
rect 388610 -20022 388666 -19966
rect 388114 -20146 388170 -20090
rect 388238 -20146 388294 -20090
rect 388362 -20146 388418 -20090
rect 388486 -20146 388542 -20090
rect 388610 -20146 388666 -20090
rect 388114 -20270 388170 -20214
rect 388238 -20270 388294 -20214
rect 388362 -20270 388418 -20214
rect 388486 -20270 388542 -20214
rect 388610 -20270 388666 -20214
rect 388114 -20394 388170 -20338
rect 388238 -20394 388294 -20338
rect 388362 -20394 388418 -20338
rect 388486 -20394 388542 -20338
rect 388610 -20394 388666 -20338
rect 388114 -20518 388170 -20462
rect 388238 -20518 388294 -20462
rect 388362 -20518 388418 -20462
rect 388486 -20518 388542 -20462
rect 388610 -20518 388666 -20462
rect 388114 -20642 388170 -20586
rect 388238 -20642 388294 -20586
rect 388362 -20642 388418 -20586
rect 388486 -20642 388542 -20586
rect 388610 -20642 388666 -20586
rect 388114 -20766 388170 -20710
rect 388238 -20766 388294 -20710
rect 388362 -20766 388418 -20710
rect 388486 -20766 388542 -20710
rect 388610 -20766 388666 -20710
rect 388114 -20890 388170 -20834
rect 388238 -20890 388294 -20834
rect 388362 -20890 388418 -20834
rect 388486 -20890 388542 -20834
rect 388610 -20890 388666 -20834
rect 388114 -21014 388170 -20958
rect 388238 -21014 388294 -20958
rect 388362 -21014 388418 -20958
rect 388486 -21014 388542 -20958
rect 388610 -21014 388666 -20958
rect 388114 -21138 388170 -21082
rect 388238 -21138 388294 -21082
rect 388362 -21138 388418 -21082
rect 388486 -21138 388542 -21082
rect 388610 -21138 388666 -21082
rect 388114 -21262 388170 -21206
rect 388238 -21262 388294 -21206
rect 388362 -21262 388418 -21206
rect 388486 -21262 388542 -21206
rect 388610 -21262 388666 -21206
rect 388114 -21386 388170 -21330
rect 388238 -21386 388294 -21330
rect 388362 -21386 388418 -21330
rect 388486 -21386 388542 -21330
rect 388610 -21386 388666 -21330
rect 388114 -21510 388170 -21454
rect 388238 -21510 388294 -21454
rect 388362 -21510 388418 -21454
rect 388486 -21510 388542 -21454
rect 388610 -21510 388666 -21454
rect 388114 -21634 388170 -21578
rect 388238 -21634 388294 -21578
rect 388362 -21634 388418 -21578
rect 388486 -21634 388542 -21578
rect 388610 -21634 388666 -21578
rect 388114 -21758 388170 -21702
rect 388238 -21758 388294 -21702
rect 388362 -21758 388418 -21702
rect 388486 -21758 388542 -21702
rect 388610 -21758 388666 -21702
rect 388114 -21882 388170 -21826
rect 388238 -21882 388294 -21826
rect 388362 -21882 388418 -21826
rect 388486 -21882 388542 -21826
rect 388610 -21882 388666 -21826
rect 388114 -22006 388170 -21950
rect 388238 -22006 388294 -21950
rect 388362 -22006 388418 -21950
rect 388486 -22006 388542 -21950
rect 388610 -22006 388666 -21950
rect 388114 -22130 388170 -22074
rect 388238 -22130 388294 -22074
rect 388362 -22130 388418 -22074
rect 388486 -22130 388542 -22074
rect 388610 -22130 388666 -22074
rect 388114 -22254 388170 -22198
rect 388238 -22254 388294 -22198
rect 388362 -22254 388418 -22198
rect 388486 -22254 388542 -22198
rect 388610 -22254 388666 -22198
rect 388114 -22378 388170 -22322
rect 388238 -22378 388294 -22322
rect 388362 -22378 388418 -22322
rect 388486 -22378 388542 -22322
rect 388610 -22378 388666 -22322
rect 388114 -22502 388170 -22446
rect 388238 -22502 388294 -22446
rect 388362 -22502 388418 -22446
rect 388486 -22502 388542 -22446
rect 388610 -22502 388666 -22446
rect 388114 -22626 388170 -22570
rect 388238 -22626 388294 -22570
rect 388362 -22626 388418 -22570
rect 388486 -22626 388542 -22570
rect 388610 -22626 388666 -22570
rect 388114 -22750 388170 -22694
rect 388238 -22750 388294 -22694
rect 388362 -22750 388418 -22694
rect 388486 -22750 388542 -22694
rect 388610 -22750 388666 -22694
rect 388114 -22874 388170 -22818
rect 388238 -22874 388294 -22818
rect 388362 -22874 388418 -22818
rect 388486 -22874 388542 -22818
rect 388610 -22874 388666 -22818
rect 388114 -22998 388170 -22942
rect 388238 -22998 388294 -22942
rect 388362 -22998 388418 -22942
rect 388486 -22998 388542 -22942
rect 388610 -22998 388666 -22942
rect 388114 -23122 388170 -23066
rect 388238 -23122 388294 -23066
rect 388362 -23122 388418 -23066
rect 388486 -23122 388542 -23066
rect 388610 -23122 388666 -23066
rect 388114 -23246 388170 -23190
rect 388238 -23246 388294 -23190
rect 388362 -23246 388418 -23190
rect 388486 -23246 388542 -23190
rect 388610 -23246 388666 -23190
rect 388114 -23370 388170 -23314
rect 388238 -23370 388294 -23314
rect 388362 -23370 388418 -23314
rect 388486 -23370 388542 -23314
rect 388610 -23370 388666 -23314
rect 388114 -23494 388170 -23438
rect 388238 -23494 388294 -23438
rect 388362 -23494 388418 -23438
rect 388486 -23494 388542 -23438
rect 388610 -23494 388666 -23438
rect 388114 -23618 388170 -23562
rect 388238 -23618 388294 -23562
rect 388362 -23618 388418 -23562
rect 388486 -23618 388542 -23562
rect 388610 -23618 388666 -23562
rect 388114 -23742 388170 -23686
rect 388238 -23742 388294 -23686
rect 388362 -23742 388418 -23686
rect 388486 -23742 388542 -23686
rect 388610 -23742 388666 -23686
rect 388114 -23866 388170 -23810
rect 388238 -23866 388294 -23810
rect 388362 -23866 388418 -23810
rect 388486 -23866 388542 -23810
rect 388610 -23866 388666 -23810
rect 388114 -23990 388170 -23934
rect 388238 -23990 388294 -23934
rect 388362 -23990 388418 -23934
rect 388486 -23990 388542 -23934
rect 388610 -23990 388666 -23934
rect 388114 -24114 388170 -24058
rect 388238 -24114 388294 -24058
rect 388362 -24114 388418 -24058
rect 388486 -24114 388542 -24058
rect 388610 -24114 388666 -24058
rect 388114 -24238 388170 -24182
rect 388238 -24238 388294 -24182
rect 388362 -24238 388418 -24182
rect 388486 -24238 388542 -24182
rect 388610 -24238 388666 -24182
rect 388114 -24362 388170 -24306
rect 388238 -24362 388294 -24306
rect 388362 -24362 388418 -24306
rect 388486 -24362 388542 -24306
rect 388610 -24362 388666 -24306
rect 388114 -24486 388170 -24430
rect 388238 -24486 388294 -24430
rect 388362 -24486 388418 -24430
rect 388486 -24486 388542 -24430
rect 388610 -24486 388666 -24430
rect 388114 -24610 388170 -24554
rect 388238 -24610 388294 -24554
rect 388362 -24610 388418 -24554
rect 388486 -24610 388542 -24554
rect 388610 -24610 388666 -24554
rect 388114 -24734 388170 -24678
rect 388238 -24734 388294 -24678
rect 388362 -24734 388418 -24678
rect 388486 -24734 388542 -24678
rect 388610 -24734 388666 -24678
rect 388114 -24858 388170 -24802
rect 388238 -24858 388294 -24802
rect 388362 -24858 388418 -24802
rect 388486 -24858 388542 -24802
rect 388610 -24858 388666 -24802
rect 388114 -24982 388170 -24926
rect 388238 -24982 388294 -24926
rect 388362 -24982 388418 -24926
rect 388486 -24982 388542 -24926
rect 388610 -24982 388666 -24926
rect 388114 -25106 388170 -25050
rect 388238 -25106 388294 -25050
rect 388362 -25106 388418 -25050
rect 388486 -25106 388542 -25050
rect 388610 -25106 388666 -25050
rect 388114 -25230 388170 -25174
rect 388238 -25230 388294 -25174
rect 388362 -25230 388418 -25174
rect 388486 -25230 388542 -25174
rect 388610 -25230 388666 -25174
rect 388114 -25354 388170 -25298
rect 388238 -25354 388294 -25298
rect 388362 -25354 388418 -25298
rect 388486 -25354 388542 -25298
rect 388610 -25354 388666 -25298
rect 388114 -25478 388170 -25422
rect 388238 -25478 388294 -25422
rect 388362 -25478 388418 -25422
rect 388486 -25478 388542 -25422
rect 388610 -25478 388666 -25422
rect 389141 -18006 389197 -17950
rect 389283 -18006 389339 -17950
rect 389141 -18148 389197 -18092
rect 389283 -18148 389339 -18092
rect 389141 -18290 389197 -18234
rect 389283 -18290 389339 -18234
rect 389141 -18432 389197 -18376
rect 389283 -18432 389339 -18376
rect 389141 -18574 389197 -18518
rect 389283 -18574 389339 -18518
rect 389141 -18716 389197 -18660
rect 389283 -18716 389339 -18660
rect 389141 -18858 389197 -18802
rect 389283 -18858 389339 -18802
rect 389141 -19000 389197 -18944
rect 389283 -19000 389339 -18944
rect 389141 -19142 389197 -19086
rect 389283 -19142 389339 -19086
rect 389141 -19284 389197 -19228
rect 389283 -19284 389339 -19228
rect 389141 -19426 389197 -19370
rect 389283 -19426 389339 -19370
rect 389141 -19568 389197 -19512
rect 389283 -19568 389339 -19512
rect 389141 -19710 389197 -19654
rect 389283 -19710 389339 -19654
rect 389141 -19852 389197 -19796
rect 389283 -19852 389339 -19796
rect 389141 -19994 389197 -19938
rect 389283 -19994 389339 -19938
rect 389141 -20136 389197 -20080
rect 389283 -20136 389339 -20080
rect 389141 -20278 389197 -20222
rect 389283 -20278 389339 -20222
rect 389141 -20420 389197 -20364
rect 389283 -20420 389339 -20364
rect 389141 -20562 389197 -20506
rect 389283 -20562 389339 -20506
rect 389141 -20704 389197 -20648
rect 389283 -20704 389339 -20648
rect 389141 -20846 389197 -20790
rect 389283 -20846 389339 -20790
rect 389141 -20988 389197 -20932
rect 389283 -20988 389339 -20932
rect 389141 -21130 389197 -21074
rect 389283 -21130 389339 -21074
rect 389141 -21272 389197 -21216
rect 389283 -21272 389339 -21216
rect 389141 -21414 389197 -21358
rect 389283 -21414 389339 -21358
rect 389141 -21556 389197 -21500
rect 389283 -21556 389339 -21500
rect 389141 -21698 389197 -21642
rect 389283 -21698 389339 -21642
rect 389141 -21840 389197 -21784
rect 389283 -21840 389339 -21784
rect 389141 -21982 389197 -21926
rect 389283 -21982 389339 -21926
rect 389141 -22124 389197 -22068
rect 389283 -22124 389339 -22068
rect 389141 -22266 389197 -22210
rect 389283 -22266 389339 -22210
rect 389141 -22408 389197 -22352
rect 389283 -22408 389339 -22352
rect 389141 -22550 389197 -22494
rect 389283 -22550 389339 -22494
rect 389141 -22692 389197 -22636
rect 389283 -22692 389339 -22636
rect 389141 -22834 389197 -22778
rect 389283 -22834 389339 -22778
rect 389141 -22976 389197 -22920
rect 389283 -22976 389339 -22920
rect 389141 -23118 389197 -23062
rect 389283 -23118 389339 -23062
rect 389141 -23260 389197 -23204
rect 389283 -23260 389339 -23204
rect 389141 -23402 389197 -23346
rect 389283 -23402 389339 -23346
rect 389141 -23544 389197 -23488
rect 389283 -23544 389339 -23488
rect 389141 -23686 389197 -23630
rect 389283 -23686 389339 -23630
rect 389141 -23828 389197 -23772
rect 389283 -23828 389339 -23772
rect 389141 -23970 389197 -23914
rect 389283 -23970 389339 -23914
rect 389141 -24112 389197 -24056
rect 389283 -24112 389339 -24056
rect 389141 -24254 389197 -24198
rect 389283 -24254 389339 -24198
rect 389141 -24396 389197 -24340
rect 389283 -24396 389339 -24340
rect 389141 -24538 389197 -24482
rect 389283 -24538 389339 -24482
rect 389141 -24680 389197 -24624
rect 389283 -24680 389339 -24624
rect 389141 -24822 389197 -24766
rect 389283 -24822 389339 -24766
rect 389141 -24964 389197 -24908
rect 389283 -24964 389339 -24908
rect 389141 -25106 389197 -25050
rect 389283 -25106 389339 -25050
rect 389141 -25248 389197 -25192
rect 389283 -25248 389339 -25192
rect 389141 -25390 389197 -25334
rect 389283 -25390 389339 -25334
rect 389141 -25532 389197 -25476
rect 389283 -25532 389339 -25476
rect 389542 -18006 389598 -17950
rect 389684 -18006 389740 -17950
rect 389542 -18148 389598 -18092
rect 389684 -18148 389740 -18092
rect 389542 -18290 389598 -18234
rect 389684 -18290 389740 -18234
rect 389542 -18432 389598 -18376
rect 389684 -18432 389740 -18376
rect 389542 -18574 389598 -18518
rect 389684 -18574 389740 -18518
rect 389542 -18716 389598 -18660
rect 389684 -18716 389740 -18660
rect 389542 -18858 389598 -18802
rect 389684 -18858 389740 -18802
rect 389542 -19000 389598 -18944
rect 389684 -19000 389740 -18944
rect 389542 -19142 389598 -19086
rect 389684 -19142 389740 -19086
rect 389542 -19284 389598 -19228
rect 389684 -19284 389740 -19228
rect 389542 -19426 389598 -19370
rect 389684 -19426 389740 -19370
rect 389542 -19568 389598 -19512
rect 389684 -19568 389740 -19512
rect 389542 -19710 389598 -19654
rect 389684 -19710 389740 -19654
rect 389542 -19852 389598 -19796
rect 389684 -19852 389740 -19796
rect 389542 -19994 389598 -19938
rect 389684 -19994 389740 -19938
rect 389542 -20136 389598 -20080
rect 389684 -20136 389740 -20080
rect 389542 -20278 389598 -20222
rect 389684 -20278 389740 -20222
rect 389542 -20420 389598 -20364
rect 389684 -20420 389740 -20364
rect 389542 -20562 389598 -20506
rect 389684 -20562 389740 -20506
rect 389542 -20704 389598 -20648
rect 389684 -20704 389740 -20648
rect 389542 -20846 389598 -20790
rect 389684 -20846 389740 -20790
rect 389542 -20988 389598 -20932
rect 389684 -20988 389740 -20932
rect 389542 -21130 389598 -21074
rect 389684 -21130 389740 -21074
rect 389542 -21272 389598 -21216
rect 389684 -21272 389740 -21216
rect 389542 -21414 389598 -21358
rect 389684 -21414 389740 -21358
rect 389542 -21556 389598 -21500
rect 389684 -21556 389740 -21500
rect 389542 -21698 389598 -21642
rect 389684 -21698 389740 -21642
rect 389542 -21840 389598 -21784
rect 389684 -21840 389740 -21784
rect 389542 -21982 389598 -21926
rect 389684 -21982 389740 -21926
rect 389542 -22124 389598 -22068
rect 389684 -22124 389740 -22068
rect 389542 -22266 389598 -22210
rect 389684 -22266 389740 -22210
rect 389542 -22408 389598 -22352
rect 389684 -22408 389740 -22352
rect 389542 -22550 389598 -22494
rect 389684 -22550 389740 -22494
rect 389542 -22692 389598 -22636
rect 389684 -22692 389740 -22636
rect 389542 -22834 389598 -22778
rect 389684 -22834 389740 -22778
rect 389542 -22976 389598 -22920
rect 389684 -22976 389740 -22920
rect 389542 -23118 389598 -23062
rect 389684 -23118 389740 -23062
rect 389542 -23260 389598 -23204
rect 389684 -23260 389740 -23204
rect 389542 -23402 389598 -23346
rect 389684 -23402 389740 -23346
rect 389542 -23544 389598 -23488
rect 389684 -23544 389740 -23488
rect 389542 -23686 389598 -23630
rect 389684 -23686 389740 -23630
rect 389542 -23828 389598 -23772
rect 389684 -23828 389740 -23772
rect 389542 -23970 389598 -23914
rect 389684 -23970 389740 -23914
rect 389542 -24112 389598 -24056
rect 389684 -24112 389740 -24056
rect 389542 -24254 389598 -24198
rect 389684 -24254 389740 -24198
rect 389542 -24396 389598 -24340
rect 389684 -24396 389740 -24340
rect 389542 -24538 389598 -24482
rect 389684 -24538 389740 -24482
rect 389542 -24680 389598 -24624
rect 389684 -24680 389740 -24624
rect 389542 -24822 389598 -24766
rect 389684 -24822 389740 -24766
rect 389542 -24964 389598 -24908
rect 389684 -24964 389740 -24908
rect 389542 -25106 389598 -25050
rect 389684 -25106 389740 -25050
rect 389542 -25248 389598 -25192
rect 389684 -25248 389740 -25192
rect 389542 -25390 389598 -25334
rect 389684 -25390 389740 -25334
rect 389542 -25532 389598 -25476
rect 389684 -25532 389740 -25476
rect 389942 -18006 389998 -17950
rect 390084 -18006 390140 -17950
rect 389942 -18148 389998 -18092
rect 390084 -18148 390140 -18092
rect 389942 -18290 389998 -18234
rect 390084 -18290 390140 -18234
rect 389942 -18432 389998 -18376
rect 390084 -18432 390140 -18376
rect 389942 -18574 389998 -18518
rect 390084 -18574 390140 -18518
rect 389942 -18716 389998 -18660
rect 390084 -18716 390140 -18660
rect 389942 -18858 389998 -18802
rect 390084 -18858 390140 -18802
rect 389942 -19000 389998 -18944
rect 390084 -19000 390140 -18944
rect 389942 -19142 389998 -19086
rect 390084 -19142 390140 -19086
rect 389942 -19284 389998 -19228
rect 390084 -19284 390140 -19228
rect 389942 -19426 389998 -19370
rect 390084 -19426 390140 -19370
rect 389942 -19568 389998 -19512
rect 390084 -19568 390140 -19512
rect 389942 -19710 389998 -19654
rect 390084 -19710 390140 -19654
rect 389942 -19852 389998 -19796
rect 390084 -19852 390140 -19796
rect 389942 -19994 389998 -19938
rect 390084 -19994 390140 -19938
rect 389942 -20136 389998 -20080
rect 390084 -20136 390140 -20080
rect 389942 -20278 389998 -20222
rect 390084 -20278 390140 -20222
rect 389942 -20420 389998 -20364
rect 390084 -20420 390140 -20364
rect 389942 -20562 389998 -20506
rect 390084 -20562 390140 -20506
rect 389942 -20704 389998 -20648
rect 390084 -20704 390140 -20648
rect 389942 -20846 389998 -20790
rect 390084 -20846 390140 -20790
rect 389942 -20988 389998 -20932
rect 390084 -20988 390140 -20932
rect 389942 -21130 389998 -21074
rect 390084 -21130 390140 -21074
rect 389942 -21272 389998 -21216
rect 390084 -21272 390140 -21216
rect 389942 -21414 389998 -21358
rect 390084 -21414 390140 -21358
rect 389942 -21556 389998 -21500
rect 390084 -21556 390140 -21500
rect 389942 -21698 389998 -21642
rect 390084 -21698 390140 -21642
rect 389942 -21840 389998 -21784
rect 390084 -21840 390140 -21784
rect 389942 -21982 389998 -21926
rect 390084 -21982 390140 -21926
rect 389942 -22124 389998 -22068
rect 390084 -22124 390140 -22068
rect 389942 -22266 389998 -22210
rect 390084 -22266 390140 -22210
rect 389942 -22408 389998 -22352
rect 390084 -22408 390140 -22352
rect 389942 -22550 389998 -22494
rect 390084 -22550 390140 -22494
rect 389942 -22692 389998 -22636
rect 390084 -22692 390140 -22636
rect 389942 -22834 389998 -22778
rect 390084 -22834 390140 -22778
rect 389942 -22976 389998 -22920
rect 390084 -22976 390140 -22920
rect 389942 -23118 389998 -23062
rect 390084 -23118 390140 -23062
rect 389942 -23260 389998 -23204
rect 390084 -23260 390140 -23204
rect 389942 -23402 389998 -23346
rect 390084 -23402 390140 -23346
rect 389942 -23544 389998 -23488
rect 390084 -23544 390140 -23488
rect 389942 -23686 389998 -23630
rect 390084 -23686 390140 -23630
rect 389942 -23828 389998 -23772
rect 390084 -23828 390140 -23772
rect 389942 -23970 389998 -23914
rect 390084 -23970 390140 -23914
rect 389942 -24112 389998 -24056
rect 390084 -24112 390140 -24056
rect 389942 -24254 389998 -24198
rect 390084 -24254 390140 -24198
rect 389942 -24396 389998 -24340
rect 390084 -24396 390140 -24340
rect 389942 -24538 389998 -24482
rect 390084 -24538 390140 -24482
rect 389942 -24680 389998 -24624
rect 390084 -24680 390140 -24624
rect 389942 -24822 389998 -24766
rect 390084 -24822 390140 -24766
rect 389942 -24964 389998 -24908
rect 390084 -24964 390140 -24908
rect 389942 -25106 389998 -25050
rect 390084 -25106 390140 -25050
rect 389942 -25248 389998 -25192
rect 390084 -25248 390140 -25192
rect 389942 -25390 389998 -25334
rect 390084 -25390 390140 -25334
rect 389942 -25532 389998 -25476
rect 390084 -25532 390140 -25476
rect 390339 -18006 390395 -17950
rect 390481 -18006 390537 -17950
rect 390339 -18148 390395 -18092
rect 390481 -18148 390537 -18092
rect 390339 -18290 390395 -18234
rect 390481 -18290 390537 -18234
rect 390339 -18432 390395 -18376
rect 390481 -18432 390537 -18376
rect 390339 -18574 390395 -18518
rect 390481 -18574 390537 -18518
rect 390339 -18716 390395 -18660
rect 390481 -18716 390537 -18660
rect 390339 -18858 390395 -18802
rect 390481 -18858 390537 -18802
rect 390339 -19000 390395 -18944
rect 390481 -19000 390537 -18944
rect 390339 -19142 390395 -19086
rect 390481 -19142 390537 -19086
rect 390339 -19284 390395 -19228
rect 390481 -19284 390537 -19228
rect 390339 -19426 390395 -19370
rect 390481 -19426 390537 -19370
rect 390339 -19568 390395 -19512
rect 390481 -19568 390537 -19512
rect 390339 -19710 390395 -19654
rect 390481 -19710 390537 -19654
rect 390339 -19852 390395 -19796
rect 390481 -19852 390537 -19796
rect 390339 -19994 390395 -19938
rect 390481 -19994 390537 -19938
rect 390339 -20136 390395 -20080
rect 390481 -20136 390537 -20080
rect 390339 -20278 390395 -20222
rect 390481 -20278 390537 -20222
rect 390339 -20420 390395 -20364
rect 390481 -20420 390537 -20364
rect 390339 -20562 390395 -20506
rect 390481 -20562 390537 -20506
rect 390339 -20704 390395 -20648
rect 390481 -20704 390537 -20648
rect 390339 -20846 390395 -20790
rect 390481 -20846 390537 -20790
rect 390339 -20988 390395 -20932
rect 390481 -20988 390537 -20932
rect 390339 -21130 390395 -21074
rect 390481 -21130 390537 -21074
rect 390339 -21272 390395 -21216
rect 390481 -21272 390537 -21216
rect 390339 -21414 390395 -21358
rect 390481 -21414 390537 -21358
rect 390339 -21556 390395 -21500
rect 390481 -21556 390537 -21500
rect 390339 -21698 390395 -21642
rect 390481 -21698 390537 -21642
rect 390339 -21840 390395 -21784
rect 390481 -21840 390537 -21784
rect 390339 -21982 390395 -21926
rect 390481 -21982 390537 -21926
rect 390339 -22124 390395 -22068
rect 390481 -22124 390537 -22068
rect 390339 -22266 390395 -22210
rect 390481 -22266 390537 -22210
rect 390339 -22408 390395 -22352
rect 390481 -22408 390537 -22352
rect 390339 -22550 390395 -22494
rect 390481 -22550 390537 -22494
rect 390339 -22692 390395 -22636
rect 390481 -22692 390537 -22636
rect 390339 -22834 390395 -22778
rect 390481 -22834 390537 -22778
rect 390339 -22976 390395 -22920
rect 390481 -22976 390537 -22920
rect 390339 -23118 390395 -23062
rect 390481 -23118 390537 -23062
rect 390339 -23260 390395 -23204
rect 390481 -23260 390537 -23204
rect 390339 -23402 390395 -23346
rect 390481 -23402 390537 -23346
rect 390339 -23544 390395 -23488
rect 390481 -23544 390537 -23488
rect 390339 -23686 390395 -23630
rect 390481 -23686 390537 -23630
rect 390339 -23828 390395 -23772
rect 390481 -23828 390537 -23772
rect 390339 -23970 390395 -23914
rect 390481 -23970 390537 -23914
rect 390339 -24112 390395 -24056
rect 390481 -24112 390537 -24056
rect 390339 -24254 390395 -24198
rect 390481 -24254 390537 -24198
rect 390339 -24396 390395 -24340
rect 390481 -24396 390537 -24340
rect 390339 -24538 390395 -24482
rect 390481 -24538 390537 -24482
rect 390339 -24680 390395 -24624
rect 390481 -24680 390537 -24624
rect 390339 -24822 390395 -24766
rect 390481 -24822 390537 -24766
rect 390339 -24964 390395 -24908
rect 390481 -24964 390537 -24908
rect 390339 -25106 390395 -25050
rect 390481 -25106 390537 -25050
rect 390339 -25248 390395 -25192
rect 390481 -25248 390537 -25192
rect 390339 -25390 390395 -25334
rect 390481 -25390 390537 -25334
rect 390339 -25532 390395 -25476
rect 390481 -25532 390537 -25476
rect 390736 -18006 390792 -17950
rect 390878 -18006 390934 -17950
rect 390736 -18148 390792 -18092
rect 390878 -18148 390934 -18092
rect 390736 -18290 390792 -18234
rect 390878 -18290 390934 -18234
rect 390736 -18432 390792 -18376
rect 390878 -18432 390934 -18376
rect 390736 -18574 390792 -18518
rect 390878 -18574 390934 -18518
rect 390736 -18716 390792 -18660
rect 390878 -18716 390934 -18660
rect 390736 -18858 390792 -18802
rect 390878 -18858 390934 -18802
rect 390736 -19000 390792 -18944
rect 390878 -19000 390934 -18944
rect 390736 -19142 390792 -19086
rect 390878 -19142 390934 -19086
rect 390736 -19284 390792 -19228
rect 390878 -19284 390934 -19228
rect 390736 -19426 390792 -19370
rect 390878 -19426 390934 -19370
rect 390736 -19568 390792 -19512
rect 390878 -19568 390934 -19512
rect 390736 -19710 390792 -19654
rect 390878 -19710 390934 -19654
rect 390736 -19852 390792 -19796
rect 390878 -19852 390934 -19796
rect 390736 -19994 390792 -19938
rect 390878 -19994 390934 -19938
rect 390736 -20136 390792 -20080
rect 390878 -20136 390934 -20080
rect 390736 -20278 390792 -20222
rect 390878 -20278 390934 -20222
rect 390736 -20420 390792 -20364
rect 390878 -20420 390934 -20364
rect 390736 -20562 390792 -20506
rect 390878 -20562 390934 -20506
rect 390736 -20704 390792 -20648
rect 390878 -20704 390934 -20648
rect 390736 -20846 390792 -20790
rect 390878 -20846 390934 -20790
rect 390736 -20988 390792 -20932
rect 390878 -20988 390934 -20932
rect 390736 -21130 390792 -21074
rect 390878 -21130 390934 -21074
rect 390736 -21272 390792 -21216
rect 390878 -21272 390934 -21216
rect 390736 -21414 390792 -21358
rect 390878 -21414 390934 -21358
rect 390736 -21556 390792 -21500
rect 390878 -21556 390934 -21500
rect 390736 -21698 390792 -21642
rect 390878 -21698 390934 -21642
rect 390736 -21840 390792 -21784
rect 390878 -21840 390934 -21784
rect 390736 -21982 390792 -21926
rect 390878 -21982 390934 -21926
rect 390736 -22124 390792 -22068
rect 390878 -22124 390934 -22068
rect 390736 -22266 390792 -22210
rect 390878 -22266 390934 -22210
rect 390736 -22408 390792 -22352
rect 390878 -22408 390934 -22352
rect 390736 -22550 390792 -22494
rect 390878 -22550 390934 -22494
rect 390736 -22692 390792 -22636
rect 390878 -22692 390934 -22636
rect 390736 -22834 390792 -22778
rect 390878 -22834 390934 -22778
rect 390736 -22976 390792 -22920
rect 390878 -22976 390934 -22920
rect 390736 -23118 390792 -23062
rect 390878 -23118 390934 -23062
rect 390736 -23260 390792 -23204
rect 390878 -23260 390934 -23204
rect 390736 -23402 390792 -23346
rect 390878 -23402 390934 -23346
rect 390736 -23544 390792 -23488
rect 390878 -23544 390934 -23488
rect 390736 -23686 390792 -23630
rect 390878 -23686 390934 -23630
rect 390736 -23828 390792 -23772
rect 390878 -23828 390934 -23772
rect 390736 -23970 390792 -23914
rect 390878 -23970 390934 -23914
rect 390736 -24112 390792 -24056
rect 390878 -24112 390934 -24056
rect 390736 -24254 390792 -24198
rect 390878 -24254 390934 -24198
rect 390736 -24396 390792 -24340
rect 390878 -24396 390934 -24340
rect 390736 -24538 390792 -24482
rect 390878 -24538 390934 -24482
rect 390736 -24680 390792 -24624
rect 390878 -24680 390934 -24624
rect 390736 -24822 390792 -24766
rect 390878 -24822 390934 -24766
rect 390736 -24964 390792 -24908
rect 390878 -24964 390934 -24908
rect 390736 -25106 390792 -25050
rect 390878 -25106 390934 -25050
rect 390736 -25248 390792 -25192
rect 390878 -25248 390934 -25192
rect 390736 -25390 390792 -25334
rect 390878 -25390 390934 -25334
rect 390736 -25532 390792 -25476
rect 390878 -25532 390934 -25476
rect 391140 -18006 391196 -17950
rect 391282 -18006 391338 -17950
rect 391140 -18148 391196 -18092
rect 391282 -18148 391338 -18092
rect 391140 -18290 391196 -18234
rect 391282 -18290 391338 -18234
rect 391140 -18432 391196 -18376
rect 391282 -18432 391338 -18376
rect 391140 -18574 391196 -18518
rect 391282 -18574 391338 -18518
rect 391140 -18716 391196 -18660
rect 391282 -18716 391338 -18660
rect 391140 -18858 391196 -18802
rect 391282 -18858 391338 -18802
rect 391140 -19000 391196 -18944
rect 391282 -19000 391338 -18944
rect 391140 -19142 391196 -19086
rect 391282 -19142 391338 -19086
rect 391140 -19284 391196 -19228
rect 391282 -19284 391338 -19228
rect 391140 -19426 391196 -19370
rect 391282 -19426 391338 -19370
rect 391140 -19568 391196 -19512
rect 391282 -19568 391338 -19512
rect 391140 -19710 391196 -19654
rect 391282 -19710 391338 -19654
rect 391140 -19852 391196 -19796
rect 391282 -19852 391338 -19796
rect 391140 -19994 391196 -19938
rect 391282 -19994 391338 -19938
rect 391140 -20136 391196 -20080
rect 391282 -20136 391338 -20080
rect 391140 -20278 391196 -20222
rect 391282 -20278 391338 -20222
rect 391140 -20420 391196 -20364
rect 391282 -20420 391338 -20364
rect 391140 -20562 391196 -20506
rect 391282 -20562 391338 -20506
rect 391140 -20704 391196 -20648
rect 391282 -20704 391338 -20648
rect 391140 -20846 391196 -20790
rect 391282 -20846 391338 -20790
rect 391140 -20988 391196 -20932
rect 391282 -20988 391338 -20932
rect 391140 -21130 391196 -21074
rect 391282 -21130 391338 -21074
rect 391140 -21272 391196 -21216
rect 391282 -21272 391338 -21216
rect 391140 -21414 391196 -21358
rect 391282 -21414 391338 -21358
rect 391140 -21556 391196 -21500
rect 391282 -21556 391338 -21500
rect 391140 -21698 391196 -21642
rect 391282 -21698 391338 -21642
rect 391140 -21840 391196 -21784
rect 391282 -21840 391338 -21784
rect 391140 -21982 391196 -21926
rect 391282 -21982 391338 -21926
rect 391140 -22124 391196 -22068
rect 391282 -22124 391338 -22068
rect 391140 -22266 391196 -22210
rect 391282 -22266 391338 -22210
rect 391140 -22408 391196 -22352
rect 391282 -22408 391338 -22352
rect 391140 -22550 391196 -22494
rect 391282 -22550 391338 -22494
rect 391140 -22692 391196 -22636
rect 391282 -22692 391338 -22636
rect 391140 -22834 391196 -22778
rect 391282 -22834 391338 -22778
rect 391140 -22976 391196 -22920
rect 391282 -22976 391338 -22920
rect 391140 -23118 391196 -23062
rect 391282 -23118 391338 -23062
rect 391140 -23260 391196 -23204
rect 391282 -23260 391338 -23204
rect 391140 -23402 391196 -23346
rect 391282 -23402 391338 -23346
rect 391140 -23544 391196 -23488
rect 391282 -23544 391338 -23488
rect 391140 -23686 391196 -23630
rect 391282 -23686 391338 -23630
rect 391140 -23828 391196 -23772
rect 391282 -23828 391338 -23772
rect 391140 -23970 391196 -23914
rect 391282 -23970 391338 -23914
rect 391140 -24112 391196 -24056
rect 391282 -24112 391338 -24056
rect 391140 -24254 391196 -24198
rect 391282 -24254 391338 -24198
rect 391140 -24396 391196 -24340
rect 391282 -24396 391338 -24340
rect 391140 -24538 391196 -24482
rect 391282 -24538 391338 -24482
rect 391140 -24680 391196 -24624
rect 391282 -24680 391338 -24624
rect 391140 -24822 391196 -24766
rect 391282 -24822 391338 -24766
rect 391140 -24964 391196 -24908
rect 391282 -24964 391338 -24908
rect 391140 -25106 391196 -25050
rect 391282 -25106 391338 -25050
rect 391140 -25248 391196 -25192
rect 391282 -25248 391338 -25192
rect 391140 -25390 391196 -25334
rect 391282 -25390 391338 -25334
rect 391140 -25532 391196 -25476
rect 391282 -25532 391338 -25476
rect 391536 -18006 391592 -17950
rect 391678 -18006 391734 -17950
rect 391536 -18148 391592 -18092
rect 391678 -18148 391734 -18092
rect 391536 -18290 391592 -18234
rect 391678 -18290 391734 -18234
rect 391536 -18432 391592 -18376
rect 391678 -18432 391734 -18376
rect 391536 -18574 391592 -18518
rect 391678 -18574 391734 -18518
rect 391536 -18716 391592 -18660
rect 391678 -18716 391734 -18660
rect 391536 -18858 391592 -18802
rect 391678 -18858 391734 -18802
rect 391536 -19000 391592 -18944
rect 391678 -19000 391734 -18944
rect 391536 -19142 391592 -19086
rect 391678 -19142 391734 -19086
rect 391536 -19284 391592 -19228
rect 391678 -19284 391734 -19228
rect 391536 -19426 391592 -19370
rect 391678 -19426 391734 -19370
rect 391536 -19568 391592 -19512
rect 391678 -19568 391734 -19512
rect 391536 -19710 391592 -19654
rect 391678 -19710 391734 -19654
rect 391536 -19852 391592 -19796
rect 391678 -19852 391734 -19796
rect 391536 -19994 391592 -19938
rect 391678 -19994 391734 -19938
rect 391536 -20136 391592 -20080
rect 391678 -20136 391734 -20080
rect 391536 -20278 391592 -20222
rect 391678 -20278 391734 -20222
rect 391536 -20420 391592 -20364
rect 391678 -20420 391734 -20364
rect 391536 -20562 391592 -20506
rect 391678 -20562 391734 -20506
rect 391536 -20704 391592 -20648
rect 391678 -20704 391734 -20648
rect 391536 -20846 391592 -20790
rect 391678 -20846 391734 -20790
rect 391536 -20988 391592 -20932
rect 391678 -20988 391734 -20932
rect 391536 -21130 391592 -21074
rect 391678 -21130 391734 -21074
rect 391536 -21272 391592 -21216
rect 391678 -21272 391734 -21216
rect 391536 -21414 391592 -21358
rect 391678 -21414 391734 -21358
rect 391536 -21556 391592 -21500
rect 391678 -21556 391734 -21500
rect 391536 -21698 391592 -21642
rect 391678 -21698 391734 -21642
rect 391536 -21840 391592 -21784
rect 391678 -21840 391734 -21784
rect 391536 -21982 391592 -21926
rect 391678 -21982 391734 -21926
rect 391536 -22124 391592 -22068
rect 391678 -22124 391734 -22068
rect 391536 -22266 391592 -22210
rect 391678 -22266 391734 -22210
rect 391536 -22408 391592 -22352
rect 391678 -22408 391734 -22352
rect 391536 -22550 391592 -22494
rect 391678 -22550 391734 -22494
rect 391536 -22692 391592 -22636
rect 391678 -22692 391734 -22636
rect 391536 -22834 391592 -22778
rect 391678 -22834 391734 -22778
rect 391536 -22976 391592 -22920
rect 391678 -22976 391734 -22920
rect 391536 -23118 391592 -23062
rect 391678 -23118 391734 -23062
rect 391536 -23260 391592 -23204
rect 391678 -23260 391734 -23204
rect 391536 -23402 391592 -23346
rect 391678 -23402 391734 -23346
rect 391536 -23544 391592 -23488
rect 391678 -23544 391734 -23488
rect 391536 -23686 391592 -23630
rect 391678 -23686 391734 -23630
rect 391536 -23828 391592 -23772
rect 391678 -23828 391734 -23772
rect 391536 -23970 391592 -23914
rect 391678 -23970 391734 -23914
rect 391536 -24112 391592 -24056
rect 391678 -24112 391734 -24056
rect 391536 -24254 391592 -24198
rect 391678 -24254 391734 -24198
rect 391536 -24396 391592 -24340
rect 391678 -24396 391734 -24340
rect 391536 -24538 391592 -24482
rect 391678 -24538 391734 -24482
rect 391536 -24680 391592 -24624
rect 391678 -24680 391734 -24624
rect 391536 -24822 391592 -24766
rect 391678 -24822 391734 -24766
rect 391536 -24964 391592 -24908
rect 391678 -24964 391734 -24908
rect 391536 -25106 391592 -25050
rect 391678 -25106 391734 -25050
rect 391536 -25248 391592 -25192
rect 391678 -25248 391734 -25192
rect 391536 -25390 391592 -25334
rect 391678 -25390 391734 -25334
rect 391536 -25532 391592 -25476
rect 391678 -25532 391734 -25476
rect 391936 -18006 391992 -17950
rect 392078 -18006 392134 -17950
rect 391936 -18148 391992 -18092
rect 392078 -18148 392134 -18092
rect 391936 -18290 391992 -18234
rect 392078 -18290 392134 -18234
rect 391936 -18432 391992 -18376
rect 392078 -18432 392134 -18376
rect 391936 -18574 391992 -18518
rect 392078 -18574 392134 -18518
rect 391936 -18716 391992 -18660
rect 392078 -18716 392134 -18660
rect 391936 -18858 391992 -18802
rect 392078 -18858 392134 -18802
rect 391936 -19000 391992 -18944
rect 392078 -19000 392134 -18944
rect 391936 -19142 391992 -19086
rect 392078 -19142 392134 -19086
rect 391936 -19284 391992 -19228
rect 392078 -19284 392134 -19228
rect 391936 -19426 391992 -19370
rect 392078 -19426 392134 -19370
rect 391936 -19568 391992 -19512
rect 392078 -19568 392134 -19512
rect 391936 -19710 391992 -19654
rect 392078 -19710 392134 -19654
rect 391936 -19852 391992 -19796
rect 392078 -19852 392134 -19796
rect 391936 -19994 391992 -19938
rect 392078 -19994 392134 -19938
rect 391936 -20136 391992 -20080
rect 392078 -20136 392134 -20080
rect 391936 -20278 391992 -20222
rect 392078 -20278 392134 -20222
rect 391936 -20420 391992 -20364
rect 392078 -20420 392134 -20364
rect 391936 -20562 391992 -20506
rect 392078 -20562 392134 -20506
rect 391936 -20704 391992 -20648
rect 392078 -20704 392134 -20648
rect 391936 -20846 391992 -20790
rect 392078 -20846 392134 -20790
rect 391936 -20988 391992 -20932
rect 392078 -20988 392134 -20932
rect 391936 -21130 391992 -21074
rect 392078 -21130 392134 -21074
rect 391936 -21272 391992 -21216
rect 392078 -21272 392134 -21216
rect 391936 -21414 391992 -21358
rect 392078 -21414 392134 -21358
rect 391936 -21556 391992 -21500
rect 392078 -21556 392134 -21500
rect 391936 -21698 391992 -21642
rect 392078 -21698 392134 -21642
rect 391936 -21840 391992 -21784
rect 392078 -21840 392134 -21784
rect 391936 -21982 391992 -21926
rect 392078 -21982 392134 -21926
rect 391936 -22124 391992 -22068
rect 392078 -22124 392134 -22068
rect 391936 -22266 391992 -22210
rect 392078 -22266 392134 -22210
rect 391936 -22408 391992 -22352
rect 392078 -22408 392134 -22352
rect 391936 -22550 391992 -22494
rect 392078 -22550 392134 -22494
rect 391936 -22692 391992 -22636
rect 392078 -22692 392134 -22636
rect 391936 -22834 391992 -22778
rect 392078 -22834 392134 -22778
rect 391936 -22976 391992 -22920
rect 392078 -22976 392134 -22920
rect 391936 -23118 391992 -23062
rect 392078 -23118 392134 -23062
rect 391936 -23260 391992 -23204
rect 392078 -23260 392134 -23204
rect 391936 -23402 391992 -23346
rect 392078 -23402 392134 -23346
rect 391936 -23544 391992 -23488
rect 392078 -23544 392134 -23488
rect 391936 -23686 391992 -23630
rect 392078 -23686 392134 -23630
rect 391936 -23828 391992 -23772
rect 392078 -23828 392134 -23772
rect 391936 -23970 391992 -23914
rect 392078 -23970 392134 -23914
rect 391936 -24112 391992 -24056
rect 392078 -24112 392134 -24056
rect 391936 -24254 391992 -24198
rect 392078 -24254 392134 -24198
rect 391936 -24396 391992 -24340
rect 392078 -24396 392134 -24340
rect 391936 -24538 391992 -24482
rect 392078 -24538 392134 -24482
rect 391936 -24680 391992 -24624
rect 392078 -24680 392134 -24624
rect 391936 -24822 391992 -24766
rect 392078 -24822 392134 -24766
rect 391936 -24964 391992 -24908
rect 392078 -24964 392134 -24908
rect 391936 -25106 391992 -25050
rect 392078 -25106 392134 -25050
rect 391936 -25248 391992 -25192
rect 392078 -25248 392134 -25192
rect 391936 -25390 391992 -25334
rect 392078 -25390 392134 -25334
rect 391936 -25532 391992 -25476
rect 392078 -25532 392134 -25476
rect 392333 -18006 392389 -17950
rect 392475 -18006 392531 -17950
rect 392333 -18148 392389 -18092
rect 392475 -18148 392531 -18092
rect 392333 -18290 392389 -18234
rect 392475 -18290 392531 -18234
rect 392333 -18432 392389 -18376
rect 392475 -18432 392531 -18376
rect 392333 -18574 392389 -18518
rect 392475 -18574 392531 -18518
rect 392333 -18716 392389 -18660
rect 392475 -18716 392531 -18660
rect 392333 -18858 392389 -18802
rect 392475 -18858 392531 -18802
rect 392333 -19000 392389 -18944
rect 392475 -19000 392531 -18944
rect 392333 -19142 392389 -19086
rect 392475 -19142 392531 -19086
rect 392333 -19284 392389 -19228
rect 392475 -19284 392531 -19228
rect 392333 -19426 392389 -19370
rect 392475 -19426 392531 -19370
rect 392333 -19568 392389 -19512
rect 392475 -19568 392531 -19512
rect 392333 -19710 392389 -19654
rect 392475 -19710 392531 -19654
rect 392333 -19852 392389 -19796
rect 392475 -19852 392531 -19796
rect 392333 -19994 392389 -19938
rect 392475 -19994 392531 -19938
rect 392333 -20136 392389 -20080
rect 392475 -20136 392531 -20080
rect 392333 -20278 392389 -20222
rect 392475 -20278 392531 -20222
rect 392333 -20420 392389 -20364
rect 392475 -20420 392531 -20364
rect 392333 -20562 392389 -20506
rect 392475 -20562 392531 -20506
rect 392333 -20704 392389 -20648
rect 392475 -20704 392531 -20648
rect 392333 -20846 392389 -20790
rect 392475 -20846 392531 -20790
rect 392333 -20988 392389 -20932
rect 392475 -20988 392531 -20932
rect 392333 -21130 392389 -21074
rect 392475 -21130 392531 -21074
rect 392333 -21272 392389 -21216
rect 392475 -21272 392531 -21216
rect 392333 -21414 392389 -21358
rect 392475 -21414 392531 -21358
rect 392333 -21556 392389 -21500
rect 392475 -21556 392531 -21500
rect 392333 -21698 392389 -21642
rect 392475 -21698 392531 -21642
rect 392333 -21840 392389 -21784
rect 392475 -21840 392531 -21784
rect 392333 -21982 392389 -21926
rect 392475 -21982 392531 -21926
rect 392333 -22124 392389 -22068
rect 392475 -22124 392531 -22068
rect 392333 -22266 392389 -22210
rect 392475 -22266 392531 -22210
rect 392333 -22408 392389 -22352
rect 392475 -22408 392531 -22352
rect 392333 -22550 392389 -22494
rect 392475 -22550 392531 -22494
rect 392333 -22692 392389 -22636
rect 392475 -22692 392531 -22636
rect 392333 -22834 392389 -22778
rect 392475 -22834 392531 -22778
rect 392333 -22976 392389 -22920
rect 392475 -22976 392531 -22920
rect 392333 -23118 392389 -23062
rect 392475 -23118 392531 -23062
rect 392333 -23260 392389 -23204
rect 392475 -23260 392531 -23204
rect 392333 -23402 392389 -23346
rect 392475 -23402 392531 -23346
rect 392333 -23544 392389 -23488
rect 392475 -23544 392531 -23488
rect 392333 -23686 392389 -23630
rect 392475 -23686 392531 -23630
rect 392333 -23828 392389 -23772
rect 392475 -23828 392531 -23772
rect 392333 -23970 392389 -23914
rect 392475 -23970 392531 -23914
rect 392333 -24112 392389 -24056
rect 392475 -24112 392531 -24056
rect 392333 -24254 392389 -24198
rect 392475 -24254 392531 -24198
rect 392333 -24396 392389 -24340
rect 392475 -24396 392531 -24340
rect 392333 -24538 392389 -24482
rect 392475 -24538 392531 -24482
rect 392333 -24680 392389 -24624
rect 392475 -24680 392531 -24624
rect 392333 -24822 392389 -24766
rect 392475 -24822 392531 -24766
rect 392333 -24964 392389 -24908
rect 392475 -24964 392531 -24908
rect 392333 -25106 392389 -25050
rect 392475 -25106 392531 -25050
rect 392333 -25248 392389 -25192
rect 392475 -25248 392531 -25192
rect 392333 -25390 392389 -25334
rect 392475 -25390 392531 -25334
rect 392333 -25532 392389 -25476
rect 392475 -25532 392531 -25476
rect 392738 -18006 392794 -17950
rect 392880 -18006 392936 -17950
rect 392738 -18148 392794 -18092
rect 392880 -18148 392936 -18092
rect 392738 -18290 392794 -18234
rect 392880 -18290 392936 -18234
rect 392738 -18432 392794 -18376
rect 392880 -18432 392936 -18376
rect 392738 -18574 392794 -18518
rect 392880 -18574 392936 -18518
rect 392738 -18716 392794 -18660
rect 392880 -18716 392936 -18660
rect 392738 -18858 392794 -18802
rect 392880 -18858 392936 -18802
rect 392738 -19000 392794 -18944
rect 392880 -19000 392936 -18944
rect 392738 -19142 392794 -19086
rect 392880 -19142 392936 -19086
rect 392738 -19284 392794 -19228
rect 392880 -19284 392936 -19228
rect 392738 -19426 392794 -19370
rect 392880 -19426 392936 -19370
rect 392738 -19568 392794 -19512
rect 392880 -19568 392936 -19512
rect 392738 -19710 392794 -19654
rect 392880 -19710 392936 -19654
rect 392738 -19852 392794 -19796
rect 392880 -19852 392936 -19796
rect 392738 -19994 392794 -19938
rect 392880 -19994 392936 -19938
rect 392738 -20136 392794 -20080
rect 392880 -20136 392936 -20080
rect 392738 -20278 392794 -20222
rect 392880 -20278 392936 -20222
rect 392738 -20420 392794 -20364
rect 392880 -20420 392936 -20364
rect 392738 -20562 392794 -20506
rect 392880 -20562 392936 -20506
rect 392738 -20704 392794 -20648
rect 392880 -20704 392936 -20648
rect 392738 -20846 392794 -20790
rect 392880 -20846 392936 -20790
rect 392738 -20988 392794 -20932
rect 392880 -20988 392936 -20932
rect 392738 -21130 392794 -21074
rect 392880 -21130 392936 -21074
rect 392738 -21272 392794 -21216
rect 392880 -21272 392936 -21216
rect 392738 -21414 392794 -21358
rect 392880 -21414 392936 -21358
rect 392738 -21556 392794 -21500
rect 392880 -21556 392936 -21500
rect 392738 -21698 392794 -21642
rect 392880 -21698 392936 -21642
rect 392738 -21840 392794 -21784
rect 392880 -21840 392936 -21784
rect 392738 -21982 392794 -21926
rect 392880 -21982 392936 -21926
rect 392738 -22124 392794 -22068
rect 392880 -22124 392936 -22068
rect 392738 -22266 392794 -22210
rect 392880 -22266 392936 -22210
rect 392738 -22408 392794 -22352
rect 392880 -22408 392936 -22352
rect 392738 -22550 392794 -22494
rect 392880 -22550 392936 -22494
rect 392738 -22692 392794 -22636
rect 392880 -22692 392936 -22636
rect 392738 -22834 392794 -22778
rect 392880 -22834 392936 -22778
rect 392738 -22976 392794 -22920
rect 392880 -22976 392936 -22920
rect 392738 -23118 392794 -23062
rect 392880 -23118 392936 -23062
rect 392738 -23260 392794 -23204
rect 392880 -23260 392936 -23204
rect 392738 -23402 392794 -23346
rect 392880 -23402 392936 -23346
rect 392738 -23544 392794 -23488
rect 392880 -23544 392936 -23488
rect 392738 -23686 392794 -23630
rect 392880 -23686 392936 -23630
rect 392738 -23828 392794 -23772
rect 392880 -23828 392936 -23772
rect 392738 -23970 392794 -23914
rect 392880 -23970 392936 -23914
rect 392738 -24112 392794 -24056
rect 392880 -24112 392936 -24056
rect 392738 -24254 392794 -24198
rect 392880 -24254 392936 -24198
rect 392738 -24396 392794 -24340
rect 392880 -24396 392936 -24340
rect 392738 -24538 392794 -24482
rect 392880 -24538 392936 -24482
rect 392738 -24680 392794 -24624
rect 392880 -24680 392936 -24624
rect 392738 -24822 392794 -24766
rect 392880 -24822 392936 -24766
rect 392738 -24964 392794 -24908
rect 392880 -24964 392936 -24908
rect 392738 -25106 392794 -25050
rect 392880 -25106 392936 -25050
rect 392738 -25248 392794 -25192
rect 392880 -25248 392936 -25192
rect 392738 -25390 392794 -25334
rect 392880 -25390 392936 -25334
rect 392738 -25532 392794 -25476
rect 392880 -25532 392936 -25476
rect 393138 -18006 393194 -17950
rect 393280 -18006 393336 -17950
rect 393138 -18148 393194 -18092
rect 393280 -18148 393336 -18092
rect 393138 -18290 393194 -18234
rect 393280 -18290 393336 -18234
rect 393138 -18432 393194 -18376
rect 393280 -18432 393336 -18376
rect 393138 -18574 393194 -18518
rect 393280 -18574 393336 -18518
rect 393138 -18716 393194 -18660
rect 393280 -18716 393336 -18660
rect 393138 -18858 393194 -18802
rect 393280 -18858 393336 -18802
rect 393138 -19000 393194 -18944
rect 393280 -19000 393336 -18944
rect 393138 -19142 393194 -19086
rect 393280 -19142 393336 -19086
rect 393138 -19284 393194 -19228
rect 393280 -19284 393336 -19228
rect 393138 -19426 393194 -19370
rect 393280 -19426 393336 -19370
rect 393138 -19568 393194 -19512
rect 393280 -19568 393336 -19512
rect 393138 -19710 393194 -19654
rect 393280 -19710 393336 -19654
rect 393138 -19852 393194 -19796
rect 393280 -19852 393336 -19796
rect 393138 -19994 393194 -19938
rect 393280 -19994 393336 -19938
rect 393138 -20136 393194 -20080
rect 393280 -20136 393336 -20080
rect 393138 -20278 393194 -20222
rect 393280 -20278 393336 -20222
rect 393138 -20420 393194 -20364
rect 393280 -20420 393336 -20364
rect 393138 -20562 393194 -20506
rect 393280 -20562 393336 -20506
rect 393138 -20704 393194 -20648
rect 393280 -20704 393336 -20648
rect 393138 -20846 393194 -20790
rect 393280 -20846 393336 -20790
rect 393138 -20988 393194 -20932
rect 393280 -20988 393336 -20932
rect 393138 -21130 393194 -21074
rect 393280 -21130 393336 -21074
rect 393138 -21272 393194 -21216
rect 393280 -21272 393336 -21216
rect 393138 -21414 393194 -21358
rect 393280 -21414 393336 -21358
rect 393138 -21556 393194 -21500
rect 393280 -21556 393336 -21500
rect 393138 -21698 393194 -21642
rect 393280 -21698 393336 -21642
rect 393138 -21840 393194 -21784
rect 393280 -21840 393336 -21784
rect 393138 -21982 393194 -21926
rect 393280 -21982 393336 -21926
rect 393138 -22124 393194 -22068
rect 393280 -22124 393336 -22068
rect 393138 -22266 393194 -22210
rect 393280 -22266 393336 -22210
rect 393138 -22408 393194 -22352
rect 393280 -22408 393336 -22352
rect 393138 -22550 393194 -22494
rect 393280 -22550 393336 -22494
rect 393138 -22692 393194 -22636
rect 393280 -22692 393336 -22636
rect 393138 -22834 393194 -22778
rect 393280 -22834 393336 -22778
rect 393138 -22976 393194 -22920
rect 393280 -22976 393336 -22920
rect 393138 -23118 393194 -23062
rect 393280 -23118 393336 -23062
rect 393138 -23260 393194 -23204
rect 393280 -23260 393336 -23204
rect 393138 -23402 393194 -23346
rect 393280 -23402 393336 -23346
rect 393138 -23544 393194 -23488
rect 393280 -23544 393336 -23488
rect 393138 -23686 393194 -23630
rect 393280 -23686 393336 -23630
rect 393138 -23828 393194 -23772
rect 393280 -23828 393336 -23772
rect 393138 -23970 393194 -23914
rect 393280 -23970 393336 -23914
rect 393138 -24112 393194 -24056
rect 393280 -24112 393336 -24056
rect 393138 -24254 393194 -24198
rect 393280 -24254 393336 -24198
rect 393138 -24396 393194 -24340
rect 393280 -24396 393336 -24340
rect 393138 -24538 393194 -24482
rect 393280 -24538 393336 -24482
rect 393138 -24680 393194 -24624
rect 393280 -24680 393336 -24624
rect 393138 -24822 393194 -24766
rect 393280 -24822 393336 -24766
rect 393138 -24964 393194 -24908
rect 393280 -24964 393336 -24908
rect 393138 -25106 393194 -25050
rect 393280 -25106 393336 -25050
rect 393138 -25248 393194 -25192
rect 393280 -25248 393336 -25192
rect 393138 -25390 393194 -25334
rect 393280 -25390 393336 -25334
rect 393138 -25532 393194 -25476
rect 393280 -25532 393336 -25476
rect 393543 -18006 393599 -17950
rect 393685 -18006 393741 -17950
rect 393543 -18148 393599 -18092
rect 393685 -18148 393741 -18092
rect 393543 -18290 393599 -18234
rect 393685 -18290 393741 -18234
rect 393543 -18432 393599 -18376
rect 393685 -18432 393741 -18376
rect 393543 -18574 393599 -18518
rect 393685 -18574 393741 -18518
rect 393543 -18716 393599 -18660
rect 393685 -18716 393741 -18660
rect 393543 -18858 393599 -18802
rect 393685 -18858 393741 -18802
rect 393543 -19000 393599 -18944
rect 393685 -19000 393741 -18944
rect 393543 -19142 393599 -19086
rect 393685 -19142 393741 -19086
rect 393543 -19284 393599 -19228
rect 393685 -19284 393741 -19228
rect 393543 -19426 393599 -19370
rect 393685 -19426 393741 -19370
rect 393543 -19568 393599 -19512
rect 393685 -19568 393741 -19512
rect 393543 -19710 393599 -19654
rect 393685 -19710 393741 -19654
rect 393543 -19852 393599 -19796
rect 393685 -19852 393741 -19796
rect 393543 -19994 393599 -19938
rect 393685 -19994 393741 -19938
rect 393543 -20136 393599 -20080
rect 393685 -20136 393741 -20080
rect 393543 -20278 393599 -20222
rect 393685 -20278 393741 -20222
rect 393543 -20420 393599 -20364
rect 393685 -20420 393741 -20364
rect 393543 -20562 393599 -20506
rect 393685 -20562 393741 -20506
rect 393543 -20704 393599 -20648
rect 393685 -20704 393741 -20648
rect 393543 -20846 393599 -20790
rect 393685 -20846 393741 -20790
rect 393543 -20988 393599 -20932
rect 393685 -20988 393741 -20932
rect 393543 -21130 393599 -21074
rect 393685 -21130 393741 -21074
rect 393543 -21272 393599 -21216
rect 393685 -21272 393741 -21216
rect 393543 -21414 393599 -21358
rect 393685 -21414 393741 -21358
rect 393543 -21556 393599 -21500
rect 393685 -21556 393741 -21500
rect 393543 -21698 393599 -21642
rect 393685 -21698 393741 -21642
rect 393543 -21840 393599 -21784
rect 393685 -21840 393741 -21784
rect 393543 -21982 393599 -21926
rect 393685 -21982 393741 -21926
rect 393543 -22124 393599 -22068
rect 393685 -22124 393741 -22068
rect 393543 -22266 393599 -22210
rect 393685 -22266 393741 -22210
rect 393543 -22408 393599 -22352
rect 393685 -22408 393741 -22352
rect 393543 -22550 393599 -22494
rect 393685 -22550 393741 -22494
rect 393543 -22692 393599 -22636
rect 393685 -22692 393741 -22636
rect 393543 -22834 393599 -22778
rect 393685 -22834 393741 -22778
rect 393543 -22976 393599 -22920
rect 393685 -22976 393741 -22920
rect 393543 -23118 393599 -23062
rect 393685 -23118 393741 -23062
rect 393543 -23260 393599 -23204
rect 393685 -23260 393741 -23204
rect 393543 -23402 393599 -23346
rect 393685 -23402 393741 -23346
rect 393543 -23544 393599 -23488
rect 393685 -23544 393741 -23488
rect 393543 -23686 393599 -23630
rect 393685 -23686 393741 -23630
rect 393543 -23828 393599 -23772
rect 393685 -23828 393741 -23772
rect 393543 -23970 393599 -23914
rect 393685 -23970 393741 -23914
rect 393543 -24112 393599 -24056
rect 393685 -24112 393741 -24056
rect 393543 -24254 393599 -24198
rect 393685 -24254 393741 -24198
rect 393543 -24396 393599 -24340
rect 393685 -24396 393741 -24340
rect 393543 -24538 393599 -24482
rect 393685 -24538 393741 -24482
rect 393543 -24680 393599 -24624
rect 393685 -24680 393741 -24624
rect 393543 -24822 393599 -24766
rect 393685 -24822 393741 -24766
rect 393543 -24964 393599 -24908
rect 393685 -24964 393741 -24908
rect 393543 -25106 393599 -25050
rect 393685 -25106 393741 -25050
rect 393543 -25248 393599 -25192
rect 393685 -25248 393741 -25192
rect 393543 -25390 393599 -25334
rect 393685 -25390 393741 -25334
rect 393543 -25532 393599 -25476
rect 393685 -25532 393741 -25476
rect 393940 -18006 393996 -17950
rect 394082 -18006 394138 -17950
rect 393940 -18148 393996 -18092
rect 394082 -18148 394138 -18092
rect 393940 -18290 393996 -18234
rect 394082 -18290 394138 -18234
rect 393940 -18432 393996 -18376
rect 394082 -18432 394138 -18376
rect 393940 -18574 393996 -18518
rect 394082 -18574 394138 -18518
rect 393940 -18716 393996 -18660
rect 394082 -18716 394138 -18660
rect 393940 -18858 393996 -18802
rect 394082 -18858 394138 -18802
rect 393940 -19000 393996 -18944
rect 394082 -19000 394138 -18944
rect 393940 -19142 393996 -19086
rect 394082 -19142 394138 -19086
rect 393940 -19284 393996 -19228
rect 394082 -19284 394138 -19228
rect 393940 -19426 393996 -19370
rect 394082 -19426 394138 -19370
rect 393940 -19568 393996 -19512
rect 394082 -19568 394138 -19512
rect 393940 -19710 393996 -19654
rect 394082 -19710 394138 -19654
rect 393940 -19852 393996 -19796
rect 394082 -19852 394138 -19796
rect 393940 -19994 393996 -19938
rect 394082 -19994 394138 -19938
rect 393940 -20136 393996 -20080
rect 394082 -20136 394138 -20080
rect 393940 -20278 393996 -20222
rect 394082 -20278 394138 -20222
rect 393940 -20420 393996 -20364
rect 394082 -20420 394138 -20364
rect 393940 -20562 393996 -20506
rect 394082 -20562 394138 -20506
rect 393940 -20704 393996 -20648
rect 394082 -20704 394138 -20648
rect 393940 -20846 393996 -20790
rect 394082 -20846 394138 -20790
rect 393940 -20988 393996 -20932
rect 394082 -20988 394138 -20932
rect 393940 -21130 393996 -21074
rect 394082 -21130 394138 -21074
rect 393940 -21272 393996 -21216
rect 394082 -21272 394138 -21216
rect 393940 -21414 393996 -21358
rect 394082 -21414 394138 -21358
rect 393940 -21556 393996 -21500
rect 394082 -21556 394138 -21500
rect 393940 -21698 393996 -21642
rect 394082 -21698 394138 -21642
rect 393940 -21840 393996 -21784
rect 394082 -21840 394138 -21784
rect 393940 -21982 393996 -21926
rect 394082 -21982 394138 -21926
rect 393940 -22124 393996 -22068
rect 394082 -22124 394138 -22068
rect 393940 -22266 393996 -22210
rect 394082 -22266 394138 -22210
rect 393940 -22408 393996 -22352
rect 394082 -22408 394138 -22352
rect 393940 -22550 393996 -22494
rect 394082 -22550 394138 -22494
rect 393940 -22692 393996 -22636
rect 394082 -22692 394138 -22636
rect 393940 -22834 393996 -22778
rect 394082 -22834 394138 -22778
rect 393940 -22976 393996 -22920
rect 394082 -22976 394138 -22920
rect 393940 -23118 393996 -23062
rect 394082 -23118 394138 -23062
rect 393940 -23260 393996 -23204
rect 394082 -23260 394138 -23204
rect 393940 -23402 393996 -23346
rect 394082 -23402 394138 -23346
rect 393940 -23544 393996 -23488
rect 394082 -23544 394138 -23488
rect 393940 -23686 393996 -23630
rect 394082 -23686 394138 -23630
rect 393940 -23828 393996 -23772
rect 394082 -23828 394138 -23772
rect 393940 -23970 393996 -23914
rect 394082 -23970 394138 -23914
rect 393940 -24112 393996 -24056
rect 394082 -24112 394138 -24056
rect 393940 -24254 393996 -24198
rect 394082 -24254 394138 -24198
rect 393940 -24396 393996 -24340
rect 394082 -24396 394138 -24340
rect 393940 -24538 393996 -24482
rect 394082 -24538 394138 -24482
rect 393940 -24680 393996 -24624
rect 394082 -24680 394138 -24624
rect 393940 -24822 393996 -24766
rect 394082 -24822 394138 -24766
rect 393940 -24964 393996 -24908
rect 394082 -24964 394138 -24908
rect 393940 -25106 393996 -25050
rect 394082 -25106 394138 -25050
rect 393940 -25248 393996 -25192
rect 394082 -25248 394138 -25192
rect 393940 -25390 393996 -25334
rect 394082 -25390 394138 -25334
rect 393940 -25532 393996 -25476
rect 394082 -25532 394138 -25476
rect 394337 -18006 394393 -17950
rect 394479 -18006 394535 -17950
rect 394337 -18148 394393 -18092
rect 394479 -18148 394535 -18092
rect 394337 -18290 394393 -18234
rect 394479 -18290 394535 -18234
rect 394337 -18432 394393 -18376
rect 394479 -18432 394535 -18376
rect 394337 -18574 394393 -18518
rect 394479 -18574 394535 -18518
rect 394337 -18716 394393 -18660
rect 394479 -18716 394535 -18660
rect 394337 -18858 394393 -18802
rect 394479 -18858 394535 -18802
rect 394337 -19000 394393 -18944
rect 394479 -19000 394535 -18944
rect 394337 -19142 394393 -19086
rect 394479 -19142 394535 -19086
rect 394337 -19284 394393 -19228
rect 394479 -19284 394535 -19228
rect 394337 -19426 394393 -19370
rect 394479 -19426 394535 -19370
rect 394337 -19568 394393 -19512
rect 394479 -19568 394535 -19512
rect 394337 -19710 394393 -19654
rect 394479 -19710 394535 -19654
rect 394337 -19852 394393 -19796
rect 394479 -19852 394535 -19796
rect 394337 -19994 394393 -19938
rect 394479 -19994 394535 -19938
rect 394337 -20136 394393 -20080
rect 394479 -20136 394535 -20080
rect 394337 -20278 394393 -20222
rect 394479 -20278 394535 -20222
rect 394337 -20420 394393 -20364
rect 394479 -20420 394535 -20364
rect 394337 -20562 394393 -20506
rect 394479 -20562 394535 -20506
rect 394337 -20704 394393 -20648
rect 394479 -20704 394535 -20648
rect 394337 -20846 394393 -20790
rect 394479 -20846 394535 -20790
rect 394337 -20988 394393 -20932
rect 394479 -20988 394535 -20932
rect 394337 -21130 394393 -21074
rect 394479 -21130 394535 -21074
rect 394337 -21272 394393 -21216
rect 394479 -21272 394535 -21216
rect 394337 -21414 394393 -21358
rect 394479 -21414 394535 -21358
rect 394337 -21556 394393 -21500
rect 394479 -21556 394535 -21500
rect 394337 -21698 394393 -21642
rect 394479 -21698 394535 -21642
rect 394337 -21840 394393 -21784
rect 394479 -21840 394535 -21784
rect 394337 -21982 394393 -21926
rect 394479 -21982 394535 -21926
rect 394337 -22124 394393 -22068
rect 394479 -22124 394535 -22068
rect 394337 -22266 394393 -22210
rect 394479 -22266 394535 -22210
rect 394337 -22408 394393 -22352
rect 394479 -22408 394535 -22352
rect 394337 -22550 394393 -22494
rect 394479 -22550 394535 -22494
rect 394337 -22692 394393 -22636
rect 394479 -22692 394535 -22636
rect 394337 -22834 394393 -22778
rect 394479 -22834 394535 -22778
rect 394337 -22976 394393 -22920
rect 394479 -22976 394535 -22920
rect 394337 -23118 394393 -23062
rect 394479 -23118 394535 -23062
rect 394337 -23260 394393 -23204
rect 394479 -23260 394535 -23204
rect 394337 -23402 394393 -23346
rect 394479 -23402 394535 -23346
rect 394337 -23544 394393 -23488
rect 394479 -23544 394535 -23488
rect 394337 -23686 394393 -23630
rect 394479 -23686 394535 -23630
rect 394337 -23828 394393 -23772
rect 394479 -23828 394535 -23772
rect 394337 -23970 394393 -23914
rect 394479 -23970 394535 -23914
rect 394337 -24112 394393 -24056
rect 394479 -24112 394535 -24056
rect 394337 -24254 394393 -24198
rect 394479 -24254 394535 -24198
rect 394337 -24396 394393 -24340
rect 394479 -24396 394535 -24340
rect 394337 -24538 394393 -24482
rect 394479 -24538 394535 -24482
rect 394337 -24680 394393 -24624
rect 394479 -24680 394535 -24624
rect 394337 -24822 394393 -24766
rect 394479 -24822 394535 -24766
rect 394337 -24964 394393 -24908
rect 394479 -24964 394535 -24908
rect 394337 -25106 394393 -25050
rect 394479 -25106 394535 -25050
rect 394337 -25248 394393 -25192
rect 394479 -25248 394535 -25192
rect 394337 -25390 394393 -25334
rect 394479 -25390 394535 -25334
rect 394337 -25532 394393 -25476
rect 394479 -25532 394535 -25476
rect 394740 -18006 394796 -17950
rect 394882 -18006 394938 -17950
rect 394740 -18148 394796 -18092
rect 394882 -18148 394938 -18092
rect 394740 -18290 394796 -18234
rect 394882 -18290 394938 -18234
rect 394740 -18432 394796 -18376
rect 394882 -18432 394938 -18376
rect 394740 -18574 394796 -18518
rect 394882 -18574 394938 -18518
rect 394740 -18716 394796 -18660
rect 394882 -18716 394938 -18660
rect 394740 -18858 394796 -18802
rect 394882 -18858 394938 -18802
rect 394740 -19000 394796 -18944
rect 394882 -19000 394938 -18944
rect 394740 -19142 394796 -19086
rect 394882 -19142 394938 -19086
rect 394740 -19284 394796 -19228
rect 394882 -19284 394938 -19228
rect 394740 -19426 394796 -19370
rect 394882 -19426 394938 -19370
rect 394740 -19568 394796 -19512
rect 394882 -19568 394938 -19512
rect 394740 -19710 394796 -19654
rect 394882 -19710 394938 -19654
rect 394740 -19852 394796 -19796
rect 394882 -19852 394938 -19796
rect 394740 -19994 394796 -19938
rect 394882 -19994 394938 -19938
rect 394740 -20136 394796 -20080
rect 394882 -20136 394938 -20080
rect 394740 -20278 394796 -20222
rect 394882 -20278 394938 -20222
rect 394740 -20420 394796 -20364
rect 394882 -20420 394938 -20364
rect 394740 -20562 394796 -20506
rect 394882 -20562 394938 -20506
rect 394740 -20704 394796 -20648
rect 394882 -20704 394938 -20648
rect 394740 -20846 394796 -20790
rect 394882 -20846 394938 -20790
rect 394740 -20988 394796 -20932
rect 394882 -20988 394938 -20932
rect 394740 -21130 394796 -21074
rect 394882 -21130 394938 -21074
rect 394740 -21272 394796 -21216
rect 394882 -21272 394938 -21216
rect 394740 -21414 394796 -21358
rect 394882 -21414 394938 -21358
rect 394740 -21556 394796 -21500
rect 394882 -21556 394938 -21500
rect 394740 -21698 394796 -21642
rect 394882 -21698 394938 -21642
rect 394740 -21840 394796 -21784
rect 394882 -21840 394938 -21784
rect 394740 -21982 394796 -21926
rect 394882 -21982 394938 -21926
rect 394740 -22124 394796 -22068
rect 394882 -22124 394938 -22068
rect 394740 -22266 394796 -22210
rect 394882 -22266 394938 -22210
rect 394740 -22408 394796 -22352
rect 394882 -22408 394938 -22352
rect 394740 -22550 394796 -22494
rect 394882 -22550 394938 -22494
rect 394740 -22692 394796 -22636
rect 394882 -22692 394938 -22636
rect 394740 -22834 394796 -22778
rect 394882 -22834 394938 -22778
rect 394740 -22976 394796 -22920
rect 394882 -22976 394938 -22920
rect 394740 -23118 394796 -23062
rect 394882 -23118 394938 -23062
rect 394740 -23260 394796 -23204
rect 394882 -23260 394938 -23204
rect 394740 -23402 394796 -23346
rect 394882 -23402 394938 -23346
rect 394740 -23544 394796 -23488
rect 394882 -23544 394938 -23488
rect 394740 -23686 394796 -23630
rect 394882 -23686 394938 -23630
rect 394740 -23828 394796 -23772
rect 394882 -23828 394938 -23772
rect 394740 -23970 394796 -23914
rect 394882 -23970 394938 -23914
rect 394740 -24112 394796 -24056
rect 394882 -24112 394938 -24056
rect 394740 -24254 394796 -24198
rect 394882 -24254 394938 -24198
rect 394740 -24396 394796 -24340
rect 394882 -24396 394938 -24340
rect 394740 -24538 394796 -24482
rect 394882 -24538 394938 -24482
rect 394740 -24680 394796 -24624
rect 394882 -24680 394938 -24624
rect 394740 -24822 394796 -24766
rect 394882 -24822 394938 -24766
rect 394740 -24964 394796 -24908
rect 394882 -24964 394938 -24908
rect 394740 -25106 394796 -25050
rect 394882 -25106 394938 -25050
rect 394740 -25248 394796 -25192
rect 394882 -25248 394938 -25192
rect 394740 -25390 394796 -25334
rect 394882 -25390 394938 -25334
rect 394740 -25532 394796 -25476
rect 394882 -25532 394938 -25476
rect 395142 -18006 395198 -17950
rect 395284 -18006 395340 -17950
rect 395142 -18148 395198 -18092
rect 395284 -18148 395340 -18092
rect 395142 -18290 395198 -18234
rect 395284 -18290 395340 -18234
rect 395142 -18432 395198 -18376
rect 395284 -18432 395340 -18376
rect 395142 -18574 395198 -18518
rect 395284 -18574 395340 -18518
rect 395142 -18716 395198 -18660
rect 395284 -18716 395340 -18660
rect 395142 -18858 395198 -18802
rect 395284 -18858 395340 -18802
rect 395142 -19000 395198 -18944
rect 395284 -19000 395340 -18944
rect 395142 -19142 395198 -19086
rect 395284 -19142 395340 -19086
rect 395142 -19284 395198 -19228
rect 395284 -19284 395340 -19228
rect 395142 -19426 395198 -19370
rect 395284 -19426 395340 -19370
rect 395142 -19568 395198 -19512
rect 395284 -19568 395340 -19512
rect 395142 -19710 395198 -19654
rect 395284 -19710 395340 -19654
rect 395142 -19852 395198 -19796
rect 395284 -19852 395340 -19796
rect 395142 -19994 395198 -19938
rect 395284 -19994 395340 -19938
rect 395142 -20136 395198 -20080
rect 395284 -20136 395340 -20080
rect 395142 -20278 395198 -20222
rect 395284 -20278 395340 -20222
rect 395142 -20420 395198 -20364
rect 395284 -20420 395340 -20364
rect 395142 -20562 395198 -20506
rect 395284 -20562 395340 -20506
rect 395142 -20704 395198 -20648
rect 395284 -20704 395340 -20648
rect 395142 -20846 395198 -20790
rect 395284 -20846 395340 -20790
rect 395142 -20988 395198 -20932
rect 395284 -20988 395340 -20932
rect 395142 -21130 395198 -21074
rect 395284 -21130 395340 -21074
rect 395142 -21272 395198 -21216
rect 395284 -21272 395340 -21216
rect 395142 -21414 395198 -21358
rect 395284 -21414 395340 -21358
rect 395142 -21556 395198 -21500
rect 395284 -21556 395340 -21500
rect 395142 -21698 395198 -21642
rect 395284 -21698 395340 -21642
rect 395142 -21840 395198 -21784
rect 395284 -21840 395340 -21784
rect 395142 -21982 395198 -21926
rect 395284 -21982 395340 -21926
rect 395142 -22124 395198 -22068
rect 395284 -22124 395340 -22068
rect 395142 -22266 395198 -22210
rect 395284 -22266 395340 -22210
rect 395142 -22408 395198 -22352
rect 395284 -22408 395340 -22352
rect 395142 -22550 395198 -22494
rect 395284 -22550 395340 -22494
rect 395142 -22692 395198 -22636
rect 395284 -22692 395340 -22636
rect 395142 -22834 395198 -22778
rect 395284 -22834 395340 -22778
rect 395142 -22976 395198 -22920
rect 395284 -22976 395340 -22920
rect 395142 -23118 395198 -23062
rect 395284 -23118 395340 -23062
rect 395142 -23260 395198 -23204
rect 395284 -23260 395340 -23204
rect 395142 -23402 395198 -23346
rect 395284 -23402 395340 -23346
rect 395142 -23544 395198 -23488
rect 395284 -23544 395340 -23488
rect 395142 -23686 395198 -23630
rect 395284 -23686 395340 -23630
rect 395142 -23828 395198 -23772
rect 395284 -23828 395340 -23772
rect 395142 -23970 395198 -23914
rect 395284 -23970 395340 -23914
rect 395142 -24112 395198 -24056
rect 395284 -24112 395340 -24056
rect 395142 -24254 395198 -24198
rect 395284 -24254 395340 -24198
rect 395142 -24396 395198 -24340
rect 395284 -24396 395340 -24340
rect 395142 -24538 395198 -24482
rect 395284 -24538 395340 -24482
rect 395142 -24680 395198 -24624
rect 395284 -24680 395340 -24624
rect 395142 -24822 395198 -24766
rect 395284 -24822 395340 -24766
rect 395142 -24964 395198 -24908
rect 395284 -24964 395340 -24908
rect 395142 -25106 395198 -25050
rect 395284 -25106 395340 -25050
rect 395142 -25248 395198 -25192
rect 395284 -25248 395340 -25192
rect 395142 -25390 395198 -25334
rect 395284 -25390 395340 -25334
rect 395142 -25532 395198 -25476
rect 395284 -25532 395340 -25476
rect 395545 -18006 395601 -17950
rect 395687 -18006 395743 -17950
rect 395545 -18148 395601 -18092
rect 395687 -18148 395743 -18092
rect 395545 -18290 395601 -18234
rect 395687 -18290 395743 -18234
rect 395545 -18432 395601 -18376
rect 395687 -18432 395743 -18376
rect 395545 -18574 395601 -18518
rect 395687 -18574 395743 -18518
rect 395545 -18716 395601 -18660
rect 395687 -18716 395743 -18660
rect 395545 -18858 395601 -18802
rect 395687 -18858 395743 -18802
rect 395545 -19000 395601 -18944
rect 395687 -19000 395743 -18944
rect 395545 -19142 395601 -19086
rect 395687 -19142 395743 -19086
rect 395545 -19284 395601 -19228
rect 395687 -19284 395743 -19228
rect 395545 -19426 395601 -19370
rect 395687 -19426 395743 -19370
rect 395545 -19568 395601 -19512
rect 395687 -19568 395743 -19512
rect 395545 -19710 395601 -19654
rect 395687 -19710 395743 -19654
rect 395545 -19852 395601 -19796
rect 395687 -19852 395743 -19796
rect 395545 -19994 395601 -19938
rect 395687 -19994 395743 -19938
rect 395545 -20136 395601 -20080
rect 395687 -20136 395743 -20080
rect 395545 -20278 395601 -20222
rect 395687 -20278 395743 -20222
rect 395545 -20420 395601 -20364
rect 395687 -20420 395743 -20364
rect 395545 -20562 395601 -20506
rect 395687 -20562 395743 -20506
rect 395545 -20704 395601 -20648
rect 395687 -20704 395743 -20648
rect 395545 -20846 395601 -20790
rect 395687 -20846 395743 -20790
rect 395545 -20988 395601 -20932
rect 395687 -20988 395743 -20932
rect 395545 -21130 395601 -21074
rect 395687 -21130 395743 -21074
rect 395545 -21272 395601 -21216
rect 395687 -21272 395743 -21216
rect 395545 -21414 395601 -21358
rect 395687 -21414 395743 -21358
rect 395545 -21556 395601 -21500
rect 395687 -21556 395743 -21500
rect 395545 -21698 395601 -21642
rect 395687 -21698 395743 -21642
rect 395545 -21840 395601 -21784
rect 395687 -21840 395743 -21784
rect 395545 -21982 395601 -21926
rect 395687 -21982 395743 -21926
rect 395545 -22124 395601 -22068
rect 395687 -22124 395743 -22068
rect 395545 -22266 395601 -22210
rect 395687 -22266 395743 -22210
rect 395545 -22408 395601 -22352
rect 395687 -22408 395743 -22352
rect 395545 -22550 395601 -22494
rect 395687 -22550 395743 -22494
rect 395545 -22692 395601 -22636
rect 395687 -22692 395743 -22636
rect 395545 -22834 395601 -22778
rect 395687 -22834 395743 -22778
rect 395545 -22976 395601 -22920
rect 395687 -22976 395743 -22920
rect 395545 -23118 395601 -23062
rect 395687 -23118 395743 -23062
rect 395545 -23260 395601 -23204
rect 395687 -23260 395743 -23204
rect 395545 -23402 395601 -23346
rect 395687 -23402 395743 -23346
rect 395545 -23544 395601 -23488
rect 395687 -23544 395743 -23488
rect 395545 -23686 395601 -23630
rect 395687 -23686 395743 -23630
rect 395545 -23828 395601 -23772
rect 395687 -23828 395743 -23772
rect 395545 -23970 395601 -23914
rect 395687 -23970 395743 -23914
rect 395545 -24112 395601 -24056
rect 395687 -24112 395743 -24056
rect 395545 -24254 395601 -24198
rect 395687 -24254 395743 -24198
rect 395545 -24396 395601 -24340
rect 395687 -24396 395743 -24340
rect 395545 -24538 395601 -24482
rect 395687 -24538 395743 -24482
rect 395545 -24680 395601 -24624
rect 395687 -24680 395743 -24624
rect 395545 -24822 395601 -24766
rect 395687 -24822 395743 -24766
rect 395545 -24964 395601 -24908
rect 395687 -24964 395743 -24908
rect 395545 -25106 395601 -25050
rect 395687 -25106 395743 -25050
rect 395545 -25248 395601 -25192
rect 395687 -25248 395743 -25192
rect 395545 -25390 395601 -25334
rect 395687 -25390 395743 -25334
rect 395545 -25532 395601 -25476
rect 395687 -25532 395743 -25476
rect 395941 -18006 395997 -17950
rect 396083 -18006 396139 -17950
rect 395941 -18148 395997 -18092
rect 396083 -18148 396139 -18092
rect 395941 -18290 395997 -18234
rect 396083 -18290 396139 -18234
rect 395941 -18432 395997 -18376
rect 396083 -18432 396139 -18376
rect 395941 -18574 395997 -18518
rect 396083 -18574 396139 -18518
rect 395941 -18716 395997 -18660
rect 396083 -18716 396139 -18660
rect 395941 -18858 395997 -18802
rect 396083 -18858 396139 -18802
rect 395941 -19000 395997 -18944
rect 396083 -19000 396139 -18944
rect 395941 -19142 395997 -19086
rect 396083 -19142 396139 -19086
rect 395941 -19284 395997 -19228
rect 396083 -19284 396139 -19228
rect 395941 -19426 395997 -19370
rect 396083 -19426 396139 -19370
rect 395941 -19568 395997 -19512
rect 396083 -19568 396139 -19512
rect 395941 -19710 395997 -19654
rect 396083 -19710 396139 -19654
rect 395941 -19852 395997 -19796
rect 396083 -19852 396139 -19796
rect 395941 -19994 395997 -19938
rect 396083 -19994 396139 -19938
rect 395941 -20136 395997 -20080
rect 396083 -20136 396139 -20080
rect 395941 -20278 395997 -20222
rect 396083 -20278 396139 -20222
rect 395941 -20420 395997 -20364
rect 396083 -20420 396139 -20364
rect 395941 -20562 395997 -20506
rect 396083 -20562 396139 -20506
rect 395941 -20704 395997 -20648
rect 396083 -20704 396139 -20648
rect 395941 -20846 395997 -20790
rect 396083 -20846 396139 -20790
rect 395941 -20988 395997 -20932
rect 396083 -20988 396139 -20932
rect 395941 -21130 395997 -21074
rect 396083 -21130 396139 -21074
rect 395941 -21272 395997 -21216
rect 396083 -21272 396139 -21216
rect 395941 -21414 395997 -21358
rect 396083 -21414 396139 -21358
rect 395941 -21556 395997 -21500
rect 396083 -21556 396139 -21500
rect 395941 -21698 395997 -21642
rect 396083 -21698 396139 -21642
rect 395941 -21840 395997 -21784
rect 396083 -21840 396139 -21784
rect 395941 -21982 395997 -21926
rect 396083 -21982 396139 -21926
rect 395941 -22124 395997 -22068
rect 396083 -22124 396139 -22068
rect 395941 -22266 395997 -22210
rect 396083 -22266 396139 -22210
rect 395941 -22408 395997 -22352
rect 396083 -22408 396139 -22352
rect 395941 -22550 395997 -22494
rect 396083 -22550 396139 -22494
rect 395941 -22692 395997 -22636
rect 396083 -22692 396139 -22636
rect 395941 -22834 395997 -22778
rect 396083 -22834 396139 -22778
rect 395941 -22976 395997 -22920
rect 396083 -22976 396139 -22920
rect 395941 -23118 395997 -23062
rect 396083 -23118 396139 -23062
rect 395941 -23260 395997 -23204
rect 396083 -23260 396139 -23204
rect 395941 -23402 395997 -23346
rect 396083 -23402 396139 -23346
rect 395941 -23544 395997 -23488
rect 396083 -23544 396139 -23488
rect 395941 -23686 395997 -23630
rect 396083 -23686 396139 -23630
rect 395941 -23828 395997 -23772
rect 396083 -23828 396139 -23772
rect 395941 -23970 395997 -23914
rect 396083 -23970 396139 -23914
rect 395941 -24112 395997 -24056
rect 396083 -24112 396139 -24056
rect 395941 -24254 395997 -24198
rect 396083 -24254 396139 -24198
rect 395941 -24396 395997 -24340
rect 396083 -24396 396139 -24340
rect 395941 -24538 395997 -24482
rect 396083 -24538 396139 -24482
rect 395941 -24680 395997 -24624
rect 396083 -24680 396139 -24624
rect 395941 -24822 395997 -24766
rect 396083 -24822 396139 -24766
rect 395941 -24964 395997 -24908
rect 396083 -24964 396139 -24908
rect 395941 -25106 395997 -25050
rect 396083 -25106 396139 -25050
rect 395941 -25248 395997 -25192
rect 396083 -25248 396139 -25192
rect 395941 -25390 395997 -25334
rect 396083 -25390 396139 -25334
rect 395941 -25532 395997 -25476
rect 396083 -25532 396139 -25476
rect 396526 -17914 396582 -17858
rect 396650 -17914 396706 -17858
rect 396774 -17914 396830 -17858
rect 396898 -17914 396954 -17858
rect 397022 -17914 397078 -17858
rect 396526 -18038 396582 -17982
rect 396650 -18038 396706 -17982
rect 396774 -18038 396830 -17982
rect 396898 -18038 396954 -17982
rect 397022 -18038 397078 -17982
rect 396526 -18162 396582 -18106
rect 396650 -18162 396706 -18106
rect 396774 -18162 396830 -18106
rect 396898 -18162 396954 -18106
rect 397022 -18162 397078 -18106
rect 396526 -18286 396582 -18230
rect 396650 -18286 396706 -18230
rect 396774 -18286 396830 -18230
rect 396898 -18286 396954 -18230
rect 397022 -18286 397078 -18230
rect 396526 -18410 396582 -18354
rect 396650 -18410 396706 -18354
rect 396774 -18410 396830 -18354
rect 396898 -18410 396954 -18354
rect 397022 -18410 397078 -18354
rect 396526 -18534 396582 -18478
rect 396650 -18534 396706 -18478
rect 396774 -18534 396830 -18478
rect 396898 -18534 396954 -18478
rect 397022 -18534 397078 -18478
rect 396526 -18658 396582 -18602
rect 396650 -18658 396706 -18602
rect 396774 -18658 396830 -18602
rect 396898 -18658 396954 -18602
rect 397022 -18658 397078 -18602
rect 396526 -18782 396582 -18726
rect 396650 -18782 396706 -18726
rect 396774 -18782 396830 -18726
rect 396898 -18782 396954 -18726
rect 397022 -18782 397078 -18726
rect 396526 -18906 396582 -18850
rect 396650 -18906 396706 -18850
rect 396774 -18906 396830 -18850
rect 396898 -18906 396954 -18850
rect 397022 -18906 397078 -18850
rect 396526 -19030 396582 -18974
rect 396650 -19030 396706 -18974
rect 396774 -19030 396830 -18974
rect 396898 -19030 396954 -18974
rect 397022 -19030 397078 -18974
rect 396526 -19154 396582 -19098
rect 396650 -19154 396706 -19098
rect 396774 -19154 396830 -19098
rect 396898 -19154 396954 -19098
rect 397022 -19154 397078 -19098
rect 396526 -19278 396582 -19222
rect 396650 -19278 396706 -19222
rect 396774 -19278 396830 -19222
rect 396898 -19278 396954 -19222
rect 397022 -19278 397078 -19222
rect 396526 -19402 396582 -19346
rect 396650 -19402 396706 -19346
rect 396774 -19402 396830 -19346
rect 396898 -19402 396954 -19346
rect 397022 -19402 397078 -19346
rect 396526 -19526 396582 -19470
rect 396650 -19526 396706 -19470
rect 396774 -19526 396830 -19470
rect 396898 -19526 396954 -19470
rect 397022 -19526 397078 -19470
rect 396526 -19650 396582 -19594
rect 396650 -19650 396706 -19594
rect 396774 -19650 396830 -19594
rect 396898 -19650 396954 -19594
rect 397022 -19650 397078 -19594
rect 396526 -19774 396582 -19718
rect 396650 -19774 396706 -19718
rect 396774 -19774 396830 -19718
rect 396898 -19774 396954 -19718
rect 397022 -19774 397078 -19718
rect 396526 -19898 396582 -19842
rect 396650 -19898 396706 -19842
rect 396774 -19898 396830 -19842
rect 396898 -19898 396954 -19842
rect 397022 -19898 397078 -19842
rect 396526 -20022 396582 -19966
rect 396650 -20022 396706 -19966
rect 396774 -20022 396830 -19966
rect 396898 -20022 396954 -19966
rect 397022 -20022 397078 -19966
rect 396526 -20146 396582 -20090
rect 396650 -20146 396706 -20090
rect 396774 -20146 396830 -20090
rect 396898 -20146 396954 -20090
rect 397022 -20146 397078 -20090
rect 396526 -20270 396582 -20214
rect 396650 -20270 396706 -20214
rect 396774 -20270 396830 -20214
rect 396898 -20270 396954 -20214
rect 397022 -20270 397078 -20214
rect 396526 -20394 396582 -20338
rect 396650 -20394 396706 -20338
rect 396774 -20394 396830 -20338
rect 396898 -20394 396954 -20338
rect 397022 -20394 397078 -20338
rect 396526 -20518 396582 -20462
rect 396650 -20518 396706 -20462
rect 396774 -20518 396830 -20462
rect 396898 -20518 396954 -20462
rect 397022 -20518 397078 -20462
rect 396526 -20642 396582 -20586
rect 396650 -20642 396706 -20586
rect 396774 -20642 396830 -20586
rect 396898 -20642 396954 -20586
rect 397022 -20642 397078 -20586
rect 396526 -20766 396582 -20710
rect 396650 -20766 396706 -20710
rect 396774 -20766 396830 -20710
rect 396898 -20766 396954 -20710
rect 397022 -20766 397078 -20710
rect 396526 -20890 396582 -20834
rect 396650 -20890 396706 -20834
rect 396774 -20890 396830 -20834
rect 396898 -20890 396954 -20834
rect 397022 -20890 397078 -20834
rect 396526 -21014 396582 -20958
rect 396650 -21014 396706 -20958
rect 396774 -21014 396830 -20958
rect 396898 -21014 396954 -20958
rect 397022 -21014 397078 -20958
rect 396526 -21138 396582 -21082
rect 396650 -21138 396706 -21082
rect 396774 -21138 396830 -21082
rect 396898 -21138 396954 -21082
rect 397022 -21138 397078 -21082
rect 396526 -21262 396582 -21206
rect 396650 -21262 396706 -21206
rect 396774 -21262 396830 -21206
rect 396898 -21262 396954 -21206
rect 397022 -21262 397078 -21206
rect 396526 -21386 396582 -21330
rect 396650 -21386 396706 -21330
rect 396774 -21386 396830 -21330
rect 396898 -21386 396954 -21330
rect 397022 -21386 397078 -21330
rect 396526 -21510 396582 -21454
rect 396650 -21510 396706 -21454
rect 396774 -21510 396830 -21454
rect 396898 -21510 396954 -21454
rect 397022 -21510 397078 -21454
rect 396526 -21634 396582 -21578
rect 396650 -21634 396706 -21578
rect 396774 -21634 396830 -21578
rect 396898 -21634 396954 -21578
rect 397022 -21634 397078 -21578
rect 396526 -21758 396582 -21702
rect 396650 -21758 396706 -21702
rect 396774 -21758 396830 -21702
rect 396898 -21758 396954 -21702
rect 397022 -21758 397078 -21702
rect 396526 -21882 396582 -21826
rect 396650 -21882 396706 -21826
rect 396774 -21882 396830 -21826
rect 396898 -21882 396954 -21826
rect 397022 -21882 397078 -21826
rect 396526 -22006 396582 -21950
rect 396650 -22006 396706 -21950
rect 396774 -22006 396830 -21950
rect 396898 -22006 396954 -21950
rect 397022 -22006 397078 -21950
rect 396526 -22130 396582 -22074
rect 396650 -22130 396706 -22074
rect 396774 -22130 396830 -22074
rect 396898 -22130 396954 -22074
rect 397022 -22130 397078 -22074
rect 396526 -22254 396582 -22198
rect 396650 -22254 396706 -22198
rect 396774 -22254 396830 -22198
rect 396898 -22254 396954 -22198
rect 397022 -22254 397078 -22198
rect 396526 -22378 396582 -22322
rect 396650 -22378 396706 -22322
rect 396774 -22378 396830 -22322
rect 396898 -22378 396954 -22322
rect 397022 -22378 397078 -22322
rect 396526 -22502 396582 -22446
rect 396650 -22502 396706 -22446
rect 396774 -22502 396830 -22446
rect 396898 -22502 396954 -22446
rect 397022 -22502 397078 -22446
rect 396526 -22626 396582 -22570
rect 396650 -22626 396706 -22570
rect 396774 -22626 396830 -22570
rect 396898 -22626 396954 -22570
rect 397022 -22626 397078 -22570
rect 396526 -22750 396582 -22694
rect 396650 -22750 396706 -22694
rect 396774 -22750 396830 -22694
rect 396898 -22750 396954 -22694
rect 397022 -22750 397078 -22694
rect 396526 -22874 396582 -22818
rect 396650 -22874 396706 -22818
rect 396774 -22874 396830 -22818
rect 396898 -22874 396954 -22818
rect 397022 -22874 397078 -22818
rect 396526 -22998 396582 -22942
rect 396650 -22998 396706 -22942
rect 396774 -22998 396830 -22942
rect 396898 -22998 396954 -22942
rect 397022 -22998 397078 -22942
rect 396526 -23122 396582 -23066
rect 396650 -23122 396706 -23066
rect 396774 -23122 396830 -23066
rect 396898 -23122 396954 -23066
rect 397022 -23122 397078 -23066
rect 396526 -23246 396582 -23190
rect 396650 -23246 396706 -23190
rect 396774 -23246 396830 -23190
rect 396898 -23246 396954 -23190
rect 397022 -23246 397078 -23190
rect 396526 -23370 396582 -23314
rect 396650 -23370 396706 -23314
rect 396774 -23370 396830 -23314
rect 396898 -23370 396954 -23314
rect 397022 -23370 397078 -23314
rect 396526 -23494 396582 -23438
rect 396650 -23494 396706 -23438
rect 396774 -23494 396830 -23438
rect 396898 -23494 396954 -23438
rect 397022 -23494 397078 -23438
rect 396526 -23618 396582 -23562
rect 396650 -23618 396706 -23562
rect 396774 -23618 396830 -23562
rect 396898 -23618 396954 -23562
rect 397022 -23618 397078 -23562
rect 396526 -23742 396582 -23686
rect 396650 -23742 396706 -23686
rect 396774 -23742 396830 -23686
rect 396898 -23742 396954 -23686
rect 397022 -23742 397078 -23686
rect 396526 -23866 396582 -23810
rect 396650 -23866 396706 -23810
rect 396774 -23866 396830 -23810
rect 396898 -23866 396954 -23810
rect 397022 -23866 397078 -23810
rect 396526 -23990 396582 -23934
rect 396650 -23990 396706 -23934
rect 396774 -23990 396830 -23934
rect 396898 -23990 396954 -23934
rect 397022 -23990 397078 -23934
rect 396526 -24114 396582 -24058
rect 396650 -24114 396706 -24058
rect 396774 -24114 396830 -24058
rect 396898 -24114 396954 -24058
rect 397022 -24114 397078 -24058
rect 396526 -24238 396582 -24182
rect 396650 -24238 396706 -24182
rect 396774 -24238 396830 -24182
rect 396898 -24238 396954 -24182
rect 397022 -24238 397078 -24182
rect 396526 -24362 396582 -24306
rect 396650 -24362 396706 -24306
rect 396774 -24362 396830 -24306
rect 396898 -24362 396954 -24306
rect 397022 -24362 397078 -24306
rect 396526 -24486 396582 -24430
rect 396650 -24486 396706 -24430
rect 396774 -24486 396830 -24430
rect 396898 -24486 396954 -24430
rect 397022 -24486 397078 -24430
rect 396526 -24610 396582 -24554
rect 396650 -24610 396706 -24554
rect 396774 -24610 396830 -24554
rect 396898 -24610 396954 -24554
rect 397022 -24610 397078 -24554
rect 396526 -24734 396582 -24678
rect 396650 -24734 396706 -24678
rect 396774 -24734 396830 -24678
rect 396898 -24734 396954 -24678
rect 397022 -24734 397078 -24678
rect 396526 -24858 396582 -24802
rect 396650 -24858 396706 -24802
rect 396774 -24858 396830 -24802
rect 396898 -24858 396954 -24802
rect 397022 -24858 397078 -24802
rect 396526 -24982 396582 -24926
rect 396650 -24982 396706 -24926
rect 396774 -24982 396830 -24926
rect 396898 -24982 396954 -24926
rect 397022 -24982 397078 -24926
rect 396526 -25106 396582 -25050
rect 396650 -25106 396706 -25050
rect 396774 -25106 396830 -25050
rect 396898 -25106 396954 -25050
rect 397022 -25106 397078 -25050
rect 396526 -25230 396582 -25174
rect 396650 -25230 396706 -25174
rect 396774 -25230 396830 -25174
rect 396898 -25230 396954 -25174
rect 397022 -25230 397078 -25174
rect 396526 -25354 396582 -25298
rect 396650 -25354 396706 -25298
rect 396774 -25354 396830 -25298
rect 396898 -25354 396954 -25298
rect 397022 -25354 397078 -25298
rect 396526 -25478 396582 -25422
rect 396650 -25478 396706 -25422
rect 396774 -25478 396830 -25422
rect 396898 -25478 396954 -25422
rect 397022 -25478 397078 -25422
rect 388146 -25777 388202 -25721
rect 388270 -25777 388326 -25721
rect 388394 -25777 388450 -25721
rect 388518 -25777 388574 -25721
rect 388642 -25777 388698 -25721
rect 388766 -25777 388822 -25721
rect 388890 -25777 388946 -25721
rect 389014 -25777 389070 -25721
rect 389138 -25777 389194 -25721
rect 389262 -25777 389318 -25721
rect 389386 -25777 389442 -25721
rect 389510 -25777 389566 -25721
rect 389634 -25777 389690 -25721
rect 389758 -25777 389814 -25721
rect 389882 -25777 389938 -25721
rect 390006 -25777 390062 -25721
rect 390130 -25777 390186 -25721
rect 390254 -25777 390310 -25721
rect 390378 -25777 390434 -25721
rect 390502 -25777 390558 -25721
rect 390626 -25777 390682 -25721
rect 390750 -25777 390806 -25721
rect 390874 -25777 390930 -25721
rect 390998 -25777 391054 -25721
rect 391122 -25777 391178 -25721
rect 391246 -25777 391302 -25721
rect 391370 -25777 391426 -25721
rect 391494 -25777 391550 -25721
rect 391618 -25777 391674 -25721
rect 391742 -25777 391798 -25721
rect 391866 -25777 391922 -25721
rect 391990 -25777 392046 -25721
rect 392114 -25777 392170 -25721
rect 392238 -25777 392294 -25721
rect 392362 -25777 392418 -25721
rect 392486 -25777 392542 -25721
rect 392610 -25777 392666 -25721
rect 392734 -25777 392790 -25721
rect 392858 -25777 392914 -25721
rect 392982 -25777 393038 -25721
rect 393106 -25777 393162 -25721
rect 393230 -25777 393286 -25721
rect 393354 -25777 393410 -25721
rect 393478 -25777 393534 -25721
rect 393602 -25777 393658 -25721
rect 393726 -25777 393782 -25721
rect 393850 -25777 393906 -25721
rect 393974 -25777 394030 -25721
rect 394098 -25777 394154 -25721
rect 394222 -25777 394278 -25721
rect 394346 -25777 394402 -25721
rect 394470 -25777 394526 -25721
rect 394594 -25777 394650 -25721
rect 394718 -25777 394774 -25721
rect 394842 -25777 394898 -25721
rect 394966 -25777 395022 -25721
rect 395090 -25777 395146 -25721
rect 395214 -25777 395270 -25721
rect 395338 -25777 395394 -25721
rect 395462 -25777 395518 -25721
rect 395586 -25777 395642 -25721
rect 395710 -25777 395766 -25721
rect 395898 -25777 395954 -25721
rect 396022 -25777 396078 -25721
rect 396146 -25777 396202 -25721
rect 396270 -25777 396326 -25721
rect 396394 -25777 396450 -25721
rect 396518 -25777 396574 -25721
rect 396642 -25777 396698 -25721
rect 396766 -25777 396822 -25721
rect 396890 -25777 396946 -25721
rect 397014 -25777 397070 -25721
rect 388146 -25901 388202 -25845
rect 388270 -25901 388326 -25845
rect 388394 -25901 388450 -25845
rect 388518 -25901 388574 -25845
rect 388642 -25901 388698 -25845
rect 388766 -25901 388822 -25845
rect 388890 -25901 388946 -25845
rect 389014 -25901 389070 -25845
rect 389138 -25901 389194 -25845
rect 389262 -25901 389318 -25845
rect 389386 -25901 389442 -25845
rect 389510 -25901 389566 -25845
rect 389634 -25901 389690 -25845
rect 389758 -25901 389814 -25845
rect 389882 -25901 389938 -25845
rect 390006 -25901 390062 -25845
rect 390130 -25901 390186 -25845
rect 390254 -25901 390310 -25845
rect 390378 -25901 390434 -25845
rect 390502 -25901 390558 -25845
rect 390626 -25901 390682 -25845
rect 390750 -25901 390806 -25845
rect 390874 -25901 390930 -25845
rect 390998 -25901 391054 -25845
rect 391122 -25901 391178 -25845
rect 391246 -25901 391302 -25845
rect 391370 -25901 391426 -25845
rect 391494 -25901 391550 -25845
rect 391618 -25901 391674 -25845
rect 391742 -25901 391798 -25845
rect 391866 -25901 391922 -25845
rect 391990 -25901 392046 -25845
rect 392114 -25901 392170 -25845
rect 392238 -25901 392294 -25845
rect 392362 -25901 392418 -25845
rect 392486 -25901 392542 -25845
rect 392610 -25901 392666 -25845
rect 392734 -25901 392790 -25845
rect 392858 -25901 392914 -25845
rect 392982 -25901 393038 -25845
rect 393106 -25901 393162 -25845
rect 393230 -25901 393286 -25845
rect 393354 -25901 393410 -25845
rect 393478 -25901 393534 -25845
rect 393602 -25901 393658 -25845
rect 393726 -25901 393782 -25845
rect 393850 -25901 393906 -25845
rect 393974 -25901 394030 -25845
rect 394098 -25901 394154 -25845
rect 394222 -25901 394278 -25845
rect 394346 -25901 394402 -25845
rect 394470 -25901 394526 -25845
rect 394594 -25901 394650 -25845
rect 394718 -25901 394774 -25845
rect 394842 -25901 394898 -25845
rect 394966 -25901 395022 -25845
rect 395090 -25901 395146 -25845
rect 395214 -25901 395270 -25845
rect 395338 -25901 395394 -25845
rect 395462 -25901 395518 -25845
rect 395586 -25901 395642 -25845
rect 395710 -25901 395766 -25845
rect 395898 -25901 395954 -25845
rect 396022 -25901 396078 -25845
rect 396146 -25901 396202 -25845
rect 396270 -25901 396326 -25845
rect 396394 -25901 396450 -25845
rect 396518 -25901 396574 -25845
rect 396642 -25901 396698 -25845
rect 396766 -25901 396822 -25845
rect 396890 -25901 396946 -25845
rect 397014 -25901 397070 -25845
rect 388146 -26025 388202 -25969
rect 388270 -26025 388326 -25969
rect 388394 -26025 388450 -25969
rect 388518 -26025 388574 -25969
rect 388642 -26025 388698 -25969
rect 388766 -26025 388822 -25969
rect 388890 -26025 388946 -25969
rect 389014 -26025 389070 -25969
rect 389138 -26025 389194 -25969
rect 389262 -26025 389318 -25969
rect 389386 -26025 389442 -25969
rect 389510 -26025 389566 -25969
rect 389634 -26025 389690 -25969
rect 389758 -26025 389814 -25969
rect 389882 -26025 389938 -25969
rect 390006 -26025 390062 -25969
rect 390130 -26025 390186 -25969
rect 390254 -26025 390310 -25969
rect 390378 -26025 390434 -25969
rect 390502 -26025 390558 -25969
rect 390626 -26025 390682 -25969
rect 390750 -26025 390806 -25969
rect 390874 -26025 390930 -25969
rect 390998 -26025 391054 -25969
rect 391122 -26025 391178 -25969
rect 391246 -26025 391302 -25969
rect 391370 -26025 391426 -25969
rect 391494 -26025 391550 -25969
rect 391618 -26025 391674 -25969
rect 391742 -26025 391798 -25969
rect 391866 -26025 391922 -25969
rect 391990 -26025 392046 -25969
rect 392114 -26025 392170 -25969
rect 392238 -26025 392294 -25969
rect 392362 -26025 392418 -25969
rect 392486 -26025 392542 -25969
rect 392610 -26025 392666 -25969
rect 392734 -26025 392790 -25969
rect 392858 -26025 392914 -25969
rect 392982 -26025 393038 -25969
rect 393106 -26025 393162 -25969
rect 393230 -26025 393286 -25969
rect 393354 -26025 393410 -25969
rect 393478 -26025 393534 -25969
rect 393602 -26025 393658 -25969
rect 393726 -26025 393782 -25969
rect 393850 -26025 393906 -25969
rect 393974 -26025 394030 -25969
rect 394098 -26025 394154 -25969
rect 394222 -26025 394278 -25969
rect 394346 -26025 394402 -25969
rect 394470 -26025 394526 -25969
rect 394594 -26025 394650 -25969
rect 394718 -26025 394774 -25969
rect 394842 -26025 394898 -25969
rect 394966 -26025 395022 -25969
rect 395090 -26025 395146 -25969
rect 395214 -26025 395270 -25969
rect 395338 -26025 395394 -25969
rect 395462 -26025 395518 -25969
rect 395586 -26025 395642 -25969
rect 395710 -26025 395766 -25969
rect 395898 -26025 395954 -25969
rect 396022 -26025 396078 -25969
rect 396146 -26025 396202 -25969
rect 396270 -26025 396326 -25969
rect 396394 -26025 396450 -25969
rect 396518 -26025 396574 -25969
rect 396642 -26025 396698 -25969
rect 396766 -26025 396822 -25969
rect 396890 -26025 396946 -25969
rect 397014 -26025 397070 -25969
rect 388146 -26149 388202 -26093
rect 388270 -26149 388326 -26093
rect 388394 -26149 388450 -26093
rect 388518 -26149 388574 -26093
rect 388642 -26149 388698 -26093
rect 388766 -26149 388822 -26093
rect 388890 -26149 388946 -26093
rect 389014 -26149 389070 -26093
rect 389138 -26149 389194 -26093
rect 389262 -26149 389318 -26093
rect 389386 -26149 389442 -26093
rect 389510 -26149 389566 -26093
rect 389634 -26149 389690 -26093
rect 389758 -26149 389814 -26093
rect 389882 -26149 389938 -26093
rect 390006 -26149 390062 -26093
rect 390130 -26149 390186 -26093
rect 390254 -26149 390310 -26093
rect 390378 -26149 390434 -26093
rect 390502 -26149 390558 -26093
rect 390626 -26149 390682 -26093
rect 390750 -26149 390806 -26093
rect 390874 -26149 390930 -26093
rect 390998 -26149 391054 -26093
rect 391122 -26149 391178 -26093
rect 391246 -26149 391302 -26093
rect 391370 -26149 391426 -26093
rect 391494 -26149 391550 -26093
rect 391618 -26149 391674 -26093
rect 391742 -26149 391798 -26093
rect 391866 -26149 391922 -26093
rect 391990 -26149 392046 -26093
rect 392114 -26149 392170 -26093
rect 392238 -26149 392294 -26093
rect 392362 -26149 392418 -26093
rect 392486 -26149 392542 -26093
rect 392610 -26149 392666 -26093
rect 392734 -26149 392790 -26093
rect 392858 -26149 392914 -26093
rect 392982 -26149 393038 -26093
rect 393106 -26149 393162 -26093
rect 393230 -26149 393286 -26093
rect 393354 -26149 393410 -26093
rect 393478 -26149 393534 -26093
rect 393602 -26149 393658 -26093
rect 393726 -26149 393782 -26093
rect 393850 -26149 393906 -26093
rect 393974 -26149 394030 -26093
rect 394098 -26149 394154 -26093
rect 394222 -26149 394278 -26093
rect 394346 -26149 394402 -26093
rect 394470 -26149 394526 -26093
rect 394594 -26149 394650 -26093
rect 394718 -26149 394774 -26093
rect 394842 -26149 394898 -26093
rect 394966 -26149 395022 -26093
rect 395090 -26149 395146 -26093
rect 395214 -26149 395270 -26093
rect 395338 -26149 395394 -26093
rect 395462 -26149 395518 -26093
rect 395586 -26149 395642 -26093
rect 395710 -26149 395766 -26093
rect 395898 -26149 395954 -26093
rect 396022 -26149 396078 -26093
rect 396146 -26149 396202 -26093
rect 396270 -26149 396326 -26093
rect 396394 -26149 396450 -26093
rect 396518 -26149 396574 -26093
rect 396642 -26149 396698 -26093
rect 396766 -26149 396822 -26093
rect 396890 -26149 396946 -26093
rect 397014 -26149 397070 -26093
<< metal5 >>
rect 388000 -17191 397200 -17070
rect 388000 -17247 388146 -17191
rect 388202 -17247 388270 -17191
rect 388326 -17247 388394 -17191
rect 388450 -17247 388518 -17191
rect 388574 -17247 388642 -17191
rect 388698 -17247 388766 -17191
rect 388822 -17247 388890 -17191
rect 388946 -17247 389014 -17191
rect 389070 -17247 389138 -17191
rect 389194 -17247 389262 -17191
rect 389318 -17247 389386 -17191
rect 389442 -17247 389510 -17191
rect 389566 -17247 389634 -17191
rect 389690 -17247 389758 -17191
rect 389814 -17247 389882 -17191
rect 389938 -17247 390006 -17191
rect 390062 -17247 390130 -17191
rect 390186 -17247 390254 -17191
rect 390310 -17247 390378 -17191
rect 390434 -17247 390502 -17191
rect 390558 -17247 390626 -17191
rect 390682 -17247 390750 -17191
rect 390806 -17247 390874 -17191
rect 390930 -17247 390998 -17191
rect 391054 -17247 391122 -17191
rect 391178 -17247 391246 -17191
rect 391302 -17247 391370 -17191
rect 391426 -17247 391494 -17191
rect 391550 -17247 391618 -17191
rect 391674 -17247 391742 -17191
rect 391798 -17247 391866 -17191
rect 391922 -17247 391990 -17191
rect 392046 -17247 392114 -17191
rect 392170 -17247 392238 -17191
rect 392294 -17247 392362 -17191
rect 392418 -17247 392486 -17191
rect 392542 -17247 392610 -17191
rect 392666 -17247 392734 -17191
rect 392790 -17247 392858 -17191
rect 392914 -17247 392982 -17191
rect 393038 -17247 393106 -17191
rect 393162 -17247 393230 -17191
rect 393286 -17247 393354 -17191
rect 393410 -17247 393478 -17191
rect 393534 -17247 393602 -17191
rect 393658 -17247 393726 -17191
rect 393782 -17247 393850 -17191
rect 393906 -17247 393974 -17191
rect 394030 -17247 394098 -17191
rect 394154 -17247 394222 -17191
rect 394278 -17247 394346 -17191
rect 394402 -17247 394470 -17191
rect 394526 -17247 394594 -17191
rect 394650 -17247 394718 -17191
rect 394774 -17247 394842 -17191
rect 394898 -17247 394966 -17191
rect 395022 -17247 395090 -17191
rect 395146 -17247 395214 -17191
rect 395270 -17247 395338 -17191
rect 395394 -17247 395462 -17191
rect 395518 -17247 395586 -17191
rect 395642 -17247 395710 -17191
rect 395766 -17247 395898 -17191
rect 395954 -17247 396022 -17191
rect 396078 -17247 396146 -17191
rect 396202 -17247 396270 -17191
rect 396326 -17247 396394 -17191
rect 396450 -17247 396518 -17191
rect 396574 -17247 396642 -17191
rect 396698 -17247 396766 -17191
rect 396822 -17247 396890 -17191
rect 396946 -17247 397014 -17191
rect 397070 -17247 397200 -17191
rect 388000 -17315 397200 -17247
rect 388000 -17371 388146 -17315
rect 388202 -17371 388270 -17315
rect 388326 -17371 388394 -17315
rect 388450 -17371 388518 -17315
rect 388574 -17371 388642 -17315
rect 388698 -17371 388766 -17315
rect 388822 -17371 388890 -17315
rect 388946 -17371 389014 -17315
rect 389070 -17371 389138 -17315
rect 389194 -17371 389262 -17315
rect 389318 -17371 389386 -17315
rect 389442 -17371 389510 -17315
rect 389566 -17371 389634 -17315
rect 389690 -17371 389758 -17315
rect 389814 -17371 389882 -17315
rect 389938 -17371 390006 -17315
rect 390062 -17371 390130 -17315
rect 390186 -17371 390254 -17315
rect 390310 -17371 390378 -17315
rect 390434 -17371 390502 -17315
rect 390558 -17371 390626 -17315
rect 390682 -17371 390750 -17315
rect 390806 -17371 390874 -17315
rect 390930 -17371 390998 -17315
rect 391054 -17371 391122 -17315
rect 391178 -17371 391246 -17315
rect 391302 -17371 391370 -17315
rect 391426 -17371 391494 -17315
rect 391550 -17371 391618 -17315
rect 391674 -17371 391742 -17315
rect 391798 -17371 391866 -17315
rect 391922 -17371 391990 -17315
rect 392046 -17371 392114 -17315
rect 392170 -17371 392238 -17315
rect 392294 -17371 392362 -17315
rect 392418 -17371 392486 -17315
rect 392542 -17371 392610 -17315
rect 392666 -17371 392734 -17315
rect 392790 -17371 392858 -17315
rect 392914 -17371 392982 -17315
rect 393038 -17371 393106 -17315
rect 393162 -17371 393230 -17315
rect 393286 -17371 393354 -17315
rect 393410 -17371 393478 -17315
rect 393534 -17371 393602 -17315
rect 393658 -17371 393726 -17315
rect 393782 -17371 393850 -17315
rect 393906 -17371 393974 -17315
rect 394030 -17371 394098 -17315
rect 394154 -17371 394222 -17315
rect 394278 -17371 394346 -17315
rect 394402 -17371 394470 -17315
rect 394526 -17371 394594 -17315
rect 394650 -17371 394718 -17315
rect 394774 -17371 394842 -17315
rect 394898 -17371 394966 -17315
rect 395022 -17371 395090 -17315
rect 395146 -17371 395214 -17315
rect 395270 -17371 395338 -17315
rect 395394 -17371 395462 -17315
rect 395518 -17371 395586 -17315
rect 395642 -17371 395710 -17315
rect 395766 -17371 395898 -17315
rect 395954 -17371 396022 -17315
rect 396078 -17371 396146 -17315
rect 396202 -17371 396270 -17315
rect 396326 -17371 396394 -17315
rect 396450 -17371 396518 -17315
rect 396574 -17371 396642 -17315
rect 396698 -17371 396766 -17315
rect 396822 -17371 396890 -17315
rect 396946 -17371 397014 -17315
rect 397070 -17371 397200 -17315
rect 388000 -17439 397200 -17371
rect 388000 -17495 388146 -17439
rect 388202 -17495 388270 -17439
rect 388326 -17495 388394 -17439
rect 388450 -17495 388518 -17439
rect 388574 -17495 388642 -17439
rect 388698 -17495 388766 -17439
rect 388822 -17495 388890 -17439
rect 388946 -17495 389014 -17439
rect 389070 -17495 389138 -17439
rect 389194 -17495 389262 -17439
rect 389318 -17495 389386 -17439
rect 389442 -17495 389510 -17439
rect 389566 -17495 389634 -17439
rect 389690 -17495 389758 -17439
rect 389814 -17495 389882 -17439
rect 389938 -17495 390006 -17439
rect 390062 -17495 390130 -17439
rect 390186 -17495 390254 -17439
rect 390310 -17495 390378 -17439
rect 390434 -17495 390502 -17439
rect 390558 -17495 390626 -17439
rect 390682 -17495 390750 -17439
rect 390806 -17495 390874 -17439
rect 390930 -17495 390998 -17439
rect 391054 -17495 391122 -17439
rect 391178 -17495 391246 -17439
rect 391302 -17495 391370 -17439
rect 391426 -17495 391494 -17439
rect 391550 -17495 391618 -17439
rect 391674 -17495 391742 -17439
rect 391798 -17495 391866 -17439
rect 391922 -17495 391990 -17439
rect 392046 -17495 392114 -17439
rect 392170 -17495 392238 -17439
rect 392294 -17495 392362 -17439
rect 392418 -17495 392486 -17439
rect 392542 -17495 392610 -17439
rect 392666 -17495 392734 -17439
rect 392790 -17495 392858 -17439
rect 392914 -17495 392982 -17439
rect 393038 -17495 393106 -17439
rect 393162 -17495 393230 -17439
rect 393286 -17495 393354 -17439
rect 393410 -17495 393478 -17439
rect 393534 -17495 393602 -17439
rect 393658 -17495 393726 -17439
rect 393782 -17495 393850 -17439
rect 393906 -17495 393974 -17439
rect 394030 -17495 394098 -17439
rect 394154 -17495 394222 -17439
rect 394278 -17495 394346 -17439
rect 394402 -17495 394470 -17439
rect 394526 -17495 394594 -17439
rect 394650 -17495 394718 -17439
rect 394774 -17495 394842 -17439
rect 394898 -17495 394966 -17439
rect 395022 -17495 395090 -17439
rect 395146 -17495 395214 -17439
rect 395270 -17495 395338 -17439
rect 395394 -17495 395462 -17439
rect 395518 -17495 395586 -17439
rect 395642 -17495 395710 -17439
rect 395766 -17495 395898 -17439
rect 395954 -17495 396022 -17439
rect 396078 -17495 396146 -17439
rect 396202 -17495 396270 -17439
rect 396326 -17495 396394 -17439
rect 396450 -17495 396518 -17439
rect 396574 -17495 396642 -17439
rect 396698 -17495 396766 -17439
rect 396822 -17495 396890 -17439
rect 396946 -17495 397014 -17439
rect 397070 -17495 397200 -17439
rect 388000 -17563 397200 -17495
rect 388000 -17619 388146 -17563
rect 388202 -17619 388270 -17563
rect 388326 -17619 388394 -17563
rect 388450 -17619 388518 -17563
rect 388574 -17619 388642 -17563
rect 388698 -17619 388766 -17563
rect 388822 -17619 388890 -17563
rect 388946 -17619 389014 -17563
rect 389070 -17619 389138 -17563
rect 389194 -17619 389262 -17563
rect 389318 -17619 389386 -17563
rect 389442 -17619 389510 -17563
rect 389566 -17619 389634 -17563
rect 389690 -17619 389758 -17563
rect 389814 -17619 389882 -17563
rect 389938 -17619 390006 -17563
rect 390062 -17619 390130 -17563
rect 390186 -17619 390254 -17563
rect 390310 -17619 390378 -17563
rect 390434 -17619 390502 -17563
rect 390558 -17619 390626 -17563
rect 390682 -17619 390750 -17563
rect 390806 -17619 390874 -17563
rect 390930 -17619 390998 -17563
rect 391054 -17619 391122 -17563
rect 391178 -17619 391246 -17563
rect 391302 -17619 391370 -17563
rect 391426 -17619 391494 -17563
rect 391550 -17619 391618 -17563
rect 391674 -17619 391742 -17563
rect 391798 -17619 391866 -17563
rect 391922 -17619 391990 -17563
rect 392046 -17619 392114 -17563
rect 392170 -17619 392238 -17563
rect 392294 -17619 392362 -17563
rect 392418 -17619 392486 -17563
rect 392542 -17619 392610 -17563
rect 392666 -17619 392734 -17563
rect 392790 -17619 392858 -17563
rect 392914 -17619 392982 -17563
rect 393038 -17619 393106 -17563
rect 393162 -17619 393230 -17563
rect 393286 -17619 393354 -17563
rect 393410 -17619 393478 -17563
rect 393534 -17619 393602 -17563
rect 393658 -17619 393726 -17563
rect 393782 -17619 393850 -17563
rect 393906 -17619 393974 -17563
rect 394030 -17619 394098 -17563
rect 394154 -17619 394222 -17563
rect 394278 -17619 394346 -17563
rect 394402 -17619 394470 -17563
rect 394526 -17619 394594 -17563
rect 394650 -17619 394718 -17563
rect 394774 -17619 394842 -17563
rect 394898 -17619 394966 -17563
rect 395022 -17619 395090 -17563
rect 395146 -17619 395214 -17563
rect 395270 -17619 395338 -17563
rect 395394 -17619 395462 -17563
rect 395518 -17619 395586 -17563
rect 395642 -17619 395710 -17563
rect 395766 -17619 395898 -17563
rect 395954 -17619 396022 -17563
rect 396078 -17619 396146 -17563
rect 396202 -17619 396270 -17563
rect 396326 -17619 396394 -17563
rect 396450 -17619 396518 -17563
rect 396574 -17619 396642 -17563
rect 396698 -17619 396766 -17563
rect 396822 -17619 396890 -17563
rect 396946 -17619 397014 -17563
rect 397070 -17619 397200 -17563
rect 388000 -17858 397200 -17619
rect 388000 -17914 388114 -17858
rect 388170 -17914 388238 -17858
rect 388294 -17914 388362 -17858
rect 388418 -17914 388486 -17858
rect 388542 -17914 388610 -17858
rect 388666 -17914 396526 -17858
rect 396582 -17914 396650 -17858
rect 396706 -17914 396774 -17858
rect 396830 -17914 396898 -17858
rect 396954 -17914 397022 -17858
rect 397078 -17914 397200 -17858
rect 388000 -17950 397200 -17914
rect 388000 -17982 389141 -17950
rect 388000 -18038 388114 -17982
rect 388170 -18038 388238 -17982
rect 388294 -18038 388362 -17982
rect 388418 -18038 388486 -17982
rect 388542 -18038 388610 -17982
rect 388666 -18006 389141 -17982
rect 389197 -18006 389283 -17950
rect 389339 -18006 389542 -17950
rect 389598 -18006 389684 -17950
rect 389740 -18006 389942 -17950
rect 389998 -18006 390084 -17950
rect 390140 -18006 390339 -17950
rect 390395 -18006 390481 -17950
rect 390537 -18006 390736 -17950
rect 390792 -18006 390878 -17950
rect 390934 -18006 391140 -17950
rect 391196 -18006 391282 -17950
rect 391338 -18006 391536 -17950
rect 391592 -18006 391678 -17950
rect 391734 -18006 391936 -17950
rect 391992 -18006 392078 -17950
rect 392134 -18006 392333 -17950
rect 392389 -18006 392475 -17950
rect 392531 -18006 392738 -17950
rect 392794 -18006 392880 -17950
rect 392936 -18006 393138 -17950
rect 393194 -18006 393280 -17950
rect 393336 -18006 393543 -17950
rect 393599 -18006 393685 -17950
rect 393741 -18006 393940 -17950
rect 393996 -18006 394082 -17950
rect 394138 -18006 394337 -17950
rect 394393 -18006 394479 -17950
rect 394535 -18006 394740 -17950
rect 394796 -18006 394882 -17950
rect 394938 -18006 395142 -17950
rect 395198 -18006 395284 -17950
rect 395340 -18006 395545 -17950
rect 395601 -18006 395687 -17950
rect 395743 -18006 395941 -17950
rect 395997 -18006 396083 -17950
rect 396139 -17982 397200 -17950
rect 396139 -18006 396526 -17982
rect 388666 -18038 396526 -18006
rect 396582 -18038 396650 -17982
rect 396706 -18038 396774 -17982
rect 396830 -18038 396898 -17982
rect 396954 -18038 397022 -17982
rect 397078 -18038 397200 -17982
rect 388000 -18092 397200 -18038
rect 388000 -18106 389141 -18092
rect 388000 -18162 388114 -18106
rect 388170 -18162 388238 -18106
rect 388294 -18162 388362 -18106
rect 388418 -18162 388486 -18106
rect 388542 -18162 388610 -18106
rect 388666 -18148 389141 -18106
rect 389197 -18148 389283 -18092
rect 389339 -18148 389542 -18092
rect 389598 -18148 389684 -18092
rect 389740 -18148 389942 -18092
rect 389998 -18148 390084 -18092
rect 390140 -18148 390339 -18092
rect 390395 -18148 390481 -18092
rect 390537 -18148 390736 -18092
rect 390792 -18148 390878 -18092
rect 390934 -18148 391140 -18092
rect 391196 -18148 391282 -18092
rect 391338 -18148 391536 -18092
rect 391592 -18148 391678 -18092
rect 391734 -18148 391936 -18092
rect 391992 -18148 392078 -18092
rect 392134 -18148 392333 -18092
rect 392389 -18148 392475 -18092
rect 392531 -18148 392738 -18092
rect 392794 -18148 392880 -18092
rect 392936 -18148 393138 -18092
rect 393194 -18148 393280 -18092
rect 393336 -18148 393543 -18092
rect 393599 -18148 393685 -18092
rect 393741 -18148 393940 -18092
rect 393996 -18148 394082 -18092
rect 394138 -18148 394337 -18092
rect 394393 -18148 394479 -18092
rect 394535 -18148 394740 -18092
rect 394796 -18148 394882 -18092
rect 394938 -18148 395142 -18092
rect 395198 -18148 395284 -18092
rect 395340 -18148 395545 -18092
rect 395601 -18148 395687 -18092
rect 395743 -18148 395941 -18092
rect 395997 -18148 396083 -18092
rect 396139 -18106 397200 -18092
rect 396139 -18148 396526 -18106
rect 388666 -18162 396526 -18148
rect 396582 -18162 396650 -18106
rect 396706 -18162 396774 -18106
rect 396830 -18162 396898 -18106
rect 396954 -18162 397022 -18106
rect 397078 -18162 397200 -18106
rect 388000 -18230 397200 -18162
rect 388000 -18286 388114 -18230
rect 388170 -18286 388238 -18230
rect 388294 -18286 388362 -18230
rect 388418 -18286 388486 -18230
rect 388542 -18286 388610 -18230
rect 388666 -18234 396526 -18230
rect 388666 -18286 389141 -18234
rect 388000 -18290 389141 -18286
rect 389197 -18290 389283 -18234
rect 389339 -18290 389542 -18234
rect 389598 -18290 389684 -18234
rect 389740 -18290 389942 -18234
rect 389998 -18290 390084 -18234
rect 390140 -18290 390339 -18234
rect 390395 -18290 390481 -18234
rect 390537 -18290 390736 -18234
rect 390792 -18290 390878 -18234
rect 390934 -18290 391140 -18234
rect 391196 -18290 391282 -18234
rect 391338 -18290 391536 -18234
rect 391592 -18290 391678 -18234
rect 391734 -18290 391936 -18234
rect 391992 -18290 392078 -18234
rect 392134 -18290 392333 -18234
rect 392389 -18290 392475 -18234
rect 392531 -18290 392738 -18234
rect 392794 -18290 392880 -18234
rect 392936 -18290 393138 -18234
rect 393194 -18290 393280 -18234
rect 393336 -18290 393543 -18234
rect 393599 -18290 393685 -18234
rect 393741 -18290 393940 -18234
rect 393996 -18290 394082 -18234
rect 394138 -18290 394337 -18234
rect 394393 -18290 394479 -18234
rect 394535 -18290 394740 -18234
rect 394796 -18290 394882 -18234
rect 394938 -18290 395142 -18234
rect 395198 -18290 395284 -18234
rect 395340 -18290 395545 -18234
rect 395601 -18290 395687 -18234
rect 395743 -18290 395941 -18234
rect 395997 -18290 396083 -18234
rect 396139 -18286 396526 -18234
rect 396582 -18286 396650 -18230
rect 396706 -18286 396774 -18230
rect 396830 -18286 396898 -18230
rect 396954 -18286 397022 -18230
rect 397078 -18286 397200 -18230
rect 396139 -18290 397200 -18286
rect 388000 -18354 397200 -18290
rect 388000 -18410 388114 -18354
rect 388170 -18410 388238 -18354
rect 388294 -18410 388362 -18354
rect 388418 -18410 388486 -18354
rect 388542 -18410 388610 -18354
rect 388666 -18376 396526 -18354
rect 388666 -18410 389141 -18376
rect 388000 -18432 389141 -18410
rect 389197 -18432 389283 -18376
rect 389339 -18432 389542 -18376
rect 389598 -18432 389684 -18376
rect 389740 -18432 389942 -18376
rect 389998 -18432 390084 -18376
rect 390140 -18432 390339 -18376
rect 390395 -18432 390481 -18376
rect 390537 -18432 390736 -18376
rect 390792 -18432 390878 -18376
rect 390934 -18432 391140 -18376
rect 391196 -18432 391282 -18376
rect 391338 -18432 391536 -18376
rect 391592 -18432 391678 -18376
rect 391734 -18432 391936 -18376
rect 391992 -18432 392078 -18376
rect 392134 -18432 392333 -18376
rect 392389 -18432 392475 -18376
rect 392531 -18432 392738 -18376
rect 392794 -18432 392880 -18376
rect 392936 -18432 393138 -18376
rect 393194 -18432 393280 -18376
rect 393336 -18432 393543 -18376
rect 393599 -18432 393685 -18376
rect 393741 -18432 393940 -18376
rect 393996 -18432 394082 -18376
rect 394138 -18432 394337 -18376
rect 394393 -18432 394479 -18376
rect 394535 -18432 394740 -18376
rect 394796 -18432 394882 -18376
rect 394938 -18432 395142 -18376
rect 395198 -18432 395284 -18376
rect 395340 -18432 395545 -18376
rect 395601 -18432 395687 -18376
rect 395743 -18432 395941 -18376
rect 395997 -18432 396083 -18376
rect 396139 -18410 396526 -18376
rect 396582 -18410 396650 -18354
rect 396706 -18410 396774 -18354
rect 396830 -18410 396898 -18354
rect 396954 -18410 397022 -18354
rect 397078 -18410 397200 -18354
rect 396139 -18432 397200 -18410
rect 388000 -18478 397200 -18432
rect 388000 -18534 388114 -18478
rect 388170 -18534 388238 -18478
rect 388294 -18534 388362 -18478
rect 388418 -18534 388486 -18478
rect 388542 -18534 388610 -18478
rect 388666 -18518 396526 -18478
rect 388666 -18534 389141 -18518
rect 388000 -18574 389141 -18534
rect 389197 -18574 389283 -18518
rect 389339 -18574 389542 -18518
rect 389598 -18574 389684 -18518
rect 389740 -18574 389942 -18518
rect 389998 -18574 390084 -18518
rect 390140 -18574 390339 -18518
rect 390395 -18574 390481 -18518
rect 390537 -18574 390736 -18518
rect 390792 -18574 390878 -18518
rect 390934 -18574 391140 -18518
rect 391196 -18574 391282 -18518
rect 391338 -18574 391536 -18518
rect 391592 -18574 391678 -18518
rect 391734 -18574 391936 -18518
rect 391992 -18574 392078 -18518
rect 392134 -18574 392333 -18518
rect 392389 -18574 392475 -18518
rect 392531 -18574 392738 -18518
rect 392794 -18574 392880 -18518
rect 392936 -18574 393138 -18518
rect 393194 -18574 393280 -18518
rect 393336 -18574 393543 -18518
rect 393599 -18574 393685 -18518
rect 393741 -18574 393940 -18518
rect 393996 -18574 394082 -18518
rect 394138 -18574 394337 -18518
rect 394393 -18574 394479 -18518
rect 394535 -18574 394740 -18518
rect 394796 -18574 394882 -18518
rect 394938 -18574 395142 -18518
rect 395198 -18574 395284 -18518
rect 395340 -18574 395545 -18518
rect 395601 -18574 395687 -18518
rect 395743 -18574 395941 -18518
rect 395997 -18574 396083 -18518
rect 396139 -18534 396526 -18518
rect 396582 -18534 396650 -18478
rect 396706 -18534 396774 -18478
rect 396830 -18534 396898 -18478
rect 396954 -18534 397022 -18478
rect 397078 -18534 397200 -18478
rect 396139 -18574 397200 -18534
rect 388000 -18602 397200 -18574
rect 388000 -18658 388114 -18602
rect 388170 -18658 388238 -18602
rect 388294 -18658 388362 -18602
rect 388418 -18658 388486 -18602
rect 388542 -18658 388610 -18602
rect 388666 -18658 396526 -18602
rect 396582 -18658 396650 -18602
rect 396706 -18658 396774 -18602
rect 396830 -18658 396898 -18602
rect 396954 -18658 397022 -18602
rect 397078 -18658 397200 -18602
rect 388000 -18660 397200 -18658
rect 388000 -18716 389141 -18660
rect 389197 -18716 389283 -18660
rect 389339 -18716 389542 -18660
rect 389598 -18716 389684 -18660
rect 389740 -18716 389942 -18660
rect 389998 -18716 390084 -18660
rect 390140 -18716 390339 -18660
rect 390395 -18716 390481 -18660
rect 390537 -18716 390736 -18660
rect 390792 -18716 390878 -18660
rect 390934 -18716 391140 -18660
rect 391196 -18716 391282 -18660
rect 391338 -18716 391536 -18660
rect 391592 -18716 391678 -18660
rect 391734 -18716 391936 -18660
rect 391992 -18716 392078 -18660
rect 392134 -18716 392333 -18660
rect 392389 -18716 392475 -18660
rect 392531 -18716 392738 -18660
rect 392794 -18716 392880 -18660
rect 392936 -18716 393138 -18660
rect 393194 -18716 393280 -18660
rect 393336 -18716 393543 -18660
rect 393599 -18716 393685 -18660
rect 393741 -18716 393940 -18660
rect 393996 -18716 394082 -18660
rect 394138 -18716 394337 -18660
rect 394393 -18716 394479 -18660
rect 394535 -18716 394740 -18660
rect 394796 -18716 394882 -18660
rect 394938 -18716 395142 -18660
rect 395198 -18716 395284 -18660
rect 395340 -18716 395545 -18660
rect 395601 -18716 395687 -18660
rect 395743 -18716 395941 -18660
rect 395997 -18716 396083 -18660
rect 396139 -18716 397200 -18660
rect 388000 -18726 397200 -18716
rect 388000 -18782 388114 -18726
rect 388170 -18782 388238 -18726
rect 388294 -18782 388362 -18726
rect 388418 -18782 388486 -18726
rect 388542 -18782 388610 -18726
rect 388666 -18782 396526 -18726
rect 396582 -18782 396650 -18726
rect 396706 -18782 396774 -18726
rect 396830 -18782 396898 -18726
rect 396954 -18782 397022 -18726
rect 397078 -18782 397200 -18726
rect 388000 -18802 397200 -18782
rect 388000 -18850 389141 -18802
rect 388000 -18906 388114 -18850
rect 388170 -18906 388238 -18850
rect 388294 -18906 388362 -18850
rect 388418 -18906 388486 -18850
rect 388542 -18906 388610 -18850
rect 388666 -18858 389141 -18850
rect 389197 -18858 389283 -18802
rect 389339 -18858 389542 -18802
rect 389598 -18858 389684 -18802
rect 389740 -18858 389942 -18802
rect 389998 -18858 390084 -18802
rect 390140 -18858 390339 -18802
rect 390395 -18858 390481 -18802
rect 390537 -18858 390736 -18802
rect 390792 -18858 390878 -18802
rect 390934 -18858 391140 -18802
rect 391196 -18858 391282 -18802
rect 391338 -18858 391536 -18802
rect 391592 -18858 391678 -18802
rect 391734 -18858 391936 -18802
rect 391992 -18858 392078 -18802
rect 392134 -18858 392333 -18802
rect 392389 -18858 392475 -18802
rect 392531 -18858 392738 -18802
rect 392794 -18858 392880 -18802
rect 392936 -18858 393138 -18802
rect 393194 -18858 393280 -18802
rect 393336 -18858 393543 -18802
rect 393599 -18858 393685 -18802
rect 393741 -18858 393940 -18802
rect 393996 -18858 394082 -18802
rect 394138 -18858 394337 -18802
rect 394393 -18858 394479 -18802
rect 394535 -18858 394740 -18802
rect 394796 -18858 394882 -18802
rect 394938 -18858 395142 -18802
rect 395198 -18858 395284 -18802
rect 395340 -18858 395545 -18802
rect 395601 -18858 395687 -18802
rect 395743 -18858 395941 -18802
rect 395997 -18858 396083 -18802
rect 396139 -18850 397200 -18802
rect 396139 -18858 396526 -18850
rect 388666 -18906 396526 -18858
rect 396582 -18906 396650 -18850
rect 396706 -18906 396774 -18850
rect 396830 -18906 396898 -18850
rect 396954 -18906 397022 -18850
rect 397078 -18906 397200 -18850
rect 388000 -18944 397200 -18906
rect 388000 -18974 389141 -18944
rect 388000 -19030 388114 -18974
rect 388170 -19030 388238 -18974
rect 388294 -19030 388362 -18974
rect 388418 -19030 388486 -18974
rect 388542 -19030 388610 -18974
rect 388666 -19000 389141 -18974
rect 389197 -19000 389283 -18944
rect 389339 -19000 389542 -18944
rect 389598 -19000 389684 -18944
rect 389740 -19000 389942 -18944
rect 389998 -19000 390084 -18944
rect 390140 -19000 390339 -18944
rect 390395 -19000 390481 -18944
rect 390537 -19000 390736 -18944
rect 390792 -19000 390878 -18944
rect 390934 -19000 391140 -18944
rect 391196 -19000 391282 -18944
rect 391338 -19000 391536 -18944
rect 391592 -19000 391678 -18944
rect 391734 -19000 391936 -18944
rect 391992 -19000 392078 -18944
rect 392134 -19000 392333 -18944
rect 392389 -19000 392475 -18944
rect 392531 -19000 392738 -18944
rect 392794 -19000 392880 -18944
rect 392936 -19000 393138 -18944
rect 393194 -19000 393280 -18944
rect 393336 -19000 393543 -18944
rect 393599 -19000 393685 -18944
rect 393741 -19000 393940 -18944
rect 393996 -19000 394082 -18944
rect 394138 -19000 394337 -18944
rect 394393 -19000 394479 -18944
rect 394535 -19000 394740 -18944
rect 394796 -19000 394882 -18944
rect 394938 -19000 395142 -18944
rect 395198 -19000 395284 -18944
rect 395340 -19000 395545 -18944
rect 395601 -19000 395687 -18944
rect 395743 -19000 395941 -18944
rect 395997 -19000 396083 -18944
rect 396139 -18974 397200 -18944
rect 396139 -19000 396526 -18974
rect 388666 -19030 396526 -19000
rect 396582 -19030 396650 -18974
rect 396706 -19030 396774 -18974
rect 396830 -19030 396898 -18974
rect 396954 -19030 397022 -18974
rect 397078 -19030 397200 -18974
rect 388000 -19086 397200 -19030
rect 388000 -19098 389141 -19086
rect 388000 -19154 388114 -19098
rect 388170 -19154 388238 -19098
rect 388294 -19154 388362 -19098
rect 388418 -19154 388486 -19098
rect 388542 -19154 388610 -19098
rect 388666 -19142 389141 -19098
rect 389197 -19142 389283 -19086
rect 389339 -19142 389542 -19086
rect 389598 -19142 389684 -19086
rect 389740 -19142 389942 -19086
rect 389998 -19142 390084 -19086
rect 390140 -19142 390339 -19086
rect 390395 -19142 390481 -19086
rect 390537 -19142 390736 -19086
rect 390792 -19142 390878 -19086
rect 390934 -19142 391140 -19086
rect 391196 -19142 391282 -19086
rect 391338 -19142 391536 -19086
rect 391592 -19142 391678 -19086
rect 391734 -19142 391936 -19086
rect 391992 -19142 392078 -19086
rect 392134 -19142 392333 -19086
rect 392389 -19142 392475 -19086
rect 392531 -19142 392738 -19086
rect 392794 -19142 392880 -19086
rect 392936 -19142 393138 -19086
rect 393194 -19142 393280 -19086
rect 393336 -19142 393543 -19086
rect 393599 -19142 393685 -19086
rect 393741 -19142 393940 -19086
rect 393996 -19142 394082 -19086
rect 394138 -19142 394337 -19086
rect 394393 -19142 394479 -19086
rect 394535 -19142 394740 -19086
rect 394796 -19142 394882 -19086
rect 394938 -19142 395142 -19086
rect 395198 -19142 395284 -19086
rect 395340 -19142 395545 -19086
rect 395601 -19142 395687 -19086
rect 395743 -19142 395941 -19086
rect 395997 -19142 396083 -19086
rect 396139 -19098 397200 -19086
rect 396139 -19142 396526 -19098
rect 388666 -19154 396526 -19142
rect 396582 -19154 396650 -19098
rect 396706 -19154 396774 -19098
rect 396830 -19154 396898 -19098
rect 396954 -19154 397022 -19098
rect 397078 -19154 397200 -19098
rect 388000 -19222 397200 -19154
rect 388000 -19278 388114 -19222
rect 388170 -19278 388238 -19222
rect 388294 -19278 388362 -19222
rect 388418 -19278 388486 -19222
rect 388542 -19278 388610 -19222
rect 388666 -19228 396526 -19222
rect 388666 -19278 389141 -19228
rect 388000 -19284 389141 -19278
rect 389197 -19284 389283 -19228
rect 389339 -19284 389542 -19228
rect 389598 -19284 389684 -19228
rect 389740 -19284 389942 -19228
rect 389998 -19284 390084 -19228
rect 390140 -19284 390339 -19228
rect 390395 -19284 390481 -19228
rect 390537 -19284 390736 -19228
rect 390792 -19284 390878 -19228
rect 390934 -19284 391140 -19228
rect 391196 -19284 391282 -19228
rect 391338 -19284 391536 -19228
rect 391592 -19284 391678 -19228
rect 391734 -19284 391936 -19228
rect 391992 -19284 392078 -19228
rect 392134 -19284 392333 -19228
rect 392389 -19284 392475 -19228
rect 392531 -19284 392738 -19228
rect 392794 -19284 392880 -19228
rect 392936 -19284 393138 -19228
rect 393194 -19284 393280 -19228
rect 393336 -19284 393543 -19228
rect 393599 -19284 393685 -19228
rect 393741 -19284 393940 -19228
rect 393996 -19284 394082 -19228
rect 394138 -19284 394337 -19228
rect 394393 -19284 394479 -19228
rect 394535 -19284 394740 -19228
rect 394796 -19284 394882 -19228
rect 394938 -19284 395142 -19228
rect 395198 -19284 395284 -19228
rect 395340 -19284 395545 -19228
rect 395601 -19284 395687 -19228
rect 395743 -19284 395941 -19228
rect 395997 -19284 396083 -19228
rect 396139 -19278 396526 -19228
rect 396582 -19278 396650 -19222
rect 396706 -19278 396774 -19222
rect 396830 -19278 396898 -19222
rect 396954 -19278 397022 -19222
rect 397078 -19278 397200 -19222
rect 396139 -19284 397200 -19278
rect 388000 -19346 397200 -19284
rect 388000 -19402 388114 -19346
rect 388170 -19402 388238 -19346
rect 388294 -19402 388362 -19346
rect 388418 -19402 388486 -19346
rect 388542 -19402 388610 -19346
rect 388666 -19370 396526 -19346
rect 388666 -19402 389141 -19370
rect 388000 -19426 389141 -19402
rect 389197 -19426 389283 -19370
rect 389339 -19426 389542 -19370
rect 389598 -19426 389684 -19370
rect 389740 -19426 389942 -19370
rect 389998 -19426 390084 -19370
rect 390140 -19426 390339 -19370
rect 390395 -19426 390481 -19370
rect 390537 -19426 390736 -19370
rect 390792 -19426 390878 -19370
rect 390934 -19426 391140 -19370
rect 391196 -19426 391282 -19370
rect 391338 -19426 391536 -19370
rect 391592 -19426 391678 -19370
rect 391734 -19426 391936 -19370
rect 391992 -19426 392078 -19370
rect 392134 -19426 392333 -19370
rect 392389 -19426 392475 -19370
rect 392531 -19426 392738 -19370
rect 392794 -19426 392880 -19370
rect 392936 -19426 393138 -19370
rect 393194 -19426 393280 -19370
rect 393336 -19426 393543 -19370
rect 393599 -19426 393685 -19370
rect 393741 -19426 393940 -19370
rect 393996 -19426 394082 -19370
rect 394138 -19426 394337 -19370
rect 394393 -19426 394479 -19370
rect 394535 -19426 394740 -19370
rect 394796 -19426 394882 -19370
rect 394938 -19426 395142 -19370
rect 395198 -19426 395284 -19370
rect 395340 -19426 395545 -19370
rect 395601 -19426 395687 -19370
rect 395743 -19426 395941 -19370
rect 395997 -19426 396083 -19370
rect 396139 -19402 396526 -19370
rect 396582 -19402 396650 -19346
rect 396706 -19402 396774 -19346
rect 396830 -19402 396898 -19346
rect 396954 -19402 397022 -19346
rect 397078 -19402 397200 -19346
rect 396139 -19426 397200 -19402
rect 388000 -19470 397200 -19426
rect 388000 -19526 388114 -19470
rect 388170 -19526 388238 -19470
rect 388294 -19526 388362 -19470
rect 388418 -19526 388486 -19470
rect 388542 -19526 388610 -19470
rect 388666 -19512 396526 -19470
rect 388666 -19526 389141 -19512
rect 388000 -19568 389141 -19526
rect 389197 -19568 389283 -19512
rect 389339 -19568 389542 -19512
rect 389598 -19568 389684 -19512
rect 389740 -19568 389942 -19512
rect 389998 -19568 390084 -19512
rect 390140 -19568 390339 -19512
rect 390395 -19568 390481 -19512
rect 390537 -19568 390736 -19512
rect 390792 -19568 390878 -19512
rect 390934 -19568 391140 -19512
rect 391196 -19568 391282 -19512
rect 391338 -19568 391536 -19512
rect 391592 -19568 391678 -19512
rect 391734 -19568 391936 -19512
rect 391992 -19568 392078 -19512
rect 392134 -19568 392333 -19512
rect 392389 -19568 392475 -19512
rect 392531 -19568 392738 -19512
rect 392794 -19568 392880 -19512
rect 392936 -19568 393138 -19512
rect 393194 -19568 393280 -19512
rect 393336 -19568 393543 -19512
rect 393599 -19568 393685 -19512
rect 393741 -19568 393940 -19512
rect 393996 -19568 394082 -19512
rect 394138 -19568 394337 -19512
rect 394393 -19568 394479 -19512
rect 394535 -19568 394740 -19512
rect 394796 -19568 394882 -19512
rect 394938 -19568 395142 -19512
rect 395198 -19568 395284 -19512
rect 395340 -19568 395545 -19512
rect 395601 -19568 395687 -19512
rect 395743 -19568 395941 -19512
rect 395997 -19568 396083 -19512
rect 396139 -19526 396526 -19512
rect 396582 -19526 396650 -19470
rect 396706 -19526 396774 -19470
rect 396830 -19526 396898 -19470
rect 396954 -19526 397022 -19470
rect 397078 -19526 397200 -19470
rect 396139 -19568 397200 -19526
rect 388000 -19594 397200 -19568
rect 388000 -19650 388114 -19594
rect 388170 -19650 388238 -19594
rect 388294 -19650 388362 -19594
rect 388418 -19650 388486 -19594
rect 388542 -19650 388610 -19594
rect 388666 -19650 396526 -19594
rect 396582 -19650 396650 -19594
rect 396706 -19650 396774 -19594
rect 396830 -19650 396898 -19594
rect 396954 -19650 397022 -19594
rect 397078 -19650 397200 -19594
rect 388000 -19654 397200 -19650
rect 388000 -19710 389141 -19654
rect 389197 -19710 389283 -19654
rect 389339 -19710 389542 -19654
rect 389598 -19710 389684 -19654
rect 389740 -19710 389942 -19654
rect 389998 -19710 390084 -19654
rect 390140 -19710 390339 -19654
rect 390395 -19710 390481 -19654
rect 390537 -19710 390736 -19654
rect 390792 -19710 390878 -19654
rect 390934 -19710 391140 -19654
rect 391196 -19710 391282 -19654
rect 391338 -19710 391536 -19654
rect 391592 -19710 391678 -19654
rect 391734 -19710 391936 -19654
rect 391992 -19710 392078 -19654
rect 392134 -19710 392333 -19654
rect 392389 -19710 392475 -19654
rect 392531 -19710 392738 -19654
rect 392794 -19710 392880 -19654
rect 392936 -19710 393138 -19654
rect 393194 -19710 393280 -19654
rect 393336 -19710 393543 -19654
rect 393599 -19710 393685 -19654
rect 393741 -19710 393940 -19654
rect 393996 -19710 394082 -19654
rect 394138 -19710 394337 -19654
rect 394393 -19710 394479 -19654
rect 394535 -19710 394740 -19654
rect 394796 -19710 394882 -19654
rect 394938 -19710 395142 -19654
rect 395198 -19710 395284 -19654
rect 395340 -19710 395545 -19654
rect 395601 -19710 395687 -19654
rect 395743 -19710 395941 -19654
rect 395997 -19710 396083 -19654
rect 396139 -19710 397200 -19654
rect 388000 -19718 397200 -19710
rect 388000 -19774 388114 -19718
rect 388170 -19774 388238 -19718
rect 388294 -19774 388362 -19718
rect 388418 -19774 388486 -19718
rect 388542 -19774 388610 -19718
rect 388666 -19774 396526 -19718
rect 396582 -19774 396650 -19718
rect 396706 -19774 396774 -19718
rect 396830 -19774 396898 -19718
rect 396954 -19774 397022 -19718
rect 397078 -19774 397200 -19718
rect 388000 -19796 397200 -19774
rect 388000 -19842 389141 -19796
rect 388000 -19898 388114 -19842
rect 388170 -19898 388238 -19842
rect 388294 -19898 388362 -19842
rect 388418 -19898 388486 -19842
rect 388542 -19898 388610 -19842
rect 388666 -19852 389141 -19842
rect 389197 -19852 389283 -19796
rect 389339 -19852 389542 -19796
rect 389598 -19852 389684 -19796
rect 389740 -19852 389942 -19796
rect 389998 -19852 390084 -19796
rect 390140 -19852 390339 -19796
rect 390395 -19852 390481 -19796
rect 390537 -19852 390736 -19796
rect 390792 -19852 390878 -19796
rect 390934 -19852 391140 -19796
rect 391196 -19852 391282 -19796
rect 391338 -19852 391536 -19796
rect 391592 -19852 391678 -19796
rect 391734 -19852 391936 -19796
rect 391992 -19852 392078 -19796
rect 392134 -19852 392333 -19796
rect 392389 -19852 392475 -19796
rect 392531 -19852 392738 -19796
rect 392794 -19852 392880 -19796
rect 392936 -19852 393138 -19796
rect 393194 -19852 393280 -19796
rect 393336 -19852 393543 -19796
rect 393599 -19852 393685 -19796
rect 393741 -19852 393940 -19796
rect 393996 -19852 394082 -19796
rect 394138 -19852 394337 -19796
rect 394393 -19852 394479 -19796
rect 394535 -19852 394740 -19796
rect 394796 -19852 394882 -19796
rect 394938 -19852 395142 -19796
rect 395198 -19852 395284 -19796
rect 395340 -19852 395545 -19796
rect 395601 -19852 395687 -19796
rect 395743 -19852 395941 -19796
rect 395997 -19852 396083 -19796
rect 396139 -19842 397200 -19796
rect 396139 -19852 396526 -19842
rect 388666 -19898 396526 -19852
rect 396582 -19898 396650 -19842
rect 396706 -19898 396774 -19842
rect 396830 -19898 396898 -19842
rect 396954 -19898 397022 -19842
rect 397078 -19898 397200 -19842
rect 388000 -19938 397200 -19898
rect 388000 -19966 389141 -19938
rect 388000 -20022 388114 -19966
rect 388170 -20022 388238 -19966
rect 388294 -20022 388362 -19966
rect 388418 -20022 388486 -19966
rect 388542 -20022 388610 -19966
rect 388666 -19994 389141 -19966
rect 389197 -19994 389283 -19938
rect 389339 -19994 389542 -19938
rect 389598 -19994 389684 -19938
rect 389740 -19994 389942 -19938
rect 389998 -19994 390084 -19938
rect 390140 -19994 390339 -19938
rect 390395 -19994 390481 -19938
rect 390537 -19994 390736 -19938
rect 390792 -19994 390878 -19938
rect 390934 -19994 391140 -19938
rect 391196 -19994 391282 -19938
rect 391338 -19994 391536 -19938
rect 391592 -19994 391678 -19938
rect 391734 -19994 391936 -19938
rect 391992 -19994 392078 -19938
rect 392134 -19994 392333 -19938
rect 392389 -19994 392475 -19938
rect 392531 -19994 392738 -19938
rect 392794 -19994 392880 -19938
rect 392936 -19994 393138 -19938
rect 393194 -19994 393280 -19938
rect 393336 -19994 393543 -19938
rect 393599 -19994 393685 -19938
rect 393741 -19994 393940 -19938
rect 393996 -19994 394082 -19938
rect 394138 -19994 394337 -19938
rect 394393 -19994 394479 -19938
rect 394535 -19994 394740 -19938
rect 394796 -19994 394882 -19938
rect 394938 -19994 395142 -19938
rect 395198 -19994 395284 -19938
rect 395340 -19994 395545 -19938
rect 395601 -19994 395687 -19938
rect 395743 -19994 395941 -19938
rect 395997 -19994 396083 -19938
rect 396139 -19966 397200 -19938
rect 396139 -19994 396526 -19966
rect 388666 -20022 396526 -19994
rect 396582 -20022 396650 -19966
rect 396706 -20022 396774 -19966
rect 396830 -20022 396898 -19966
rect 396954 -20022 397022 -19966
rect 397078 -20022 397200 -19966
rect 388000 -20080 397200 -20022
rect 388000 -20090 389141 -20080
rect 388000 -20146 388114 -20090
rect 388170 -20146 388238 -20090
rect 388294 -20146 388362 -20090
rect 388418 -20146 388486 -20090
rect 388542 -20146 388610 -20090
rect 388666 -20136 389141 -20090
rect 389197 -20136 389283 -20080
rect 389339 -20136 389542 -20080
rect 389598 -20136 389684 -20080
rect 389740 -20136 389942 -20080
rect 389998 -20136 390084 -20080
rect 390140 -20136 390339 -20080
rect 390395 -20136 390481 -20080
rect 390537 -20136 390736 -20080
rect 390792 -20136 390878 -20080
rect 390934 -20136 391140 -20080
rect 391196 -20136 391282 -20080
rect 391338 -20136 391536 -20080
rect 391592 -20136 391678 -20080
rect 391734 -20136 391936 -20080
rect 391992 -20136 392078 -20080
rect 392134 -20136 392333 -20080
rect 392389 -20136 392475 -20080
rect 392531 -20136 392738 -20080
rect 392794 -20136 392880 -20080
rect 392936 -20136 393138 -20080
rect 393194 -20136 393280 -20080
rect 393336 -20136 393543 -20080
rect 393599 -20136 393685 -20080
rect 393741 -20136 393940 -20080
rect 393996 -20136 394082 -20080
rect 394138 -20136 394337 -20080
rect 394393 -20136 394479 -20080
rect 394535 -20136 394740 -20080
rect 394796 -20136 394882 -20080
rect 394938 -20136 395142 -20080
rect 395198 -20136 395284 -20080
rect 395340 -20136 395545 -20080
rect 395601 -20136 395687 -20080
rect 395743 -20136 395941 -20080
rect 395997 -20136 396083 -20080
rect 396139 -20090 397200 -20080
rect 396139 -20136 396526 -20090
rect 388666 -20146 396526 -20136
rect 396582 -20146 396650 -20090
rect 396706 -20146 396774 -20090
rect 396830 -20146 396898 -20090
rect 396954 -20146 397022 -20090
rect 397078 -20146 397200 -20090
rect 388000 -20214 397200 -20146
rect 388000 -20270 388114 -20214
rect 388170 -20270 388238 -20214
rect 388294 -20270 388362 -20214
rect 388418 -20270 388486 -20214
rect 388542 -20270 388610 -20214
rect 388666 -20222 396526 -20214
rect 388666 -20270 389141 -20222
rect 388000 -20278 389141 -20270
rect 389197 -20278 389283 -20222
rect 389339 -20278 389542 -20222
rect 389598 -20278 389684 -20222
rect 389740 -20278 389942 -20222
rect 389998 -20278 390084 -20222
rect 390140 -20278 390339 -20222
rect 390395 -20278 390481 -20222
rect 390537 -20278 390736 -20222
rect 390792 -20278 390878 -20222
rect 390934 -20278 391140 -20222
rect 391196 -20278 391282 -20222
rect 391338 -20278 391536 -20222
rect 391592 -20278 391678 -20222
rect 391734 -20278 391936 -20222
rect 391992 -20278 392078 -20222
rect 392134 -20278 392333 -20222
rect 392389 -20278 392475 -20222
rect 392531 -20278 392738 -20222
rect 392794 -20278 392880 -20222
rect 392936 -20278 393138 -20222
rect 393194 -20278 393280 -20222
rect 393336 -20278 393543 -20222
rect 393599 -20278 393685 -20222
rect 393741 -20278 393940 -20222
rect 393996 -20278 394082 -20222
rect 394138 -20278 394337 -20222
rect 394393 -20278 394479 -20222
rect 394535 -20278 394740 -20222
rect 394796 -20278 394882 -20222
rect 394938 -20278 395142 -20222
rect 395198 -20278 395284 -20222
rect 395340 -20278 395545 -20222
rect 395601 -20278 395687 -20222
rect 395743 -20278 395941 -20222
rect 395997 -20278 396083 -20222
rect 396139 -20270 396526 -20222
rect 396582 -20270 396650 -20214
rect 396706 -20270 396774 -20214
rect 396830 -20270 396898 -20214
rect 396954 -20270 397022 -20214
rect 397078 -20270 397200 -20214
rect 396139 -20278 397200 -20270
rect 388000 -20338 397200 -20278
rect 388000 -20394 388114 -20338
rect 388170 -20394 388238 -20338
rect 388294 -20394 388362 -20338
rect 388418 -20394 388486 -20338
rect 388542 -20394 388610 -20338
rect 388666 -20364 396526 -20338
rect 388666 -20394 389141 -20364
rect 388000 -20420 389141 -20394
rect 389197 -20420 389283 -20364
rect 389339 -20420 389542 -20364
rect 389598 -20420 389684 -20364
rect 389740 -20420 389942 -20364
rect 389998 -20420 390084 -20364
rect 390140 -20420 390339 -20364
rect 390395 -20420 390481 -20364
rect 390537 -20420 390736 -20364
rect 390792 -20420 390878 -20364
rect 390934 -20420 391140 -20364
rect 391196 -20420 391282 -20364
rect 391338 -20420 391536 -20364
rect 391592 -20420 391678 -20364
rect 391734 -20420 391936 -20364
rect 391992 -20420 392078 -20364
rect 392134 -20420 392333 -20364
rect 392389 -20420 392475 -20364
rect 392531 -20420 392738 -20364
rect 392794 -20420 392880 -20364
rect 392936 -20420 393138 -20364
rect 393194 -20420 393280 -20364
rect 393336 -20420 393543 -20364
rect 393599 -20420 393685 -20364
rect 393741 -20420 393940 -20364
rect 393996 -20420 394082 -20364
rect 394138 -20420 394337 -20364
rect 394393 -20420 394479 -20364
rect 394535 -20420 394740 -20364
rect 394796 -20420 394882 -20364
rect 394938 -20420 395142 -20364
rect 395198 -20420 395284 -20364
rect 395340 -20420 395545 -20364
rect 395601 -20420 395687 -20364
rect 395743 -20420 395941 -20364
rect 395997 -20420 396083 -20364
rect 396139 -20394 396526 -20364
rect 396582 -20394 396650 -20338
rect 396706 -20394 396774 -20338
rect 396830 -20394 396898 -20338
rect 396954 -20394 397022 -20338
rect 397078 -20394 397200 -20338
rect 396139 -20420 397200 -20394
rect 388000 -20462 397200 -20420
rect 388000 -20518 388114 -20462
rect 388170 -20518 388238 -20462
rect 388294 -20518 388362 -20462
rect 388418 -20518 388486 -20462
rect 388542 -20518 388610 -20462
rect 388666 -20506 396526 -20462
rect 388666 -20518 389141 -20506
rect 388000 -20562 389141 -20518
rect 389197 -20562 389283 -20506
rect 389339 -20562 389542 -20506
rect 389598 -20562 389684 -20506
rect 389740 -20562 389942 -20506
rect 389998 -20562 390084 -20506
rect 390140 -20562 390339 -20506
rect 390395 -20562 390481 -20506
rect 390537 -20562 390736 -20506
rect 390792 -20562 390878 -20506
rect 390934 -20562 391140 -20506
rect 391196 -20562 391282 -20506
rect 391338 -20562 391536 -20506
rect 391592 -20562 391678 -20506
rect 391734 -20562 391936 -20506
rect 391992 -20562 392078 -20506
rect 392134 -20562 392333 -20506
rect 392389 -20562 392475 -20506
rect 392531 -20562 392738 -20506
rect 392794 -20562 392880 -20506
rect 392936 -20562 393138 -20506
rect 393194 -20562 393280 -20506
rect 393336 -20562 393543 -20506
rect 393599 -20562 393685 -20506
rect 393741 -20562 393940 -20506
rect 393996 -20562 394082 -20506
rect 394138 -20562 394337 -20506
rect 394393 -20562 394479 -20506
rect 394535 -20562 394740 -20506
rect 394796 -20562 394882 -20506
rect 394938 -20562 395142 -20506
rect 395198 -20562 395284 -20506
rect 395340 -20562 395545 -20506
rect 395601 -20562 395687 -20506
rect 395743 -20562 395941 -20506
rect 395997 -20562 396083 -20506
rect 396139 -20518 396526 -20506
rect 396582 -20518 396650 -20462
rect 396706 -20518 396774 -20462
rect 396830 -20518 396898 -20462
rect 396954 -20518 397022 -20462
rect 397078 -20518 397200 -20462
rect 396139 -20562 397200 -20518
rect 388000 -20586 397200 -20562
rect 388000 -20642 388114 -20586
rect 388170 -20642 388238 -20586
rect 388294 -20642 388362 -20586
rect 388418 -20642 388486 -20586
rect 388542 -20642 388610 -20586
rect 388666 -20642 396526 -20586
rect 396582 -20642 396650 -20586
rect 396706 -20642 396774 -20586
rect 396830 -20642 396898 -20586
rect 396954 -20642 397022 -20586
rect 397078 -20642 397200 -20586
rect 388000 -20648 397200 -20642
rect 388000 -20704 389141 -20648
rect 389197 -20704 389283 -20648
rect 389339 -20704 389542 -20648
rect 389598 -20704 389684 -20648
rect 389740 -20704 389942 -20648
rect 389998 -20704 390084 -20648
rect 390140 -20704 390339 -20648
rect 390395 -20704 390481 -20648
rect 390537 -20704 390736 -20648
rect 390792 -20704 390878 -20648
rect 390934 -20704 391140 -20648
rect 391196 -20704 391282 -20648
rect 391338 -20704 391536 -20648
rect 391592 -20704 391678 -20648
rect 391734 -20704 391936 -20648
rect 391992 -20704 392078 -20648
rect 392134 -20704 392333 -20648
rect 392389 -20704 392475 -20648
rect 392531 -20704 392738 -20648
rect 392794 -20704 392880 -20648
rect 392936 -20704 393138 -20648
rect 393194 -20704 393280 -20648
rect 393336 -20704 393543 -20648
rect 393599 -20704 393685 -20648
rect 393741 -20704 393940 -20648
rect 393996 -20704 394082 -20648
rect 394138 -20704 394337 -20648
rect 394393 -20704 394479 -20648
rect 394535 -20704 394740 -20648
rect 394796 -20704 394882 -20648
rect 394938 -20704 395142 -20648
rect 395198 -20704 395284 -20648
rect 395340 -20704 395545 -20648
rect 395601 -20704 395687 -20648
rect 395743 -20704 395941 -20648
rect 395997 -20704 396083 -20648
rect 396139 -20704 397200 -20648
rect 388000 -20710 397200 -20704
rect 388000 -20766 388114 -20710
rect 388170 -20766 388238 -20710
rect 388294 -20766 388362 -20710
rect 388418 -20766 388486 -20710
rect 388542 -20766 388610 -20710
rect 388666 -20766 396526 -20710
rect 396582 -20766 396650 -20710
rect 396706 -20766 396774 -20710
rect 396830 -20766 396898 -20710
rect 396954 -20766 397022 -20710
rect 397078 -20766 397200 -20710
rect 388000 -20790 397200 -20766
rect 388000 -20834 389141 -20790
rect 388000 -20890 388114 -20834
rect 388170 -20890 388238 -20834
rect 388294 -20890 388362 -20834
rect 388418 -20890 388486 -20834
rect 388542 -20890 388610 -20834
rect 388666 -20846 389141 -20834
rect 389197 -20846 389283 -20790
rect 389339 -20846 389542 -20790
rect 389598 -20846 389684 -20790
rect 389740 -20846 389942 -20790
rect 389998 -20846 390084 -20790
rect 390140 -20846 390339 -20790
rect 390395 -20846 390481 -20790
rect 390537 -20846 390736 -20790
rect 390792 -20846 390878 -20790
rect 390934 -20846 391140 -20790
rect 391196 -20846 391282 -20790
rect 391338 -20846 391536 -20790
rect 391592 -20846 391678 -20790
rect 391734 -20846 391936 -20790
rect 391992 -20846 392078 -20790
rect 392134 -20846 392333 -20790
rect 392389 -20846 392475 -20790
rect 392531 -20846 392738 -20790
rect 392794 -20846 392880 -20790
rect 392936 -20846 393138 -20790
rect 393194 -20846 393280 -20790
rect 393336 -20846 393543 -20790
rect 393599 -20846 393685 -20790
rect 393741 -20846 393940 -20790
rect 393996 -20846 394082 -20790
rect 394138 -20846 394337 -20790
rect 394393 -20846 394479 -20790
rect 394535 -20846 394740 -20790
rect 394796 -20846 394882 -20790
rect 394938 -20846 395142 -20790
rect 395198 -20846 395284 -20790
rect 395340 -20846 395545 -20790
rect 395601 -20846 395687 -20790
rect 395743 -20846 395941 -20790
rect 395997 -20846 396083 -20790
rect 396139 -20834 397200 -20790
rect 396139 -20846 396526 -20834
rect 388666 -20890 396526 -20846
rect 396582 -20890 396650 -20834
rect 396706 -20890 396774 -20834
rect 396830 -20890 396898 -20834
rect 396954 -20890 397022 -20834
rect 397078 -20890 397200 -20834
rect 388000 -20932 397200 -20890
rect 388000 -20958 389141 -20932
rect 388000 -21014 388114 -20958
rect 388170 -21014 388238 -20958
rect 388294 -21014 388362 -20958
rect 388418 -21014 388486 -20958
rect 388542 -21014 388610 -20958
rect 388666 -20988 389141 -20958
rect 389197 -20988 389283 -20932
rect 389339 -20988 389542 -20932
rect 389598 -20988 389684 -20932
rect 389740 -20988 389942 -20932
rect 389998 -20988 390084 -20932
rect 390140 -20988 390339 -20932
rect 390395 -20988 390481 -20932
rect 390537 -20988 390736 -20932
rect 390792 -20988 390878 -20932
rect 390934 -20988 391140 -20932
rect 391196 -20988 391282 -20932
rect 391338 -20988 391536 -20932
rect 391592 -20988 391678 -20932
rect 391734 -20988 391936 -20932
rect 391992 -20988 392078 -20932
rect 392134 -20988 392333 -20932
rect 392389 -20988 392475 -20932
rect 392531 -20988 392738 -20932
rect 392794 -20988 392880 -20932
rect 392936 -20988 393138 -20932
rect 393194 -20988 393280 -20932
rect 393336 -20988 393543 -20932
rect 393599 -20988 393685 -20932
rect 393741 -20988 393940 -20932
rect 393996 -20988 394082 -20932
rect 394138 -20988 394337 -20932
rect 394393 -20988 394479 -20932
rect 394535 -20988 394740 -20932
rect 394796 -20988 394882 -20932
rect 394938 -20988 395142 -20932
rect 395198 -20988 395284 -20932
rect 395340 -20988 395545 -20932
rect 395601 -20988 395687 -20932
rect 395743 -20988 395941 -20932
rect 395997 -20988 396083 -20932
rect 396139 -20958 397200 -20932
rect 396139 -20988 396526 -20958
rect 388666 -21014 396526 -20988
rect 396582 -21014 396650 -20958
rect 396706 -21014 396774 -20958
rect 396830 -21014 396898 -20958
rect 396954 -21014 397022 -20958
rect 397078 -21014 397200 -20958
rect 388000 -21074 397200 -21014
rect 388000 -21082 389141 -21074
rect 388000 -21138 388114 -21082
rect 388170 -21138 388238 -21082
rect 388294 -21138 388362 -21082
rect 388418 -21138 388486 -21082
rect 388542 -21138 388610 -21082
rect 388666 -21130 389141 -21082
rect 389197 -21130 389283 -21074
rect 389339 -21130 389542 -21074
rect 389598 -21130 389684 -21074
rect 389740 -21130 389942 -21074
rect 389998 -21130 390084 -21074
rect 390140 -21130 390339 -21074
rect 390395 -21130 390481 -21074
rect 390537 -21130 390736 -21074
rect 390792 -21130 390878 -21074
rect 390934 -21130 391140 -21074
rect 391196 -21130 391282 -21074
rect 391338 -21130 391536 -21074
rect 391592 -21130 391678 -21074
rect 391734 -21130 391936 -21074
rect 391992 -21130 392078 -21074
rect 392134 -21130 392333 -21074
rect 392389 -21130 392475 -21074
rect 392531 -21130 392738 -21074
rect 392794 -21130 392880 -21074
rect 392936 -21130 393138 -21074
rect 393194 -21130 393280 -21074
rect 393336 -21130 393543 -21074
rect 393599 -21130 393685 -21074
rect 393741 -21130 393940 -21074
rect 393996 -21130 394082 -21074
rect 394138 -21130 394337 -21074
rect 394393 -21130 394479 -21074
rect 394535 -21130 394740 -21074
rect 394796 -21130 394882 -21074
rect 394938 -21130 395142 -21074
rect 395198 -21130 395284 -21074
rect 395340 -21130 395545 -21074
rect 395601 -21130 395687 -21074
rect 395743 -21130 395941 -21074
rect 395997 -21130 396083 -21074
rect 396139 -21082 397200 -21074
rect 396139 -21130 396526 -21082
rect 388666 -21138 396526 -21130
rect 396582 -21138 396650 -21082
rect 396706 -21138 396774 -21082
rect 396830 -21138 396898 -21082
rect 396954 -21138 397022 -21082
rect 397078 -21138 397200 -21082
rect 388000 -21206 397200 -21138
rect 388000 -21262 388114 -21206
rect 388170 -21262 388238 -21206
rect 388294 -21262 388362 -21206
rect 388418 -21262 388486 -21206
rect 388542 -21262 388610 -21206
rect 388666 -21216 396526 -21206
rect 388666 -21262 389141 -21216
rect 388000 -21272 389141 -21262
rect 389197 -21272 389283 -21216
rect 389339 -21272 389542 -21216
rect 389598 -21272 389684 -21216
rect 389740 -21272 389942 -21216
rect 389998 -21272 390084 -21216
rect 390140 -21272 390339 -21216
rect 390395 -21272 390481 -21216
rect 390537 -21272 390736 -21216
rect 390792 -21272 390878 -21216
rect 390934 -21272 391140 -21216
rect 391196 -21272 391282 -21216
rect 391338 -21272 391536 -21216
rect 391592 -21272 391678 -21216
rect 391734 -21272 391936 -21216
rect 391992 -21272 392078 -21216
rect 392134 -21272 392333 -21216
rect 392389 -21272 392475 -21216
rect 392531 -21272 392738 -21216
rect 392794 -21272 392880 -21216
rect 392936 -21272 393138 -21216
rect 393194 -21272 393280 -21216
rect 393336 -21272 393543 -21216
rect 393599 -21272 393685 -21216
rect 393741 -21272 393940 -21216
rect 393996 -21272 394082 -21216
rect 394138 -21272 394337 -21216
rect 394393 -21272 394479 -21216
rect 394535 -21272 394740 -21216
rect 394796 -21272 394882 -21216
rect 394938 -21272 395142 -21216
rect 395198 -21272 395284 -21216
rect 395340 -21272 395545 -21216
rect 395601 -21272 395687 -21216
rect 395743 -21272 395941 -21216
rect 395997 -21272 396083 -21216
rect 396139 -21262 396526 -21216
rect 396582 -21262 396650 -21206
rect 396706 -21262 396774 -21206
rect 396830 -21262 396898 -21206
rect 396954 -21262 397022 -21206
rect 397078 -21262 397200 -21206
rect 396139 -21272 397200 -21262
rect 388000 -21330 397200 -21272
rect 388000 -21386 388114 -21330
rect 388170 -21386 388238 -21330
rect 388294 -21386 388362 -21330
rect 388418 -21386 388486 -21330
rect 388542 -21386 388610 -21330
rect 388666 -21358 396526 -21330
rect 388666 -21386 389141 -21358
rect 388000 -21414 389141 -21386
rect 389197 -21414 389283 -21358
rect 389339 -21414 389542 -21358
rect 389598 -21414 389684 -21358
rect 389740 -21414 389942 -21358
rect 389998 -21414 390084 -21358
rect 390140 -21414 390339 -21358
rect 390395 -21414 390481 -21358
rect 390537 -21414 390736 -21358
rect 390792 -21414 390878 -21358
rect 390934 -21414 391140 -21358
rect 391196 -21414 391282 -21358
rect 391338 -21414 391536 -21358
rect 391592 -21414 391678 -21358
rect 391734 -21414 391936 -21358
rect 391992 -21414 392078 -21358
rect 392134 -21414 392333 -21358
rect 392389 -21414 392475 -21358
rect 392531 -21414 392738 -21358
rect 392794 -21414 392880 -21358
rect 392936 -21414 393138 -21358
rect 393194 -21414 393280 -21358
rect 393336 -21414 393543 -21358
rect 393599 -21414 393685 -21358
rect 393741 -21414 393940 -21358
rect 393996 -21414 394082 -21358
rect 394138 -21414 394337 -21358
rect 394393 -21414 394479 -21358
rect 394535 -21414 394740 -21358
rect 394796 -21414 394882 -21358
rect 394938 -21414 395142 -21358
rect 395198 -21414 395284 -21358
rect 395340 -21414 395545 -21358
rect 395601 -21414 395687 -21358
rect 395743 -21414 395941 -21358
rect 395997 -21414 396083 -21358
rect 396139 -21386 396526 -21358
rect 396582 -21386 396650 -21330
rect 396706 -21386 396774 -21330
rect 396830 -21386 396898 -21330
rect 396954 -21386 397022 -21330
rect 397078 -21386 397200 -21330
rect 396139 -21414 397200 -21386
rect 388000 -21454 397200 -21414
rect 388000 -21510 388114 -21454
rect 388170 -21510 388238 -21454
rect 388294 -21510 388362 -21454
rect 388418 -21510 388486 -21454
rect 388542 -21510 388610 -21454
rect 388666 -21500 396526 -21454
rect 388666 -21510 389141 -21500
rect 388000 -21556 389141 -21510
rect 389197 -21556 389283 -21500
rect 389339 -21556 389542 -21500
rect 389598 -21556 389684 -21500
rect 389740 -21556 389942 -21500
rect 389998 -21556 390084 -21500
rect 390140 -21556 390339 -21500
rect 390395 -21556 390481 -21500
rect 390537 -21556 390736 -21500
rect 390792 -21556 390878 -21500
rect 390934 -21556 391140 -21500
rect 391196 -21556 391282 -21500
rect 391338 -21556 391536 -21500
rect 391592 -21556 391678 -21500
rect 391734 -21556 391936 -21500
rect 391992 -21556 392078 -21500
rect 392134 -21556 392333 -21500
rect 392389 -21556 392475 -21500
rect 392531 -21556 392738 -21500
rect 392794 -21556 392880 -21500
rect 392936 -21556 393138 -21500
rect 393194 -21556 393280 -21500
rect 393336 -21556 393543 -21500
rect 393599 -21556 393685 -21500
rect 393741 -21556 393940 -21500
rect 393996 -21556 394082 -21500
rect 394138 -21556 394337 -21500
rect 394393 -21556 394479 -21500
rect 394535 -21556 394740 -21500
rect 394796 -21556 394882 -21500
rect 394938 -21556 395142 -21500
rect 395198 -21556 395284 -21500
rect 395340 -21556 395545 -21500
rect 395601 -21556 395687 -21500
rect 395743 -21556 395941 -21500
rect 395997 -21556 396083 -21500
rect 396139 -21510 396526 -21500
rect 396582 -21510 396650 -21454
rect 396706 -21510 396774 -21454
rect 396830 -21510 396898 -21454
rect 396954 -21510 397022 -21454
rect 397078 -21510 397200 -21454
rect 396139 -21556 397200 -21510
rect 388000 -21578 397200 -21556
rect 388000 -21634 388114 -21578
rect 388170 -21634 388238 -21578
rect 388294 -21634 388362 -21578
rect 388418 -21634 388486 -21578
rect 388542 -21634 388610 -21578
rect 388666 -21634 396526 -21578
rect 396582 -21634 396650 -21578
rect 396706 -21634 396774 -21578
rect 396830 -21634 396898 -21578
rect 396954 -21634 397022 -21578
rect 397078 -21634 397200 -21578
rect 388000 -21642 397200 -21634
rect 388000 -21698 389141 -21642
rect 389197 -21698 389283 -21642
rect 389339 -21698 389542 -21642
rect 389598 -21698 389684 -21642
rect 389740 -21698 389942 -21642
rect 389998 -21698 390084 -21642
rect 390140 -21698 390339 -21642
rect 390395 -21698 390481 -21642
rect 390537 -21698 390736 -21642
rect 390792 -21698 390878 -21642
rect 390934 -21698 391140 -21642
rect 391196 -21698 391282 -21642
rect 391338 -21698 391536 -21642
rect 391592 -21698 391678 -21642
rect 391734 -21698 391936 -21642
rect 391992 -21698 392078 -21642
rect 392134 -21698 392333 -21642
rect 392389 -21698 392475 -21642
rect 392531 -21698 392738 -21642
rect 392794 -21698 392880 -21642
rect 392936 -21698 393138 -21642
rect 393194 -21698 393280 -21642
rect 393336 -21698 393543 -21642
rect 393599 -21698 393685 -21642
rect 393741 -21698 393940 -21642
rect 393996 -21698 394082 -21642
rect 394138 -21698 394337 -21642
rect 394393 -21698 394479 -21642
rect 394535 -21698 394740 -21642
rect 394796 -21698 394882 -21642
rect 394938 -21698 395142 -21642
rect 395198 -21698 395284 -21642
rect 395340 -21698 395545 -21642
rect 395601 -21698 395687 -21642
rect 395743 -21698 395941 -21642
rect 395997 -21698 396083 -21642
rect 396139 -21698 397200 -21642
rect 388000 -21702 397200 -21698
rect 388000 -21758 388114 -21702
rect 388170 -21758 388238 -21702
rect 388294 -21758 388362 -21702
rect 388418 -21758 388486 -21702
rect 388542 -21758 388610 -21702
rect 388666 -21758 396526 -21702
rect 396582 -21758 396650 -21702
rect 396706 -21758 396774 -21702
rect 396830 -21758 396898 -21702
rect 396954 -21758 397022 -21702
rect 397078 -21758 397200 -21702
rect 388000 -21784 397200 -21758
rect 388000 -21826 389141 -21784
rect 388000 -21882 388114 -21826
rect 388170 -21882 388238 -21826
rect 388294 -21882 388362 -21826
rect 388418 -21882 388486 -21826
rect 388542 -21882 388610 -21826
rect 388666 -21840 389141 -21826
rect 389197 -21840 389283 -21784
rect 389339 -21840 389542 -21784
rect 389598 -21840 389684 -21784
rect 389740 -21840 389942 -21784
rect 389998 -21840 390084 -21784
rect 390140 -21840 390339 -21784
rect 390395 -21840 390481 -21784
rect 390537 -21840 390736 -21784
rect 390792 -21840 390878 -21784
rect 390934 -21840 391140 -21784
rect 391196 -21840 391282 -21784
rect 391338 -21840 391536 -21784
rect 391592 -21840 391678 -21784
rect 391734 -21840 391936 -21784
rect 391992 -21840 392078 -21784
rect 392134 -21840 392333 -21784
rect 392389 -21840 392475 -21784
rect 392531 -21840 392738 -21784
rect 392794 -21840 392880 -21784
rect 392936 -21840 393138 -21784
rect 393194 -21840 393280 -21784
rect 393336 -21840 393543 -21784
rect 393599 -21840 393685 -21784
rect 393741 -21840 393940 -21784
rect 393996 -21840 394082 -21784
rect 394138 -21840 394337 -21784
rect 394393 -21840 394479 -21784
rect 394535 -21840 394740 -21784
rect 394796 -21840 394882 -21784
rect 394938 -21840 395142 -21784
rect 395198 -21840 395284 -21784
rect 395340 -21840 395545 -21784
rect 395601 -21840 395687 -21784
rect 395743 -21840 395941 -21784
rect 395997 -21840 396083 -21784
rect 396139 -21826 397200 -21784
rect 396139 -21840 396526 -21826
rect 388666 -21882 396526 -21840
rect 396582 -21882 396650 -21826
rect 396706 -21882 396774 -21826
rect 396830 -21882 396898 -21826
rect 396954 -21882 397022 -21826
rect 397078 -21882 397200 -21826
rect 388000 -21926 397200 -21882
rect 388000 -21950 389141 -21926
rect 388000 -22006 388114 -21950
rect 388170 -22006 388238 -21950
rect 388294 -22006 388362 -21950
rect 388418 -22006 388486 -21950
rect 388542 -22006 388610 -21950
rect 388666 -21982 389141 -21950
rect 389197 -21982 389283 -21926
rect 389339 -21982 389542 -21926
rect 389598 -21982 389684 -21926
rect 389740 -21982 389942 -21926
rect 389998 -21982 390084 -21926
rect 390140 -21982 390339 -21926
rect 390395 -21982 390481 -21926
rect 390537 -21982 390736 -21926
rect 390792 -21982 390878 -21926
rect 390934 -21982 391140 -21926
rect 391196 -21982 391282 -21926
rect 391338 -21982 391536 -21926
rect 391592 -21982 391678 -21926
rect 391734 -21982 391936 -21926
rect 391992 -21982 392078 -21926
rect 392134 -21982 392333 -21926
rect 392389 -21982 392475 -21926
rect 392531 -21982 392738 -21926
rect 392794 -21982 392880 -21926
rect 392936 -21982 393138 -21926
rect 393194 -21982 393280 -21926
rect 393336 -21982 393543 -21926
rect 393599 -21982 393685 -21926
rect 393741 -21982 393940 -21926
rect 393996 -21982 394082 -21926
rect 394138 -21982 394337 -21926
rect 394393 -21982 394479 -21926
rect 394535 -21982 394740 -21926
rect 394796 -21982 394882 -21926
rect 394938 -21982 395142 -21926
rect 395198 -21982 395284 -21926
rect 395340 -21982 395545 -21926
rect 395601 -21982 395687 -21926
rect 395743 -21982 395941 -21926
rect 395997 -21982 396083 -21926
rect 396139 -21950 397200 -21926
rect 396139 -21982 396526 -21950
rect 388666 -22006 396526 -21982
rect 396582 -22006 396650 -21950
rect 396706 -22006 396774 -21950
rect 396830 -22006 396898 -21950
rect 396954 -22006 397022 -21950
rect 397078 -22006 397200 -21950
rect 388000 -22068 397200 -22006
rect 388000 -22074 389141 -22068
rect 388000 -22130 388114 -22074
rect 388170 -22130 388238 -22074
rect 388294 -22130 388362 -22074
rect 388418 -22130 388486 -22074
rect 388542 -22130 388610 -22074
rect 388666 -22124 389141 -22074
rect 389197 -22124 389283 -22068
rect 389339 -22124 389542 -22068
rect 389598 -22124 389684 -22068
rect 389740 -22124 389942 -22068
rect 389998 -22124 390084 -22068
rect 390140 -22124 390339 -22068
rect 390395 -22124 390481 -22068
rect 390537 -22124 390736 -22068
rect 390792 -22124 390878 -22068
rect 390934 -22124 391140 -22068
rect 391196 -22124 391282 -22068
rect 391338 -22124 391536 -22068
rect 391592 -22124 391678 -22068
rect 391734 -22124 391936 -22068
rect 391992 -22124 392078 -22068
rect 392134 -22124 392333 -22068
rect 392389 -22124 392475 -22068
rect 392531 -22124 392738 -22068
rect 392794 -22124 392880 -22068
rect 392936 -22124 393138 -22068
rect 393194 -22124 393280 -22068
rect 393336 -22124 393543 -22068
rect 393599 -22124 393685 -22068
rect 393741 -22124 393940 -22068
rect 393996 -22124 394082 -22068
rect 394138 -22124 394337 -22068
rect 394393 -22124 394479 -22068
rect 394535 -22124 394740 -22068
rect 394796 -22124 394882 -22068
rect 394938 -22124 395142 -22068
rect 395198 -22124 395284 -22068
rect 395340 -22124 395545 -22068
rect 395601 -22124 395687 -22068
rect 395743 -22124 395941 -22068
rect 395997 -22124 396083 -22068
rect 396139 -22074 397200 -22068
rect 396139 -22124 396526 -22074
rect 388666 -22130 396526 -22124
rect 396582 -22130 396650 -22074
rect 396706 -22130 396774 -22074
rect 396830 -22130 396898 -22074
rect 396954 -22130 397022 -22074
rect 397078 -22130 397200 -22074
rect 388000 -22198 397200 -22130
rect 388000 -22254 388114 -22198
rect 388170 -22254 388238 -22198
rect 388294 -22254 388362 -22198
rect 388418 -22254 388486 -22198
rect 388542 -22254 388610 -22198
rect 388666 -22210 396526 -22198
rect 388666 -22254 389141 -22210
rect 388000 -22266 389141 -22254
rect 389197 -22266 389283 -22210
rect 389339 -22266 389542 -22210
rect 389598 -22266 389684 -22210
rect 389740 -22266 389942 -22210
rect 389998 -22266 390084 -22210
rect 390140 -22266 390339 -22210
rect 390395 -22266 390481 -22210
rect 390537 -22266 390736 -22210
rect 390792 -22266 390878 -22210
rect 390934 -22266 391140 -22210
rect 391196 -22266 391282 -22210
rect 391338 -22266 391536 -22210
rect 391592 -22266 391678 -22210
rect 391734 -22266 391936 -22210
rect 391992 -22266 392078 -22210
rect 392134 -22266 392333 -22210
rect 392389 -22266 392475 -22210
rect 392531 -22266 392738 -22210
rect 392794 -22266 392880 -22210
rect 392936 -22266 393138 -22210
rect 393194 -22266 393280 -22210
rect 393336 -22266 393543 -22210
rect 393599 -22266 393685 -22210
rect 393741 -22266 393940 -22210
rect 393996 -22266 394082 -22210
rect 394138 -22266 394337 -22210
rect 394393 -22266 394479 -22210
rect 394535 -22266 394740 -22210
rect 394796 -22266 394882 -22210
rect 394938 -22266 395142 -22210
rect 395198 -22266 395284 -22210
rect 395340 -22266 395545 -22210
rect 395601 -22266 395687 -22210
rect 395743 -22266 395941 -22210
rect 395997 -22266 396083 -22210
rect 396139 -22254 396526 -22210
rect 396582 -22254 396650 -22198
rect 396706 -22254 396774 -22198
rect 396830 -22254 396898 -22198
rect 396954 -22254 397022 -22198
rect 397078 -22254 397200 -22198
rect 396139 -22266 397200 -22254
rect 388000 -22322 397200 -22266
rect 388000 -22378 388114 -22322
rect 388170 -22378 388238 -22322
rect 388294 -22378 388362 -22322
rect 388418 -22378 388486 -22322
rect 388542 -22378 388610 -22322
rect 388666 -22352 396526 -22322
rect 388666 -22378 389141 -22352
rect 388000 -22408 389141 -22378
rect 389197 -22408 389283 -22352
rect 389339 -22408 389542 -22352
rect 389598 -22408 389684 -22352
rect 389740 -22408 389942 -22352
rect 389998 -22408 390084 -22352
rect 390140 -22408 390339 -22352
rect 390395 -22408 390481 -22352
rect 390537 -22408 390736 -22352
rect 390792 -22408 390878 -22352
rect 390934 -22408 391140 -22352
rect 391196 -22408 391282 -22352
rect 391338 -22408 391536 -22352
rect 391592 -22408 391678 -22352
rect 391734 -22408 391936 -22352
rect 391992 -22408 392078 -22352
rect 392134 -22408 392333 -22352
rect 392389 -22408 392475 -22352
rect 392531 -22408 392738 -22352
rect 392794 -22408 392880 -22352
rect 392936 -22408 393138 -22352
rect 393194 -22408 393280 -22352
rect 393336 -22408 393543 -22352
rect 393599 -22408 393685 -22352
rect 393741 -22408 393940 -22352
rect 393996 -22408 394082 -22352
rect 394138 -22408 394337 -22352
rect 394393 -22408 394479 -22352
rect 394535 -22408 394740 -22352
rect 394796 -22408 394882 -22352
rect 394938 -22408 395142 -22352
rect 395198 -22408 395284 -22352
rect 395340 -22408 395545 -22352
rect 395601 -22408 395687 -22352
rect 395743 -22408 395941 -22352
rect 395997 -22408 396083 -22352
rect 396139 -22378 396526 -22352
rect 396582 -22378 396650 -22322
rect 396706 -22378 396774 -22322
rect 396830 -22378 396898 -22322
rect 396954 -22378 397022 -22322
rect 397078 -22378 397200 -22322
rect 396139 -22408 397200 -22378
rect 388000 -22446 397200 -22408
rect 388000 -22502 388114 -22446
rect 388170 -22502 388238 -22446
rect 388294 -22502 388362 -22446
rect 388418 -22502 388486 -22446
rect 388542 -22502 388610 -22446
rect 388666 -22494 396526 -22446
rect 388666 -22502 389141 -22494
rect 388000 -22550 389141 -22502
rect 389197 -22550 389283 -22494
rect 389339 -22550 389542 -22494
rect 389598 -22550 389684 -22494
rect 389740 -22550 389942 -22494
rect 389998 -22550 390084 -22494
rect 390140 -22550 390339 -22494
rect 390395 -22550 390481 -22494
rect 390537 -22550 390736 -22494
rect 390792 -22550 390878 -22494
rect 390934 -22550 391140 -22494
rect 391196 -22550 391282 -22494
rect 391338 -22550 391536 -22494
rect 391592 -22550 391678 -22494
rect 391734 -22550 391936 -22494
rect 391992 -22550 392078 -22494
rect 392134 -22550 392333 -22494
rect 392389 -22550 392475 -22494
rect 392531 -22550 392738 -22494
rect 392794 -22550 392880 -22494
rect 392936 -22550 393138 -22494
rect 393194 -22550 393280 -22494
rect 393336 -22550 393543 -22494
rect 393599 -22550 393685 -22494
rect 393741 -22550 393940 -22494
rect 393996 -22550 394082 -22494
rect 394138 -22550 394337 -22494
rect 394393 -22550 394479 -22494
rect 394535 -22550 394740 -22494
rect 394796 -22550 394882 -22494
rect 394938 -22550 395142 -22494
rect 395198 -22550 395284 -22494
rect 395340 -22550 395545 -22494
rect 395601 -22550 395687 -22494
rect 395743 -22550 395941 -22494
rect 395997 -22550 396083 -22494
rect 396139 -22502 396526 -22494
rect 396582 -22502 396650 -22446
rect 396706 -22502 396774 -22446
rect 396830 -22502 396898 -22446
rect 396954 -22502 397022 -22446
rect 397078 -22502 397200 -22446
rect 396139 -22550 397200 -22502
rect 388000 -22570 397200 -22550
rect 388000 -22626 388114 -22570
rect 388170 -22626 388238 -22570
rect 388294 -22626 388362 -22570
rect 388418 -22626 388486 -22570
rect 388542 -22626 388610 -22570
rect 388666 -22626 396526 -22570
rect 396582 -22626 396650 -22570
rect 396706 -22626 396774 -22570
rect 396830 -22626 396898 -22570
rect 396954 -22626 397022 -22570
rect 397078 -22626 397200 -22570
rect 388000 -22636 397200 -22626
rect 388000 -22692 389141 -22636
rect 389197 -22692 389283 -22636
rect 389339 -22692 389542 -22636
rect 389598 -22692 389684 -22636
rect 389740 -22692 389942 -22636
rect 389998 -22692 390084 -22636
rect 390140 -22692 390339 -22636
rect 390395 -22692 390481 -22636
rect 390537 -22692 390736 -22636
rect 390792 -22692 390878 -22636
rect 390934 -22692 391140 -22636
rect 391196 -22692 391282 -22636
rect 391338 -22692 391536 -22636
rect 391592 -22692 391678 -22636
rect 391734 -22692 391936 -22636
rect 391992 -22692 392078 -22636
rect 392134 -22692 392333 -22636
rect 392389 -22692 392475 -22636
rect 392531 -22692 392738 -22636
rect 392794 -22692 392880 -22636
rect 392936 -22692 393138 -22636
rect 393194 -22692 393280 -22636
rect 393336 -22692 393543 -22636
rect 393599 -22692 393685 -22636
rect 393741 -22692 393940 -22636
rect 393996 -22692 394082 -22636
rect 394138 -22692 394337 -22636
rect 394393 -22692 394479 -22636
rect 394535 -22692 394740 -22636
rect 394796 -22692 394882 -22636
rect 394938 -22692 395142 -22636
rect 395198 -22692 395284 -22636
rect 395340 -22692 395545 -22636
rect 395601 -22692 395687 -22636
rect 395743 -22692 395941 -22636
rect 395997 -22692 396083 -22636
rect 396139 -22692 397200 -22636
rect 388000 -22694 397200 -22692
rect 388000 -22750 388114 -22694
rect 388170 -22750 388238 -22694
rect 388294 -22750 388362 -22694
rect 388418 -22750 388486 -22694
rect 388542 -22750 388610 -22694
rect 388666 -22750 396526 -22694
rect 396582 -22750 396650 -22694
rect 396706 -22750 396774 -22694
rect 396830 -22750 396898 -22694
rect 396954 -22750 397022 -22694
rect 397078 -22750 397200 -22694
rect 388000 -22778 397200 -22750
rect 388000 -22818 389141 -22778
rect 388000 -22874 388114 -22818
rect 388170 -22874 388238 -22818
rect 388294 -22874 388362 -22818
rect 388418 -22874 388486 -22818
rect 388542 -22874 388610 -22818
rect 388666 -22834 389141 -22818
rect 389197 -22834 389283 -22778
rect 389339 -22834 389542 -22778
rect 389598 -22834 389684 -22778
rect 389740 -22834 389942 -22778
rect 389998 -22834 390084 -22778
rect 390140 -22834 390339 -22778
rect 390395 -22834 390481 -22778
rect 390537 -22834 390736 -22778
rect 390792 -22834 390878 -22778
rect 390934 -22834 391140 -22778
rect 391196 -22834 391282 -22778
rect 391338 -22834 391536 -22778
rect 391592 -22834 391678 -22778
rect 391734 -22834 391936 -22778
rect 391992 -22834 392078 -22778
rect 392134 -22834 392333 -22778
rect 392389 -22834 392475 -22778
rect 392531 -22834 392738 -22778
rect 392794 -22834 392880 -22778
rect 392936 -22834 393138 -22778
rect 393194 -22834 393280 -22778
rect 393336 -22834 393543 -22778
rect 393599 -22834 393685 -22778
rect 393741 -22834 393940 -22778
rect 393996 -22834 394082 -22778
rect 394138 -22834 394337 -22778
rect 394393 -22834 394479 -22778
rect 394535 -22834 394740 -22778
rect 394796 -22834 394882 -22778
rect 394938 -22834 395142 -22778
rect 395198 -22834 395284 -22778
rect 395340 -22834 395545 -22778
rect 395601 -22834 395687 -22778
rect 395743 -22834 395941 -22778
rect 395997 -22834 396083 -22778
rect 396139 -22818 397200 -22778
rect 396139 -22834 396526 -22818
rect 388666 -22874 396526 -22834
rect 396582 -22874 396650 -22818
rect 396706 -22874 396774 -22818
rect 396830 -22874 396898 -22818
rect 396954 -22874 397022 -22818
rect 397078 -22874 397200 -22818
rect 388000 -22920 397200 -22874
rect 388000 -22942 389141 -22920
rect 388000 -22998 388114 -22942
rect 388170 -22998 388238 -22942
rect 388294 -22998 388362 -22942
rect 388418 -22998 388486 -22942
rect 388542 -22998 388610 -22942
rect 388666 -22976 389141 -22942
rect 389197 -22976 389283 -22920
rect 389339 -22976 389542 -22920
rect 389598 -22976 389684 -22920
rect 389740 -22976 389942 -22920
rect 389998 -22976 390084 -22920
rect 390140 -22976 390339 -22920
rect 390395 -22976 390481 -22920
rect 390537 -22976 390736 -22920
rect 390792 -22976 390878 -22920
rect 390934 -22976 391140 -22920
rect 391196 -22976 391282 -22920
rect 391338 -22976 391536 -22920
rect 391592 -22976 391678 -22920
rect 391734 -22976 391936 -22920
rect 391992 -22976 392078 -22920
rect 392134 -22976 392333 -22920
rect 392389 -22976 392475 -22920
rect 392531 -22976 392738 -22920
rect 392794 -22976 392880 -22920
rect 392936 -22976 393138 -22920
rect 393194 -22976 393280 -22920
rect 393336 -22976 393543 -22920
rect 393599 -22976 393685 -22920
rect 393741 -22976 393940 -22920
rect 393996 -22976 394082 -22920
rect 394138 -22976 394337 -22920
rect 394393 -22976 394479 -22920
rect 394535 -22976 394740 -22920
rect 394796 -22976 394882 -22920
rect 394938 -22976 395142 -22920
rect 395198 -22976 395284 -22920
rect 395340 -22976 395545 -22920
rect 395601 -22976 395687 -22920
rect 395743 -22976 395941 -22920
rect 395997 -22976 396083 -22920
rect 396139 -22942 397200 -22920
rect 396139 -22976 396526 -22942
rect 388666 -22998 396526 -22976
rect 396582 -22998 396650 -22942
rect 396706 -22998 396774 -22942
rect 396830 -22998 396898 -22942
rect 396954 -22998 397022 -22942
rect 397078 -22998 397200 -22942
rect 388000 -23062 397200 -22998
rect 388000 -23066 389141 -23062
rect 388000 -23122 388114 -23066
rect 388170 -23122 388238 -23066
rect 388294 -23122 388362 -23066
rect 388418 -23122 388486 -23066
rect 388542 -23122 388610 -23066
rect 388666 -23118 389141 -23066
rect 389197 -23118 389283 -23062
rect 389339 -23118 389542 -23062
rect 389598 -23118 389684 -23062
rect 389740 -23118 389942 -23062
rect 389998 -23118 390084 -23062
rect 390140 -23118 390339 -23062
rect 390395 -23118 390481 -23062
rect 390537 -23118 390736 -23062
rect 390792 -23118 390878 -23062
rect 390934 -23118 391140 -23062
rect 391196 -23118 391282 -23062
rect 391338 -23118 391536 -23062
rect 391592 -23118 391678 -23062
rect 391734 -23118 391936 -23062
rect 391992 -23118 392078 -23062
rect 392134 -23118 392333 -23062
rect 392389 -23118 392475 -23062
rect 392531 -23118 392738 -23062
rect 392794 -23118 392880 -23062
rect 392936 -23118 393138 -23062
rect 393194 -23118 393280 -23062
rect 393336 -23118 393543 -23062
rect 393599 -23118 393685 -23062
rect 393741 -23118 393940 -23062
rect 393996 -23118 394082 -23062
rect 394138 -23118 394337 -23062
rect 394393 -23118 394479 -23062
rect 394535 -23118 394740 -23062
rect 394796 -23118 394882 -23062
rect 394938 -23118 395142 -23062
rect 395198 -23118 395284 -23062
rect 395340 -23118 395545 -23062
rect 395601 -23118 395687 -23062
rect 395743 -23118 395941 -23062
rect 395997 -23118 396083 -23062
rect 396139 -23066 397200 -23062
rect 396139 -23118 396526 -23066
rect 388666 -23122 396526 -23118
rect 396582 -23122 396650 -23066
rect 396706 -23122 396774 -23066
rect 396830 -23122 396898 -23066
rect 396954 -23122 397022 -23066
rect 397078 -23122 397200 -23066
rect 388000 -23190 397200 -23122
rect 388000 -23246 388114 -23190
rect 388170 -23246 388238 -23190
rect 388294 -23246 388362 -23190
rect 388418 -23246 388486 -23190
rect 388542 -23246 388610 -23190
rect 388666 -23204 396526 -23190
rect 388666 -23246 389141 -23204
rect 388000 -23260 389141 -23246
rect 389197 -23260 389283 -23204
rect 389339 -23260 389542 -23204
rect 389598 -23260 389684 -23204
rect 389740 -23260 389942 -23204
rect 389998 -23260 390084 -23204
rect 390140 -23260 390339 -23204
rect 390395 -23260 390481 -23204
rect 390537 -23260 390736 -23204
rect 390792 -23260 390878 -23204
rect 390934 -23260 391140 -23204
rect 391196 -23260 391282 -23204
rect 391338 -23260 391536 -23204
rect 391592 -23260 391678 -23204
rect 391734 -23260 391936 -23204
rect 391992 -23260 392078 -23204
rect 392134 -23260 392333 -23204
rect 392389 -23260 392475 -23204
rect 392531 -23260 392738 -23204
rect 392794 -23260 392880 -23204
rect 392936 -23260 393138 -23204
rect 393194 -23260 393280 -23204
rect 393336 -23260 393543 -23204
rect 393599 -23260 393685 -23204
rect 393741 -23260 393940 -23204
rect 393996 -23260 394082 -23204
rect 394138 -23260 394337 -23204
rect 394393 -23260 394479 -23204
rect 394535 -23260 394740 -23204
rect 394796 -23260 394882 -23204
rect 394938 -23260 395142 -23204
rect 395198 -23260 395284 -23204
rect 395340 -23260 395545 -23204
rect 395601 -23260 395687 -23204
rect 395743 -23260 395941 -23204
rect 395997 -23260 396083 -23204
rect 396139 -23246 396526 -23204
rect 396582 -23246 396650 -23190
rect 396706 -23246 396774 -23190
rect 396830 -23246 396898 -23190
rect 396954 -23246 397022 -23190
rect 397078 -23246 397200 -23190
rect 396139 -23260 397200 -23246
rect 388000 -23314 397200 -23260
rect 388000 -23370 388114 -23314
rect 388170 -23370 388238 -23314
rect 388294 -23370 388362 -23314
rect 388418 -23370 388486 -23314
rect 388542 -23370 388610 -23314
rect 388666 -23346 396526 -23314
rect 388666 -23370 389141 -23346
rect 388000 -23402 389141 -23370
rect 389197 -23402 389283 -23346
rect 389339 -23402 389542 -23346
rect 389598 -23402 389684 -23346
rect 389740 -23402 389942 -23346
rect 389998 -23402 390084 -23346
rect 390140 -23402 390339 -23346
rect 390395 -23402 390481 -23346
rect 390537 -23402 390736 -23346
rect 390792 -23402 390878 -23346
rect 390934 -23402 391140 -23346
rect 391196 -23402 391282 -23346
rect 391338 -23402 391536 -23346
rect 391592 -23402 391678 -23346
rect 391734 -23402 391936 -23346
rect 391992 -23402 392078 -23346
rect 392134 -23402 392333 -23346
rect 392389 -23402 392475 -23346
rect 392531 -23402 392738 -23346
rect 392794 -23402 392880 -23346
rect 392936 -23402 393138 -23346
rect 393194 -23402 393280 -23346
rect 393336 -23402 393543 -23346
rect 393599 -23402 393685 -23346
rect 393741 -23402 393940 -23346
rect 393996 -23402 394082 -23346
rect 394138 -23402 394337 -23346
rect 394393 -23402 394479 -23346
rect 394535 -23402 394740 -23346
rect 394796 -23402 394882 -23346
rect 394938 -23402 395142 -23346
rect 395198 -23402 395284 -23346
rect 395340 -23402 395545 -23346
rect 395601 -23402 395687 -23346
rect 395743 -23402 395941 -23346
rect 395997 -23402 396083 -23346
rect 396139 -23370 396526 -23346
rect 396582 -23370 396650 -23314
rect 396706 -23370 396774 -23314
rect 396830 -23370 396898 -23314
rect 396954 -23370 397022 -23314
rect 397078 -23370 397200 -23314
rect 396139 -23402 397200 -23370
rect 388000 -23438 397200 -23402
rect 388000 -23494 388114 -23438
rect 388170 -23494 388238 -23438
rect 388294 -23494 388362 -23438
rect 388418 -23494 388486 -23438
rect 388542 -23494 388610 -23438
rect 388666 -23488 396526 -23438
rect 388666 -23494 389141 -23488
rect 388000 -23544 389141 -23494
rect 389197 -23544 389283 -23488
rect 389339 -23544 389542 -23488
rect 389598 -23544 389684 -23488
rect 389740 -23544 389942 -23488
rect 389998 -23544 390084 -23488
rect 390140 -23544 390339 -23488
rect 390395 -23544 390481 -23488
rect 390537 -23544 390736 -23488
rect 390792 -23544 390878 -23488
rect 390934 -23544 391140 -23488
rect 391196 -23544 391282 -23488
rect 391338 -23544 391536 -23488
rect 391592 -23544 391678 -23488
rect 391734 -23544 391936 -23488
rect 391992 -23544 392078 -23488
rect 392134 -23544 392333 -23488
rect 392389 -23544 392475 -23488
rect 392531 -23544 392738 -23488
rect 392794 -23544 392880 -23488
rect 392936 -23544 393138 -23488
rect 393194 -23544 393280 -23488
rect 393336 -23544 393543 -23488
rect 393599 -23544 393685 -23488
rect 393741 -23544 393940 -23488
rect 393996 -23544 394082 -23488
rect 394138 -23544 394337 -23488
rect 394393 -23544 394479 -23488
rect 394535 -23544 394740 -23488
rect 394796 -23544 394882 -23488
rect 394938 -23544 395142 -23488
rect 395198 -23544 395284 -23488
rect 395340 -23544 395545 -23488
rect 395601 -23544 395687 -23488
rect 395743 -23544 395941 -23488
rect 395997 -23544 396083 -23488
rect 396139 -23494 396526 -23488
rect 396582 -23494 396650 -23438
rect 396706 -23494 396774 -23438
rect 396830 -23494 396898 -23438
rect 396954 -23494 397022 -23438
rect 397078 -23494 397200 -23438
rect 396139 -23544 397200 -23494
rect 388000 -23562 397200 -23544
rect 388000 -23618 388114 -23562
rect 388170 -23618 388238 -23562
rect 388294 -23618 388362 -23562
rect 388418 -23618 388486 -23562
rect 388542 -23618 388610 -23562
rect 388666 -23618 396526 -23562
rect 396582 -23618 396650 -23562
rect 396706 -23618 396774 -23562
rect 396830 -23618 396898 -23562
rect 396954 -23618 397022 -23562
rect 397078 -23618 397200 -23562
rect 388000 -23630 397200 -23618
rect 388000 -23686 389141 -23630
rect 389197 -23686 389283 -23630
rect 389339 -23686 389542 -23630
rect 389598 -23686 389684 -23630
rect 389740 -23686 389942 -23630
rect 389998 -23686 390084 -23630
rect 390140 -23686 390339 -23630
rect 390395 -23686 390481 -23630
rect 390537 -23686 390736 -23630
rect 390792 -23686 390878 -23630
rect 390934 -23686 391140 -23630
rect 391196 -23686 391282 -23630
rect 391338 -23686 391536 -23630
rect 391592 -23686 391678 -23630
rect 391734 -23686 391936 -23630
rect 391992 -23686 392078 -23630
rect 392134 -23686 392333 -23630
rect 392389 -23686 392475 -23630
rect 392531 -23686 392738 -23630
rect 392794 -23686 392880 -23630
rect 392936 -23686 393138 -23630
rect 393194 -23686 393280 -23630
rect 393336 -23686 393543 -23630
rect 393599 -23686 393685 -23630
rect 393741 -23686 393940 -23630
rect 393996 -23686 394082 -23630
rect 394138 -23686 394337 -23630
rect 394393 -23686 394479 -23630
rect 394535 -23686 394740 -23630
rect 394796 -23686 394882 -23630
rect 394938 -23686 395142 -23630
rect 395198 -23686 395284 -23630
rect 395340 -23686 395545 -23630
rect 395601 -23686 395687 -23630
rect 395743 -23686 395941 -23630
rect 395997 -23686 396083 -23630
rect 396139 -23686 397200 -23630
rect 388000 -23742 388114 -23686
rect 388170 -23742 388238 -23686
rect 388294 -23742 388362 -23686
rect 388418 -23742 388486 -23686
rect 388542 -23742 388610 -23686
rect 388666 -23742 396526 -23686
rect 396582 -23742 396650 -23686
rect 396706 -23742 396774 -23686
rect 396830 -23742 396898 -23686
rect 396954 -23742 397022 -23686
rect 397078 -23742 397200 -23686
rect 388000 -23772 397200 -23742
rect 388000 -23810 389141 -23772
rect 388000 -23866 388114 -23810
rect 388170 -23866 388238 -23810
rect 388294 -23866 388362 -23810
rect 388418 -23866 388486 -23810
rect 388542 -23866 388610 -23810
rect 388666 -23828 389141 -23810
rect 389197 -23828 389283 -23772
rect 389339 -23828 389542 -23772
rect 389598 -23828 389684 -23772
rect 389740 -23828 389942 -23772
rect 389998 -23828 390084 -23772
rect 390140 -23828 390339 -23772
rect 390395 -23828 390481 -23772
rect 390537 -23828 390736 -23772
rect 390792 -23828 390878 -23772
rect 390934 -23828 391140 -23772
rect 391196 -23828 391282 -23772
rect 391338 -23828 391536 -23772
rect 391592 -23828 391678 -23772
rect 391734 -23828 391936 -23772
rect 391992 -23828 392078 -23772
rect 392134 -23828 392333 -23772
rect 392389 -23828 392475 -23772
rect 392531 -23828 392738 -23772
rect 392794 -23828 392880 -23772
rect 392936 -23828 393138 -23772
rect 393194 -23828 393280 -23772
rect 393336 -23828 393543 -23772
rect 393599 -23828 393685 -23772
rect 393741 -23828 393940 -23772
rect 393996 -23828 394082 -23772
rect 394138 -23828 394337 -23772
rect 394393 -23828 394479 -23772
rect 394535 -23828 394740 -23772
rect 394796 -23828 394882 -23772
rect 394938 -23828 395142 -23772
rect 395198 -23828 395284 -23772
rect 395340 -23828 395545 -23772
rect 395601 -23828 395687 -23772
rect 395743 -23828 395941 -23772
rect 395997 -23828 396083 -23772
rect 396139 -23810 397200 -23772
rect 396139 -23828 396526 -23810
rect 388666 -23866 396526 -23828
rect 396582 -23866 396650 -23810
rect 396706 -23866 396774 -23810
rect 396830 -23866 396898 -23810
rect 396954 -23866 397022 -23810
rect 397078 -23866 397200 -23810
rect 388000 -23914 397200 -23866
rect 388000 -23934 389141 -23914
rect 388000 -23990 388114 -23934
rect 388170 -23990 388238 -23934
rect 388294 -23990 388362 -23934
rect 388418 -23990 388486 -23934
rect 388542 -23990 388610 -23934
rect 388666 -23970 389141 -23934
rect 389197 -23970 389283 -23914
rect 389339 -23970 389542 -23914
rect 389598 -23970 389684 -23914
rect 389740 -23970 389942 -23914
rect 389998 -23970 390084 -23914
rect 390140 -23970 390339 -23914
rect 390395 -23970 390481 -23914
rect 390537 -23970 390736 -23914
rect 390792 -23970 390878 -23914
rect 390934 -23970 391140 -23914
rect 391196 -23970 391282 -23914
rect 391338 -23970 391536 -23914
rect 391592 -23970 391678 -23914
rect 391734 -23970 391936 -23914
rect 391992 -23970 392078 -23914
rect 392134 -23970 392333 -23914
rect 392389 -23970 392475 -23914
rect 392531 -23970 392738 -23914
rect 392794 -23970 392880 -23914
rect 392936 -23970 393138 -23914
rect 393194 -23970 393280 -23914
rect 393336 -23970 393543 -23914
rect 393599 -23970 393685 -23914
rect 393741 -23970 393940 -23914
rect 393996 -23970 394082 -23914
rect 394138 -23970 394337 -23914
rect 394393 -23970 394479 -23914
rect 394535 -23970 394740 -23914
rect 394796 -23970 394882 -23914
rect 394938 -23970 395142 -23914
rect 395198 -23970 395284 -23914
rect 395340 -23970 395545 -23914
rect 395601 -23970 395687 -23914
rect 395743 -23970 395941 -23914
rect 395997 -23970 396083 -23914
rect 396139 -23934 397200 -23914
rect 396139 -23970 396526 -23934
rect 388666 -23990 396526 -23970
rect 396582 -23990 396650 -23934
rect 396706 -23990 396774 -23934
rect 396830 -23990 396898 -23934
rect 396954 -23990 397022 -23934
rect 397078 -23990 397200 -23934
rect 388000 -24056 397200 -23990
rect 388000 -24058 389141 -24056
rect 388000 -24114 388114 -24058
rect 388170 -24114 388238 -24058
rect 388294 -24114 388362 -24058
rect 388418 -24114 388486 -24058
rect 388542 -24114 388610 -24058
rect 388666 -24112 389141 -24058
rect 389197 -24112 389283 -24056
rect 389339 -24112 389542 -24056
rect 389598 -24112 389684 -24056
rect 389740 -24112 389942 -24056
rect 389998 -24112 390084 -24056
rect 390140 -24112 390339 -24056
rect 390395 -24112 390481 -24056
rect 390537 -24112 390736 -24056
rect 390792 -24112 390878 -24056
rect 390934 -24112 391140 -24056
rect 391196 -24112 391282 -24056
rect 391338 -24112 391536 -24056
rect 391592 -24112 391678 -24056
rect 391734 -24112 391936 -24056
rect 391992 -24112 392078 -24056
rect 392134 -24112 392333 -24056
rect 392389 -24112 392475 -24056
rect 392531 -24112 392738 -24056
rect 392794 -24112 392880 -24056
rect 392936 -24112 393138 -24056
rect 393194 -24112 393280 -24056
rect 393336 -24112 393543 -24056
rect 393599 -24112 393685 -24056
rect 393741 -24112 393940 -24056
rect 393996 -24112 394082 -24056
rect 394138 -24112 394337 -24056
rect 394393 -24112 394479 -24056
rect 394535 -24112 394740 -24056
rect 394796 -24112 394882 -24056
rect 394938 -24112 395142 -24056
rect 395198 -24112 395284 -24056
rect 395340 -24112 395545 -24056
rect 395601 -24112 395687 -24056
rect 395743 -24112 395941 -24056
rect 395997 -24112 396083 -24056
rect 396139 -24058 397200 -24056
rect 396139 -24112 396526 -24058
rect 388666 -24114 396526 -24112
rect 396582 -24114 396650 -24058
rect 396706 -24114 396774 -24058
rect 396830 -24114 396898 -24058
rect 396954 -24114 397022 -24058
rect 397078 -24114 397200 -24058
rect 388000 -24182 397200 -24114
rect 388000 -24238 388114 -24182
rect 388170 -24238 388238 -24182
rect 388294 -24238 388362 -24182
rect 388418 -24238 388486 -24182
rect 388542 -24238 388610 -24182
rect 388666 -24198 396526 -24182
rect 388666 -24238 389141 -24198
rect 388000 -24254 389141 -24238
rect 389197 -24254 389283 -24198
rect 389339 -24254 389542 -24198
rect 389598 -24254 389684 -24198
rect 389740 -24254 389942 -24198
rect 389998 -24254 390084 -24198
rect 390140 -24254 390339 -24198
rect 390395 -24254 390481 -24198
rect 390537 -24254 390736 -24198
rect 390792 -24254 390878 -24198
rect 390934 -24254 391140 -24198
rect 391196 -24254 391282 -24198
rect 391338 -24254 391536 -24198
rect 391592 -24254 391678 -24198
rect 391734 -24254 391936 -24198
rect 391992 -24254 392078 -24198
rect 392134 -24254 392333 -24198
rect 392389 -24254 392475 -24198
rect 392531 -24254 392738 -24198
rect 392794 -24254 392880 -24198
rect 392936 -24254 393138 -24198
rect 393194 -24254 393280 -24198
rect 393336 -24254 393543 -24198
rect 393599 -24254 393685 -24198
rect 393741 -24254 393940 -24198
rect 393996 -24254 394082 -24198
rect 394138 -24254 394337 -24198
rect 394393 -24254 394479 -24198
rect 394535 -24254 394740 -24198
rect 394796 -24254 394882 -24198
rect 394938 -24254 395142 -24198
rect 395198 -24254 395284 -24198
rect 395340 -24254 395545 -24198
rect 395601 -24254 395687 -24198
rect 395743 -24254 395941 -24198
rect 395997 -24254 396083 -24198
rect 396139 -24238 396526 -24198
rect 396582 -24238 396650 -24182
rect 396706 -24238 396774 -24182
rect 396830 -24238 396898 -24182
rect 396954 -24238 397022 -24182
rect 397078 -24238 397200 -24182
rect 396139 -24254 397200 -24238
rect 388000 -24306 397200 -24254
rect 388000 -24362 388114 -24306
rect 388170 -24362 388238 -24306
rect 388294 -24362 388362 -24306
rect 388418 -24362 388486 -24306
rect 388542 -24362 388610 -24306
rect 388666 -24340 396526 -24306
rect 388666 -24362 389141 -24340
rect 388000 -24396 389141 -24362
rect 389197 -24396 389283 -24340
rect 389339 -24396 389542 -24340
rect 389598 -24396 389684 -24340
rect 389740 -24396 389942 -24340
rect 389998 -24396 390084 -24340
rect 390140 -24396 390339 -24340
rect 390395 -24396 390481 -24340
rect 390537 -24396 390736 -24340
rect 390792 -24396 390878 -24340
rect 390934 -24396 391140 -24340
rect 391196 -24396 391282 -24340
rect 391338 -24396 391536 -24340
rect 391592 -24396 391678 -24340
rect 391734 -24396 391936 -24340
rect 391992 -24396 392078 -24340
rect 392134 -24396 392333 -24340
rect 392389 -24396 392475 -24340
rect 392531 -24396 392738 -24340
rect 392794 -24396 392880 -24340
rect 392936 -24396 393138 -24340
rect 393194 -24396 393280 -24340
rect 393336 -24396 393543 -24340
rect 393599 -24396 393685 -24340
rect 393741 -24396 393940 -24340
rect 393996 -24396 394082 -24340
rect 394138 -24396 394337 -24340
rect 394393 -24396 394479 -24340
rect 394535 -24396 394740 -24340
rect 394796 -24396 394882 -24340
rect 394938 -24396 395142 -24340
rect 395198 -24396 395284 -24340
rect 395340 -24396 395545 -24340
rect 395601 -24396 395687 -24340
rect 395743 -24396 395941 -24340
rect 395997 -24396 396083 -24340
rect 396139 -24362 396526 -24340
rect 396582 -24362 396650 -24306
rect 396706 -24362 396774 -24306
rect 396830 -24362 396898 -24306
rect 396954 -24362 397022 -24306
rect 397078 -24362 397200 -24306
rect 396139 -24396 397200 -24362
rect 388000 -24430 397200 -24396
rect 388000 -24486 388114 -24430
rect 388170 -24486 388238 -24430
rect 388294 -24486 388362 -24430
rect 388418 -24486 388486 -24430
rect 388542 -24486 388610 -24430
rect 388666 -24482 396526 -24430
rect 388666 -24486 389141 -24482
rect 388000 -24538 389141 -24486
rect 389197 -24538 389283 -24482
rect 389339 -24538 389542 -24482
rect 389598 -24538 389684 -24482
rect 389740 -24538 389942 -24482
rect 389998 -24538 390084 -24482
rect 390140 -24538 390339 -24482
rect 390395 -24538 390481 -24482
rect 390537 -24538 390736 -24482
rect 390792 -24538 390878 -24482
rect 390934 -24538 391140 -24482
rect 391196 -24538 391282 -24482
rect 391338 -24538 391536 -24482
rect 391592 -24538 391678 -24482
rect 391734 -24538 391936 -24482
rect 391992 -24538 392078 -24482
rect 392134 -24538 392333 -24482
rect 392389 -24538 392475 -24482
rect 392531 -24538 392738 -24482
rect 392794 -24538 392880 -24482
rect 392936 -24538 393138 -24482
rect 393194 -24538 393280 -24482
rect 393336 -24538 393543 -24482
rect 393599 -24538 393685 -24482
rect 393741 -24538 393940 -24482
rect 393996 -24538 394082 -24482
rect 394138 -24538 394337 -24482
rect 394393 -24538 394479 -24482
rect 394535 -24538 394740 -24482
rect 394796 -24538 394882 -24482
rect 394938 -24538 395142 -24482
rect 395198 -24538 395284 -24482
rect 395340 -24538 395545 -24482
rect 395601 -24538 395687 -24482
rect 395743 -24538 395941 -24482
rect 395997 -24538 396083 -24482
rect 396139 -24486 396526 -24482
rect 396582 -24486 396650 -24430
rect 396706 -24486 396774 -24430
rect 396830 -24486 396898 -24430
rect 396954 -24486 397022 -24430
rect 397078 -24486 397200 -24430
rect 396139 -24538 397200 -24486
rect 388000 -24554 397200 -24538
rect 388000 -24610 388114 -24554
rect 388170 -24610 388238 -24554
rect 388294 -24610 388362 -24554
rect 388418 -24610 388486 -24554
rect 388542 -24610 388610 -24554
rect 388666 -24610 396526 -24554
rect 396582 -24610 396650 -24554
rect 396706 -24610 396774 -24554
rect 396830 -24610 396898 -24554
rect 396954 -24610 397022 -24554
rect 397078 -24610 397200 -24554
rect 388000 -24624 397200 -24610
rect 388000 -24678 389141 -24624
rect 388000 -24734 388114 -24678
rect 388170 -24734 388238 -24678
rect 388294 -24734 388362 -24678
rect 388418 -24734 388486 -24678
rect 388542 -24734 388610 -24678
rect 388666 -24680 389141 -24678
rect 389197 -24680 389283 -24624
rect 389339 -24680 389542 -24624
rect 389598 -24680 389684 -24624
rect 389740 -24680 389942 -24624
rect 389998 -24680 390084 -24624
rect 390140 -24680 390339 -24624
rect 390395 -24680 390481 -24624
rect 390537 -24680 390736 -24624
rect 390792 -24680 390878 -24624
rect 390934 -24680 391140 -24624
rect 391196 -24680 391282 -24624
rect 391338 -24680 391536 -24624
rect 391592 -24680 391678 -24624
rect 391734 -24680 391936 -24624
rect 391992 -24680 392078 -24624
rect 392134 -24680 392333 -24624
rect 392389 -24680 392475 -24624
rect 392531 -24680 392738 -24624
rect 392794 -24680 392880 -24624
rect 392936 -24680 393138 -24624
rect 393194 -24680 393280 -24624
rect 393336 -24680 393543 -24624
rect 393599 -24680 393685 -24624
rect 393741 -24680 393940 -24624
rect 393996 -24680 394082 -24624
rect 394138 -24680 394337 -24624
rect 394393 -24680 394479 -24624
rect 394535 -24680 394740 -24624
rect 394796 -24680 394882 -24624
rect 394938 -24680 395142 -24624
rect 395198 -24680 395284 -24624
rect 395340 -24680 395545 -24624
rect 395601 -24680 395687 -24624
rect 395743 -24680 395941 -24624
rect 395997 -24680 396083 -24624
rect 396139 -24678 397200 -24624
rect 396139 -24680 396526 -24678
rect 388666 -24734 396526 -24680
rect 396582 -24734 396650 -24678
rect 396706 -24734 396774 -24678
rect 396830 -24734 396898 -24678
rect 396954 -24734 397022 -24678
rect 397078 -24734 397200 -24678
rect 388000 -24766 397200 -24734
rect 388000 -24802 389141 -24766
rect 388000 -24858 388114 -24802
rect 388170 -24858 388238 -24802
rect 388294 -24858 388362 -24802
rect 388418 -24858 388486 -24802
rect 388542 -24858 388610 -24802
rect 388666 -24822 389141 -24802
rect 389197 -24822 389283 -24766
rect 389339 -24822 389542 -24766
rect 389598 -24822 389684 -24766
rect 389740 -24822 389942 -24766
rect 389998 -24822 390084 -24766
rect 390140 -24822 390339 -24766
rect 390395 -24822 390481 -24766
rect 390537 -24822 390736 -24766
rect 390792 -24822 390878 -24766
rect 390934 -24822 391140 -24766
rect 391196 -24822 391282 -24766
rect 391338 -24822 391536 -24766
rect 391592 -24822 391678 -24766
rect 391734 -24822 391936 -24766
rect 391992 -24822 392078 -24766
rect 392134 -24822 392333 -24766
rect 392389 -24822 392475 -24766
rect 392531 -24822 392738 -24766
rect 392794 -24822 392880 -24766
rect 392936 -24822 393138 -24766
rect 393194 -24822 393280 -24766
rect 393336 -24822 393543 -24766
rect 393599 -24822 393685 -24766
rect 393741 -24822 393940 -24766
rect 393996 -24822 394082 -24766
rect 394138 -24822 394337 -24766
rect 394393 -24822 394479 -24766
rect 394535 -24822 394740 -24766
rect 394796 -24822 394882 -24766
rect 394938 -24822 395142 -24766
rect 395198 -24822 395284 -24766
rect 395340 -24822 395545 -24766
rect 395601 -24822 395687 -24766
rect 395743 -24822 395941 -24766
rect 395997 -24822 396083 -24766
rect 396139 -24802 397200 -24766
rect 396139 -24822 396526 -24802
rect 388666 -24858 396526 -24822
rect 396582 -24858 396650 -24802
rect 396706 -24858 396774 -24802
rect 396830 -24858 396898 -24802
rect 396954 -24858 397022 -24802
rect 397078 -24858 397200 -24802
rect 388000 -24908 397200 -24858
rect 388000 -24926 389141 -24908
rect 388000 -24982 388114 -24926
rect 388170 -24982 388238 -24926
rect 388294 -24982 388362 -24926
rect 388418 -24982 388486 -24926
rect 388542 -24982 388610 -24926
rect 388666 -24964 389141 -24926
rect 389197 -24964 389283 -24908
rect 389339 -24964 389542 -24908
rect 389598 -24964 389684 -24908
rect 389740 -24964 389942 -24908
rect 389998 -24964 390084 -24908
rect 390140 -24964 390339 -24908
rect 390395 -24964 390481 -24908
rect 390537 -24964 390736 -24908
rect 390792 -24964 390878 -24908
rect 390934 -24964 391140 -24908
rect 391196 -24964 391282 -24908
rect 391338 -24964 391536 -24908
rect 391592 -24964 391678 -24908
rect 391734 -24964 391936 -24908
rect 391992 -24964 392078 -24908
rect 392134 -24964 392333 -24908
rect 392389 -24964 392475 -24908
rect 392531 -24964 392738 -24908
rect 392794 -24964 392880 -24908
rect 392936 -24964 393138 -24908
rect 393194 -24964 393280 -24908
rect 393336 -24964 393543 -24908
rect 393599 -24964 393685 -24908
rect 393741 -24964 393940 -24908
rect 393996 -24964 394082 -24908
rect 394138 -24964 394337 -24908
rect 394393 -24964 394479 -24908
rect 394535 -24964 394740 -24908
rect 394796 -24964 394882 -24908
rect 394938 -24964 395142 -24908
rect 395198 -24964 395284 -24908
rect 395340 -24964 395545 -24908
rect 395601 -24964 395687 -24908
rect 395743 -24964 395941 -24908
rect 395997 -24964 396083 -24908
rect 396139 -24926 397200 -24908
rect 396139 -24964 396526 -24926
rect 388666 -24982 396526 -24964
rect 396582 -24982 396650 -24926
rect 396706 -24982 396774 -24926
rect 396830 -24982 396898 -24926
rect 396954 -24982 397022 -24926
rect 397078 -24982 397200 -24926
rect 388000 -25050 397200 -24982
rect 388000 -25106 388114 -25050
rect 388170 -25106 388238 -25050
rect 388294 -25106 388362 -25050
rect 388418 -25106 388486 -25050
rect 388542 -25106 388610 -25050
rect 388666 -25106 389141 -25050
rect 389197 -25106 389283 -25050
rect 389339 -25106 389542 -25050
rect 389598 -25106 389684 -25050
rect 389740 -25106 389942 -25050
rect 389998 -25106 390084 -25050
rect 390140 -25106 390339 -25050
rect 390395 -25106 390481 -25050
rect 390537 -25106 390736 -25050
rect 390792 -25106 390878 -25050
rect 390934 -25106 391140 -25050
rect 391196 -25106 391282 -25050
rect 391338 -25106 391536 -25050
rect 391592 -25106 391678 -25050
rect 391734 -25106 391936 -25050
rect 391992 -25106 392078 -25050
rect 392134 -25106 392333 -25050
rect 392389 -25106 392475 -25050
rect 392531 -25106 392738 -25050
rect 392794 -25106 392880 -25050
rect 392936 -25106 393138 -25050
rect 393194 -25106 393280 -25050
rect 393336 -25106 393543 -25050
rect 393599 -25106 393685 -25050
rect 393741 -25106 393940 -25050
rect 393996 -25106 394082 -25050
rect 394138 -25106 394337 -25050
rect 394393 -25106 394479 -25050
rect 394535 -25106 394740 -25050
rect 394796 -25106 394882 -25050
rect 394938 -25106 395142 -25050
rect 395198 -25106 395284 -25050
rect 395340 -25106 395545 -25050
rect 395601 -25106 395687 -25050
rect 395743 -25106 395941 -25050
rect 395997 -25106 396083 -25050
rect 396139 -25106 396526 -25050
rect 396582 -25106 396650 -25050
rect 396706 -25106 396774 -25050
rect 396830 -25106 396898 -25050
rect 396954 -25106 397022 -25050
rect 397078 -25106 397200 -25050
rect 388000 -25174 397200 -25106
rect 388000 -25230 388114 -25174
rect 388170 -25230 388238 -25174
rect 388294 -25230 388362 -25174
rect 388418 -25230 388486 -25174
rect 388542 -25230 388610 -25174
rect 388666 -25192 396526 -25174
rect 388666 -25230 389141 -25192
rect 388000 -25248 389141 -25230
rect 389197 -25248 389283 -25192
rect 389339 -25248 389542 -25192
rect 389598 -25248 389684 -25192
rect 389740 -25248 389942 -25192
rect 389998 -25248 390084 -25192
rect 390140 -25248 390339 -25192
rect 390395 -25248 390481 -25192
rect 390537 -25248 390736 -25192
rect 390792 -25248 390878 -25192
rect 390934 -25248 391140 -25192
rect 391196 -25248 391282 -25192
rect 391338 -25248 391536 -25192
rect 391592 -25248 391678 -25192
rect 391734 -25248 391936 -25192
rect 391992 -25248 392078 -25192
rect 392134 -25248 392333 -25192
rect 392389 -25248 392475 -25192
rect 392531 -25248 392738 -25192
rect 392794 -25248 392880 -25192
rect 392936 -25248 393138 -25192
rect 393194 -25248 393280 -25192
rect 393336 -25248 393543 -25192
rect 393599 -25248 393685 -25192
rect 393741 -25248 393940 -25192
rect 393996 -25248 394082 -25192
rect 394138 -25248 394337 -25192
rect 394393 -25248 394479 -25192
rect 394535 -25248 394740 -25192
rect 394796 -25248 394882 -25192
rect 394938 -25248 395142 -25192
rect 395198 -25248 395284 -25192
rect 395340 -25248 395545 -25192
rect 395601 -25248 395687 -25192
rect 395743 -25248 395941 -25192
rect 395997 -25248 396083 -25192
rect 396139 -25230 396526 -25192
rect 396582 -25230 396650 -25174
rect 396706 -25230 396774 -25174
rect 396830 -25230 396898 -25174
rect 396954 -25230 397022 -25174
rect 397078 -25230 397200 -25174
rect 396139 -25248 397200 -25230
rect 388000 -25298 397200 -25248
rect 388000 -25354 388114 -25298
rect 388170 -25354 388238 -25298
rect 388294 -25354 388362 -25298
rect 388418 -25354 388486 -25298
rect 388542 -25354 388610 -25298
rect 388666 -25334 396526 -25298
rect 388666 -25354 389141 -25334
rect 388000 -25390 389141 -25354
rect 389197 -25390 389283 -25334
rect 389339 -25390 389542 -25334
rect 389598 -25390 389684 -25334
rect 389740 -25390 389942 -25334
rect 389998 -25390 390084 -25334
rect 390140 -25390 390339 -25334
rect 390395 -25390 390481 -25334
rect 390537 -25390 390736 -25334
rect 390792 -25390 390878 -25334
rect 390934 -25390 391140 -25334
rect 391196 -25390 391282 -25334
rect 391338 -25390 391536 -25334
rect 391592 -25390 391678 -25334
rect 391734 -25390 391936 -25334
rect 391992 -25390 392078 -25334
rect 392134 -25390 392333 -25334
rect 392389 -25390 392475 -25334
rect 392531 -25390 392738 -25334
rect 392794 -25390 392880 -25334
rect 392936 -25390 393138 -25334
rect 393194 -25390 393280 -25334
rect 393336 -25390 393543 -25334
rect 393599 -25390 393685 -25334
rect 393741 -25390 393940 -25334
rect 393996 -25390 394082 -25334
rect 394138 -25390 394337 -25334
rect 394393 -25390 394479 -25334
rect 394535 -25390 394740 -25334
rect 394796 -25390 394882 -25334
rect 394938 -25390 395142 -25334
rect 395198 -25390 395284 -25334
rect 395340 -25390 395545 -25334
rect 395601 -25390 395687 -25334
rect 395743 -25390 395941 -25334
rect 395997 -25390 396083 -25334
rect 396139 -25354 396526 -25334
rect 396582 -25354 396650 -25298
rect 396706 -25354 396774 -25298
rect 396830 -25354 396898 -25298
rect 396954 -25354 397022 -25298
rect 397078 -25354 397200 -25298
rect 396139 -25390 397200 -25354
rect 388000 -25422 397200 -25390
rect 388000 -25478 388114 -25422
rect 388170 -25478 388238 -25422
rect 388294 -25478 388362 -25422
rect 388418 -25478 388486 -25422
rect 388542 -25478 388610 -25422
rect 388666 -25476 396526 -25422
rect 388666 -25478 389141 -25476
rect 388000 -25532 389141 -25478
rect 389197 -25532 389283 -25476
rect 389339 -25532 389542 -25476
rect 389598 -25532 389684 -25476
rect 389740 -25532 389942 -25476
rect 389998 -25532 390084 -25476
rect 390140 -25532 390339 -25476
rect 390395 -25532 390481 -25476
rect 390537 -25532 390736 -25476
rect 390792 -25532 390878 -25476
rect 390934 -25532 391140 -25476
rect 391196 -25532 391282 -25476
rect 391338 -25532 391536 -25476
rect 391592 -25532 391678 -25476
rect 391734 -25532 391936 -25476
rect 391992 -25532 392078 -25476
rect 392134 -25532 392333 -25476
rect 392389 -25532 392475 -25476
rect 392531 -25532 392738 -25476
rect 392794 -25532 392880 -25476
rect 392936 -25532 393138 -25476
rect 393194 -25532 393280 -25476
rect 393336 -25532 393543 -25476
rect 393599 -25532 393685 -25476
rect 393741 -25532 393940 -25476
rect 393996 -25532 394082 -25476
rect 394138 -25532 394337 -25476
rect 394393 -25532 394479 -25476
rect 394535 -25532 394740 -25476
rect 394796 -25532 394882 -25476
rect 394938 -25532 395142 -25476
rect 395198 -25532 395284 -25476
rect 395340 -25532 395545 -25476
rect 395601 -25532 395687 -25476
rect 395743 -25532 395941 -25476
rect 395997 -25532 396083 -25476
rect 396139 -25478 396526 -25476
rect 396582 -25478 396650 -25422
rect 396706 -25478 396774 -25422
rect 396830 -25478 396898 -25422
rect 396954 -25478 397022 -25422
rect 397078 -25478 397200 -25422
rect 396139 -25532 397200 -25478
rect 388000 -25721 397200 -25532
rect 388000 -25777 388146 -25721
rect 388202 -25777 388270 -25721
rect 388326 -25777 388394 -25721
rect 388450 -25777 388518 -25721
rect 388574 -25777 388642 -25721
rect 388698 -25777 388766 -25721
rect 388822 -25777 388890 -25721
rect 388946 -25777 389014 -25721
rect 389070 -25777 389138 -25721
rect 389194 -25777 389262 -25721
rect 389318 -25777 389386 -25721
rect 389442 -25777 389510 -25721
rect 389566 -25777 389634 -25721
rect 389690 -25777 389758 -25721
rect 389814 -25777 389882 -25721
rect 389938 -25777 390006 -25721
rect 390062 -25777 390130 -25721
rect 390186 -25777 390254 -25721
rect 390310 -25777 390378 -25721
rect 390434 -25777 390502 -25721
rect 390558 -25777 390626 -25721
rect 390682 -25777 390750 -25721
rect 390806 -25777 390874 -25721
rect 390930 -25777 390998 -25721
rect 391054 -25777 391122 -25721
rect 391178 -25777 391246 -25721
rect 391302 -25777 391370 -25721
rect 391426 -25777 391494 -25721
rect 391550 -25777 391618 -25721
rect 391674 -25777 391742 -25721
rect 391798 -25777 391866 -25721
rect 391922 -25777 391990 -25721
rect 392046 -25777 392114 -25721
rect 392170 -25777 392238 -25721
rect 392294 -25777 392362 -25721
rect 392418 -25777 392486 -25721
rect 392542 -25777 392610 -25721
rect 392666 -25777 392734 -25721
rect 392790 -25777 392858 -25721
rect 392914 -25777 392982 -25721
rect 393038 -25777 393106 -25721
rect 393162 -25777 393230 -25721
rect 393286 -25777 393354 -25721
rect 393410 -25777 393478 -25721
rect 393534 -25777 393602 -25721
rect 393658 -25777 393726 -25721
rect 393782 -25777 393850 -25721
rect 393906 -25777 393974 -25721
rect 394030 -25777 394098 -25721
rect 394154 -25777 394222 -25721
rect 394278 -25777 394346 -25721
rect 394402 -25777 394470 -25721
rect 394526 -25777 394594 -25721
rect 394650 -25777 394718 -25721
rect 394774 -25777 394842 -25721
rect 394898 -25777 394966 -25721
rect 395022 -25777 395090 -25721
rect 395146 -25777 395214 -25721
rect 395270 -25777 395338 -25721
rect 395394 -25777 395462 -25721
rect 395518 -25777 395586 -25721
rect 395642 -25777 395710 -25721
rect 395766 -25777 395898 -25721
rect 395954 -25777 396022 -25721
rect 396078 -25777 396146 -25721
rect 396202 -25777 396270 -25721
rect 396326 -25777 396394 -25721
rect 396450 -25777 396518 -25721
rect 396574 -25777 396642 -25721
rect 396698 -25777 396766 -25721
rect 396822 -25777 396890 -25721
rect 396946 -25777 397014 -25721
rect 397070 -25777 397200 -25721
rect 388000 -25845 397200 -25777
rect 388000 -25901 388146 -25845
rect 388202 -25901 388270 -25845
rect 388326 -25901 388394 -25845
rect 388450 -25901 388518 -25845
rect 388574 -25901 388642 -25845
rect 388698 -25901 388766 -25845
rect 388822 -25901 388890 -25845
rect 388946 -25901 389014 -25845
rect 389070 -25901 389138 -25845
rect 389194 -25901 389262 -25845
rect 389318 -25901 389386 -25845
rect 389442 -25901 389510 -25845
rect 389566 -25901 389634 -25845
rect 389690 -25901 389758 -25845
rect 389814 -25901 389882 -25845
rect 389938 -25901 390006 -25845
rect 390062 -25901 390130 -25845
rect 390186 -25901 390254 -25845
rect 390310 -25901 390378 -25845
rect 390434 -25901 390502 -25845
rect 390558 -25901 390626 -25845
rect 390682 -25901 390750 -25845
rect 390806 -25901 390874 -25845
rect 390930 -25901 390998 -25845
rect 391054 -25901 391122 -25845
rect 391178 -25901 391246 -25845
rect 391302 -25901 391370 -25845
rect 391426 -25901 391494 -25845
rect 391550 -25901 391618 -25845
rect 391674 -25901 391742 -25845
rect 391798 -25901 391866 -25845
rect 391922 -25901 391990 -25845
rect 392046 -25901 392114 -25845
rect 392170 -25901 392238 -25845
rect 392294 -25901 392362 -25845
rect 392418 -25901 392486 -25845
rect 392542 -25901 392610 -25845
rect 392666 -25901 392734 -25845
rect 392790 -25901 392858 -25845
rect 392914 -25901 392982 -25845
rect 393038 -25901 393106 -25845
rect 393162 -25901 393230 -25845
rect 393286 -25901 393354 -25845
rect 393410 -25901 393478 -25845
rect 393534 -25901 393602 -25845
rect 393658 -25901 393726 -25845
rect 393782 -25901 393850 -25845
rect 393906 -25901 393974 -25845
rect 394030 -25901 394098 -25845
rect 394154 -25901 394222 -25845
rect 394278 -25901 394346 -25845
rect 394402 -25901 394470 -25845
rect 394526 -25901 394594 -25845
rect 394650 -25901 394718 -25845
rect 394774 -25901 394842 -25845
rect 394898 -25901 394966 -25845
rect 395022 -25901 395090 -25845
rect 395146 -25901 395214 -25845
rect 395270 -25901 395338 -25845
rect 395394 -25901 395462 -25845
rect 395518 -25901 395586 -25845
rect 395642 -25901 395710 -25845
rect 395766 -25901 395898 -25845
rect 395954 -25901 396022 -25845
rect 396078 -25901 396146 -25845
rect 396202 -25901 396270 -25845
rect 396326 -25901 396394 -25845
rect 396450 -25901 396518 -25845
rect 396574 -25901 396642 -25845
rect 396698 -25901 396766 -25845
rect 396822 -25901 396890 -25845
rect 396946 -25901 397014 -25845
rect 397070 -25901 397200 -25845
rect 388000 -25969 397200 -25901
rect 388000 -26025 388146 -25969
rect 388202 -26025 388270 -25969
rect 388326 -26025 388394 -25969
rect 388450 -26025 388518 -25969
rect 388574 -26025 388642 -25969
rect 388698 -26025 388766 -25969
rect 388822 -26025 388890 -25969
rect 388946 -26025 389014 -25969
rect 389070 -26025 389138 -25969
rect 389194 -26025 389262 -25969
rect 389318 -26025 389386 -25969
rect 389442 -26025 389510 -25969
rect 389566 -26025 389634 -25969
rect 389690 -26025 389758 -25969
rect 389814 -26025 389882 -25969
rect 389938 -26025 390006 -25969
rect 390062 -26025 390130 -25969
rect 390186 -26025 390254 -25969
rect 390310 -26025 390378 -25969
rect 390434 -26025 390502 -25969
rect 390558 -26025 390626 -25969
rect 390682 -26025 390750 -25969
rect 390806 -26025 390874 -25969
rect 390930 -26025 390998 -25969
rect 391054 -26025 391122 -25969
rect 391178 -26025 391246 -25969
rect 391302 -26025 391370 -25969
rect 391426 -26025 391494 -25969
rect 391550 -26025 391618 -25969
rect 391674 -26025 391742 -25969
rect 391798 -26025 391866 -25969
rect 391922 -26025 391990 -25969
rect 392046 -26025 392114 -25969
rect 392170 -26025 392238 -25969
rect 392294 -26025 392362 -25969
rect 392418 -26025 392486 -25969
rect 392542 -26025 392610 -25969
rect 392666 -26025 392734 -25969
rect 392790 -26025 392858 -25969
rect 392914 -26025 392982 -25969
rect 393038 -26025 393106 -25969
rect 393162 -26025 393230 -25969
rect 393286 -26025 393354 -25969
rect 393410 -26025 393478 -25969
rect 393534 -26025 393602 -25969
rect 393658 -26025 393726 -25969
rect 393782 -26025 393850 -25969
rect 393906 -26025 393974 -25969
rect 394030 -26025 394098 -25969
rect 394154 -26025 394222 -25969
rect 394278 -26025 394346 -25969
rect 394402 -26025 394470 -25969
rect 394526 -26025 394594 -25969
rect 394650 -26025 394718 -25969
rect 394774 -26025 394842 -25969
rect 394898 -26025 394966 -25969
rect 395022 -26025 395090 -25969
rect 395146 -26025 395214 -25969
rect 395270 -26025 395338 -25969
rect 395394 -26025 395462 -25969
rect 395518 -26025 395586 -25969
rect 395642 -26025 395710 -25969
rect 395766 -26025 395898 -25969
rect 395954 -26025 396022 -25969
rect 396078 -26025 396146 -25969
rect 396202 -26025 396270 -25969
rect 396326 -26025 396394 -25969
rect 396450 -26025 396518 -25969
rect 396574 -26025 396642 -25969
rect 396698 -26025 396766 -25969
rect 396822 -26025 396890 -25969
rect 396946 -26025 397014 -25969
rect 397070 -26025 397200 -25969
rect 388000 -26093 397200 -26025
rect 388000 -26149 388146 -26093
rect 388202 -26149 388270 -26093
rect 388326 -26149 388394 -26093
rect 388450 -26149 388518 -26093
rect 388574 -26149 388642 -26093
rect 388698 -26149 388766 -26093
rect 388822 -26149 388890 -26093
rect 388946 -26149 389014 -26093
rect 389070 -26149 389138 -26093
rect 389194 -26149 389262 -26093
rect 389318 -26149 389386 -26093
rect 389442 -26149 389510 -26093
rect 389566 -26149 389634 -26093
rect 389690 -26149 389758 -26093
rect 389814 -26149 389882 -26093
rect 389938 -26149 390006 -26093
rect 390062 -26149 390130 -26093
rect 390186 -26149 390254 -26093
rect 390310 -26149 390378 -26093
rect 390434 -26149 390502 -26093
rect 390558 -26149 390626 -26093
rect 390682 -26149 390750 -26093
rect 390806 -26149 390874 -26093
rect 390930 -26149 390998 -26093
rect 391054 -26149 391122 -26093
rect 391178 -26149 391246 -26093
rect 391302 -26149 391370 -26093
rect 391426 -26149 391494 -26093
rect 391550 -26149 391618 -26093
rect 391674 -26149 391742 -26093
rect 391798 -26149 391866 -26093
rect 391922 -26149 391990 -26093
rect 392046 -26149 392114 -26093
rect 392170 -26149 392238 -26093
rect 392294 -26149 392362 -26093
rect 392418 -26149 392486 -26093
rect 392542 -26149 392610 -26093
rect 392666 -26149 392734 -26093
rect 392790 -26149 392858 -26093
rect 392914 -26149 392982 -26093
rect 393038 -26149 393106 -26093
rect 393162 -26149 393230 -26093
rect 393286 -26149 393354 -26093
rect 393410 -26149 393478 -26093
rect 393534 -26149 393602 -26093
rect 393658 -26149 393726 -26093
rect 393782 -26149 393850 -26093
rect 393906 -26149 393974 -26093
rect 394030 -26149 394098 -26093
rect 394154 -26149 394222 -26093
rect 394278 -26149 394346 -26093
rect 394402 -26149 394470 -26093
rect 394526 -26149 394594 -26093
rect 394650 -26149 394718 -26093
rect 394774 -26149 394842 -26093
rect 394898 -26149 394966 -26093
rect 395022 -26149 395090 -26093
rect 395146 -26149 395214 -26093
rect 395270 -26149 395338 -26093
rect 395394 -26149 395462 -26093
rect 395518 -26149 395586 -26093
rect 395642 -26149 395710 -26093
rect 395766 -26149 395898 -26093
rect 395954 -26149 396022 -26093
rect 396078 -26149 396146 -26093
rect 396202 -26149 396270 -26093
rect 396326 -26149 396394 -26093
rect 396450 -26149 396518 -26093
rect 396574 -26149 396642 -26093
rect 396698 -26149 396766 -26093
rect 396822 -26149 396890 -26093
rect 396946 -26149 397014 -26093
rect 397070 -26149 397200 -26093
rect 388000 -26270 397200 -26149
<< glass >>
rect 388800 -25600 396400 -17740
<< comment >>
rect 397220 -26270 397230 -17070
rect 388000 -26300 397200 -26290
rect 397110 -26330 397120 -26310
rect 397130 -26330 397140 -26310
rect 397110 -26340 397140 -26330
rect 397130 -26360 397140 -26340
rect 397150 -26320 397180 -26310
rect 397150 -26330 397160 -26320
rect 397150 -26340 397180 -26330
rect 397150 -26350 397160 -26340
rect 397170 -26350 397180 -26340
rect 397150 -26360 397180 -26350
rect 388800 -26400 396400 -26390
rect 396330 -26420 396360 -26410
rect 396350 -26430 396360 -26420
rect 396340 -26440 396360 -26430
rect 396350 -26450 396360 -26440
rect 396330 -26460 396360 -26450
rect 396370 -26420 396400 -26410
rect 396370 -26430 396380 -26420
rect 396390 -26430 396400 -26420
rect 396370 -26440 396400 -26430
rect 396370 -26450 396380 -26440
rect 396390 -26450 396400 -26440
rect 396370 -26460 396400 -26450
<< labels >>
rlabel metal5 s 392300 -22000 397300 -17000 4 PAD
port 7 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 778000 1020000
<< end >>
