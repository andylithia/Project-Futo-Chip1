VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO filterstage
  CLASS BLOCK ;
  FOREIGN filterstage ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 100.000 ;
  PIN nbusin_nshunt
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.480 4.000 75.040 ;
    END
  END nbusin_nshunt
  PIN nbusout
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 74.480 120.000 75.040 ;
    END
  END nbusout
  PIN nseries_gy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END nseries_gy
  PIN nseries_gygy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.640 0.000 109.200 4.000 ;
    END
  END nseries_gygy
  PIN nshunt_gy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END nshunt_gy
  PIN pbusin_pshunt
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 4.000 25.200 ;
    END
  END pbusin_pshunt
  PIN pbusout
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 116.000 24.640 120.000 25.200 ;
    END
  END pbusout
  PIN pseries_gy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.840 0.000 50.400 4.000 ;
    END
  END pseries_gy
  PIN pseries_gygy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.040 0.000 89.600 4.000 ;
    END
  END pseries_gygy
  PIN pshunt_gy
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.640 0.000 11.200 4.000 ;
    END
  END pshunt_gy
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.220 15.380 20.820 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 45.820 15.380 47.420 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 72.420 15.380 74.020 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.020 15.380 100.620 82.620 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 32.520 15.380 34.120 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 59.120 15.380 60.720 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 85.720 15.380 87.320 82.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 112.320 15.380 113.920 82.620 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 113.920 82.620 ;
      LAYER Metal2 ;
        RECT 10.220 4.300 113.780 82.510 ;
        RECT 10.220 4.000 10.340 4.300 ;
        RECT 11.500 4.000 29.940 4.300 ;
        RECT 31.100 4.000 49.540 4.300 ;
        RECT 50.700 4.000 69.140 4.300 ;
        RECT 70.300 4.000 88.740 4.300 ;
        RECT 89.900 4.000 108.340 4.300 ;
        RECT 109.500 4.000 113.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 75.340 116.000 82.460 ;
        RECT 4.300 74.180 115.700 75.340 ;
        RECT 4.000 25.500 116.000 74.180 ;
        RECT 4.300 24.340 115.700 25.500 ;
        RECT 4.000 15.540 116.000 24.340 ;
  END
END filterstage
END LIBRARY

