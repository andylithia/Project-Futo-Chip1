* NGSPICE file created from shiftreg.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

.subckt shiftreg latch sclk sdin sr_out tune_s1_series_gy[0] tune_s1_series_gy[1]
+ tune_s1_series_gy[2] tune_s1_series_gy[3] tune_s1_series_gy[4] tune_s1_series_gy[5]
+ tune_s1_series_gygy[0] tune_s1_series_gygy[1] tune_s1_series_gygy[2] tune_s1_series_gygy[3]
+ tune_s1_series_gygy[4] tune_s1_series_gygy[5] tune_s1_shunt[0] tune_s1_shunt[1]
+ tune_s1_shunt[2] tune_s1_shunt[3] tune_s1_shunt[4] tune_s1_shunt[5] tune_s1_shunt[6]
+ tune_s1_shunt[7] tune_s1_shunt_gy[0] tune_s1_shunt_gy[1] tune_s1_shunt_gy[2] tune_s1_shunt_gy[3]
+ tune_s1_shunt_gy[4] tune_s1_shunt_gy[5] tune_s1_shunt_gy[6] tune_s2_series_gy[0]
+ tune_s2_series_gy[1] tune_s2_series_gy[2] tune_s2_series_gy[3] tune_s2_series_gy[4]
+ tune_s2_series_gy[5] tune_s2_series_gy[6] tune_s2_series_gy[7] tune_s2_series_gygy[0]
+ tune_s2_series_gygy[1] tune_s2_series_gygy[2] tune_s2_series_gygy[3] tune_s2_series_gygy[4]
+ tune_s2_series_gygy[5] tune_s2_series_gygy[6] tune_s2_series_gygy[7] tune_s2_shunt[0]
+ tune_s2_shunt[10] tune_s2_shunt[1] tune_s2_shunt[2] tune_s2_shunt[3] tune_s2_shunt[4]
+ tune_s2_shunt[5] tune_s2_shunt[6] tune_s2_shunt[7] tune_s2_shunt[8] tune_s2_shunt[9]
+ tune_s2_shunt_gy[0] tune_s2_shunt_gy[1] tune_s2_shunt_gy[2] tune_s2_shunt_gy[3]
+ tune_s2_shunt_gy[4] vdd vss
XFILLER_3_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_062_ sr\[20\] clknet_3_3__leaf_sclk sr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_114_ sr\[14\] latch tune_s1_shunt_gy[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_045_ sr\[3\] clknet_3_3__leaf_sclk sr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_028_ sr\[46\] latch tune_s2_series_gy[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_061_ sr\[19\] clknet_3_3__leaf_sclk sr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_044_ sr\[2\] clknet_3_0__leaf_sclk sr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_113_ sr\[13\] latch tune_s1_shunt_gy[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_027_ sr\[45\] latch tune_s2_series_gy[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_060_ sr\[18\] clknet_3_3__leaf_sclk sr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_112_ sr\[12\] latch tune_s1_shunt_gy[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_043_ sr\[1\] clknet_3_2__leaf_sclk sr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_026_ sr\[44\] latch tune_s2_series_gy[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_009_ sr\[27\] latch tune_s2_shunt[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_042_ sr\[0\] clknet_3_0__leaf_sclk sr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_111_ sr\[11\] latch tune_s1_shunt_gy[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_025_ sr\[43\] latch tune_s2_series_gy[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_008_ sr\[26\] latch tune_s1_series_gygy[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_041_ sdin clknet_3_0__leaf_sclk sr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_110_ sr\[10\] latch tune_s1_shunt_gy[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_024_ sr\[42\] latch tune_s2_shunt_gy[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_007_ sr\[25\] latch tune_s1_series_gygy[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_6__f_sclk clknet_0_sclk clknet_3_6__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_040_ sr_out latch tune_s2_series_gygy[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_023_ sr\[41\] latch tune_s2_shunt_gy[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_006_ sr\[24\] latch tune_s1_series_gygy[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_2__f_sclk clknet_0_sclk clknet_3_2__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_099_ sr\[57\] clknet_3_7__leaf_sclk sr_out vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_022_ sr\[40\] latch tune_s2_shunt_gy[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_005_ sr\[23\] latch tune_s1_series_gygy[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_098_ sr\[56\] clknet_3_5__leaf_sclk sr\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_021_ sr\[39\] latch tune_s2_shunt_gy[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_004_ sr\[22\] latch tune_s1_series_gygy[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_097_ sr\[55\] clknet_3_6__leaf_sclk sr\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_020_ sr\[38\] latch tune_s2_shunt_gy[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_003_ sr\[21\] latch tune_s1_series_gygy[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_096_ sr\[54\] clknet_3_4__leaf_sclk sr\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_079_ sr\[37\] clknet_3_6__leaf_sclk sr\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_002_ sr\[20\] latch tune_s1_series_gy[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_095_ sr\[53\] clknet_3_6__leaf_sclk sr\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_078_ sr\[36\] clknet_3_5__leaf_sclk sr\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_001_ sr\[19\] latch tune_s1_series_gy[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_094_ sr\[52\] clknet_3_7__leaf_sclk sr\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_077_ sr\[35\] clknet_3_6__leaf_sclk sr\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_000_ sr\[18\] latch tune_s1_series_gy[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_093_ sr\[51\] clknet_3_4__leaf_sclk sr\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_076_ sr\[34\] clknet_3_5__leaf_sclk sr\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_059_ sr\[17\] clknet_3_0__leaf_sclk sr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_092_ sr\[50\] clknet_3_4__leaf_sclk sr\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_075_ sr\[33\] clknet_3_4__leaf_sclk sr\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_058_ sr\[16\] clknet_3_3__leaf_sclk sr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_sclk clknet_0_sclk clknet_3_5__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_091_ sr\[49\] clknet_3_5__leaf_sclk sr\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_074_ sr\[32\] clknet_3_7__leaf_sclk sr\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_057_ sr\[15\] clknet_3_0__leaf_sclk sr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_109_ sr\[9\] latch tune_s1_shunt_gy[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_1__f_sclk clknet_0_sclk clknet_3_1__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_090_ sr\[48\] clknet_3_7__leaf_sclk sr\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_073_ sr\[31\] clknet_3_7__leaf_sclk sr\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_056_ sr\[14\] clknet_3_1__leaf_sclk sr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_039_ sr\[57\] latch tune_s2_series_gygy[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_108_ sr\[8\] latch tune_s1_shunt_gy[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_072_ sr\[30\] clknet_3_7__leaf_sclk sr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_055_ sr\[13\] clknet_3_1__leaf_sclk sr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_107_ sr\[7\] latch tune_s1_shunt[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_038_ sr\[56\] latch tune_s2_series_gygy[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_071_ sr\[29\] clknet_3_6__leaf_sclk sr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_054_ sr\[12\] clknet_3_1__leaf_sclk sr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_106_ sr\[6\] latch tune_s1_shunt[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_037_ sr\[55\] latch tune_s2_series_gygy[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_070_ sr\[28\] clknet_3_7__leaf_sclk sr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_053_ sr\[11\] clknet_3_2__leaf_sclk sr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_105_ sr\[5\] latch tune_s1_shunt[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_036_ sr\[54\] latch tune_s2_series_gygy[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_019_ sr\[37\] latch tune_s2_shunt[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_052_ sr\[10\] clknet_3_1__leaf_sclk sr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_035_ sr\[53\] latch tune_s2_series_gygy[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_104_ sr\[4\] latch tune_s1_shunt[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_018_ sr\[36\] latch tune_s2_shunt[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_051_ sr\[9\] clknet_3_2__leaf_sclk sr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_034_ sr\[52\] latch tune_s2_series_gygy[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_103_ sr\[3\] latch tune_s1_shunt[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_017_ sr\[35\] latch tune_s2_shunt[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_050_ sr\[8\] clknet_3_2__leaf_sclk sr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_033_ sr\[51\] latch tune_s2_series_gygy[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_102_ sr\[2\] latch tune_s1_shunt[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_016_ sr\[34\] latch tune_s2_shunt[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_032_ sr\[50\] latch tune_s2_series_gy[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_101_ sr\[1\] latch tune_s1_shunt[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_015_ sr\[33\] latch tune_s2_shunt[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_4__f_sclk clknet_0_sclk clknet_3_4__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_100_ sr\[0\] latch tune_s1_shunt[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_031_ sr\[49\] latch tune_s2_series_gy[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_014_ sr\[32\] latch tune_s2_shunt[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_0__f_sclk clknet_0_sclk clknet_3_0__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_030_ sr\[48\] latch tune_s2_series_gy[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_013_ sr\[31\] latch tune_s2_shunt[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_sclk sclk clknet_0_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_089_ sr\[47\] clknet_3_7__leaf_sclk sr\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_012_ sr\[30\] latch tune_s2_shunt[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_088_ sr\[46\] clknet_3_4__leaf_sclk sr\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_011_ sr\[29\] latch tune_s2_shunt[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_087_ sr\[45\] clknet_3_5__leaf_sclk sr\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_010_ sr\[28\] latch tune_s2_shunt[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_086_ sr\[44\] clknet_3_5__leaf_sclk sr\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_069_ sr\[27\] clknet_3_1__leaf_sclk sr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_085_ sr\[43\] clknet_3_7__leaf_sclk sr\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_068_ sr\[26\] clknet_3_3__leaf_sclk sr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_084_ sr\[42\] clknet_3_5__leaf_sclk sr\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_067_ sr\[25\] clknet_3_2__leaf_sclk sr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7__f_sclk clknet_0_sclk clknet_3_7__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_083_ sr\[41\] clknet_3_7__leaf_sclk sr\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_066_ sr\[24\] clknet_3_0__leaf_sclk sr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_049_ sr\[7\] clknet_3_3__leaf_sclk sr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_3__f_sclk clknet_0_sclk clknet_3_3__leaf_sclk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_082_ sr\[40\] clknet_3_6__leaf_sclk sr\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_065_ sr\[23\] clknet_3_3__leaf_sclk sr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_117_ sr\[17\] latch tune_s1_series_gy[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_048_ sr\[6\] clknet_3_3__leaf_sclk sr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_081_ sr\[39\] clknet_3_6__leaf_sclk sr\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_064_ sr\[22\] clknet_3_2__leaf_sclk sr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_116_ sr\[16\] latch tune_s1_series_gy[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_047_ sr\[5\] clknet_3_3__leaf_sclk sr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_080_ sr\[38\] clknet_3_6__leaf_sclk sr\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_063_ sr\[21\] clknet_3_0__leaf_sclk sr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_046_ sr\[4\] clknet_3_2__leaf_sclk sr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_115_ sr\[15\] latch tune_s1_series_gy[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_029_ sr\[47\] latch tune_s2_series_gy[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

