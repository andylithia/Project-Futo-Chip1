// This is the unpowered netlist.
module ringosc (Y);
 output Y;

 wire \con[0] ;
 wire \con[100] ;
 wire \con[101] ;
 wire \con[102] ;
 wire \con[103] ;
 wire \con[104] ;
 wire \con[105] ;
 wire \con[106] ;
 wire \con[107] ;
 wire \con[108] ;
 wire \con[109] ;
 wire \con[10] ;
 wire \con[110] ;
 wire \con[111] ;
 wire \con[112] ;
 wire \con[113] ;
 wire \con[114] ;
 wire \con[115] ;
 wire \con[116] ;
 wire \con[117] ;
 wire \con[118] ;
 wire \con[119] ;
 wire \con[11] ;
 wire \con[120] ;
 wire \con[121] ;
 wire \con[122] ;
 wire \con[123] ;
 wire \con[124] ;
 wire \con[125] ;
 wire \con[126] ;
 wire \con[12] ;
 wire \con[13] ;
 wire \con[14] ;
 wire \con[15] ;
 wire \con[16] ;
 wire \con[17] ;
 wire \con[18] ;
 wire \con[19] ;
 wire \con[1] ;
 wire \con[20] ;
 wire \con[21] ;
 wire \con[22] ;
 wire \con[23] ;
 wire \con[24] ;
 wire \con[25] ;
 wire \con[26] ;
 wire \con[27] ;
 wire \con[28] ;
 wire \con[29] ;
 wire \con[2] ;
 wire \con[30] ;
 wire \con[31] ;
 wire \con[32] ;
 wire \con[33] ;
 wire \con[34] ;
 wire \con[35] ;
 wire \con[36] ;
 wire \con[37] ;
 wire \con[38] ;
 wire \con[39] ;
 wire \con[3] ;
 wire \con[40] ;
 wire \con[41] ;
 wire \con[42] ;
 wire \con[43] ;
 wire \con[44] ;
 wire \con[45] ;
 wire \con[46] ;
 wire \con[47] ;
 wire \con[48] ;
 wire \con[49] ;
 wire \con[4] ;
 wire \con[50] ;
 wire \con[51] ;
 wire \con[52] ;
 wire \con[53] ;
 wire \con[54] ;
 wire \con[55] ;
 wire \con[56] ;
 wire \con[57] ;
 wire \con[58] ;
 wire \con[59] ;
 wire \con[5] ;
 wire \con[60] ;
 wire \con[61] ;
 wire \con[62] ;
 wire \con[63] ;
 wire \con[64] ;
 wire \con[65] ;
 wire \con[66] ;
 wire \con[67] ;
 wire \con[68] ;
 wire \con[69] ;
 wire \con[6] ;
 wire \con[70] ;
 wire \con[71] ;
 wire \con[72] ;
 wire \con[73] ;
 wire \con[74] ;
 wire \con[75] ;
 wire \con[76] ;
 wire \con[77] ;
 wire \con[78] ;
 wire \con[79] ;
 wire \con[7] ;
 wire \con[80] ;
 wire \con[81] ;
 wire \con[82] ;
 wire \con[83] ;
 wire \con[84] ;
 wire \con[85] ;
 wire \con[86] ;
 wire \con[87] ;
 wire \con[88] ;
 wire \con[89] ;
 wire \con[8] ;
 wire \con[90] ;
 wire \con[91] ;
 wire \con[92] ;
 wire \con[93] ;
 wire \con[94] ;
 wire \con[95] ;
 wire \con[96] ;
 wire \con[97] ;
 wire \con[98] ;
 wire \con[99] ;
 wire \con[9] ;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0_ (.I(Y),
    .Z(\con[125] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[0].u_uinv  (.I(\con[0] ),
    .ZN(\con[1] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[100].u_uinv  (.I(\con[100] ),
    .ZN(\con[101] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[101].u_uinv  (.I(\con[101] ),
    .ZN(\con[102] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[102].u_uinv  (.I(\con[102] ),
    .ZN(\con[103] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[103].u_uinv  (.I(\con[103] ),
    .ZN(\con[104] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[104].u_uinv  (.I(\con[104] ),
    .ZN(\con[105] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[105].u_uinv  (.I(\con[105] ),
    .ZN(\con[106] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[106].u_uinv  (.I(\con[106] ),
    .ZN(\con[107] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[107].u_uinv  (.I(\con[107] ),
    .ZN(\con[108] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[108].u_uinv  (.I(\con[108] ),
    .ZN(\con[109] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[109].u_uinv  (.I(\con[109] ),
    .ZN(\con[110] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[10].u_uinv  (.I(\con[10] ),
    .ZN(\con[11] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[110].u_uinv  (.I(\con[110] ),
    .ZN(\con[111] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[111].u_uinv  (.I(\con[111] ),
    .ZN(\con[112] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[112].u_uinv  (.I(\con[112] ),
    .ZN(\con[113] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[113].u_uinv  (.I(\con[113] ),
    .ZN(\con[114] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[114].u_uinv  (.I(\con[114] ),
    .ZN(\con[115] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[115].u_uinv  (.I(\con[115] ),
    .ZN(\con[116] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[116].u_uinv  (.I(\con[116] ),
    .ZN(\con[117] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[117].u_uinv  (.I(\con[117] ),
    .ZN(\con[118] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[118].u_uinv  (.I(\con[118] ),
    .ZN(\con[119] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[119].u_uinv  (.I(\con[119] ),
    .ZN(\con[120] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[11].u_uinv  (.I(\con[11] ),
    .ZN(\con[12] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[120].u_uinv  (.I(\con[120] ),
    .ZN(\con[121] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[121].u_uinv  (.I(\con[121] ),
    .ZN(\con[122] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[122].u_uinv  (.I(\con[122] ),
    .ZN(\con[123] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[123].u_uinv  (.I(\con[123] ),
    .ZN(\con[124] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[124].u_uinv  (.I(\con[124] ),
    .ZN(Y));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[125].u_uinv  (.I(Y),
    .ZN(\con[126] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[12].u_uinv  (.I(\con[12] ),
    .ZN(\con[13] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[13].u_uinv  (.I(\con[13] ),
    .ZN(\con[14] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[14].u_uinv  (.I(\con[14] ),
    .ZN(\con[15] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[15].u_uinv  (.I(\con[15] ),
    .ZN(\con[16] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[16].u_uinv  (.I(\con[16] ),
    .ZN(\con[17] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[17].u_uinv  (.I(\con[17] ),
    .ZN(\con[18] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[18].u_uinv  (.I(\con[18] ),
    .ZN(\con[19] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[19].u_uinv  (.I(\con[19] ),
    .ZN(\con[20] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[1].u_uinv  (.I(\con[1] ),
    .ZN(\con[2] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[20].u_uinv  (.I(\con[20] ),
    .ZN(\con[21] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[21].u_uinv  (.I(\con[21] ),
    .ZN(\con[22] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[22].u_uinv  (.I(\con[22] ),
    .ZN(\con[23] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[23].u_uinv  (.I(\con[23] ),
    .ZN(\con[24] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[24].u_uinv  (.I(\con[24] ),
    .ZN(\con[25] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[25].u_uinv  (.I(\con[25] ),
    .ZN(\con[26] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[26].u_uinv  (.I(\con[26] ),
    .ZN(\con[27] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[27].u_uinv  (.I(\con[27] ),
    .ZN(\con[28] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[28].u_uinv  (.I(\con[28] ),
    .ZN(\con[29] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[29].u_uinv  (.I(\con[29] ),
    .ZN(\con[30] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[2].u_uinv  (.I(\con[2] ),
    .ZN(\con[3] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[30].u_uinv  (.I(\con[30] ),
    .ZN(\con[31] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[31].u_uinv  (.I(\con[31] ),
    .ZN(\con[32] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[32].u_uinv  (.I(\con[32] ),
    .ZN(\con[33] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[33].u_uinv  (.I(\con[33] ),
    .ZN(\con[34] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[34].u_uinv  (.I(\con[34] ),
    .ZN(\con[35] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[35].u_uinv  (.I(\con[35] ),
    .ZN(\con[36] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[36].u_uinv  (.I(\con[36] ),
    .ZN(\con[37] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[37].u_uinv  (.I(\con[37] ),
    .ZN(\con[38] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[38].u_uinv  (.I(\con[38] ),
    .ZN(\con[39] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[39].u_uinv  (.I(\con[39] ),
    .ZN(\con[40] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[3].u_uinv  (.I(\con[3] ),
    .ZN(\con[4] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[40].u_uinv  (.I(\con[40] ),
    .ZN(\con[41] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[41].u_uinv  (.I(\con[41] ),
    .ZN(\con[42] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[42].u_uinv  (.I(\con[42] ),
    .ZN(\con[43] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[43].u_uinv  (.I(\con[43] ),
    .ZN(\con[44] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[44].u_uinv  (.I(\con[44] ),
    .ZN(\con[45] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[45].u_uinv  (.I(\con[45] ),
    .ZN(\con[46] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[46].u_uinv  (.I(\con[46] ),
    .ZN(\con[47] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[47].u_uinv  (.I(\con[47] ),
    .ZN(\con[48] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[48].u_uinv  (.I(\con[48] ),
    .ZN(\con[49] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[49].u_uinv  (.I(\con[49] ),
    .ZN(\con[50] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[4].u_uinv  (.I(\con[4] ),
    .ZN(\con[5] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[50].u_uinv  (.I(\con[50] ),
    .ZN(\con[51] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[51].u_uinv  (.I(\con[51] ),
    .ZN(\con[52] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[52].u_uinv  (.I(\con[52] ),
    .ZN(\con[53] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[53].u_uinv  (.I(\con[53] ),
    .ZN(\con[54] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[54].u_uinv  (.I(\con[54] ),
    .ZN(\con[55] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[55].u_uinv  (.I(\con[55] ),
    .ZN(\con[56] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[56].u_uinv  (.I(\con[56] ),
    .ZN(\con[57] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[57].u_uinv  (.I(\con[57] ),
    .ZN(\con[58] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[58].u_uinv  (.I(\con[58] ),
    .ZN(\con[59] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[59].u_uinv  (.I(\con[59] ),
    .ZN(\con[60] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[5].u_uinv  (.I(\con[5] ),
    .ZN(\con[6] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[60].u_uinv  (.I(\con[60] ),
    .ZN(\con[61] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[61].u_uinv  (.I(\con[61] ),
    .ZN(\con[62] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[62].u_uinv  (.I(\con[62] ),
    .ZN(\con[63] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[63].u_uinv  (.I(\con[63] ),
    .ZN(\con[64] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[64].u_uinv  (.I(\con[64] ),
    .ZN(\con[65] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[65].u_uinv  (.I(\con[65] ),
    .ZN(\con[66] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[66].u_uinv  (.I(\con[66] ),
    .ZN(\con[67] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[67].u_uinv  (.I(\con[67] ),
    .ZN(\con[68] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[68].u_uinv  (.I(\con[68] ),
    .ZN(\con[69] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[69].u_uinv  (.I(\con[69] ),
    .ZN(\con[70] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[6].u_uinv  (.I(\con[6] ),
    .ZN(\con[7] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[70].u_uinv  (.I(\con[70] ),
    .ZN(\con[71] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[71].u_uinv  (.I(\con[71] ),
    .ZN(\con[72] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[72].u_uinv  (.I(\con[72] ),
    .ZN(\con[73] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[73].u_uinv  (.I(\con[73] ),
    .ZN(\con[74] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[74].u_uinv  (.I(\con[74] ),
    .ZN(\con[75] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[75].u_uinv  (.I(\con[75] ),
    .ZN(\con[76] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[76].u_uinv  (.I(\con[76] ),
    .ZN(\con[77] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[77].u_uinv  (.I(\con[77] ),
    .ZN(\con[78] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[78].u_uinv  (.I(\con[78] ),
    .ZN(\con[79] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[79].u_uinv  (.I(\con[79] ),
    .ZN(\con[80] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[7].u_uinv  (.I(\con[7] ),
    .ZN(\con[8] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[80].u_uinv  (.I(\con[80] ),
    .ZN(\con[81] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[81].u_uinv  (.I(\con[81] ),
    .ZN(\con[82] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[82].u_uinv  (.I(\con[82] ),
    .ZN(\con[83] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[83].u_uinv  (.I(\con[83] ),
    .ZN(\con[84] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[84].u_uinv  (.I(\con[84] ),
    .ZN(\con[85] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[85].u_uinv  (.I(\con[85] ),
    .ZN(\con[86] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[86].u_uinv  (.I(\con[86] ),
    .ZN(\con[87] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[87].u_uinv  (.I(\con[87] ),
    .ZN(\con[88] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[88].u_uinv  (.I(\con[88] ),
    .ZN(\con[89] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[89].u_uinv  (.I(\con[89] ),
    .ZN(\con[90] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[8].u_uinv  (.I(\con[8] ),
    .ZN(\con[9] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[90].u_uinv  (.I(\con[90] ),
    .ZN(\con[91] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[91].u_uinv  (.I(\con[91] ),
    .ZN(\con[92] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[92].u_uinv  (.I(\con[92] ),
    .ZN(\con[93] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[93].u_uinv  (.I(\con[93] ),
    .ZN(\con[94] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[94].u_uinv  (.I(\con[94] ),
    .ZN(\con[95] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[95].u_uinv  (.I(\con[95] ),
    .ZN(\con[96] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[96].u_uinv  (.I(\con[96] ),
    .ZN(\con[97] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[97].u_uinv  (.I(\con[97] ),
    .ZN(\con[98] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[98].u_uinv  (.I(\con[98] ),
    .ZN(\con[99] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[99].u_uinv  (.I(\con[99] ),
    .ZN(\con[100] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \gen_ring[9].u_uinv  (.I(\con[9] ),
    .ZN(\con[10] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 u_uinv_init (.I(\con[126] ),
    .ZN(\con[0] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_98 ();
endmodule

