magic
tech gf180mcuC
magscale 1 5
timestamp 1669701303
<< obsm1 >>
rect 672 1538 9376 4342
<< metal2 >>
rect 4928 5600 4984 6000
rect 1400 0 1456 400
rect 1512 0 1568 400
rect 1624 0 1680 400
rect 1736 0 1792 400
rect 1848 0 1904 400
rect 1960 0 2016 400
rect 2072 0 2128 400
rect 2184 0 2240 400
rect 2296 0 2352 400
rect 2408 0 2464 400
rect 2520 0 2576 400
rect 2632 0 2688 400
rect 2744 0 2800 400
rect 2856 0 2912 400
rect 2968 0 3024 400
rect 3080 0 3136 400
rect 3192 0 3248 400
rect 3304 0 3360 400
rect 3416 0 3472 400
rect 3528 0 3584 400
rect 3640 0 3696 400
rect 3752 0 3808 400
rect 3864 0 3920 400
rect 3976 0 4032 400
rect 4088 0 4144 400
rect 4200 0 4256 400
rect 4312 0 4368 400
rect 4424 0 4480 400
rect 4536 0 4592 400
rect 4648 0 4704 400
rect 4760 0 4816 400
rect 4872 0 4928 400
rect 4984 0 5040 400
rect 5096 0 5152 400
rect 5208 0 5264 400
rect 5320 0 5376 400
rect 5432 0 5488 400
rect 5544 0 5600 400
rect 5656 0 5712 400
rect 5768 0 5824 400
rect 5880 0 5936 400
rect 5992 0 6048 400
rect 6104 0 6160 400
rect 6216 0 6272 400
rect 6328 0 6384 400
rect 6440 0 6496 400
rect 6552 0 6608 400
rect 6664 0 6720 400
rect 6776 0 6832 400
rect 6888 0 6944 400
rect 7000 0 7056 400
rect 7112 0 7168 400
rect 7224 0 7280 400
rect 7336 0 7392 400
rect 7448 0 7504 400
rect 7560 0 7616 400
rect 7672 0 7728 400
rect 7784 0 7840 400
rect 7896 0 7952 400
rect 8008 0 8064 400
rect 8120 0 8176 400
rect 8232 0 8288 400
rect 8344 0 8400 400
rect 8456 0 8512 400
<< obsm2 >>
rect 1078 5570 4898 5600
rect 5014 5570 9362 5600
rect 1078 430 9362 5570
rect 1078 400 1370 430
rect 8542 400 9362 430
<< obsm3 >>
rect 1073 1022 9367 4326
<< metal4 >>
rect 1670 1538 1830 4342
rect 2748 1538 2908 4342
rect 3826 1538 3986 4342
rect 4904 1538 5064 4342
rect 5982 1538 6142 4342
rect 7060 1538 7220 4342
rect 8138 1538 8298 4342
rect 9216 1538 9376 4342
<< obsm4 >>
rect 2086 1577 2718 3351
rect 2938 1577 3796 3351
rect 4016 1577 4874 3351
rect 5094 1577 5952 3351
rect 6172 1577 7030 3351
rect 7250 1577 7378 3351
<< labels >>
rlabel metal2 s 4928 5600 4984 6000 6 cap
port 1 nsew signal bidirectional
rlabel metal2 s 1400 0 1456 400 6 tune[0]
port 2 nsew signal input
rlabel metal2 s 2520 0 2576 400 6 tune[10]
port 3 nsew signal input
rlabel metal2 s 2632 0 2688 400 6 tune[11]
port 4 nsew signal input
rlabel metal2 s 2744 0 2800 400 6 tune[12]
port 5 nsew signal input
rlabel metal2 s 2856 0 2912 400 6 tune[13]
port 6 nsew signal input
rlabel metal2 s 2968 0 3024 400 6 tune[14]
port 7 nsew signal input
rlabel metal2 s 3080 0 3136 400 6 tune[15]
port 8 nsew signal input
rlabel metal2 s 3192 0 3248 400 6 tune[16]
port 9 nsew signal input
rlabel metal2 s 3304 0 3360 400 6 tune[17]
port 10 nsew signal input
rlabel metal2 s 3416 0 3472 400 6 tune[18]
port 11 nsew signal input
rlabel metal2 s 3528 0 3584 400 6 tune[19]
port 12 nsew signal input
rlabel metal2 s 1512 0 1568 400 6 tune[1]
port 13 nsew signal input
rlabel metal2 s 3640 0 3696 400 6 tune[20]
port 14 nsew signal input
rlabel metal2 s 3752 0 3808 400 6 tune[21]
port 15 nsew signal input
rlabel metal2 s 3864 0 3920 400 6 tune[22]
port 16 nsew signal input
rlabel metal2 s 3976 0 4032 400 6 tune[23]
port 17 nsew signal input
rlabel metal2 s 4088 0 4144 400 6 tune[24]
port 18 nsew signal input
rlabel metal2 s 4200 0 4256 400 6 tune[25]
port 19 nsew signal input
rlabel metal2 s 4312 0 4368 400 6 tune[26]
port 20 nsew signal input
rlabel metal2 s 4424 0 4480 400 6 tune[27]
port 21 nsew signal input
rlabel metal2 s 4536 0 4592 400 6 tune[28]
port 22 nsew signal input
rlabel metal2 s 4648 0 4704 400 6 tune[29]
port 23 nsew signal input
rlabel metal2 s 1624 0 1680 400 6 tune[2]
port 24 nsew signal input
rlabel metal2 s 4760 0 4816 400 6 tune[30]
port 25 nsew signal input
rlabel metal2 s 4872 0 4928 400 6 tune[31]
port 26 nsew signal input
rlabel metal2 s 4984 0 5040 400 6 tune[32]
port 27 nsew signal input
rlabel metal2 s 5096 0 5152 400 6 tune[33]
port 28 nsew signal input
rlabel metal2 s 5208 0 5264 400 6 tune[34]
port 29 nsew signal input
rlabel metal2 s 5320 0 5376 400 6 tune[35]
port 30 nsew signal input
rlabel metal2 s 5432 0 5488 400 6 tune[36]
port 31 nsew signal input
rlabel metal2 s 5544 0 5600 400 6 tune[37]
port 32 nsew signal input
rlabel metal2 s 5656 0 5712 400 6 tune[38]
port 33 nsew signal input
rlabel metal2 s 5768 0 5824 400 6 tune[39]
port 34 nsew signal input
rlabel metal2 s 1736 0 1792 400 6 tune[3]
port 35 nsew signal input
rlabel metal2 s 5880 0 5936 400 6 tune[40]
port 36 nsew signal input
rlabel metal2 s 5992 0 6048 400 6 tune[41]
port 37 nsew signal input
rlabel metal2 s 6104 0 6160 400 6 tune[42]
port 38 nsew signal input
rlabel metal2 s 6216 0 6272 400 6 tune[43]
port 39 nsew signal input
rlabel metal2 s 6328 0 6384 400 6 tune[44]
port 40 nsew signal input
rlabel metal2 s 6440 0 6496 400 6 tune[45]
port 41 nsew signal input
rlabel metal2 s 6552 0 6608 400 6 tune[46]
port 42 nsew signal input
rlabel metal2 s 6664 0 6720 400 6 tune[47]
port 43 nsew signal input
rlabel metal2 s 6776 0 6832 400 6 tune[48]
port 44 nsew signal input
rlabel metal2 s 6888 0 6944 400 6 tune[49]
port 45 nsew signal input
rlabel metal2 s 1848 0 1904 400 6 tune[4]
port 46 nsew signal input
rlabel metal2 s 7000 0 7056 400 6 tune[50]
port 47 nsew signal input
rlabel metal2 s 7112 0 7168 400 6 tune[51]
port 48 nsew signal input
rlabel metal2 s 7224 0 7280 400 6 tune[52]
port 49 nsew signal input
rlabel metal2 s 7336 0 7392 400 6 tune[53]
port 50 nsew signal input
rlabel metal2 s 7448 0 7504 400 6 tune[54]
port 51 nsew signal input
rlabel metal2 s 7560 0 7616 400 6 tune[55]
port 52 nsew signal input
rlabel metal2 s 7672 0 7728 400 6 tune[56]
port 53 nsew signal input
rlabel metal2 s 7784 0 7840 400 6 tune[57]
port 54 nsew signal input
rlabel metal2 s 7896 0 7952 400 6 tune[58]
port 55 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 tune[59]
port 56 nsew signal input
rlabel metal2 s 1960 0 2016 400 6 tune[5]
port 57 nsew signal input
rlabel metal2 s 8120 0 8176 400 6 tune[60]
port 58 nsew signal input
rlabel metal2 s 8232 0 8288 400 6 tune[61]
port 59 nsew signal input
rlabel metal2 s 8344 0 8400 400 6 tune[62]
port 60 nsew signal input
rlabel metal2 s 8456 0 8512 400 6 tune[63]
port 61 nsew signal input
rlabel metal2 s 2072 0 2128 400 6 tune[6]
port 62 nsew signal input
rlabel metal2 s 2184 0 2240 400 6 tune[7]
port 63 nsew signal input
rlabel metal2 s 2296 0 2352 400 6 tune[8]
port 64 nsew signal input
rlabel metal2 s 2408 0 2464 400 6 tune[9]
port 65 nsew signal input
rlabel metal4 s 1670 1538 1830 4342 6 vdd
port 66 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 4342 6 vdd
port 66 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 4342 6 vdd
port 66 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 4342 6 vdd
port 66 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 4342 6 vss
port 67 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 4342 6 vss
port 67 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 4342 6 vss
port 67 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 4342 6 vss
port 67 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10000 6000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 162932
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/captune_1p/runs/22_11_29_00_54/results/signoff/captune_1p.magic.gds
string GDS_START 30122
<< end >>

