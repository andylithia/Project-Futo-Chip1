magic
tech gf180mcuC
magscale 1 10
timestamp 1669699727
<< metal1 >>
rect 1344 16490 22624 16524
rect 1344 16438 3874 16490
rect 3926 16438 3978 16490
rect 4030 16438 4082 16490
rect 4134 16438 9194 16490
rect 9246 16438 9298 16490
rect 9350 16438 9402 16490
rect 9454 16438 14514 16490
rect 14566 16438 14618 16490
rect 14670 16438 14722 16490
rect 14774 16438 19834 16490
rect 19886 16438 19938 16490
rect 19990 16438 20042 16490
rect 20094 16438 22624 16490
rect 1344 16404 22624 16438
rect 1344 15706 22784 15740
rect 1344 15654 6534 15706
rect 6586 15654 6638 15706
rect 6690 15654 6742 15706
rect 6794 15654 11854 15706
rect 11906 15654 11958 15706
rect 12010 15654 12062 15706
rect 12114 15654 17174 15706
rect 17226 15654 17278 15706
rect 17330 15654 17382 15706
rect 17434 15654 22494 15706
rect 22546 15654 22598 15706
rect 22650 15654 22702 15706
rect 22754 15654 22784 15706
rect 1344 15620 22784 15654
rect 1344 14922 22624 14956
rect 1344 14870 3874 14922
rect 3926 14870 3978 14922
rect 4030 14870 4082 14922
rect 4134 14870 9194 14922
rect 9246 14870 9298 14922
rect 9350 14870 9402 14922
rect 9454 14870 14514 14922
rect 14566 14870 14618 14922
rect 14670 14870 14722 14922
rect 14774 14870 19834 14922
rect 19886 14870 19938 14922
rect 19990 14870 20042 14922
rect 20094 14870 22624 14922
rect 1344 14836 22624 14870
rect 16830 14642 16882 14654
rect 16830 14578 16882 14590
rect 16942 14418 16994 14430
rect 16942 14354 16994 14366
rect 17614 14418 17666 14430
rect 17614 14354 17666 14366
rect 17502 14306 17554 14318
rect 17502 14242 17554 14254
rect 1344 14138 22784 14172
rect 1344 14086 6534 14138
rect 6586 14086 6638 14138
rect 6690 14086 6742 14138
rect 6794 14086 11854 14138
rect 11906 14086 11958 14138
rect 12010 14086 12062 14138
rect 12114 14086 17174 14138
rect 17226 14086 17278 14138
rect 17330 14086 17382 14138
rect 17434 14086 22494 14138
rect 22546 14086 22598 14138
rect 22650 14086 22702 14138
rect 22754 14086 22784 14138
rect 1344 14052 22784 14086
rect 16158 13746 16210 13758
rect 16158 13682 16210 13694
rect 16830 13746 16882 13758
rect 16830 13682 16882 13694
rect 17726 13746 17778 13758
rect 17726 13682 17778 13694
rect 18398 13746 18450 13758
rect 18398 13682 18450 13694
rect 16270 13522 16322 13534
rect 16270 13458 16322 13470
rect 16942 13522 16994 13534
rect 16942 13458 16994 13470
rect 17838 13522 17890 13534
rect 17838 13458 17890 13470
rect 18510 13522 18562 13534
rect 18510 13458 18562 13470
rect 1344 13354 22624 13388
rect 1344 13302 3874 13354
rect 3926 13302 3978 13354
rect 4030 13302 4082 13354
rect 4134 13302 9194 13354
rect 9246 13302 9298 13354
rect 9350 13302 9402 13354
rect 9454 13302 14514 13354
rect 14566 13302 14618 13354
rect 14670 13302 14722 13354
rect 14774 13302 19834 13354
rect 19886 13302 19938 13354
rect 19990 13302 20042 13354
rect 20094 13302 22624 13354
rect 1344 13268 22624 13302
rect 14926 13186 14978 13198
rect 14926 13122 14978 13134
rect 18286 13186 18338 13198
rect 18286 13122 18338 13134
rect 18958 13186 19010 13198
rect 18958 13122 19010 13134
rect 17502 12962 17554 12974
rect 17502 12898 17554 12910
rect 18846 12962 18898 12974
rect 18846 12898 18898 12910
rect 14814 12850 14866 12862
rect 14814 12786 14866 12798
rect 15486 12850 15538 12862
rect 15486 12786 15538 12798
rect 16158 12850 16210 12862
rect 16158 12786 16210 12798
rect 16830 12850 16882 12862
rect 16830 12786 16882 12798
rect 18174 12850 18226 12862
rect 18174 12786 18226 12798
rect 19518 12850 19570 12862
rect 19518 12786 19570 12798
rect 15598 12738 15650 12750
rect 15598 12674 15650 12686
rect 16270 12738 16322 12750
rect 16270 12674 16322 12686
rect 16942 12738 16994 12750
rect 16942 12674 16994 12686
rect 17614 12738 17666 12750
rect 17614 12674 17666 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 1344 12570 22784 12604
rect 1344 12518 6534 12570
rect 6586 12518 6638 12570
rect 6690 12518 6742 12570
rect 6794 12518 11854 12570
rect 11906 12518 11958 12570
rect 12010 12518 12062 12570
rect 12114 12518 17174 12570
rect 17226 12518 17278 12570
rect 17330 12518 17382 12570
rect 17434 12518 22494 12570
rect 22546 12518 22598 12570
rect 22650 12518 22702 12570
rect 22754 12518 22784 12570
rect 1344 12484 22784 12518
rect 19182 12402 19234 12414
rect 19182 12338 19234 12350
rect 19854 12402 19906 12414
rect 19854 12338 19906 12350
rect 17726 12290 17778 12302
rect 17726 12226 17778 12238
rect 17838 12290 17890 12302
rect 17838 12226 17890 12238
rect 18398 12290 18450 12302
rect 18398 12226 18450 12238
rect 19070 12290 19122 12302
rect 19070 12226 19122 12238
rect 19742 12290 19794 12302
rect 19742 12226 19794 12238
rect 20414 12290 20466 12302
rect 20414 12226 20466 12238
rect 20526 12290 20578 12302
rect 20526 12226 20578 12238
rect 14142 12178 14194 12190
rect 14142 12114 14194 12126
rect 14814 12178 14866 12190
rect 14814 12114 14866 12126
rect 15486 12178 15538 12190
rect 15486 12114 15538 12126
rect 16158 12178 16210 12190
rect 16158 12114 16210 12126
rect 16830 12178 16882 12190
rect 16830 12114 16882 12126
rect 14254 11954 14306 11966
rect 14254 11890 14306 11902
rect 14926 11954 14978 11966
rect 14926 11890 14978 11902
rect 15598 11954 15650 11966
rect 15598 11890 15650 11902
rect 16270 11954 16322 11966
rect 16270 11890 16322 11902
rect 16942 11954 16994 11966
rect 16942 11890 16994 11902
rect 18510 11954 18562 11966
rect 18510 11890 18562 11902
rect 1344 11786 22624 11820
rect 1344 11734 3874 11786
rect 3926 11734 3978 11786
rect 4030 11734 4082 11786
rect 4134 11734 9194 11786
rect 9246 11734 9298 11786
rect 9350 11734 9402 11786
rect 9454 11734 14514 11786
rect 14566 11734 14618 11786
rect 14670 11734 14722 11786
rect 14774 11734 19834 11786
rect 19886 11734 19938 11786
rect 19990 11734 20042 11786
rect 20094 11734 22624 11786
rect 1344 11700 22624 11734
rect 17614 11618 17666 11630
rect 17614 11554 17666 11566
rect 19630 11618 19682 11630
rect 19630 11554 19682 11566
rect 10670 11506 10722 11518
rect 10670 11442 10722 11454
rect 14926 11394 14978 11406
rect 14926 11330 14978 11342
rect 15598 11394 15650 11406
rect 15598 11330 15650 11342
rect 16270 11394 16322 11406
rect 16270 11330 16322 11342
rect 16830 11394 16882 11406
rect 16830 11330 16882 11342
rect 16942 11394 16994 11406
rect 16942 11330 16994 11342
rect 17502 11394 17554 11406
rect 17502 11330 17554 11342
rect 18174 11394 18226 11406
rect 18174 11330 18226 11342
rect 18846 11394 18898 11406
rect 18846 11330 18898 11342
rect 19518 11394 19570 11406
rect 19518 11330 19570 11342
rect 6078 11282 6130 11294
rect 6078 11218 6130 11230
rect 6190 11282 6242 11294
rect 6190 11218 6242 11230
rect 6974 11282 7026 11294
rect 6974 11218 7026 11230
rect 7646 11282 7698 11294
rect 7646 11218 7698 11230
rect 8318 11282 8370 11294
rect 8318 11218 8370 11230
rect 9214 11282 9266 11294
rect 9214 11218 9266 11230
rect 9886 11282 9938 11294
rect 9886 11218 9938 11230
rect 10558 11282 10610 11294
rect 10558 11218 10610 11230
rect 12126 11282 12178 11294
rect 12126 11218 12178 11230
rect 12238 11282 12290 11294
rect 12238 11218 12290 11230
rect 12798 11282 12850 11294
rect 12798 11218 12850 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 14814 11282 14866 11294
rect 14814 11218 14866 11230
rect 15486 11282 15538 11294
rect 15486 11218 15538 11230
rect 16158 11282 16210 11294
rect 16158 11218 16210 11230
rect 20190 11282 20242 11294
rect 20190 11218 20242 11230
rect 6862 11170 6914 11182
rect 6862 11106 6914 11118
rect 7534 11170 7586 11182
rect 7534 11106 7586 11118
rect 8206 11170 8258 11182
rect 8206 11106 8258 11118
rect 9326 11170 9378 11182
rect 9326 11106 9378 11118
rect 9998 11170 10050 11182
rect 9998 11106 10050 11118
rect 12910 11170 12962 11182
rect 12910 11106 12962 11118
rect 13806 11170 13858 11182
rect 13806 11106 13858 11118
rect 18286 11170 18338 11182
rect 18286 11106 18338 11118
rect 18958 11170 19010 11182
rect 18958 11106 19010 11118
rect 20302 11170 20354 11182
rect 20302 11106 20354 11118
rect 1344 11002 22784 11036
rect 1344 10950 6534 11002
rect 6586 10950 6638 11002
rect 6690 10950 6742 11002
rect 6794 10950 11854 11002
rect 11906 10950 11958 11002
rect 12010 10950 12062 11002
rect 12114 10950 17174 11002
rect 17226 10950 17278 11002
rect 17330 10950 17382 11002
rect 17434 10950 22494 11002
rect 22546 10950 22598 11002
rect 22650 10950 22702 11002
rect 22754 10950 22784 11002
rect 1344 10916 22784 10950
rect 6862 10834 6914 10846
rect 6862 10770 6914 10782
rect 19182 10834 19234 10846
rect 19182 10770 19234 10782
rect 19854 10834 19906 10846
rect 19854 10770 19906 10782
rect 5406 10722 5458 10734
rect 5406 10658 5458 10670
rect 5518 10722 5570 10734
rect 5518 10658 5570 10670
rect 6078 10722 6130 10734
rect 6078 10658 6130 10670
rect 8094 10722 8146 10734
rect 8094 10658 8146 10670
rect 16718 10722 16770 10734
rect 16718 10658 16770 10670
rect 17726 10722 17778 10734
rect 17726 10658 17778 10670
rect 18398 10722 18450 10734
rect 18398 10658 18450 10670
rect 19070 10722 19122 10734
rect 19070 10658 19122 10670
rect 19742 10722 19794 10734
rect 19742 10658 19794 10670
rect 20414 10722 20466 10734
rect 20414 10658 20466 10670
rect 21086 10722 21138 10734
rect 21086 10658 21138 10670
rect 21758 10722 21810 10734
rect 21758 10658 21810 10670
rect 21870 10722 21922 10734
rect 21870 10658 21922 10670
rect 6750 10610 6802 10622
rect 6750 10546 6802 10558
rect 7422 10610 7474 10622
rect 7422 10546 7474 10558
rect 7534 10610 7586 10622
rect 7534 10546 7586 10558
rect 8878 10610 8930 10622
rect 8878 10546 8930 10558
rect 9886 10610 9938 10622
rect 9886 10546 9938 10558
rect 10558 10610 10610 10622
rect 10558 10546 10610 10558
rect 11230 10610 11282 10622
rect 11230 10546 11282 10558
rect 12014 10610 12066 10622
rect 12014 10546 12066 10558
rect 12686 10610 12738 10622
rect 12686 10546 12738 10558
rect 12798 10610 12850 10622
rect 12798 10546 12850 10558
rect 13358 10610 13410 10622
rect 13358 10546 13410 10558
rect 13470 10610 13522 10622
rect 13470 10546 13522 10558
rect 14030 10610 14082 10622
rect 14030 10546 14082 10558
rect 14142 10610 14194 10622
rect 14142 10546 14194 10558
rect 14702 10610 14754 10622
rect 14702 10546 14754 10558
rect 14814 10610 14866 10622
rect 14814 10546 14866 10558
rect 15374 10610 15426 10622
rect 15374 10546 15426 10558
rect 15486 10610 15538 10622
rect 15486 10546 15538 10558
rect 16046 10610 16098 10622
rect 16046 10546 16098 10558
rect 6190 10386 6242 10398
rect 6190 10322 6242 10334
rect 8206 10386 8258 10398
rect 8206 10322 8258 10334
rect 8990 10386 9042 10398
rect 8990 10322 9042 10334
rect 9998 10386 10050 10398
rect 9998 10322 10050 10334
rect 10670 10386 10722 10398
rect 10670 10322 10722 10334
rect 11342 10386 11394 10398
rect 11342 10322 11394 10334
rect 12126 10386 12178 10398
rect 12126 10322 12178 10334
rect 16158 10386 16210 10398
rect 16158 10322 16210 10334
rect 16830 10386 16882 10398
rect 16830 10322 16882 10334
rect 17838 10386 17890 10398
rect 17838 10322 17890 10334
rect 18510 10386 18562 10398
rect 18510 10322 18562 10334
rect 20526 10386 20578 10398
rect 20526 10322 20578 10334
rect 21198 10386 21250 10398
rect 21198 10322 21250 10334
rect 1344 10218 22624 10252
rect 1344 10166 3874 10218
rect 3926 10166 3978 10218
rect 4030 10166 4082 10218
rect 4134 10166 9194 10218
rect 9246 10166 9298 10218
rect 9350 10166 9402 10218
rect 9454 10166 14514 10218
rect 14566 10166 14618 10218
rect 14670 10166 14722 10218
rect 14774 10166 19834 10218
rect 19886 10166 19938 10218
rect 19990 10166 20042 10218
rect 20094 10166 22624 10218
rect 1344 10132 22624 10166
rect 11566 10050 11618 10062
rect 11566 9986 11618 9998
rect 18510 10050 18562 10062
rect 18510 9986 18562 9998
rect 20526 10050 20578 10062
rect 20526 9986 20578 9998
rect 21758 10050 21810 10062
rect 21758 9986 21810 9998
rect 4174 9826 4226 9838
rect 4174 9762 4226 9774
rect 4286 9826 4338 9838
rect 4286 9762 4338 9774
rect 4846 9826 4898 9838
rect 4846 9762 4898 9774
rect 7870 9826 7922 9838
rect 7870 9762 7922 9774
rect 8542 9826 8594 9838
rect 8542 9762 8594 9774
rect 9214 9826 9266 9838
rect 9214 9762 9266 9774
rect 10558 9826 10610 9838
rect 10558 9762 10610 9774
rect 12126 9826 12178 9838
rect 12126 9762 12178 9774
rect 12238 9826 12290 9838
rect 12238 9762 12290 9774
rect 14478 9826 14530 9838
rect 14478 9762 14530 9774
rect 15038 9826 15090 9838
rect 15038 9762 15090 9774
rect 15710 9826 15762 9838
rect 15710 9762 15762 9774
rect 17838 9826 17890 9838
rect 17838 9762 17890 9774
rect 19070 9826 19122 9838
rect 19070 9762 19122 9774
rect 19742 9826 19794 9838
rect 19742 9762 19794 9774
rect 20414 9826 20466 9838
rect 20414 9762 20466 9774
rect 21646 9826 21698 9838
rect 21646 9762 21698 9774
rect 5854 9714 5906 9726
rect 5854 9650 5906 9662
rect 6526 9714 6578 9726
rect 6526 9650 6578 9662
rect 6638 9714 6690 9726
rect 6638 9650 6690 9662
rect 7198 9714 7250 9726
rect 7198 9650 7250 9662
rect 7310 9714 7362 9726
rect 7310 9650 7362 9662
rect 9886 9714 9938 9726
rect 9886 9650 9938 9662
rect 11454 9714 11506 9726
rect 11454 9650 11506 9662
rect 12798 9714 12850 9726
rect 12798 9650 12850 9662
rect 12910 9714 12962 9726
rect 12910 9650 12962 9662
rect 13694 9714 13746 9726
rect 13694 9650 13746 9662
rect 13806 9714 13858 9726
rect 13806 9650 13858 9662
rect 14366 9714 14418 9726
rect 14366 9650 14418 9662
rect 16382 9714 16434 9726
rect 16382 9650 16434 9662
rect 17054 9714 17106 9726
rect 17054 9650 17106 9662
rect 18398 9714 18450 9726
rect 18398 9650 18450 9662
rect 4958 9602 5010 9614
rect 4958 9538 5010 9550
rect 5966 9602 6018 9614
rect 5966 9538 6018 9550
rect 7982 9602 8034 9614
rect 7982 9538 8034 9550
rect 8654 9602 8706 9614
rect 8654 9538 8706 9550
rect 9326 9602 9378 9614
rect 9326 9538 9378 9550
rect 9998 9602 10050 9614
rect 9998 9538 10050 9550
rect 10670 9602 10722 9614
rect 10670 9538 10722 9550
rect 15150 9602 15202 9614
rect 15150 9538 15202 9550
rect 15822 9602 15874 9614
rect 15822 9538 15874 9550
rect 16494 9602 16546 9614
rect 16494 9538 16546 9550
rect 17166 9602 17218 9614
rect 17166 9538 17218 9550
rect 17726 9602 17778 9614
rect 17726 9538 17778 9550
rect 19182 9602 19234 9614
rect 19182 9538 19234 9550
rect 19854 9602 19906 9614
rect 19854 9538 19906 9550
rect 1344 9434 22784 9468
rect 1344 9382 6534 9434
rect 6586 9382 6638 9434
rect 6690 9382 6742 9434
rect 6794 9382 11854 9434
rect 11906 9382 11958 9434
rect 12010 9382 12062 9434
rect 12114 9382 17174 9434
rect 17226 9382 17278 9434
rect 17330 9382 17382 9434
rect 17434 9382 22494 9434
rect 22546 9382 22598 9434
rect 22650 9382 22702 9434
rect 22754 9382 22784 9434
rect 1344 9348 22784 9382
rect 4846 9266 4898 9278
rect 4846 9202 4898 9214
rect 8990 9266 9042 9278
rect 8990 9202 9042 9214
rect 14478 9266 14530 9278
rect 14478 9202 14530 9214
rect 15150 9266 15202 9278
rect 15150 9202 15202 9214
rect 19854 9266 19906 9278
rect 19854 9202 19906 9214
rect 20526 9266 20578 9278
rect 20526 9202 20578 9214
rect 3390 9154 3442 9166
rect 3390 9090 3442 9102
rect 3502 9154 3554 9166
rect 3502 9090 3554 9102
rect 4062 9154 4114 9166
rect 4062 9090 4114 9102
rect 7422 9154 7474 9166
rect 7422 9090 7474 9102
rect 7534 9154 7586 9166
rect 7534 9090 7586 9102
rect 8206 9154 8258 9166
rect 8206 9090 8258 9102
rect 10334 9154 10386 9166
rect 10334 9090 10386 9102
rect 12350 9154 12402 9166
rect 12350 9090 12402 9102
rect 13022 9154 13074 9166
rect 13022 9090 13074 9102
rect 15710 9154 15762 9166
rect 15710 9090 15762 9102
rect 17726 9154 17778 9166
rect 17726 9090 17778 9102
rect 19070 9154 19122 9166
rect 19070 9090 19122 9102
rect 20414 9154 20466 9166
rect 20414 9090 20466 9102
rect 4734 9042 4786 9054
rect 4734 8978 4786 8990
rect 5406 9042 5458 9054
rect 5406 8978 5458 8990
rect 6078 9042 6130 9054
rect 6078 8978 6130 8990
rect 6190 9042 6242 9054
rect 6190 8978 6242 8990
rect 6750 9042 6802 9054
rect 6750 8978 6802 8990
rect 6862 9042 6914 9054
rect 6862 8978 6914 8990
rect 8878 9042 8930 9054
rect 8878 8978 8930 8990
rect 11006 9042 11058 9054
rect 11006 8978 11058 8990
rect 11678 9042 11730 9054
rect 11678 8978 11730 8990
rect 13694 9042 13746 9054
rect 13694 8978 13746 8990
rect 14366 9042 14418 9054
rect 14366 8978 14418 8990
rect 15038 9042 15090 9054
rect 15038 8978 15090 8990
rect 16382 9042 16434 9054
rect 16382 8978 16434 8990
rect 18398 9042 18450 9054
rect 18398 8978 18450 8990
rect 19742 9042 19794 9054
rect 19742 8978 19794 8990
rect 10446 8930 10498 8942
rect 10446 8866 10498 8878
rect 4174 8818 4226 8830
rect 4174 8754 4226 8766
rect 5518 8818 5570 8830
rect 5518 8754 5570 8766
rect 8318 8818 8370 8830
rect 8318 8754 8370 8766
rect 11118 8818 11170 8830
rect 11118 8754 11170 8766
rect 11790 8818 11842 8830
rect 11790 8754 11842 8766
rect 12462 8818 12514 8830
rect 12462 8754 12514 8766
rect 13134 8818 13186 8830
rect 13134 8754 13186 8766
rect 13806 8818 13858 8830
rect 13806 8754 13858 8766
rect 15822 8818 15874 8830
rect 15822 8754 15874 8766
rect 16494 8818 16546 8830
rect 16494 8754 16546 8766
rect 17838 8818 17890 8830
rect 17838 8754 17890 8766
rect 18510 8818 18562 8830
rect 18510 8754 18562 8766
rect 19182 8818 19234 8830
rect 19182 8754 19234 8766
rect 1344 8650 22624 8684
rect 1344 8598 3874 8650
rect 3926 8598 3978 8650
rect 4030 8598 4082 8650
rect 4134 8598 9194 8650
rect 9246 8598 9298 8650
rect 9350 8598 9402 8650
rect 9454 8598 14514 8650
rect 14566 8598 14618 8650
rect 14670 8598 14722 8650
rect 14774 8598 19834 8650
rect 19886 8598 19938 8650
rect 19990 8598 20042 8650
rect 20094 8598 22624 8650
rect 1344 8564 22624 8598
rect 4958 8482 5010 8494
rect 4958 8418 5010 8430
rect 5966 8482 6018 8494
rect 5966 8418 6018 8430
rect 6638 8482 6690 8494
rect 6638 8418 6690 8430
rect 9326 8482 9378 8494
rect 9326 8418 9378 8430
rect 9998 8482 10050 8494
rect 9998 8418 10050 8430
rect 10670 8482 10722 8494
rect 10670 8418 10722 8430
rect 15150 8482 15202 8494
rect 15150 8418 15202 8430
rect 17166 8482 17218 8494
rect 17166 8418 17218 8430
rect 17838 8482 17890 8494
rect 17838 8418 17890 8430
rect 18510 8482 18562 8494
rect 18510 8418 18562 8430
rect 19182 8482 19234 8494
rect 19182 8418 19234 8430
rect 11230 8370 11282 8382
rect 11230 8306 11282 8318
rect 6526 8258 6578 8270
rect 6526 8194 6578 8206
rect 7198 8258 7250 8270
rect 7198 8194 7250 8206
rect 7870 8258 7922 8270
rect 7870 8194 7922 8206
rect 9214 8258 9266 8270
rect 9214 8194 9266 8206
rect 9886 8258 9938 8270
rect 9886 8194 9938 8206
rect 10558 8258 10610 8270
rect 10558 8194 10610 8206
rect 12126 8258 12178 8270
rect 12126 8194 12178 8206
rect 12238 8258 12290 8270
rect 12238 8194 12290 8206
rect 12910 8258 12962 8270
rect 12910 8194 12962 8206
rect 13694 8258 13746 8270
rect 13694 8194 13746 8206
rect 13806 8258 13858 8270
rect 13806 8194 13858 8206
rect 14366 8258 14418 8270
rect 14366 8194 14418 8206
rect 14478 8258 14530 8270
rect 14478 8194 14530 8206
rect 15038 8258 15090 8270
rect 15038 8194 15090 8206
rect 15822 8258 15874 8270
rect 15822 8194 15874 8206
rect 16494 8258 16546 8270
rect 16494 8194 16546 8206
rect 17054 8258 17106 8270
rect 17054 8194 17106 8206
rect 18398 8258 18450 8270
rect 18398 8194 18450 8206
rect 19070 8258 19122 8270
rect 19070 8194 19122 8206
rect 19742 8258 19794 8270
rect 19742 8194 19794 8206
rect 19854 8258 19906 8270
rect 19854 8194 19906 8206
rect 2942 8146 2994 8158
rect 2942 8082 2994 8094
rect 3502 8146 3554 8158
rect 3502 8082 3554 8094
rect 4174 8146 4226 8158
rect 4174 8082 4226 8094
rect 4846 8146 4898 8158
rect 4846 8082 4898 8094
rect 5854 8146 5906 8158
rect 5854 8082 5906 8094
rect 8542 8146 8594 8158
rect 8542 8082 8594 8094
rect 11342 8146 11394 8158
rect 11342 8082 11394 8094
rect 12798 8146 12850 8158
rect 12798 8082 12850 8094
rect 15710 8146 15762 8158
rect 15710 8082 15762 8094
rect 16382 8146 16434 8158
rect 16382 8082 16434 8094
rect 17726 8146 17778 8158
rect 17726 8082 17778 8094
rect 20526 8146 20578 8158
rect 20526 8082 20578 8094
rect 2830 8034 2882 8046
rect 2830 7970 2882 7982
rect 3614 8034 3666 8046
rect 3614 7970 3666 7982
rect 4286 8034 4338 8046
rect 4286 7970 4338 7982
rect 7310 8034 7362 8046
rect 7310 7970 7362 7982
rect 7982 8034 8034 8046
rect 7982 7970 8034 7982
rect 8654 8034 8706 8046
rect 8654 7970 8706 7982
rect 20414 8034 20466 8046
rect 20414 7970 20466 7982
rect 1344 7866 22784 7900
rect 1344 7814 6534 7866
rect 6586 7814 6638 7866
rect 6690 7814 6742 7866
rect 6794 7814 11854 7866
rect 11906 7814 11958 7866
rect 12010 7814 12062 7866
rect 12114 7814 17174 7866
rect 17226 7814 17278 7866
rect 17330 7814 17382 7866
rect 17434 7814 22494 7866
rect 22546 7814 22598 7866
rect 22650 7814 22702 7866
rect 22754 7814 22784 7866
rect 1344 7780 22784 7814
rect 6190 7698 6242 7710
rect 6190 7634 6242 7646
rect 6862 7698 6914 7710
rect 6862 7634 6914 7646
rect 8990 7698 9042 7710
rect 8990 7634 9042 7646
rect 9998 7698 10050 7710
rect 9998 7634 10050 7646
rect 10670 7698 10722 7710
rect 10670 7634 10722 7646
rect 11230 7698 11282 7710
rect 11230 7634 11282 7646
rect 13358 7698 13410 7710
rect 13358 7634 13410 7646
rect 14702 7698 14754 7710
rect 14702 7634 14754 7646
rect 16718 7698 16770 7710
rect 16718 7634 16770 7646
rect 17838 7698 17890 7710
rect 17838 7634 17890 7646
rect 18510 7698 18562 7710
rect 18510 7634 18562 7646
rect 4734 7586 4786 7598
rect 4734 7522 4786 7534
rect 10558 7586 10610 7598
rect 10558 7522 10610 7534
rect 13918 7586 13970 7598
rect 13918 7522 13970 7534
rect 15262 7586 15314 7598
rect 15262 7522 15314 7534
rect 15934 7586 15986 7598
rect 15934 7522 15986 7534
rect 2158 7474 2210 7486
rect 2158 7410 2210 7422
rect 2718 7474 2770 7486
rect 2718 7410 2770 7422
rect 3390 7474 3442 7486
rect 3390 7410 3442 7422
rect 4062 7474 4114 7486
rect 4062 7410 4114 7422
rect 4846 7474 4898 7486
rect 4846 7410 4898 7422
rect 5406 7474 5458 7486
rect 5406 7410 5458 7422
rect 6078 7474 6130 7486
rect 6078 7410 6130 7422
rect 6750 7474 6802 7486
rect 6750 7410 6802 7422
rect 7422 7474 7474 7486
rect 7422 7410 7474 7422
rect 8206 7474 8258 7486
rect 8206 7410 8258 7422
rect 8878 7474 8930 7486
rect 8878 7410 8930 7422
rect 9886 7474 9938 7486
rect 9886 7410 9938 7422
rect 11342 7474 11394 7486
rect 11342 7410 11394 7422
rect 11902 7474 11954 7486
rect 11902 7410 11954 7422
rect 12574 7474 12626 7486
rect 12574 7410 12626 7422
rect 13246 7474 13298 7486
rect 13246 7410 13298 7422
rect 14590 7474 14642 7486
rect 14590 7410 14642 7422
rect 16606 7474 16658 7486
rect 16606 7410 16658 7422
rect 17726 7474 17778 7486
rect 17726 7410 17778 7422
rect 18398 7474 18450 7486
rect 18398 7410 18450 7422
rect 19070 7474 19122 7486
rect 19070 7410 19122 7422
rect 19742 7474 19794 7486
rect 19742 7410 19794 7422
rect 20414 7474 20466 7486
rect 20414 7410 20466 7422
rect 21086 7474 21138 7486
rect 21086 7410 21138 7422
rect 14030 7362 14082 7374
rect 14030 7298 14082 7310
rect 2046 7250 2098 7262
rect 2046 7186 2098 7198
rect 2830 7250 2882 7262
rect 2830 7186 2882 7198
rect 3502 7250 3554 7262
rect 3502 7186 3554 7198
rect 4174 7250 4226 7262
rect 4174 7186 4226 7198
rect 5518 7250 5570 7262
rect 5518 7186 5570 7198
rect 7534 7250 7586 7262
rect 7534 7186 7586 7198
rect 8318 7250 8370 7262
rect 8318 7186 8370 7198
rect 12014 7250 12066 7262
rect 12014 7186 12066 7198
rect 12686 7250 12738 7262
rect 12686 7186 12738 7198
rect 15374 7250 15426 7262
rect 15374 7186 15426 7198
rect 16046 7250 16098 7262
rect 16046 7186 16098 7198
rect 19182 7250 19234 7262
rect 19182 7186 19234 7198
rect 19854 7250 19906 7262
rect 19854 7186 19906 7198
rect 20526 7250 20578 7262
rect 20526 7186 20578 7198
rect 21198 7250 21250 7262
rect 21198 7186 21250 7198
rect 1344 7082 22624 7116
rect 1344 7030 3874 7082
rect 3926 7030 3978 7082
rect 4030 7030 4082 7082
rect 4134 7030 9194 7082
rect 9246 7030 9298 7082
rect 9350 7030 9402 7082
rect 9454 7030 14514 7082
rect 14566 7030 14618 7082
rect 14670 7030 14722 7082
rect 14774 7030 19834 7082
rect 19886 7030 19938 7082
rect 19990 7030 20042 7082
rect 20094 7030 22624 7082
rect 1344 6996 22624 7030
rect 4286 6914 4338 6926
rect 4286 6850 4338 6862
rect 4958 6914 5010 6926
rect 4958 6850 5010 6862
rect 10558 6914 10610 6926
rect 10558 6850 10610 6862
rect 11230 6914 11282 6926
rect 11230 6850 11282 6862
rect 14254 6914 14306 6926
rect 14254 6850 14306 6862
rect 14926 6914 14978 6926
rect 14926 6850 14978 6862
rect 15598 6914 15650 6926
rect 15598 6850 15650 6862
rect 17614 6914 17666 6926
rect 17614 6850 17666 6862
rect 19630 6914 19682 6926
rect 19630 6850 19682 6862
rect 5742 6690 5794 6702
rect 5742 6626 5794 6638
rect 5854 6690 5906 6702
rect 5854 6626 5906 6638
rect 6414 6690 6466 6702
rect 6414 6626 6466 6638
rect 6526 6690 6578 6702
rect 6526 6626 6578 6638
rect 8542 6690 8594 6702
rect 8542 6626 8594 6638
rect 9214 6690 9266 6702
rect 9214 6626 9266 6638
rect 9774 6690 9826 6702
rect 9774 6626 9826 6638
rect 10446 6690 10498 6702
rect 10446 6626 10498 6638
rect 11118 6690 11170 6702
rect 11118 6626 11170 6638
rect 11790 6690 11842 6702
rect 11790 6626 11842 6638
rect 12462 6690 12514 6702
rect 12462 6626 12514 6638
rect 14142 6690 14194 6702
rect 14142 6626 14194 6638
rect 14814 6690 14866 6702
rect 14814 6626 14866 6638
rect 15486 6690 15538 6702
rect 15486 6626 15538 6638
rect 18958 6690 19010 6702
rect 18958 6626 19010 6638
rect 21646 6690 21698 6702
rect 21646 6626 21698 6638
rect 2158 6578 2210 6590
rect 2158 6514 2210 6526
rect 2830 6578 2882 6590
rect 2830 6514 2882 6526
rect 3502 6578 3554 6590
rect 3502 6514 3554 6526
rect 4174 6578 4226 6590
rect 4174 6514 4226 6526
rect 4846 6578 4898 6590
rect 4846 6514 4898 6526
rect 7086 6578 7138 6590
rect 7086 6514 7138 6526
rect 7758 6578 7810 6590
rect 7758 6514 7810 6526
rect 8430 6578 8482 6590
rect 8430 6514 8482 6526
rect 9102 6578 9154 6590
rect 9102 6514 9154 6526
rect 16158 6578 16210 6590
rect 16158 6514 16210 6526
rect 16270 6578 16322 6590
rect 16270 6514 16322 6526
rect 16830 6578 16882 6590
rect 16830 6514 16882 6526
rect 16942 6578 16994 6590
rect 16942 6514 16994 6526
rect 17502 6578 17554 6590
rect 17502 6514 17554 6526
rect 18174 6578 18226 6590
rect 18174 6514 18226 6526
rect 18846 6578 18898 6590
rect 18846 6514 18898 6526
rect 19518 6578 19570 6590
rect 19518 6514 19570 6526
rect 20302 6578 20354 6590
rect 20302 6514 20354 6526
rect 2270 6466 2322 6478
rect 2270 6402 2322 6414
rect 2942 6466 2994 6478
rect 2942 6402 2994 6414
rect 3614 6466 3666 6478
rect 3614 6402 3666 6414
rect 7198 6466 7250 6478
rect 7198 6402 7250 6414
rect 7870 6466 7922 6478
rect 7870 6402 7922 6414
rect 9886 6466 9938 6478
rect 9886 6402 9938 6414
rect 11902 6466 11954 6478
rect 11902 6402 11954 6414
rect 12574 6466 12626 6478
rect 12574 6402 12626 6414
rect 18286 6466 18338 6478
rect 18286 6402 18338 6414
rect 20190 6466 20242 6478
rect 20190 6402 20242 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 1344 6298 22784 6332
rect 1344 6246 6534 6298
rect 6586 6246 6638 6298
rect 6690 6246 6742 6298
rect 6794 6246 11854 6298
rect 11906 6246 11958 6298
rect 12010 6246 12062 6298
rect 12114 6246 17174 6298
rect 17226 6246 17278 6298
rect 17330 6246 17382 6298
rect 17434 6246 22494 6298
rect 22546 6246 22598 6298
rect 22650 6246 22702 6298
rect 22754 6246 22784 6298
rect 1344 6212 22784 6246
rect 5518 6130 5570 6142
rect 5518 6066 5570 6078
rect 6190 6130 6242 6142
rect 6190 6066 6242 6078
rect 8878 6130 8930 6142
rect 8878 6066 8930 6078
rect 9886 6130 9938 6142
rect 9886 6066 9938 6078
rect 10558 6130 10610 6142
rect 10558 6066 10610 6078
rect 11230 6130 11282 6142
rect 11230 6066 11282 6078
rect 11902 6130 11954 6142
rect 11902 6066 11954 6078
rect 13358 6130 13410 6142
rect 13358 6066 13410 6078
rect 14030 6130 14082 6142
rect 14030 6066 14082 6078
rect 14702 6130 14754 6142
rect 14702 6066 14754 6078
rect 15374 6130 15426 6142
rect 15374 6066 15426 6078
rect 16046 6130 16098 6142
rect 16046 6066 16098 6078
rect 16718 6130 16770 6142
rect 16718 6066 16770 6078
rect 6750 6018 6802 6030
rect 6750 5954 6802 5966
rect 6862 6018 6914 6030
rect 6862 5954 6914 5966
rect 7422 6018 7474 6030
rect 7422 5954 7474 5966
rect 8094 6018 8146 6030
rect 8094 5954 8146 5966
rect 8766 6018 8818 6030
rect 8766 5954 8818 5966
rect 11118 6018 11170 6030
rect 11118 5954 11170 5966
rect 11790 6018 11842 6030
rect 11790 5954 11842 5966
rect 12574 6018 12626 6030
rect 12574 5954 12626 5966
rect 14590 6018 14642 6030
rect 14590 5954 14642 5966
rect 15262 6018 15314 6030
rect 15262 5954 15314 5966
rect 15934 6018 15986 6030
rect 15934 5954 15986 5966
rect 16606 6018 16658 6030
rect 16606 5954 16658 5966
rect 19070 6018 19122 6030
rect 19070 5954 19122 5966
rect 19742 6018 19794 6030
rect 19742 5954 19794 5966
rect 2046 5906 2098 5918
rect 2046 5842 2098 5854
rect 2718 5906 2770 5918
rect 2718 5842 2770 5854
rect 3390 5906 3442 5918
rect 3390 5842 3442 5854
rect 4062 5906 4114 5918
rect 4062 5842 4114 5854
rect 4734 5906 4786 5918
rect 4734 5842 4786 5854
rect 5406 5906 5458 5918
rect 5406 5842 5458 5854
rect 6078 5906 6130 5918
rect 6078 5842 6130 5854
rect 9774 5906 9826 5918
rect 9774 5842 9826 5854
rect 10446 5906 10498 5918
rect 10446 5842 10498 5854
rect 13246 5906 13298 5918
rect 13246 5842 13298 5854
rect 13918 5906 13970 5918
rect 13918 5842 13970 5854
rect 17726 5906 17778 5918
rect 17726 5842 17778 5854
rect 18398 5906 18450 5918
rect 18398 5842 18450 5854
rect 20414 5906 20466 5918
rect 20414 5842 20466 5854
rect 21086 5906 21138 5918
rect 21086 5842 21138 5854
rect 21870 5906 21922 5918
rect 21870 5842 21922 5854
rect 18510 5794 18562 5806
rect 18510 5730 18562 5742
rect 19182 5794 19234 5806
rect 19182 5730 19234 5742
rect 2158 5682 2210 5694
rect 2158 5618 2210 5630
rect 2830 5682 2882 5694
rect 2830 5618 2882 5630
rect 3502 5682 3554 5694
rect 3502 5618 3554 5630
rect 4174 5682 4226 5694
rect 4174 5618 4226 5630
rect 4846 5682 4898 5694
rect 4846 5618 4898 5630
rect 7534 5682 7586 5694
rect 7534 5618 7586 5630
rect 8206 5682 8258 5694
rect 8206 5618 8258 5630
rect 12686 5682 12738 5694
rect 12686 5618 12738 5630
rect 17838 5682 17890 5694
rect 17838 5618 17890 5630
rect 19854 5682 19906 5694
rect 19854 5618 19906 5630
rect 20526 5682 20578 5694
rect 20526 5618 20578 5630
rect 21198 5682 21250 5694
rect 21198 5618 21250 5630
rect 21758 5682 21810 5694
rect 21758 5618 21810 5630
rect 1344 5514 22624 5548
rect 1344 5462 3874 5514
rect 3926 5462 3978 5514
rect 4030 5462 4082 5514
rect 4134 5462 9194 5514
rect 9246 5462 9298 5514
rect 9350 5462 9402 5514
rect 9454 5462 14514 5514
rect 14566 5462 14618 5514
rect 14670 5462 14722 5514
rect 14774 5462 19834 5514
rect 19886 5462 19938 5514
rect 19990 5462 20042 5514
rect 20094 5462 22624 5514
rect 1344 5428 22624 5462
rect 5854 5346 5906 5358
rect 5854 5282 5906 5294
rect 6526 5346 6578 5358
rect 6526 5282 6578 5294
rect 7198 5346 7250 5358
rect 7198 5282 7250 5294
rect 8542 5346 8594 5358
rect 8542 5282 8594 5294
rect 9886 5346 9938 5358
rect 9886 5282 9938 5294
rect 10558 5346 10610 5358
rect 10558 5282 10610 5294
rect 14142 5346 14194 5358
rect 14142 5282 14194 5294
rect 14814 5346 14866 5358
rect 14814 5282 14866 5294
rect 15486 5346 15538 5358
rect 15486 5282 15538 5294
rect 18174 5346 18226 5358
rect 18174 5282 18226 5294
rect 20190 5346 20242 5358
rect 20190 5282 20242 5294
rect 19518 5234 19570 5246
rect 19518 5170 19570 5182
rect 4174 5122 4226 5134
rect 4174 5058 4226 5070
rect 4846 5122 4898 5134
rect 4846 5058 4898 5070
rect 7086 5122 7138 5134
rect 7086 5058 7138 5070
rect 7758 5122 7810 5134
rect 7758 5058 7810 5070
rect 7870 5122 7922 5134
rect 7870 5058 7922 5070
rect 8430 5122 8482 5134
rect 8430 5058 8482 5070
rect 9102 5122 9154 5134
rect 9102 5058 9154 5070
rect 9214 5122 9266 5134
rect 9214 5058 9266 5070
rect 10446 5122 10498 5134
rect 10446 5058 10498 5070
rect 11454 5122 11506 5134
rect 11454 5058 11506 5070
rect 11566 5122 11618 5134
rect 11566 5058 11618 5070
rect 15374 5122 15426 5134
rect 15374 5058 15426 5070
rect 16830 5122 16882 5134
rect 16830 5058 16882 5070
rect 17390 5122 17442 5134
rect 17390 5058 17442 5070
rect 18062 5122 18114 5134
rect 18062 5058 18114 5070
rect 18734 5122 18786 5134
rect 18734 5058 18786 5070
rect 18846 5122 18898 5134
rect 18846 5058 18898 5070
rect 19406 5122 19458 5134
rect 19406 5058 19458 5070
rect 20078 5122 20130 5134
rect 20078 5058 20130 5070
rect 2158 5010 2210 5022
rect 2158 4946 2210 4958
rect 2830 5010 2882 5022
rect 2830 4946 2882 4958
rect 3502 5010 3554 5022
rect 3502 4946 3554 4958
rect 3614 5010 3666 5022
rect 3614 4946 3666 4958
rect 5742 5010 5794 5022
rect 5742 4946 5794 4958
rect 6414 5010 6466 5022
rect 6414 4946 6466 4958
rect 9774 5010 9826 5022
rect 9774 4946 9826 4958
rect 12126 5010 12178 5022
rect 12126 4946 12178 4958
rect 12798 5010 12850 5022
rect 12798 4946 12850 4958
rect 14030 5010 14082 5022
rect 14030 4946 14082 4958
rect 14702 5010 14754 5022
rect 14702 4946 14754 4958
rect 16046 5010 16098 5022
rect 16046 4946 16098 4958
rect 16718 5010 16770 5022
rect 16718 4946 16770 4958
rect 20750 5010 20802 5022
rect 20750 4946 20802 4958
rect 21646 5010 21698 5022
rect 21646 4946 21698 4958
rect 2270 4898 2322 4910
rect 2270 4834 2322 4846
rect 2942 4898 2994 4910
rect 2942 4834 2994 4846
rect 4286 4898 4338 4910
rect 4286 4834 4338 4846
rect 4958 4898 5010 4910
rect 4958 4834 5010 4846
rect 12238 4898 12290 4910
rect 12238 4834 12290 4846
rect 12910 4898 12962 4910
rect 12910 4834 12962 4846
rect 16158 4898 16210 4910
rect 16158 4834 16210 4846
rect 17502 4898 17554 4910
rect 17502 4834 17554 4846
rect 20862 4898 20914 4910
rect 20862 4834 20914 4846
rect 21758 4898 21810 4910
rect 21758 4834 21810 4846
rect 1344 4730 22784 4764
rect 1344 4678 6534 4730
rect 6586 4678 6638 4730
rect 6690 4678 6742 4730
rect 6794 4678 11854 4730
rect 11906 4678 11958 4730
rect 12010 4678 12062 4730
rect 12114 4678 17174 4730
rect 17226 4678 17278 4730
rect 17330 4678 17382 4730
rect 17434 4678 22494 4730
rect 22546 4678 22598 4730
rect 22650 4678 22702 4730
rect 22754 4678 22784 4730
rect 1344 4644 22784 4678
rect 3838 4562 3890 4574
rect 3838 4498 3890 4510
rect 4510 4562 4562 4574
rect 4510 4498 4562 4510
rect 7198 4562 7250 4574
rect 7198 4498 7250 4510
rect 8542 4562 8594 4574
rect 8542 4498 8594 4510
rect 15150 4562 15202 4574
rect 15150 4498 15202 4510
rect 15822 4562 15874 4574
rect 15822 4498 15874 4510
rect 17838 4562 17890 4574
rect 17838 4498 17890 4510
rect 18510 4562 18562 4574
rect 18510 4498 18562 4510
rect 19854 4562 19906 4574
rect 19854 4498 19906 4510
rect 20526 4562 20578 4574
rect 20526 4498 20578 4510
rect 21198 4562 21250 4574
rect 21198 4498 21250 4510
rect 2382 4450 2434 4462
rect 2382 4386 2434 4398
rect 5070 4450 5122 4462
rect 5070 4386 5122 4398
rect 5742 4450 5794 4462
rect 5742 4386 5794 4398
rect 8430 4450 8482 4462
rect 8430 4386 8482 4398
rect 9774 4450 9826 4462
rect 9774 4386 9826 4398
rect 10446 4450 10498 4462
rect 10446 4386 10498 4398
rect 14366 4450 14418 4462
rect 14366 4386 14418 4398
rect 16382 4450 16434 4462
rect 16382 4386 16434 4398
rect 16494 4450 16546 4462
rect 16494 4386 16546 4398
rect 17726 4450 17778 4462
rect 17726 4386 17778 4398
rect 18398 4450 18450 4462
rect 18398 4386 18450 4398
rect 19070 4450 19122 4462
rect 19070 4386 19122 4398
rect 20414 4450 20466 4462
rect 20414 4386 20466 4398
rect 21086 4450 21138 4462
rect 21086 4386 21138 4398
rect 2494 4338 2546 4350
rect 2494 4274 2546 4286
rect 3054 4338 3106 4350
rect 3054 4274 3106 4286
rect 3166 4338 3218 4350
rect 3166 4274 3218 4286
rect 3726 4338 3778 4350
rect 3726 4274 3778 4286
rect 4398 4338 4450 4350
rect 4398 4274 4450 4286
rect 6414 4338 6466 4350
rect 6414 4274 6466 4286
rect 7086 4338 7138 4350
rect 7086 4274 7138 4286
rect 7758 4338 7810 4350
rect 7758 4274 7810 4286
rect 11118 4338 11170 4350
rect 11118 4274 11170 4286
rect 12350 4338 12402 4350
rect 12350 4274 12402 4286
rect 13022 4338 13074 4350
rect 13022 4274 13074 4286
rect 13694 4338 13746 4350
rect 13694 4274 13746 4286
rect 14478 4338 14530 4350
rect 14478 4274 14530 4286
rect 15038 4338 15090 4350
rect 15038 4274 15090 4286
rect 15710 4338 15762 4350
rect 15710 4274 15762 4286
rect 19742 4338 19794 4350
rect 19742 4274 19794 4286
rect 21870 4338 21922 4350
rect 21870 4274 21922 4286
rect 5182 4114 5234 4126
rect 5182 4050 5234 4062
rect 5854 4114 5906 4126
rect 5854 4050 5906 4062
rect 6526 4114 6578 4126
rect 6526 4050 6578 4062
rect 7870 4114 7922 4126
rect 7870 4050 7922 4062
rect 9886 4114 9938 4126
rect 9886 4050 9938 4062
rect 10558 4114 10610 4126
rect 10558 4050 10610 4062
rect 11230 4114 11282 4126
rect 11230 4050 11282 4062
rect 12462 4114 12514 4126
rect 12462 4050 12514 4062
rect 13134 4114 13186 4126
rect 13134 4050 13186 4062
rect 13806 4114 13858 4126
rect 13806 4050 13858 4062
rect 19182 4114 19234 4126
rect 19182 4050 19234 4062
rect 21758 4114 21810 4126
rect 21758 4050 21810 4062
rect 1344 3946 22624 3980
rect 1344 3894 3874 3946
rect 3926 3894 3978 3946
rect 4030 3894 4082 3946
rect 4134 3894 9194 3946
rect 9246 3894 9298 3946
rect 9350 3894 9402 3946
rect 9454 3894 14514 3946
rect 14566 3894 14618 3946
rect 14670 3894 14722 3946
rect 14774 3894 19834 3946
rect 19886 3894 19938 3946
rect 19990 3894 20042 3946
rect 20094 3894 22624 3946
rect 1344 3860 22624 3894
rect 2942 3778 2994 3790
rect 2942 3714 2994 3726
rect 3614 3778 3666 3790
rect 3614 3714 3666 3726
rect 4286 3778 4338 3790
rect 4286 3714 4338 3726
rect 4958 3778 5010 3790
rect 4958 3714 5010 3726
rect 6414 3778 6466 3790
rect 6414 3714 6466 3726
rect 7086 3778 7138 3790
rect 7086 3714 7138 3726
rect 7870 3778 7922 3790
rect 7870 3714 7922 3726
rect 17614 3778 17666 3790
rect 17614 3714 17666 3726
rect 19630 3778 19682 3790
rect 19630 3714 19682 3726
rect 20302 3778 20354 3790
rect 20302 3714 20354 3726
rect 2830 3554 2882 3566
rect 2830 3490 2882 3502
rect 3502 3554 3554 3566
rect 3502 3490 3554 3502
rect 4174 3554 4226 3566
rect 4174 3490 4226 3502
rect 5854 3554 5906 3566
rect 5854 3490 5906 3502
rect 6526 3554 6578 3566
rect 6526 3490 6578 3502
rect 7198 3554 7250 3566
rect 7198 3490 7250 3502
rect 7758 3554 7810 3566
rect 7758 3490 7810 3502
rect 8430 3554 8482 3566
rect 8430 3490 8482 3502
rect 8542 3554 8594 3566
rect 8542 3490 8594 3502
rect 9662 3554 9714 3566
rect 9662 3490 9714 3502
rect 9774 3554 9826 3566
rect 9774 3490 9826 3502
rect 10334 3554 10386 3566
rect 10334 3490 10386 3502
rect 10446 3554 10498 3566
rect 10446 3490 10498 3502
rect 11118 3554 11170 3566
rect 11118 3490 11170 3502
rect 11678 3554 11730 3566
rect 11678 3490 11730 3502
rect 14590 3554 14642 3566
rect 14590 3490 14642 3502
rect 15262 3554 15314 3566
rect 16606 3554 16658 3566
rect 15586 3502 15598 3554
rect 15650 3551 15662 3554
rect 15810 3551 15822 3554
rect 15650 3505 15822 3551
rect 15650 3502 15662 3505
rect 15810 3502 15822 3505
rect 15874 3502 15886 3554
rect 15262 3490 15314 3502
rect 16606 3490 16658 3502
rect 17502 3554 17554 3566
rect 17502 3490 17554 3502
rect 18174 3554 18226 3566
rect 18174 3490 18226 3502
rect 18846 3554 18898 3566
rect 18846 3490 18898 3502
rect 20190 3554 20242 3566
rect 20190 3490 20242 3502
rect 4846 3442 4898 3454
rect 4846 3378 4898 3390
rect 5742 3442 5794 3454
rect 5742 3378 5794 3390
rect 11006 3442 11058 3454
rect 11006 3378 11058 3390
rect 11790 3442 11842 3454
rect 11790 3378 11842 3390
rect 13918 3442 13970 3454
rect 13918 3378 13970 3390
rect 14030 3442 14082 3454
rect 14030 3378 14082 3390
rect 14702 3442 14754 3454
rect 14702 3378 14754 3390
rect 15374 3442 15426 3454
rect 15374 3378 15426 3390
rect 15934 3442 15986 3454
rect 15934 3378 15986 3390
rect 16046 3442 16098 3454
rect 16046 3378 16098 3390
rect 16718 3442 16770 3454
rect 16718 3378 16770 3390
rect 18286 3442 18338 3454
rect 18286 3378 18338 3390
rect 18958 3442 19010 3454
rect 18958 3378 19010 3390
rect 19518 3442 19570 3454
rect 19518 3378 19570 3390
rect 1344 3162 22784 3196
rect 1344 3110 6534 3162
rect 6586 3110 6638 3162
rect 6690 3110 6742 3162
rect 6794 3110 11854 3162
rect 11906 3110 11958 3162
rect 12010 3110 12062 3162
rect 12114 3110 17174 3162
rect 17226 3110 17278 3162
rect 17330 3110 17382 3162
rect 17434 3110 22494 3162
rect 22546 3110 22598 3162
rect 22650 3110 22702 3162
rect 22754 3110 22784 3162
rect 1344 3076 22784 3110
<< via1 >>
rect 3874 16438 3926 16490
rect 3978 16438 4030 16490
rect 4082 16438 4134 16490
rect 9194 16438 9246 16490
rect 9298 16438 9350 16490
rect 9402 16438 9454 16490
rect 14514 16438 14566 16490
rect 14618 16438 14670 16490
rect 14722 16438 14774 16490
rect 19834 16438 19886 16490
rect 19938 16438 19990 16490
rect 20042 16438 20094 16490
rect 6534 15654 6586 15706
rect 6638 15654 6690 15706
rect 6742 15654 6794 15706
rect 11854 15654 11906 15706
rect 11958 15654 12010 15706
rect 12062 15654 12114 15706
rect 17174 15654 17226 15706
rect 17278 15654 17330 15706
rect 17382 15654 17434 15706
rect 22494 15654 22546 15706
rect 22598 15654 22650 15706
rect 22702 15654 22754 15706
rect 3874 14870 3926 14922
rect 3978 14870 4030 14922
rect 4082 14870 4134 14922
rect 9194 14870 9246 14922
rect 9298 14870 9350 14922
rect 9402 14870 9454 14922
rect 14514 14870 14566 14922
rect 14618 14870 14670 14922
rect 14722 14870 14774 14922
rect 19834 14870 19886 14922
rect 19938 14870 19990 14922
rect 20042 14870 20094 14922
rect 16830 14590 16882 14642
rect 16942 14366 16994 14418
rect 17614 14366 17666 14418
rect 17502 14254 17554 14306
rect 6534 14086 6586 14138
rect 6638 14086 6690 14138
rect 6742 14086 6794 14138
rect 11854 14086 11906 14138
rect 11958 14086 12010 14138
rect 12062 14086 12114 14138
rect 17174 14086 17226 14138
rect 17278 14086 17330 14138
rect 17382 14086 17434 14138
rect 22494 14086 22546 14138
rect 22598 14086 22650 14138
rect 22702 14086 22754 14138
rect 16158 13694 16210 13746
rect 16830 13694 16882 13746
rect 17726 13694 17778 13746
rect 18398 13694 18450 13746
rect 16270 13470 16322 13522
rect 16942 13470 16994 13522
rect 17838 13470 17890 13522
rect 18510 13470 18562 13522
rect 3874 13302 3926 13354
rect 3978 13302 4030 13354
rect 4082 13302 4134 13354
rect 9194 13302 9246 13354
rect 9298 13302 9350 13354
rect 9402 13302 9454 13354
rect 14514 13302 14566 13354
rect 14618 13302 14670 13354
rect 14722 13302 14774 13354
rect 19834 13302 19886 13354
rect 19938 13302 19990 13354
rect 20042 13302 20094 13354
rect 14926 13134 14978 13186
rect 18286 13134 18338 13186
rect 18958 13134 19010 13186
rect 17502 12910 17554 12962
rect 18846 12910 18898 12962
rect 14814 12798 14866 12850
rect 15486 12798 15538 12850
rect 16158 12798 16210 12850
rect 16830 12798 16882 12850
rect 18174 12798 18226 12850
rect 19518 12798 19570 12850
rect 15598 12686 15650 12738
rect 16270 12686 16322 12738
rect 16942 12686 16994 12738
rect 17614 12686 17666 12738
rect 19630 12686 19682 12738
rect 6534 12518 6586 12570
rect 6638 12518 6690 12570
rect 6742 12518 6794 12570
rect 11854 12518 11906 12570
rect 11958 12518 12010 12570
rect 12062 12518 12114 12570
rect 17174 12518 17226 12570
rect 17278 12518 17330 12570
rect 17382 12518 17434 12570
rect 22494 12518 22546 12570
rect 22598 12518 22650 12570
rect 22702 12518 22754 12570
rect 19182 12350 19234 12402
rect 19854 12350 19906 12402
rect 17726 12238 17778 12290
rect 17838 12238 17890 12290
rect 18398 12238 18450 12290
rect 19070 12238 19122 12290
rect 19742 12238 19794 12290
rect 20414 12238 20466 12290
rect 20526 12238 20578 12290
rect 14142 12126 14194 12178
rect 14814 12126 14866 12178
rect 15486 12126 15538 12178
rect 16158 12126 16210 12178
rect 16830 12126 16882 12178
rect 14254 11902 14306 11954
rect 14926 11902 14978 11954
rect 15598 11902 15650 11954
rect 16270 11902 16322 11954
rect 16942 11902 16994 11954
rect 18510 11902 18562 11954
rect 3874 11734 3926 11786
rect 3978 11734 4030 11786
rect 4082 11734 4134 11786
rect 9194 11734 9246 11786
rect 9298 11734 9350 11786
rect 9402 11734 9454 11786
rect 14514 11734 14566 11786
rect 14618 11734 14670 11786
rect 14722 11734 14774 11786
rect 19834 11734 19886 11786
rect 19938 11734 19990 11786
rect 20042 11734 20094 11786
rect 17614 11566 17666 11618
rect 19630 11566 19682 11618
rect 10670 11454 10722 11506
rect 14926 11342 14978 11394
rect 15598 11342 15650 11394
rect 16270 11342 16322 11394
rect 16830 11342 16882 11394
rect 16942 11342 16994 11394
rect 17502 11342 17554 11394
rect 18174 11342 18226 11394
rect 18846 11342 18898 11394
rect 19518 11342 19570 11394
rect 6078 11230 6130 11282
rect 6190 11230 6242 11282
rect 6974 11230 7026 11282
rect 7646 11230 7698 11282
rect 8318 11230 8370 11282
rect 9214 11230 9266 11282
rect 9886 11230 9938 11282
rect 10558 11230 10610 11282
rect 12126 11230 12178 11282
rect 12238 11230 12290 11282
rect 12798 11230 12850 11282
rect 13694 11230 13746 11282
rect 14814 11230 14866 11282
rect 15486 11230 15538 11282
rect 16158 11230 16210 11282
rect 20190 11230 20242 11282
rect 6862 11118 6914 11170
rect 7534 11118 7586 11170
rect 8206 11118 8258 11170
rect 9326 11118 9378 11170
rect 9998 11118 10050 11170
rect 12910 11118 12962 11170
rect 13806 11118 13858 11170
rect 18286 11118 18338 11170
rect 18958 11118 19010 11170
rect 20302 11118 20354 11170
rect 6534 10950 6586 11002
rect 6638 10950 6690 11002
rect 6742 10950 6794 11002
rect 11854 10950 11906 11002
rect 11958 10950 12010 11002
rect 12062 10950 12114 11002
rect 17174 10950 17226 11002
rect 17278 10950 17330 11002
rect 17382 10950 17434 11002
rect 22494 10950 22546 11002
rect 22598 10950 22650 11002
rect 22702 10950 22754 11002
rect 6862 10782 6914 10834
rect 19182 10782 19234 10834
rect 19854 10782 19906 10834
rect 5406 10670 5458 10722
rect 5518 10670 5570 10722
rect 6078 10670 6130 10722
rect 8094 10670 8146 10722
rect 16718 10670 16770 10722
rect 17726 10670 17778 10722
rect 18398 10670 18450 10722
rect 19070 10670 19122 10722
rect 19742 10670 19794 10722
rect 20414 10670 20466 10722
rect 21086 10670 21138 10722
rect 21758 10670 21810 10722
rect 21870 10670 21922 10722
rect 6750 10558 6802 10610
rect 7422 10558 7474 10610
rect 7534 10558 7586 10610
rect 8878 10558 8930 10610
rect 9886 10558 9938 10610
rect 10558 10558 10610 10610
rect 11230 10558 11282 10610
rect 12014 10558 12066 10610
rect 12686 10558 12738 10610
rect 12798 10558 12850 10610
rect 13358 10558 13410 10610
rect 13470 10558 13522 10610
rect 14030 10558 14082 10610
rect 14142 10558 14194 10610
rect 14702 10558 14754 10610
rect 14814 10558 14866 10610
rect 15374 10558 15426 10610
rect 15486 10558 15538 10610
rect 16046 10558 16098 10610
rect 6190 10334 6242 10386
rect 8206 10334 8258 10386
rect 8990 10334 9042 10386
rect 9998 10334 10050 10386
rect 10670 10334 10722 10386
rect 11342 10334 11394 10386
rect 12126 10334 12178 10386
rect 16158 10334 16210 10386
rect 16830 10334 16882 10386
rect 17838 10334 17890 10386
rect 18510 10334 18562 10386
rect 20526 10334 20578 10386
rect 21198 10334 21250 10386
rect 3874 10166 3926 10218
rect 3978 10166 4030 10218
rect 4082 10166 4134 10218
rect 9194 10166 9246 10218
rect 9298 10166 9350 10218
rect 9402 10166 9454 10218
rect 14514 10166 14566 10218
rect 14618 10166 14670 10218
rect 14722 10166 14774 10218
rect 19834 10166 19886 10218
rect 19938 10166 19990 10218
rect 20042 10166 20094 10218
rect 11566 9998 11618 10050
rect 18510 9998 18562 10050
rect 20526 9998 20578 10050
rect 21758 9998 21810 10050
rect 4174 9774 4226 9826
rect 4286 9774 4338 9826
rect 4846 9774 4898 9826
rect 7870 9774 7922 9826
rect 8542 9774 8594 9826
rect 9214 9774 9266 9826
rect 10558 9774 10610 9826
rect 12126 9774 12178 9826
rect 12238 9774 12290 9826
rect 14478 9774 14530 9826
rect 15038 9774 15090 9826
rect 15710 9774 15762 9826
rect 17838 9774 17890 9826
rect 19070 9774 19122 9826
rect 19742 9774 19794 9826
rect 20414 9774 20466 9826
rect 21646 9774 21698 9826
rect 5854 9662 5906 9714
rect 6526 9662 6578 9714
rect 6638 9662 6690 9714
rect 7198 9662 7250 9714
rect 7310 9662 7362 9714
rect 9886 9662 9938 9714
rect 11454 9662 11506 9714
rect 12798 9662 12850 9714
rect 12910 9662 12962 9714
rect 13694 9662 13746 9714
rect 13806 9662 13858 9714
rect 14366 9662 14418 9714
rect 16382 9662 16434 9714
rect 17054 9662 17106 9714
rect 18398 9662 18450 9714
rect 4958 9550 5010 9602
rect 5966 9550 6018 9602
rect 7982 9550 8034 9602
rect 8654 9550 8706 9602
rect 9326 9550 9378 9602
rect 9998 9550 10050 9602
rect 10670 9550 10722 9602
rect 15150 9550 15202 9602
rect 15822 9550 15874 9602
rect 16494 9550 16546 9602
rect 17166 9550 17218 9602
rect 17726 9550 17778 9602
rect 19182 9550 19234 9602
rect 19854 9550 19906 9602
rect 6534 9382 6586 9434
rect 6638 9382 6690 9434
rect 6742 9382 6794 9434
rect 11854 9382 11906 9434
rect 11958 9382 12010 9434
rect 12062 9382 12114 9434
rect 17174 9382 17226 9434
rect 17278 9382 17330 9434
rect 17382 9382 17434 9434
rect 22494 9382 22546 9434
rect 22598 9382 22650 9434
rect 22702 9382 22754 9434
rect 4846 9214 4898 9266
rect 8990 9214 9042 9266
rect 14478 9214 14530 9266
rect 15150 9214 15202 9266
rect 19854 9214 19906 9266
rect 20526 9214 20578 9266
rect 3390 9102 3442 9154
rect 3502 9102 3554 9154
rect 4062 9102 4114 9154
rect 7422 9102 7474 9154
rect 7534 9102 7586 9154
rect 8206 9102 8258 9154
rect 10334 9102 10386 9154
rect 12350 9102 12402 9154
rect 13022 9102 13074 9154
rect 15710 9102 15762 9154
rect 17726 9102 17778 9154
rect 19070 9102 19122 9154
rect 20414 9102 20466 9154
rect 4734 8990 4786 9042
rect 5406 8990 5458 9042
rect 6078 8990 6130 9042
rect 6190 8990 6242 9042
rect 6750 8990 6802 9042
rect 6862 8990 6914 9042
rect 8878 8990 8930 9042
rect 11006 8990 11058 9042
rect 11678 8990 11730 9042
rect 13694 8990 13746 9042
rect 14366 8990 14418 9042
rect 15038 8990 15090 9042
rect 16382 8990 16434 9042
rect 18398 8990 18450 9042
rect 19742 8990 19794 9042
rect 10446 8878 10498 8930
rect 4174 8766 4226 8818
rect 5518 8766 5570 8818
rect 8318 8766 8370 8818
rect 11118 8766 11170 8818
rect 11790 8766 11842 8818
rect 12462 8766 12514 8818
rect 13134 8766 13186 8818
rect 13806 8766 13858 8818
rect 15822 8766 15874 8818
rect 16494 8766 16546 8818
rect 17838 8766 17890 8818
rect 18510 8766 18562 8818
rect 19182 8766 19234 8818
rect 3874 8598 3926 8650
rect 3978 8598 4030 8650
rect 4082 8598 4134 8650
rect 9194 8598 9246 8650
rect 9298 8598 9350 8650
rect 9402 8598 9454 8650
rect 14514 8598 14566 8650
rect 14618 8598 14670 8650
rect 14722 8598 14774 8650
rect 19834 8598 19886 8650
rect 19938 8598 19990 8650
rect 20042 8598 20094 8650
rect 4958 8430 5010 8482
rect 5966 8430 6018 8482
rect 6638 8430 6690 8482
rect 9326 8430 9378 8482
rect 9998 8430 10050 8482
rect 10670 8430 10722 8482
rect 15150 8430 15202 8482
rect 17166 8430 17218 8482
rect 17838 8430 17890 8482
rect 18510 8430 18562 8482
rect 19182 8430 19234 8482
rect 11230 8318 11282 8370
rect 6526 8206 6578 8258
rect 7198 8206 7250 8258
rect 7870 8206 7922 8258
rect 9214 8206 9266 8258
rect 9886 8206 9938 8258
rect 10558 8206 10610 8258
rect 12126 8206 12178 8258
rect 12238 8206 12290 8258
rect 12910 8206 12962 8258
rect 13694 8206 13746 8258
rect 13806 8206 13858 8258
rect 14366 8206 14418 8258
rect 14478 8206 14530 8258
rect 15038 8206 15090 8258
rect 15822 8206 15874 8258
rect 16494 8206 16546 8258
rect 17054 8206 17106 8258
rect 18398 8206 18450 8258
rect 19070 8206 19122 8258
rect 19742 8206 19794 8258
rect 19854 8206 19906 8258
rect 2942 8094 2994 8146
rect 3502 8094 3554 8146
rect 4174 8094 4226 8146
rect 4846 8094 4898 8146
rect 5854 8094 5906 8146
rect 8542 8094 8594 8146
rect 11342 8094 11394 8146
rect 12798 8094 12850 8146
rect 15710 8094 15762 8146
rect 16382 8094 16434 8146
rect 17726 8094 17778 8146
rect 20526 8094 20578 8146
rect 2830 7982 2882 8034
rect 3614 7982 3666 8034
rect 4286 7982 4338 8034
rect 7310 7982 7362 8034
rect 7982 7982 8034 8034
rect 8654 7982 8706 8034
rect 20414 7982 20466 8034
rect 6534 7814 6586 7866
rect 6638 7814 6690 7866
rect 6742 7814 6794 7866
rect 11854 7814 11906 7866
rect 11958 7814 12010 7866
rect 12062 7814 12114 7866
rect 17174 7814 17226 7866
rect 17278 7814 17330 7866
rect 17382 7814 17434 7866
rect 22494 7814 22546 7866
rect 22598 7814 22650 7866
rect 22702 7814 22754 7866
rect 6190 7646 6242 7698
rect 6862 7646 6914 7698
rect 8990 7646 9042 7698
rect 9998 7646 10050 7698
rect 10670 7646 10722 7698
rect 11230 7646 11282 7698
rect 13358 7646 13410 7698
rect 14702 7646 14754 7698
rect 16718 7646 16770 7698
rect 17838 7646 17890 7698
rect 18510 7646 18562 7698
rect 4734 7534 4786 7586
rect 10558 7534 10610 7586
rect 13918 7534 13970 7586
rect 15262 7534 15314 7586
rect 15934 7534 15986 7586
rect 2158 7422 2210 7474
rect 2718 7422 2770 7474
rect 3390 7422 3442 7474
rect 4062 7422 4114 7474
rect 4846 7422 4898 7474
rect 5406 7422 5458 7474
rect 6078 7422 6130 7474
rect 6750 7422 6802 7474
rect 7422 7422 7474 7474
rect 8206 7422 8258 7474
rect 8878 7422 8930 7474
rect 9886 7422 9938 7474
rect 11342 7422 11394 7474
rect 11902 7422 11954 7474
rect 12574 7422 12626 7474
rect 13246 7422 13298 7474
rect 14590 7422 14642 7474
rect 16606 7422 16658 7474
rect 17726 7422 17778 7474
rect 18398 7422 18450 7474
rect 19070 7422 19122 7474
rect 19742 7422 19794 7474
rect 20414 7422 20466 7474
rect 21086 7422 21138 7474
rect 14030 7310 14082 7362
rect 2046 7198 2098 7250
rect 2830 7198 2882 7250
rect 3502 7198 3554 7250
rect 4174 7198 4226 7250
rect 5518 7198 5570 7250
rect 7534 7198 7586 7250
rect 8318 7198 8370 7250
rect 12014 7198 12066 7250
rect 12686 7198 12738 7250
rect 15374 7198 15426 7250
rect 16046 7198 16098 7250
rect 19182 7198 19234 7250
rect 19854 7198 19906 7250
rect 20526 7198 20578 7250
rect 21198 7198 21250 7250
rect 3874 7030 3926 7082
rect 3978 7030 4030 7082
rect 4082 7030 4134 7082
rect 9194 7030 9246 7082
rect 9298 7030 9350 7082
rect 9402 7030 9454 7082
rect 14514 7030 14566 7082
rect 14618 7030 14670 7082
rect 14722 7030 14774 7082
rect 19834 7030 19886 7082
rect 19938 7030 19990 7082
rect 20042 7030 20094 7082
rect 4286 6862 4338 6914
rect 4958 6862 5010 6914
rect 10558 6862 10610 6914
rect 11230 6862 11282 6914
rect 14254 6862 14306 6914
rect 14926 6862 14978 6914
rect 15598 6862 15650 6914
rect 17614 6862 17666 6914
rect 19630 6862 19682 6914
rect 5742 6638 5794 6690
rect 5854 6638 5906 6690
rect 6414 6638 6466 6690
rect 6526 6638 6578 6690
rect 8542 6638 8594 6690
rect 9214 6638 9266 6690
rect 9774 6638 9826 6690
rect 10446 6638 10498 6690
rect 11118 6638 11170 6690
rect 11790 6638 11842 6690
rect 12462 6638 12514 6690
rect 14142 6638 14194 6690
rect 14814 6638 14866 6690
rect 15486 6638 15538 6690
rect 18958 6638 19010 6690
rect 21646 6638 21698 6690
rect 2158 6526 2210 6578
rect 2830 6526 2882 6578
rect 3502 6526 3554 6578
rect 4174 6526 4226 6578
rect 4846 6526 4898 6578
rect 7086 6526 7138 6578
rect 7758 6526 7810 6578
rect 8430 6526 8482 6578
rect 9102 6526 9154 6578
rect 16158 6526 16210 6578
rect 16270 6526 16322 6578
rect 16830 6526 16882 6578
rect 16942 6526 16994 6578
rect 17502 6526 17554 6578
rect 18174 6526 18226 6578
rect 18846 6526 18898 6578
rect 19518 6526 19570 6578
rect 20302 6526 20354 6578
rect 2270 6414 2322 6466
rect 2942 6414 2994 6466
rect 3614 6414 3666 6466
rect 7198 6414 7250 6466
rect 7870 6414 7922 6466
rect 9886 6414 9938 6466
rect 11902 6414 11954 6466
rect 12574 6414 12626 6466
rect 18286 6414 18338 6466
rect 20190 6414 20242 6466
rect 21758 6414 21810 6466
rect 6534 6246 6586 6298
rect 6638 6246 6690 6298
rect 6742 6246 6794 6298
rect 11854 6246 11906 6298
rect 11958 6246 12010 6298
rect 12062 6246 12114 6298
rect 17174 6246 17226 6298
rect 17278 6246 17330 6298
rect 17382 6246 17434 6298
rect 22494 6246 22546 6298
rect 22598 6246 22650 6298
rect 22702 6246 22754 6298
rect 5518 6078 5570 6130
rect 6190 6078 6242 6130
rect 8878 6078 8930 6130
rect 9886 6078 9938 6130
rect 10558 6078 10610 6130
rect 11230 6078 11282 6130
rect 11902 6078 11954 6130
rect 13358 6078 13410 6130
rect 14030 6078 14082 6130
rect 14702 6078 14754 6130
rect 15374 6078 15426 6130
rect 16046 6078 16098 6130
rect 16718 6078 16770 6130
rect 6750 5966 6802 6018
rect 6862 5966 6914 6018
rect 7422 5966 7474 6018
rect 8094 5966 8146 6018
rect 8766 5966 8818 6018
rect 11118 5966 11170 6018
rect 11790 5966 11842 6018
rect 12574 5966 12626 6018
rect 14590 5966 14642 6018
rect 15262 5966 15314 6018
rect 15934 5966 15986 6018
rect 16606 5966 16658 6018
rect 19070 5966 19122 6018
rect 19742 5966 19794 6018
rect 2046 5854 2098 5906
rect 2718 5854 2770 5906
rect 3390 5854 3442 5906
rect 4062 5854 4114 5906
rect 4734 5854 4786 5906
rect 5406 5854 5458 5906
rect 6078 5854 6130 5906
rect 9774 5854 9826 5906
rect 10446 5854 10498 5906
rect 13246 5854 13298 5906
rect 13918 5854 13970 5906
rect 17726 5854 17778 5906
rect 18398 5854 18450 5906
rect 20414 5854 20466 5906
rect 21086 5854 21138 5906
rect 21870 5854 21922 5906
rect 18510 5742 18562 5794
rect 19182 5742 19234 5794
rect 2158 5630 2210 5682
rect 2830 5630 2882 5682
rect 3502 5630 3554 5682
rect 4174 5630 4226 5682
rect 4846 5630 4898 5682
rect 7534 5630 7586 5682
rect 8206 5630 8258 5682
rect 12686 5630 12738 5682
rect 17838 5630 17890 5682
rect 19854 5630 19906 5682
rect 20526 5630 20578 5682
rect 21198 5630 21250 5682
rect 21758 5630 21810 5682
rect 3874 5462 3926 5514
rect 3978 5462 4030 5514
rect 4082 5462 4134 5514
rect 9194 5462 9246 5514
rect 9298 5462 9350 5514
rect 9402 5462 9454 5514
rect 14514 5462 14566 5514
rect 14618 5462 14670 5514
rect 14722 5462 14774 5514
rect 19834 5462 19886 5514
rect 19938 5462 19990 5514
rect 20042 5462 20094 5514
rect 5854 5294 5906 5346
rect 6526 5294 6578 5346
rect 7198 5294 7250 5346
rect 8542 5294 8594 5346
rect 9886 5294 9938 5346
rect 10558 5294 10610 5346
rect 14142 5294 14194 5346
rect 14814 5294 14866 5346
rect 15486 5294 15538 5346
rect 18174 5294 18226 5346
rect 20190 5294 20242 5346
rect 19518 5182 19570 5234
rect 4174 5070 4226 5122
rect 4846 5070 4898 5122
rect 7086 5070 7138 5122
rect 7758 5070 7810 5122
rect 7870 5070 7922 5122
rect 8430 5070 8482 5122
rect 9102 5070 9154 5122
rect 9214 5070 9266 5122
rect 10446 5070 10498 5122
rect 11454 5070 11506 5122
rect 11566 5070 11618 5122
rect 15374 5070 15426 5122
rect 16830 5070 16882 5122
rect 17390 5070 17442 5122
rect 18062 5070 18114 5122
rect 18734 5070 18786 5122
rect 18846 5070 18898 5122
rect 19406 5070 19458 5122
rect 20078 5070 20130 5122
rect 2158 4958 2210 5010
rect 2830 4958 2882 5010
rect 3502 4958 3554 5010
rect 3614 4958 3666 5010
rect 5742 4958 5794 5010
rect 6414 4958 6466 5010
rect 9774 4958 9826 5010
rect 12126 4958 12178 5010
rect 12798 4958 12850 5010
rect 14030 4958 14082 5010
rect 14702 4958 14754 5010
rect 16046 4958 16098 5010
rect 16718 4958 16770 5010
rect 20750 4958 20802 5010
rect 21646 4958 21698 5010
rect 2270 4846 2322 4898
rect 2942 4846 2994 4898
rect 4286 4846 4338 4898
rect 4958 4846 5010 4898
rect 12238 4846 12290 4898
rect 12910 4846 12962 4898
rect 16158 4846 16210 4898
rect 17502 4846 17554 4898
rect 20862 4846 20914 4898
rect 21758 4846 21810 4898
rect 6534 4678 6586 4730
rect 6638 4678 6690 4730
rect 6742 4678 6794 4730
rect 11854 4678 11906 4730
rect 11958 4678 12010 4730
rect 12062 4678 12114 4730
rect 17174 4678 17226 4730
rect 17278 4678 17330 4730
rect 17382 4678 17434 4730
rect 22494 4678 22546 4730
rect 22598 4678 22650 4730
rect 22702 4678 22754 4730
rect 3838 4510 3890 4562
rect 4510 4510 4562 4562
rect 7198 4510 7250 4562
rect 8542 4510 8594 4562
rect 15150 4510 15202 4562
rect 15822 4510 15874 4562
rect 17838 4510 17890 4562
rect 18510 4510 18562 4562
rect 19854 4510 19906 4562
rect 20526 4510 20578 4562
rect 21198 4510 21250 4562
rect 2382 4398 2434 4450
rect 5070 4398 5122 4450
rect 5742 4398 5794 4450
rect 8430 4398 8482 4450
rect 9774 4398 9826 4450
rect 10446 4398 10498 4450
rect 14366 4398 14418 4450
rect 16382 4398 16434 4450
rect 16494 4398 16546 4450
rect 17726 4398 17778 4450
rect 18398 4398 18450 4450
rect 19070 4398 19122 4450
rect 20414 4398 20466 4450
rect 21086 4398 21138 4450
rect 2494 4286 2546 4338
rect 3054 4286 3106 4338
rect 3166 4286 3218 4338
rect 3726 4286 3778 4338
rect 4398 4286 4450 4338
rect 6414 4286 6466 4338
rect 7086 4286 7138 4338
rect 7758 4286 7810 4338
rect 11118 4286 11170 4338
rect 12350 4286 12402 4338
rect 13022 4286 13074 4338
rect 13694 4286 13746 4338
rect 14478 4286 14530 4338
rect 15038 4286 15090 4338
rect 15710 4286 15762 4338
rect 19742 4286 19794 4338
rect 21870 4286 21922 4338
rect 5182 4062 5234 4114
rect 5854 4062 5906 4114
rect 6526 4062 6578 4114
rect 7870 4062 7922 4114
rect 9886 4062 9938 4114
rect 10558 4062 10610 4114
rect 11230 4062 11282 4114
rect 12462 4062 12514 4114
rect 13134 4062 13186 4114
rect 13806 4062 13858 4114
rect 19182 4062 19234 4114
rect 21758 4062 21810 4114
rect 3874 3894 3926 3946
rect 3978 3894 4030 3946
rect 4082 3894 4134 3946
rect 9194 3894 9246 3946
rect 9298 3894 9350 3946
rect 9402 3894 9454 3946
rect 14514 3894 14566 3946
rect 14618 3894 14670 3946
rect 14722 3894 14774 3946
rect 19834 3894 19886 3946
rect 19938 3894 19990 3946
rect 20042 3894 20094 3946
rect 2942 3726 2994 3778
rect 3614 3726 3666 3778
rect 4286 3726 4338 3778
rect 4958 3726 5010 3778
rect 6414 3726 6466 3778
rect 7086 3726 7138 3778
rect 7870 3726 7922 3778
rect 17614 3726 17666 3778
rect 19630 3726 19682 3778
rect 20302 3726 20354 3778
rect 2830 3502 2882 3554
rect 3502 3502 3554 3554
rect 4174 3502 4226 3554
rect 5854 3502 5906 3554
rect 6526 3502 6578 3554
rect 7198 3502 7250 3554
rect 7758 3502 7810 3554
rect 8430 3502 8482 3554
rect 8542 3502 8594 3554
rect 9662 3502 9714 3554
rect 9774 3502 9826 3554
rect 10334 3502 10386 3554
rect 10446 3502 10498 3554
rect 11118 3502 11170 3554
rect 11678 3502 11730 3554
rect 14590 3502 14642 3554
rect 15262 3502 15314 3554
rect 15598 3502 15650 3554
rect 15822 3502 15874 3554
rect 16606 3502 16658 3554
rect 17502 3502 17554 3554
rect 18174 3502 18226 3554
rect 18846 3502 18898 3554
rect 20190 3502 20242 3554
rect 4846 3390 4898 3442
rect 5742 3390 5794 3442
rect 11006 3390 11058 3442
rect 11790 3390 11842 3442
rect 13918 3390 13970 3442
rect 14030 3390 14082 3442
rect 14702 3390 14754 3442
rect 15374 3390 15426 3442
rect 15934 3390 15986 3442
rect 16046 3390 16098 3442
rect 16718 3390 16770 3442
rect 18286 3390 18338 3442
rect 18958 3390 19010 3442
rect 19518 3390 19570 3442
rect 6534 3110 6586 3162
rect 6638 3110 6690 3162
rect 6742 3110 6794 3162
rect 11854 3110 11906 3162
rect 11958 3110 12010 3162
rect 12062 3110 12114 3162
rect 17174 3110 17226 3162
rect 17278 3110 17330 3162
rect 17382 3110 17434 3162
rect 22494 3110 22546 3162
rect 22598 3110 22650 3162
rect 22702 3110 22754 3162
<< metal2 >>
rect 3872 16492 4136 16502
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 3872 16426 4136 16436
rect 9192 16492 9456 16502
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9192 16426 9456 16436
rect 14512 16492 14776 16502
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14512 16426 14776 16436
rect 19832 16492 20096 16502
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 19832 16426 20096 16436
rect 6532 15708 6796 15718
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6532 15642 6796 15652
rect 11852 15708 12116 15718
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 11852 15642 12116 15652
rect 17172 15708 17436 15718
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17172 15642 17436 15652
rect 22492 15708 22756 15718
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22492 15642 22756 15652
rect 3612 14980 3668 14990
rect 3388 9156 3444 9166
rect 3500 9156 3556 9166
rect 3388 9154 3500 9156
rect 3388 9102 3390 9154
rect 3442 9102 3500 9154
rect 3388 9100 3500 9102
rect 2940 8148 2996 8158
rect 3388 8148 3444 9100
rect 3500 9062 3556 9100
rect 3612 8484 3668 14924
rect 3872 14924 4136 14934
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 3872 14858 4136 14868
rect 9192 14924 9456 14934
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9192 14858 9456 14868
rect 14512 14924 14776 14934
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14512 14858 14776 14868
rect 19832 14924 20096 14934
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 19832 14858 20096 14868
rect 19628 14756 19684 14766
rect 16828 14644 16884 14654
rect 16828 14642 17108 14644
rect 16828 14590 16830 14642
rect 16882 14590 17108 14642
rect 16828 14588 17108 14590
rect 16828 14578 16884 14588
rect 16940 14418 16996 14430
rect 16940 14366 16942 14418
rect 16994 14366 16996 14418
rect 6532 14140 6796 14150
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6532 14074 6796 14084
rect 11852 14140 12116 14150
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 11852 14074 12116 14084
rect 16156 13746 16212 13758
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 3872 13356 4136 13366
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 3872 13290 4136 13300
rect 9192 13356 9456 13366
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9192 13290 9456 13300
rect 14512 13356 14776 13366
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14512 13290 14776 13300
rect 14924 13188 14980 13198
rect 14924 13094 14980 13132
rect 16156 13076 16212 13694
rect 16828 13746 16884 13758
rect 16828 13694 16830 13746
rect 16882 13694 16884 13746
rect 16268 13524 16324 13534
rect 16268 13430 16324 13468
rect 16156 13020 16324 13076
rect 14812 12852 14868 12862
rect 14812 12850 15092 12852
rect 14812 12798 14814 12850
rect 14866 12798 15092 12850
rect 14812 12796 15092 12798
rect 14812 12786 14868 12796
rect 6532 12572 6796 12582
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6532 12506 6796 12516
rect 11852 12572 12116 12582
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 11852 12506 12116 12516
rect 14140 12178 14196 12190
rect 14140 12126 14142 12178
rect 14194 12126 14196 12178
rect 3872 11788 4136 11798
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 3872 11722 4136 11732
rect 9192 11788 9456 11798
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9192 11722 9456 11732
rect 10668 11508 10724 11518
rect 7532 11452 8148 11508
rect 6076 11284 6132 11294
rect 6188 11284 6244 11294
rect 6076 11282 6188 11284
rect 6076 11230 6078 11282
rect 6130 11230 6188 11282
rect 6076 11228 6188 11230
rect 5404 10724 5460 10734
rect 5516 10724 5572 10734
rect 5404 10722 5516 10724
rect 5404 10670 5406 10722
rect 5458 10670 5516 10722
rect 5404 10668 5516 10670
rect 3872 10220 4136 10230
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 3872 10154 4136 10164
rect 4172 9828 4228 9838
rect 4284 9828 4340 9838
rect 4172 9826 4284 9828
rect 4172 9774 4174 9826
rect 4226 9774 4284 9826
rect 4172 9772 4284 9774
rect 4060 9156 4116 9166
rect 4172 9156 4228 9772
rect 4284 9734 4340 9772
rect 4844 9828 4900 9838
rect 4844 9734 4900 9772
rect 5404 9828 5460 10668
rect 5516 10630 5572 10668
rect 6076 10724 6132 11228
rect 6188 11190 6244 11228
rect 6972 11284 7028 11294
rect 6972 11190 7028 11228
rect 6860 11170 6916 11182
rect 7532 11172 7588 11452
rect 7644 11284 7700 11294
rect 7644 11282 7812 11284
rect 7644 11230 7646 11282
rect 7698 11230 7812 11282
rect 7644 11228 7812 11230
rect 7644 11218 7700 11228
rect 6860 11118 6862 11170
rect 6914 11118 6916 11170
rect 6860 11060 6916 11118
rect 7420 11170 7588 11172
rect 7420 11118 7534 11170
rect 7586 11118 7588 11170
rect 7420 11116 7588 11118
rect 7756 11172 7812 11228
rect 8092 11172 8148 11452
rect 10444 11506 10724 11508
rect 10444 11454 10670 11506
rect 10722 11454 10724 11506
rect 10444 11452 10724 11454
rect 8316 11282 8372 11294
rect 8316 11230 8318 11282
rect 8370 11230 8372 11282
rect 8204 11172 8260 11182
rect 7756 11116 7924 11172
rect 7420 11060 7476 11116
rect 7532 11106 7588 11116
rect 6532 11004 6796 11014
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6532 10938 6796 10948
rect 6860 11004 7476 11060
rect 6860 10836 6916 11004
rect 6076 10592 6132 10668
rect 6188 10834 6916 10836
rect 6188 10782 6862 10834
rect 6914 10782 6916 10834
rect 6188 10780 6916 10782
rect 5404 9762 5460 9772
rect 6188 10386 6244 10780
rect 6860 10770 6916 10780
rect 6748 10612 6804 10622
rect 7420 10612 7476 10622
rect 7532 10612 7588 10622
rect 7868 10612 7924 11116
rect 8092 11170 8260 11172
rect 8092 11118 8206 11170
rect 8258 11118 8260 11170
rect 8092 11116 8260 11118
rect 8092 10722 8148 11116
rect 8204 11106 8260 11116
rect 8092 10670 8094 10722
rect 8146 10670 8148 10722
rect 8092 10658 8148 10670
rect 6636 10610 6804 10612
rect 6636 10558 6750 10610
rect 6802 10558 6804 10610
rect 6636 10556 6804 10558
rect 6636 10500 6692 10556
rect 6748 10546 6804 10556
rect 7308 10610 7924 10612
rect 7308 10558 7422 10610
rect 7474 10558 7534 10610
rect 7586 10558 7924 10610
rect 7308 10556 7924 10558
rect 6188 10334 6190 10386
rect 6242 10334 6244 10386
rect 5852 9716 5908 9726
rect 5740 9660 5852 9716
rect 4956 9602 5012 9614
rect 4956 9550 4958 9602
rect 5010 9550 5012 9602
rect 4116 9100 4228 9156
rect 4844 9268 4900 9278
rect 4956 9268 5012 9550
rect 4844 9266 5012 9268
rect 4844 9214 4846 9266
rect 4898 9214 5012 9266
rect 4844 9212 5012 9214
rect 4060 9024 4116 9100
rect 4732 9042 4788 9054
rect 4732 8990 4734 9042
rect 4786 8990 4788 9042
rect 4172 8820 4228 8830
rect 4172 8818 4340 8820
rect 4172 8766 4174 8818
rect 4226 8766 4340 8818
rect 4172 8764 4340 8766
rect 4172 8754 4228 8764
rect 3872 8652 4136 8662
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 3872 8586 4136 8596
rect 2940 8146 3444 8148
rect 2940 8094 2942 8146
rect 2994 8094 3444 8146
rect 2940 8092 3444 8094
rect 3500 8372 3668 8428
rect 4172 8484 4228 8494
rect 3500 8146 3556 8372
rect 3500 8094 3502 8146
rect 3554 8094 3556 8146
rect 2828 8034 2884 8046
rect 2828 7982 2830 8034
rect 2882 7982 2884 8034
rect 2828 7700 2884 7982
rect 2604 7644 2884 7700
rect 2156 7476 2212 7486
rect 2156 7382 2212 7420
rect 2044 7252 2100 7262
rect 2604 7252 2660 7644
rect 2044 7250 2660 7252
rect 2044 7198 2046 7250
rect 2098 7198 2660 7250
rect 2044 7196 2660 7198
rect 2716 7476 2772 7486
rect 2940 7476 2996 8092
rect 2772 7420 2996 7476
rect 3388 7476 3444 7486
rect 3500 7476 3556 8094
rect 4172 8146 4228 8428
rect 4172 8094 4174 8146
rect 4226 8094 4228 8146
rect 3612 8036 3668 8046
rect 3612 8034 3780 8036
rect 3612 7982 3614 8034
rect 3666 7982 3780 8034
rect 3612 7980 3780 7982
rect 3612 7970 3668 7980
rect 3388 7474 3556 7476
rect 3388 7422 3390 7474
rect 3442 7422 3556 7474
rect 3388 7420 3556 7422
rect 2044 5906 2100 7196
rect 2156 6580 2212 6590
rect 2156 6486 2212 6524
rect 2044 5854 2046 5906
rect 2098 5854 2100 5906
rect 2044 5012 2100 5854
rect 2268 6466 2324 6478
rect 2268 6414 2270 6466
rect 2322 6414 2324 6466
rect 2156 5684 2212 5694
rect 2268 5684 2324 6414
rect 2716 5908 2772 7420
rect 2828 7250 2884 7262
rect 2828 7198 2830 7250
rect 2882 7198 2884 7250
rect 2828 6804 2884 7198
rect 2828 6738 2884 6748
rect 2828 6580 2884 6590
rect 2828 6486 2884 6524
rect 3388 6580 3444 7420
rect 3500 7252 3556 7262
rect 3612 7252 3668 7262
rect 3500 7250 3612 7252
rect 3500 7198 3502 7250
rect 3554 7198 3612 7250
rect 3500 7196 3612 7198
rect 3500 7186 3556 7196
rect 3500 6580 3556 6590
rect 3444 6578 3556 6580
rect 3444 6526 3502 6578
rect 3554 6526 3556 6578
rect 3444 6524 3556 6526
rect 2940 6466 2996 6478
rect 2940 6414 2942 6466
rect 2994 6414 2996 6466
rect 2940 5908 2996 6414
rect 2716 5906 2996 5908
rect 2716 5854 2718 5906
rect 2770 5854 2996 5906
rect 2716 5852 2996 5854
rect 3388 5906 3444 6524
rect 3500 6514 3556 6524
rect 3388 5854 3390 5906
rect 3442 5854 3444 5906
rect 2716 5684 2772 5852
rect 2156 5682 2772 5684
rect 2156 5630 2158 5682
rect 2210 5630 2772 5682
rect 2156 5628 2772 5630
rect 2828 5682 2884 5694
rect 2828 5630 2830 5682
rect 2882 5630 2884 5682
rect 2156 5618 2212 5628
rect 2156 5012 2212 5022
rect 2044 5010 2212 5012
rect 2044 4958 2158 5010
rect 2210 4958 2212 5010
rect 2044 4956 2212 4958
rect 2156 4452 2212 4956
rect 2268 4898 2324 5628
rect 2828 5572 2884 5630
rect 2716 5516 2884 5572
rect 2716 5124 2772 5516
rect 2716 5058 2772 5068
rect 3388 5124 3444 5854
rect 3612 6466 3668 7196
rect 3724 6804 3780 7980
rect 4060 7476 4116 7486
rect 4172 7476 4228 8094
rect 4284 8036 4340 8764
rect 4284 7942 4340 7980
rect 4732 8484 4788 8990
rect 4732 7586 4788 8428
rect 4732 7534 4734 7586
rect 4786 7534 4788 7586
rect 4060 7474 4340 7476
rect 4060 7422 4062 7474
rect 4114 7422 4340 7474
rect 4060 7420 4340 7422
rect 4060 7410 4116 7420
rect 4172 7252 4228 7290
rect 4172 7186 4228 7196
rect 3872 7084 4136 7094
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 3872 7018 4136 7028
rect 4284 6914 4340 7420
rect 4284 6862 4286 6914
rect 4338 6862 4340 6914
rect 4284 6850 4340 6862
rect 4732 6916 4788 7534
rect 4844 8146 4900 9212
rect 5404 9044 5460 9054
rect 5740 9044 5796 9660
rect 5852 9584 5908 9660
rect 5964 9604 6020 9614
rect 6188 9604 6244 10334
rect 6524 10444 6692 10500
rect 6524 9716 6580 10444
rect 6636 9716 6692 9726
rect 6580 9714 6692 9716
rect 6580 9662 6638 9714
rect 6690 9662 6692 9714
rect 6580 9660 6692 9662
rect 6524 9622 6580 9660
rect 6636 9650 6692 9660
rect 7196 9716 7252 9726
rect 7308 9716 7364 10556
rect 7420 10546 7476 10556
rect 7532 10546 7588 10556
rect 7868 10388 7924 10556
rect 8204 10388 8260 10398
rect 8316 10388 8372 11230
rect 9212 11282 9268 11294
rect 9212 11230 9214 11282
rect 9266 11230 9268 11282
rect 7868 10386 8372 10388
rect 7868 10334 8206 10386
rect 8258 10334 8372 10386
rect 7868 10332 8372 10334
rect 7868 9826 7924 10332
rect 8204 10322 8260 10332
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9762 7924 9774
rect 8316 9828 8372 10332
rect 8876 10612 8932 10622
rect 9212 10612 9268 11230
rect 9884 11282 9940 11294
rect 9884 11230 9886 11282
rect 9938 11230 9940 11282
rect 8876 10610 9268 10612
rect 8876 10558 8878 10610
rect 8930 10558 9268 10610
rect 8876 10556 9268 10558
rect 9324 11170 9380 11182
rect 9324 11118 9326 11170
rect 9378 11118 9380 11170
rect 8540 9828 8596 9838
rect 8876 9828 8932 10556
rect 8988 10388 9044 10398
rect 9324 10388 9380 11118
rect 8988 10386 9380 10388
rect 8988 10334 8990 10386
rect 9042 10334 9380 10386
rect 8988 10332 9380 10334
rect 9884 10610 9940 11230
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 8988 10052 9044 10332
rect 9192 10220 9456 10230
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9192 10154 9456 10164
rect 8988 9986 9044 9996
rect 9884 9940 9940 10558
rect 9996 11172 10052 11182
rect 10444 11172 10500 11452
rect 10668 11442 10724 11452
rect 10556 11284 10612 11294
rect 12124 11284 12180 11294
rect 12236 11284 12292 11294
rect 10556 11282 10724 11284
rect 10556 11230 10558 11282
rect 10610 11230 10724 11282
rect 10556 11228 10724 11230
rect 10556 11218 10612 11228
rect 9996 11170 10500 11172
rect 9996 11118 9998 11170
rect 10050 11118 10500 11170
rect 9996 11116 10500 11118
rect 9996 10386 10052 11116
rect 9996 10334 9998 10386
rect 10050 10334 10052 10386
rect 9996 10164 10052 10334
rect 9996 10098 10052 10108
rect 10556 10610 10612 10622
rect 10556 10558 10558 10610
rect 10610 10558 10612 10610
rect 9212 9884 10052 9940
rect 9212 9828 9268 9884
rect 8316 9826 9268 9828
rect 8316 9774 8542 9826
rect 8594 9774 9214 9826
rect 9266 9774 9268 9826
rect 8316 9772 9268 9774
rect 8540 9762 8596 9772
rect 7252 9714 7364 9716
rect 7252 9662 7310 9714
rect 7362 9662 7364 9714
rect 7252 9660 7364 9662
rect 7196 9622 7252 9660
rect 5964 9602 6244 9604
rect 5964 9550 5966 9602
rect 6018 9550 6244 9602
rect 5964 9548 6244 9550
rect 5964 9492 6020 9548
rect 5404 9042 5796 9044
rect 5404 8990 5406 9042
rect 5458 8990 5796 9042
rect 5404 8988 5796 8990
rect 5852 9436 6020 9492
rect 6532 9436 6796 9446
rect 4956 8484 5012 8522
rect 4956 8418 5012 8428
rect 5404 8484 5460 8988
rect 5404 8418 5460 8428
rect 5516 8818 5572 8830
rect 5516 8766 5518 8818
rect 5570 8766 5572 8818
rect 4844 8094 4846 8146
rect 4898 8094 4900 8146
rect 4844 8036 4900 8094
rect 4844 7476 4900 7980
rect 5516 8148 5572 8766
rect 5852 8148 5908 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6532 9370 6796 9380
rect 7308 9156 7364 9660
rect 7980 9604 8036 9614
rect 8652 9604 8708 9614
rect 7980 9602 8260 9604
rect 7980 9550 7982 9602
rect 8034 9550 8260 9602
rect 7980 9548 8260 9550
rect 7420 9156 7476 9166
rect 7532 9156 7588 9166
rect 7308 9154 7588 9156
rect 7308 9102 7422 9154
rect 7474 9102 7534 9154
rect 7586 9102 7588 9154
rect 7308 9100 7588 9102
rect 6076 9044 6132 9054
rect 6188 9044 6244 9054
rect 6748 9044 6804 9054
rect 6860 9044 6916 9054
rect 6076 9042 6244 9044
rect 6076 8990 6078 9042
rect 6130 8990 6190 9042
rect 6242 8990 6244 9042
rect 6076 8988 6244 8990
rect 5964 8484 6020 8522
rect 6076 8428 6132 8988
rect 6188 8978 6244 8988
rect 6636 9042 6916 9044
rect 6636 8990 6750 9042
rect 6802 8990 6862 9042
rect 6914 8990 6916 9042
rect 6636 8988 6916 8990
rect 5964 8372 6132 8428
rect 5516 8146 5908 8148
rect 5516 8094 5854 8146
rect 5906 8094 5908 8146
rect 5516 8092 5908 8094
rect 4844 7382 4900 7420
rect 5404 7476 5460 7486
rect 5516 7476 5572 8092
rect 5852 8082 5908 8092
rect 6076 7700 6132 8372
rect 6524 8484 6580 8494
rect 6636 8484 6692 8988
rect 6748 8978 6804 8988
rect 6580 8482 6692 8484
rect 6580 8430 6638 8482
rect 6690 8430 6692 8482
rect 6580 8428 6692 8430
rect 6524 8258 6580 8428
rect 6636 8418 6692 8428
rect 6524 8206 6526 8258
rect 6578 8206 6580 8258
rect 6524 8194 6580 8206
rect 6532 7868 6796 7878
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6532 7802 6796 7812
rect 6188 7700 6244 7710
rect 6076 7698 6244 7700
rect 6076 7646 6190 7698
rect 6242 7646 6244 7698
rect 6076 7644 6244 7646
rect 5460 7420 5572 7476
rect 5404 7344 5460 7420
rect 5516 7250 5572 7420
rect 6076 7476 6132 7486
rect 6076 7382 6132 7420
rect 5516 7198 5518 7250
rect 5570 7198 5572 7250
rect 4956 6916 5012 6926
rect 4732 6914 5012 6916
rect 4732 6862 4958 6914
rect 5010 6862 5012 6914
rect 4732 6860 5012 6862
rect 4956 6850 5012 6860
rect 3724 6738 3780 6748
rect 4620 6804 4676 6814
rect 5516 6804 5572 7198
rect 4676 6748 4788 6804
rect 4620 6738 4676 6748
rect 3612 6414 3614 6466
rect 3666 6414 3668 6466
rect 3388 5058 3444 5068
rect 3500 5684 3556 5694
rect 3612 5684 3668 6414
rect 4172 6578 4228 6590
rect 4172 6526 4174 6578
rect 4226 6526 4228 6578
rect 4060 5908 4116 5918
rect 4060 5796 4116 5852
rect 3500 5682 3668 5684
rect 3500 5630 3502 5682
rect 3554 5630 3668 5682
rect 3500 5628 3668 5630
rect 3724 5740 4116 5796
rect 2828 5012 2884 5022
rect 2828 5010 2996 5012
rect 2828 4958 2830 5010
rect 2882 4958 2996 5010
rect 2828 4956 2996 4958
rect 2828 4946 2884 4956
rect 2268 4846 2270 4898
rect 2322 4846 2324 4898
rect 2268 4788 2324 4846
rect 2940 4900 2996 4956
rect 3500 5010 3556 5628
rect 3500 4958 3502 5010
rect 3554 4958 3556 5010
rect 2940 4898 3108 4900
rect 2940 4846 2942 4898
rect 2994 4846 3108 4898
rect 2940 4844 3108 4846
rect 2940 4834 2996 4844
rect 2268 4732 2548 4788
rect 2380 4452 2436 4462
rect 2156 4396 2380 4452
rect 2380 4358 2436 4396
rect 2492 4340 2548 4732
rect 3052 4452 3108 4844
rect 2492 4246 2548 4284
rect 2828 4340 2884 4350
rect 2156 3556 2212 3566
rect 2156 800 2212 3500
rect 2828 3556 2884 4284
rect 3052 4338 3108 4396
rect 3052 4286 3054 4338
rect 3106 4286 3108 4338
rect 2940 3780 2996 3790
rect 3052 3780 3108 4286
rect 3164 4340 3220 4350
rect 3164 4246 3220 4284
rect 3500 4340 3556 4958
rect 3612 5012 3668 5022
rect 3724 5012 3780 5740
rect 4172 5684 4228 6526
rect 4732 5908 4788 6748
rect 5516 6738 5572 6748
rect 5740 6804 5796 6814
rect 5740 6692 5796 6748
rect 5852 6692 5908 6702
rect 5740 6690 5908 6692
rect 5740 6638 5742 6690
rect 5794 6638 5854 6690
rect 5906 6638 5908 6690
rect 5740 6636 5908 6638
rect 5740 6626 5796 6636
rect 5852 6626 5908 6636
rect 4732 5814 4788 5852
rect 4844 6578 4900 6590
rect 4844 6526 4846 6578
rect 4898 6526 4900 6578
rect 4844 5684 4900 6526
rect 5516 6132 5572 6142
rect 6188 6132 6244 7644
rect 6860 7698 6916 8988
rect 7196 8484 7252 8494
rect 7196 8258 7252 8428
rect 7420 8428 7476 9100
rect 7532 9090 7588 9100
rect 7980 8484 8036 9548
rect 8204 9154 8260 9548
rect 8204 9102 8206 9154
rect 8258 9102 8260 9154
rect 8204 9090 8260 9102
rect 8540 9548 8652 9604
rect 7420 8372 7588 8428
rect 7196 8206 7198 8258
rect 7250 8206 7252 8258
rect 7196 8194 7252 8206
rect 6860 7646 6862 7698
rect 6914 7646 6916 7698
rect 6860 7634 6916 7646
rect 7308 8036 7364 8046
rect 6748 7476 6804 7486
rect 6412 6804 6468 6814
rect 6412 6692 6468 6748
rect 6524 6692 6580 6702
rect 6748 6692 6804 7420
rect 7308 7476 7364 7980
rect 7308 7410 7364 7420
rect 7420 7474 7476 7486
rect 7420 7422 7422 7474
rect 7474 7422 7476 7474
rect 7420 7252 7476 7422
rect 7532 7252 7588 8372
rect 7868 8372 8036 8428
rect 8316 8818 8372 8830
rect 8316 8766 8318 8818
rect 8370 8766 8372 8818
rect 7868 8258 7924 8372
rect 7868 8206 7870 8258
rect 7922 8206 7924 8258
rect 7868 8194 7924 8206
rect 7980 8036 8036 8046
rect 7980 7942 8036 7980
rect 8316 8036 8372 8766
rect 8540 8484 8596 9548
rect 8652 9472 8708 9548
rect 8988 9266 9044 9772
rect 9212 9762 9268 9772
rect 9884 9714 9940 9726
rect 9884 9662 9886 9714
rect 9938 9662 9940 9714
rect 9324 9604 9380 9614
rect 9324 9510 9380 9548
rect 8988 9214 8990 9266
rect 9042 9214 9044 9266
rect 8988 9202 9044 9214
rect 8540 8148 8596 8428
rect 8876 9042 8932 9054
rect 8876 8990 8878 9042
rect 8930 8990 8932 9042
rect 8876 8428 8932 8990
rect 9192 8652 9456 8662
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9192 8586 9456 8596
rect 9324 8484 9380 8522
rect 8876 8372 9044 8428
rect 9324 8418 9380 8428
rect 8316 7970 8372 7980
rect 8428 8146 8596 8148
rect 8428 8094 8542 8146
rect 8594 8094 8596 8146
rect 8428 8092 8596 8094
rect 8204 7476 8260 7486
rect 8428 7476 8484 8092
rect 8540 8082 8596 8092
rect 8652 8036 8708 8046
rect 8652 8034 8820 8036
rect 8652 7982 8654 8034
rect 8706 7982 8820 8034
rect 8652 7980 8820 7982
rect 8652 7970 8708 7980
rect 8204 7474 8484 7476
rect 8204 7422 8206 7474
rect 8258 7422 8484 7474
rect 8204 7420 8484 7422
rect 8204 7410 8260 7420
rect 7420 7250 7588 7252
rect 7420 7198 7534 7250
rect 7586 7198 7588 7250
rect 7420 7196 7588 7198
rect 7532 6916 7588 7196
rect 6412 6690 6916 6692
rect 6412 6638 6414 6690
rect 6466 6638 6526 6690
rect 6578 6638 6916 6690
rect 6412 6636 6916 6638
rect 6412 6626 6468 6636
rect 6524 6626 6580 6636
rect 6860 6580 6916 6636
rect 7084 6580 7140 6590
rect 6860 6578 7140 6580
rect 6860 6526 7086 6578
rect 7138 6526 7140 6578
rect 6860 6524 7140 6526
rect 6532 6300 6796 6310
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6532 6234 6796 6244
rect 5516 6130 6580 6132
rect 5516 6078 5518 6130
rect 5570 6078 6190 6130
rect 6242 6078 6580 6130
rect 5516 6076 6580 6078
rect 5516 6066 5572 6076
rect 4172 5682 4900 5684
rect 4172 5630 4174 5682
rect 4226 5630 4846 5682
rect 4898 5630 4900 5682
rect 4172 5628 4900 5630
rect 4172 5618 4228 5628
rect 3872 5516 4136 5526
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 3872 5450 4136 5460
rect 4172 5124 4228 5134
rect 4172 5030 4228 5068
rect 3668 4956 3780 5012
rect 3612 4564 3668 4956
rect 4284 4900 4340 4910
rect 4732 4900 4788 5628
rect 4844 5618 4900 5628
rect 5404 5906 5460 5918
rect 5404 5854 5406 5906
rect 5458 5854 5460 5906
rect 4284 4898 4452 4900
rect 4284 4846 4286 4898
rect 4338 4846 4452 4898
rect 4284 4844 4452 4846
rect 4284 4834 4340 4844
rect 3836 4564 3892 4574
rect 3612 4508 3836 4564
rect 3836 4432 3892 4508
rect 3500 4274 3556 4284
rect 3724 4340 3780 4350
rect 2940 3778 3108 3780
rect 2940 3726 2942 3778
rect 2994 3726 3108 3778
rect 2940 3724 3108 3726
rect 2940 3714 2996 3724
rect 2828 3424 2884 3500
rect 3052 3556 3108 3724
rect 3612 3780 3668 3790
rect 3724 3780 3780 4284
rect 4396 4340 4452 4844
rect 4732 4834 4788 4844
rect 4844 5122 4900 5134
rect 4844 5070 4846 5122
rect 4898 5070 4900 5122
rect 4508 4564 4564 4574
rect 4508 4470 4564 4508
rect 4844 4564 4900 5070
rect 4956 5124 5012 5134
rect 5012 5068 5124 5124
rect 4956 5058 5012 5068
rect 4956 4900 5012 4910
rect 4956 4806 5012 4844
rect 4284 4116 4340 4126
rect 3872 3948 4136 3958
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 3872 3882 4136 3892
rect 3612 3778 3780 3780
rect 3612 3726 3614 3778
rect 3666 3726 3780 3778
rect 3612 3724 3780 3726
rect 4284 3778 4340 4060
rect 4284 3726 4286 3778
rect 4338 3726 4340 3778
rect 3612 3714 3668 3724
rect 3052 3490 3108 3500
rect 3500 3556 3556 3566
rect 3500 3462 3556 3500
rect 4172 3556 4228 3566
rect 4284 3556 4340 3726
rect 4228 3500 4340 3556
rect 4172 3424 4228 3500
rect 4396 3444 4452 4284
rect 4844 3780 4900 4508
rect 5068 4450 5124 5068
rect 5404 4900 5460 5854
rect 5852 5348 5908 6076
rect 6188 6066 6244 6076
rect 6076 5906 6132 5918
rect 6076 5854 6078 5906
rect 6130 5854 6132 5906
rect 5852 5346 6020 5348
rect 5852 5294 5854 5346
rect 5906 5294 6020 5346
rect 5852 5292 6020 5294
rect 5852 5282 5908 5292
rect 5740 5012 5796 5022
rect 5740 5010 5908 5012
rect 5740 4958 5742 5010
rect 5794 4958 5908 5010
rect 5740 4956 5908 4958
rect 5740 4946 5796 4956
rect 5404 4834 5460 4844
rect 5852 4900 5908 4956
rect 5068 4398 5070 4450
rect 5122 4398 5124 4450
rect 5068 4386 5124 4398
rect 5740 4564 5796 4574
rect 5740 4450 5796 4508
rect 5740 4398 5742 4450
rect 5794 4398 5796 4450
rect 5740 4386 5796 4398
rect 5180 4114 5236 4126
rect 5180 4062 5182 4114
rect 5234 4062 5236 4114
rect 4956 3780 5012 3790
rect 4844 3778 5012 3780
rect 4844 3726 4958 3778
rect 5010 3726 5012 3778
rect 4844 3724 5012 3726
rect 4956 3714 5012 3724
rect 4396 3378 4452 3388
rect 4844 3444 4900 3454
rect 4844 3350 4900 3388
rect 5180 3444 5236 4062
rect 5852 4116 5908 4844
rect 5852 4022 5908 4060
rect 5964 4340 6020 5292
rect 6076 4900 6132 5854
rect 6524 5348 6580 6076
rect 6748 6020 6804 6030
rect 6860 6020 6916 6524
rect 6748 6018 6916 6020
rect 6748 5966 6750 6018
rect 6802 5966 6862 6018
rect 6914 5966 6916 6018
rect 6748 5964 6916 5966
rect 6748 5954 6804 5964
rect 6860 5954 6916 5964
rect 7084 6020 7140 6524
rect 7084 5572 7140 5964
rect 7196 6466 7252 6478
rect 7196 6414 7198 6466
rect 7250 6414 7252 6466
rect 7196 5684 7252 6414
rect 7420 6020 7476 6030
rect 7420 5926 7476 5964
rect 7532 5684 7588 6860
rect 8316 7250 8372 7262
rect 8316 7198 8318 7250
rect 8370 7198 8372 7250
rect 7756 6578 7812 6590
rect 7756 6526 7758 6578
rect 7810 6526 7812 6578
rect 7756 6020 7812 6526
rect 7756 5954 7812 5964
rect 7868 6466 7924 6478
rect 7868 6414 7870 6466
rect 7922 6414 7924 6466
rect 7868 5684 7924 6414
rect 8092 6020 8148 6030
rect 8316 6020 8372 7198
rect 8428 6580 8484 7420
rect 8764 7476 8820 7980
rect 8988 7698 9044 8316
rect 9884 8372 9940 9662
rect 9212 8260 9268 8270
rect 9212 8166 9268 8204
rect 9884 8258 9940 8316
rect 9884 8206 9886 8258
rect 9938 8206 9940 8258
rect 8988 7646 8990 7698
rect 9042 7646 9044 7698
rect 8988 7634 9044 7646
rect 9884 7700 9940 8206
rect 9996 9602 10052 9884
rect 10556 9828 10612 10558
rect 9996 9550 9998 9602
rect 10050 9550 10052 9602
rect 9996 8596 10052 9550
rect 10332 9826 10612 9828
rect 10332 9774 10558 9826
rect 10610 9774 10612 9826
rect 10332 9772 10612 9774
rect 10332 9156 10388 9772
rect 10556 9762 10612 9772
rect 10668 10388 10724 11228
rect 12124 11282 12292 11284
rect 12124 11230 12126 11282
rect 12178 11230 12238 11282
rect 12290 11230 12292 11282
rect 12124 11228 12292 11230
rect 12124 11218 12180 11228
rect 11852 11004 12116 11014
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 11852 10938 12116 10948
rect 11228 10610 11284 10622
rect 11228 10558 11230 10610
rect 11282 10558 11284 10610
rect 11228 10388 11284 10558
rect 12012 10610 12068 10622
rect 12012 10558 12014 10610
rect 12066 10558 12068 10610
rect 10668 10386 11284 10388
rect 10668 10334 10670 10386
rect 10722 10334 11284 10386
rect 10668 10332 11284 10334
rect 11340 10386 11396 10398
rect 11340 10334 11342 10386
rect 11394 10334 11396 10386
rect 10668 9604 10724 10332
rect 11340 10052 11396 10334
rect 12012 10388 12068 10558
rect 12236 10612 12292 11228
rect 12796 11282 12852 11294
rect 12796 11230 12798 11282
rect 12850 11230 12852 11282
rect 12796 11172 12852 11230
rect 13692 11282 13748 11294
rect 13692 11230 13694 11282
rect 13746 11230 13748 11282
rect 12908 11172 12964 11182
rect 12796 11170 12964 11172
rect 12796 11118 12910 11170
rect 12962 11118 12964 11170
rect 12796 11116 12964 11118
rect 12684 10612 12740 10622
rect 12796 10612 12852 11116
rect 12908 11106 12964 11116
rect 13692 11172 13748 11230
rect 13804 11172 13860 11182
rect 13692 11170 13860 11172
rect 13692 11118 13806 11170
rect 13858 11118 13860 11170
rect 13692 11116 13860 11118
rect 13356 10612 13412 10622
rect 13468 10612 13524 10622
rect 13692 10612 13748 11116
rect 13804 11106 13860 11116
rect 14028 10612 14084 10622
rect 14140 10612 14196 12126
rect 14812 12180 14868 12190
rect 14812 12086 14868 12124
rect 14252 11956 14308 11966
rect 14252 11862 14308 11900
rect 14924 11956 14980 11966
rect 14512 11788 14776 11798
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14512 11722 14776 11732
rect 14924 11396 14980 11900
rect 14924 11302 14980 11340
rect 14812 11282 14868 11294
rect 14812 11230 14814 11282
rect 14866 11230 14868 11282
rect 14700 10612 14756 10622
rect 14812 10612 14868 11230
rect 12236 10610 14868 10612
rect 12236 10558 12686 10610
rect 12738 10558 12798 10610
rect 12850 10558 13358 10610
rect 13410 10558 13470 10610
rect 13522 10558 14030 10610
rect 14082 10558 14142 10610
rect 14194 10558 14702 10610
rect 14754 10558 14814 10610
rect 14866 10558 14868 10610
rect 12236 10556 14868 10558
rect 12124 10388 12180 10398
rect 12236 10388 12292 10556
rect 12684 10546 12740 10556
rect 12796 10546 12852 10556
rect 13356 10546 13412 10556
rect 13468 10546 13524 10556
rect 14028 10546 14084 10556
rect 14140 10546 14196 10556
rect 14700 10546 14756 10556
rect 14812 10546 14868 10556
rect 12012 10386 12292 10388
rect 12012 10334 12126 10386
rect 12178 10334 12292 10386
rect 12012 10332 12292 10334
rect 11564 10052 11620 10062
rect 11396 10050 11620 10052
rect 11396 9998 11566 10050
rect 11618 9998 11620 10050
rect 11396 9996 11620 9998
rect 11340 9986 11396 9996
rect 11564 9986 11620 9996
rect 12012 10052 12068 10332
rect 12124 10322 12180 10332
rect 14512 10220 14776 10230
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14512 10154 14776 10164
rect 12012 9828 12068 9996
rect 12124 9828 12180 9838
rect 12236 9828 12292 9838
rect 14476 9828 14532 9838
rect 15036 9828 15092 12796
rect 15484 12850 15540 12862
rect 15484 12798 15486 12850
rect 15538 12798 15540 12850
rect 15484 12180 15540 12798
rect 16156 12850 16212 12862
rect 16156 12798 16158 12850
rect 16210 12798 16212 12850
rect 15484 11282 15540 12124
rect 15596 12738 15652 12750
rect 15596 12686 15598 12738
rect 15650 12686 15652 12738
rect 15596 11954 15652 12686
rect 15596 11902 15598 11954
rect 15650 11902 15652 11954
rect 15596 11396 15652 11902
rect 15596 11302 15652 11340
rect 16156 12180 16212 12798
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15372 10612 15428 10622
rect 15484 10612 15540 11230
rect 16156 11282 16212 12124
rect 16268 12738 16324 13020
rect 16828 12852 16884 13694
rect 16940 13524 16996 14366
rect 16940 13430 16996 13468
rect 17052 14308 17108 14588
rect 17612 14418 17668 14430
rect 17612 14366 17614 14418
rect 17666 14366 17668 14418
rect 17500 14308 17556 14318
rect 17052 14306 17556 14308
rect 17052 14254 17502 14306
rect 17554 14254 17556 14306
rect 17052 14252 17556 14254
rect 17052 13188 17108 14252
rect 17500 14242 17556 14252
rect 17172 14140 17436 14150
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17172 14074 17436 14084
rect 17052 13122 17108 13132
rect 17388 13524 17444 13534
rect 16828 12850 16996 12852
rect 16828 12798 16830 12850
rect 16882 12798 16996 12850
rect 16828 12796 16996 12798
rect 16828 12786 16884 12796
rect 16268 12686 16270 12738
rect 16322 12686 16324 12738
rect 16268 11954 16324 12686
rect 16940 12738 16996 12796
rect 16940 12686 16942 12738
rect 16994 12686 16996 12738
rect 16828 12180 16884 12190
rect 16828 12086 16884 12124
rect 16268 11902 16270 11954
rect 16322 11902 16324 11954
rect 16268 11396 16324 11902
rect 16940 11954 16996 12686
rect 17388 12740 17444 13468
rect 17612 13524 17668 14366
rect 17612 13458 17668 13468
rect 17724 13746 17780 13758
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13188 17780 13694
rect 18396 13746 18452 13758
rect 18396 13694 18398 13746
rect 18450 13694 18452 13746
rect 17724 13122 17780 13132
rect 17836 13522 17892 13534
rect 17836 13470 17838 13522
rect 17890 13470 17892 13522
rect 17500 12964 17556 12974
rect 17836 12964 17892 13470
rect 18396 13524 18452 13694
rect 18396 13458 18452 13468
rect 18508 13522 18564 13534
rect 18508 13470 18510 13522
rect 18562 13470 18564 13522
rect 18508 13300 18564 13470
rect 18508 13234 18564 13244
rect 18956 13524 19012 13534
rect 18284 13188 18340 13198
rect 18284 13094 18340 13132
rect 18844 13188 18900 13198
rect 17500 12962 17892 12964
rect 17500 12910 17502 12962
rect 17554 12910 17892 12962
rect 17500 12908 17892 12910
rect 17500 12898 17556 12908
rect 17612 12740 17668 12750
rect 17388 12738 17668 12740
rect 17388 12686 17614 12738
rect 17666 12686 17668 12738
rect 17388 12684 17668 12686
rect 17172 12572 17436 12582
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17172 12506 17436 12516
rect 16940 11902 16942 11954
rect 16994 11902 16996 11954
rect 16268 11302 16324 11340
rect 16828 11396 16884 11406
rect 16940 11396 16996 11902
rect 17612 11844 17668 12684
rect 17612 11778 17668 11788
rect 17724 12292 17780 12302
rect 17836 12292 17892 12908
rect 18844 12962 18900 13132
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 12898 18900 12910
rect 18956 13186 19012 13468
rect 19628 13524 19684 14700
rect 22492 14140 22756 14150
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22492 14074 22756 14084
rect 18956 13134 18958 13186
rect 19010 13134 19012 13186
rect 18172 12850 18228 12862
rect 18172 12798 18174 12850
rect 18226 12798 18228 12850
rect 18172 12292 18228 12798
rect 18396 12292 18452 12302
rect 17724 12290 18396 12292
rect 17724 12238 17726 12290
rect 17778 12238 17838 12290
rect 17890 12238 18396 12290
rect 17724 12236 18396 12238
rect 17612 11620 17668 11630
rect 17724 11620 17780 12236
rect 17836 12226 17892 12236
rect 17612 11618 17780 11620
rect 17612 11566 17614 11618
rect 17666 11566 17780 11618
rect 17612 11564 17780 11566
rect 16828 11394 16940 11396
rect 16828 11342 16830 11394
rect 16882 11342 16940 11394
rect 16828 11340 16940 11342
rect 16156 11230 16158 11282
rect 16210 11230 16212 11282
rect 16044 10612 16100 10622
rect 12012 9826 12404 9828
rect 12012 9774 12126 9826
rect 12178 9774 12238 9826
rect 12290 9774 12404 9826
rect 12012 9772 12404 9774
rect 12124 9762 12180 9772
rect 12236 9762 12292 9772
rect 11452 9716 11508 9726
rect 9996 8482 10052 8540
rect 9996 8430 9998 8482
rect 10050 8430 10052 8482
rect 9996 8260 10052 8430
rect 10108 9154 10388 9156
rect 10108 9102 10334 9154
rect 10386 9102 10388 9154
rect 10108 9100 10388 9102
rect 10108 8428 10164 9100
rect 10332 9090 10388 9100
rect 10556 9602 10724 9604
rect 10556 9550 10670 9602
rect 10722 9550 10724 9602
rect 10556 9548 10724 9550
rect 10444 8932 10500 8942
rect 10556 8932 10612 9548
rect 10668 9538 10724 9548
rect 11340 9714 11508 9716
rect 11340 9662 11454 9714
rect 11506 9662 11508 9714
rect 11340 9660 11508 9662
rect 11004 9044 11060 9054
rect 11004 9042 11172 9044
rect 11004 8990 11006 9042
rect 11058 8990 11172 9042
rect 11004 8988 11172 8990
rect 11004 8978 11060 8988
rect 10444 8930 10612 8932
rect 10444 8878 10446 8930
rect 10498 8878 10612 8930
rect 10444 8876 10612 8878
rect 10444 8866 10500 8876
rect 10556 8596 10612 8876
rect 11116 8820 11172 8988
rect 11340 8820 11396 9660
rect 11452 9650 11508 9660
rect 11852 9436 12116 9446
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 11852 9370 12116 9380
rect 12348 9156 12404 9772
rect 14476 9826 15092 9828
rect 14476 9774 14478 9826
rect 14530 9774 15038 9826
rect 15090 9774 15092 9826
rect 14476 9772 15092 9774
rect 12796 9716 12852 9726
rect 12908 9716 12964 9726
rect 12796 9714 12964 9716
rect 12796 9662 12798 9714
rect 12850 9662 12910 9714
rect 12962 9662 12964 9714
rect 12796 9660 12964 9662
rect 12796 9156 12852 9660
rect 12908 9650 12964 9660
rect 13692 9716 13748 9726
rect 13804 9716 13860 9726
rect 13692 9714 13860 9716
rect 13692 9662 13694 9714
rect 13746 9662 13806 9714
rect 13858 9662 13860 9714
rect 13692 9660 13860 9662
rect 13020 9156 13076 9166
rect 12348 9154 13076 9156
rect 12348 9102 12350 9154
rect 12402 9102 13022 9154
rect 13074 9102 13076 9154
rect 12348 9100 13076 9102
rect 12348 9090 12404 9100
rect 11116 8818 11396 8820
rect 11116 8766 11118 8818
rect 11170 8766 11396 8818
rect 11116 8764 11396 8766
rect 11676 9042 11732 9054
rect 11676 8990 11678 9042
rect 11730 8990 11732 9042
rect 11676 8820 11732 8990
rect 11788 8820 11844 8830
rect 11676 8818 11844 8820
rect 11676 8766 11790 8818
rect 11842 8766 11844 8818
rect 11676 8764 11844 8766
rect 11116 8754 11172 8764
rect 10556 8484 10612 8540
rect 10668 8484 10724 8494
rect 10556 8482 10836 8484
rect 10556 8430 10670 8482
rect 10722 8430 10836 8482
rect 10556 8428 10836 8430
rect 11340 8428 11396 8764
rect 11788 8428 11844 8764
rect 12460 8818 12516 8830
rect 12460 8766 12462 8818
rect 12514 8766 12516 8818
rect 10108 8372 10388 8428
rect 10668 8418 10724 8428
rect 10780 8372 11284 8428
rect 10388 8316 10612 8372
rect 10332 8306 10388 8316
rect 9996 8194 10052 8204
rect 10556 8258 10612 8316
rect 10556 8206 10558 8258
rect 10610 8206 10612 8258
rect 9996 7700 10052 7710
rect 9884 7698 10052 7700
rect 9884 7646 9998 7698
rect 10050 7646 10052 7698
rect 9884 7644 10052 7646
rect 9996 7634 10052 7644
rect 10556 7586 10612 8206
rect 10668 7700 10724 7710
rect 10780 7700 10836 8372
rect 10668 7698 10836 7700
rect 10668 7646 10670 7698
rect 10722 7646 10836 7698
rect 10668 7644 10836 7646
rect 11228 8370 11284 8372
rect 11228 8318 11230 8370
rect 11282 8318 11284 8370
rect 11228 7698 11284 8318
rect 11228 7646 11230 7698
rect 11282 7646 11284 7698
rect 10668 7634 10724 7644
rect 11228 7634 11284 7646
rect 11340 8372 12180 8428
rect 11340 8146 11396 8372
rect 12124 8260 12180 8372
rect 12236 8260 12292 8270
rect 12460 8260 12516 8766
rect 12124 8258 12460 8260
rect 12124 8206 12126 8258
rect 12178 8206 12238 8258
rect 12290 8206 12460 8258
rect 12124 8204 12460 8206
rect 12124 8194 12180 8204
rect 12236 8194 12292 8204
rect 11340 8094 11342 8146
rect 11394 8094 11396 8146
rect 12460 8128 12516 8204
rect 12796 8484 12852 9100
rect 13020 9090 13076 9100
rect 13692 9042 13748 9660
rect 13804 9650 13860 9660
rect 14364 9714 14420 9726
rect 14364 9662 14366 9714
rect 14418 9662 14420 9714
rect 13692 8990 13694 9042
rect 13746 8990 13748 9042
rect 12796 8146 12852 8428
rect 13132 8818 13188 8830
rect 13132 8766 13134 8818
rect 13186 8766 13188 8818
rect 13132 8428 13188 8766
rect 13692 8484 13748 8990
rect 14364 9044 14420 9662
rect 14476 9266 14532 9772
rect 14476 9214 14478 9266
rect 14530 9214 14532 9266
rect 14476 9202 14532 9214
rect 15036 9268 15092 9772
rect 15260 10610 15540 10612
rect 15260 10558 15374 10610
rect 15426 10558 15486 10610
rect 15538 10558 15540 10610
rect 15260 10556 15540 10558
rect 15148 9604 15204 9614
rect 15260 9604 15316 10556
rect 15372 10546 15428 10556
rect 15484 10546 15540 10556
rect 15708 10610 16100 10612
rect 15708 10558 16046 10610
rect 16098 10558 16100 10610
rect 15708 10556 16100 10558
rect 15148 9602 15316 9604
rect 15148 9550 15150 9602
rect 15202 9550 15316 9602
rect 15148 9548 15316 9550
rect 15148 9538 15204 9548
rect 15148 9268 15204 9278
rect 15036 9266 15204 9268
rect 15036 9214 15150 9266
rect 15202 9214 15204 9266
rect 15036 9212 15204 9214
rect 13132 8372 13412 8428
rect 12908 8260 12964 8270
rect 12908 8166 12964 8204
rect 13356 8260 13412 8372
rect 10556 7534 10558 7586
rect 10610 7534 10612 7586
rect 8876 7476 8932 7486
rect 8764 7474 8932 7476
rect 8764 7422 8878 7474
rect 8930 7422 8932 7474
rect 8764 7420 8932 7422
rect 8428 6486 8484 6524
rect 8540 6692 8596 6702
rect 8148 5964 8372 6020
rect 8092 5926 8148 5964
rect 8204 5684 8260 5694
rect 7196 5682 8260 5684
rect 7196 5630 7534 5682
rect 7586 5630 8206 5682
rect 8258 5630 8260 5682
rect 7196 5628 8260 5630
rect 7084 5516 7252 5572
rect 7196 5348 7252 5516
rect 6524 5346 7140 5348
rect 6524 5294 6526 5346
rect 6578 5294 7140 5346
rect 6524 5292 7140 5294
rect 6524 5282 6580 5292
rect 7084 5124 7140 5292
rect 7196 5346 7364 5348
rect 7196 5294 7198 5346
rect 7250 5294 7364 5346
rect 7196 5292 7364 5294
rect 7196 5282 7252 5292
rect 7308 5124 7364 5292
rect 7084 5122 7252 5124
rect 7084 5070 7086 5122
rect 7138 5070 7252 5122
rect 7084 5068 7252 5070
rect 7084 5058 7140 5068
rect 6076 4834 6132 4844
rect 6412 5010 6468 5022
rect 6412 4958 6414 5010
rect 6466 4958 6468 5010
rect 6300 4564 6356 4574
rect 6412 4564 6468 4958
rect 6532 4732 6796 4742
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6532 4666 6796 4676
rect 6412 4508 6580 4564
rect 6300 4340 6356 4508
rect 6412 4340 6468 4350
rect 5964 4284 6244 4340
rect 6300 4338 6468 4340
rect 6300 4286 6414 4338
rect 6466 4286 6468 4338
rect 6300 4284 6468 4286
rect 5964 3892 6020 4284
rect 5852 3836 6020 3892
rect 6076 4116 6132 4126
rect 5852 3554 5908 3836
rect 5852 3502 5854 3554
rect 5906 3502 5908 3554
rect 5852 3490 5908 3502
rect 5180 3378 5236 3388
rect 5740 3444 5796 3454
rect 5740 3350 5796 3388
rect 6076 800 6132 4060
rect 6188 3668 6244 4284
rect 6412 4274 6468 4284
rect 6524 4116 6580 4508
rect 7196 4562 7252 5068
rect 7196 4510 7198 4562
rect 7250 4510 7252 4562
rect 7196 4498 7252 4510
rect 6524 4022 6580 4060
rect 7084 4340 7140 4350
rect 7084 4116 7140 4284
rect 6412 3780 6468 3790
rect 6412 3778 6692 3780
rect 6412 3726 6414 3778
rect 6466 3726 6692 3778
rect 6412 3724 6692 3726
rect 6412 3714 6468 3724
rect 6188 3612 6356 3668
rect 6300 3556 6356 3612
rect 6524 3556 6580 3566
rect 6300 3554 6580 3556
rect 6300 3502 6526 3554
rect 6578 3502 6580 3554
rect 6300 3500 6580 3502
rect 6524 3490 6580 3500
rect 6636 3444 6692 3724
rect 7084 3778 7140 4060
rect 7084 3726 7086 3778
rect 7138 3726 7140 3778
rect 7084 3556 7140 3726
rect 7084 3490 7140 3500
rect 7196 3556 7252 3566
rect 7308 3556 7364 5068
rect 7532 4116 7588 5628
rect 8204 5618 8260 5628
rect 8540 5346 8596 6636
rect 8764 6692 8820 7420
rect 8876 7410 8932 7420
rect 9884 7474 9940 7486
rect 9884 7422 9886 7474
rect 9938 7422 9940 7474
rect 9192 7084 9456 7094
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9192 7018 9456 7028
rect 8764 6018 8820 6636
rect 8876 6916 8932 6926
rect 8876 6130 8932 6860
rect 9212 6692 9268 6702
rect 9212 6598 9268 6636
rect 9772 6692 9828 6702
rect 9884 6692 9940 7422
rect 9772 6690 9884 6692
rect 9772 6638 9774 6690
rect 9826 6638 9884 6690
rect 9772 6636 9884 6638
rect 8876 6078 8878 6130
rect 8930 6078 8932 6130
rect 8876 6066 8932 6078
rect 9100 6580 9156 6590
rect 8764 5966 8766 6018
rect 8818 5966 8820 6018
rect 8764 5954 8820 5966
rect 9100 5908 9156 6524
rect 9772 6132 9828 6636
rect 9884 6626 9940 6636
rect 9996 6916 10052 6926
rect 9884 6468 9940 6478
rect 9884 6374 9940 6412
rect 9884 6132 9940 6142
rect 9772 6130 9940 6132
rect 9772 6078 9886 6130
rect 9938 6078 9940 6130
rect 9772 6076 9940 6078
rect 9884 6066 9940 6076
rect 9100 5842 9156 5852
rect 9772 5908 9828 5918
rect 9772 5814 9828 5852
rect 9192 5516 9456 5526
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9192 5450 9456 5460
rect 8540 5294 8542 5346
rect 8594 5294 8596 5346
rect 7756 5124 7812 5134
rect 7868 5124 7924 5134
rect 7812 5122 7924 5124
rect 7812 5070 7870 5122
rect 7922 5070 7924 5122
rect 7812 5068 7924 5070
rect 7756 5030 7812 5068
rect 7868 5058 7924 5068
rect 8428 5124 8484 5134
rect 8540 5124 8596 5294
rect 9884 5348 9940 5358
rect 9996 5348 10052 6860
rect 10556 6916 10612 7534
rect 11340 7476 11396 8094
rect 12796 8094 12798 8146
rect 12850 8094 12852 8146
rect 11852 7868 12116 7878
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 11852 7802 12116 7812
rect 10444 6692 10500 6702
rect 10444 6132 10500 6636
rect 10556 6468 10612 6860
rect 11228 7474 11396 7476
rect 11228 7422 11342 7474
rect 11394 7422 11396 7474
rect 11228 7420 11396 7422
rect 11228 6916 11284 7420
rect 11340 7410 11396 7420
rect 11900 7474 11956 7486
rect 11900 7422 11902 7474
rect 11954 7422 11956 7474
rect 10556 6402 10612 6412
rect 11116 6692 11172 6702
rect 10556 6132 10612 6142
rect 10444 6130 10612 6132
rect 10444 6078 10558 6130
rect 10610 6078 10612 6130
rect 10444 6076 10612 6078
rect 9884 5346 10052 5348
rect 9884 5294 9886 5346
rect 9938 5294 10052 5346
rect 9884 5292 10052 5294
rect 10444 5908 10500 5918
rect 9884 5282 9940 5292
rect 8428 5122 8540 5124
rect 8428 5070 8430 5122
rect 8482 5070 8540 5122
rect 8428 5068 8540 5070
rect 8428 5058 8484 5068
rect 8540 4564 8596 5068
rect 9100 5124 9156 5134
rect 9212 5124 9268 5134
rect 9156 5122 9268 5124
rect 9156 5070 9214 5122
rect 9266 5070 9268 5122
rect 9156 5068 9268 5070
rect 9100 5030 9156 5068
rect 9212 5058 9268 5068
rect 9660 5124 9716 5134
rect 10444 5124 10500 5852
rect 8428 4562 8596 4564
rect 8428 4510 8542 4562
rect 8594 4510 8596 4562
rect 8428 4508 8596 4510
rect 8428 4450 8484 4508
rect 8428 4398 8430 4450
rect 8482 4398 8484 4450
rect 8428 4386 8484 4398
rect 7756 4340 7812 4350
rect 7756 4246 7812 4284
rect 7868 4116 7924 4126
rect 7532 4114 7924 4116
rect 7532 4062 7870 4114
rect 7922 4062 7924 4114
rect 7532 4060 7924 4062
rect 7868 3778 7924 4060
rect 7868 3726 7870 3778
rect 7922 3726 7924 3778
rect 7868 3714 7924 3726
rect 7196 3554 7364 3556
rect 7196 3502 7198 3554
rect 7250 3502 7364 3554
rect 7196 3500 7364 3502
rect 7756 3556 7812 3566
rect 7196 3490 7252 3500
rect 7756 3462 7812 3500
rect 8428 3556 8484 3566
rect 8428 3462 8484 3500
rect 8540 3554 8596 4508
rect 9660 4452 9716 5068
rect 9996 5122 10500 5124
rect 9996 5070 10446 5122
rect 10498 5070 10500 5122
rect 9996 5068 10500 5070
rect 9772 5012 9828 5022
rect 9772 5010 9940 5012
rect 9772 4958 9774 5010
rect 9826 4958 9940 5010
rect 9772 4956 9940 4958
rect 9772 4946 9828 4956
rect 9772 4452 9828 4462
rect 9660 4450 9828 4452
rect 9660 4398 9774 4450
rect 9826 4398 9828 4450
rect 9660 4396 9828 4398
rect 9192 3948 9456 3958
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9192 3882 9456 3892
rect 8540 3502 8542 3554
rect 8594 3502 8596 3554
rect 8540 3490 8596 3502
rect 9660 3556 9716 3566
rect 9660 3462 9716 3500
rect 9772 3554 9828 4396
rect 9772 3502 9774 3554
rect 9826 3502 9828 3554
rect 9772 3490 9828 3502
rect 9884 4114 9940 4956
rect 9884 4062 9886 4114
rect 9938 4062 9940 4114
rect 9884 3556 9940 4062
rect 9884 3490 9940 3500
rect 6636 3378 6692 3388
rect 6532 3164 6796 3174
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6532 3098 6796 3108
rect 9996 800 10052 5068
rect 10444 5058 10500 5068
rect 10556 5346 10612 6076
rect 11116 6018 11172 6636
rect 11228 6130 11284 6860
rect 11788 6692 11844 6702
rect 11900 6692 11956 7422
rect 12572 7474 12628 7486
rect 12572 7422 12574 7474
rect 12626 7422 12628 7474
rect 11228 6078 11230 6130
rect 11282 6078 11284 6130
rect 11228 6066 11284 6078
rect 11676 6690 11900 6692
rect 11676 6638 11790 6690
rect 11842 6638 11900 6690
rect 11676 6636 11900 6638
rect 11116 5966 11118 6018
rect 11170 5966 11172 6018
rect 11116 5954 11172 5966
rect 11676 6020 11732 6636
rect 11788 6626 11844 6636
rect 11900 6626 11956 6636
rect 12012 7250 12068 7262
rect 12012 7198 12014 7250
rect 12066 7198 12068 7250
rect 12012 6916 12068 7198
rect 11900 6468 11956 6478
rect 12012 6468 12068 6860
rect 12572 7252 12628 7422
rect 12796 7476 12852 8094
rect 13356 7698 13412 8204
rect 13692 8258 13748 8428
rect 13692 8206 13694 8258
rect 13746 8206 13748 8258
rect 13692 8194 13748 8206
rect 13804 8818 13860 8830
rect 13804 8766 13806 8818
rect 13858 8766 13860 8818
rect 13804 8260 13860 8766
rect 13356 7646 13358 7698
rect 13410 7646 13412 7698
rect 13356 7634 13412 7646
rect 13244 7476 13300 7486
rect 12796 7474 13300 7476
rect 12796 7422 13246 7474
rect 13298 7422 13300 7474
rect 12796 7420 13300 7422
rect 12684 7252 12740 7262
rect 12572 7250 12740 7252
rect 12572 7198 12686 7250
rect 12738 7198 12740 7250
rect 12572 7196 12740 7198
rect 12460 6692 12516 6702
rect 12460 6598 12516 6636
rect 12572 6468 12628 7196
rect 12684 7186 12740 7196
rect 11900 6466 12628 6468
rect 11900 6414 11902 6466
rect 11954 6414 12574 6466
rect 12626 6414 12628 6466
rect 11900 6412 12628 6414
rect 11900 6402 11956 6412
rect 11852 6300 12116 6310
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 11852 6234 12116 6244
rect 11900 6132 11956 6142
rect 12236 6132 12292 6412
rect 11900 6130 12292 6132
rect 11900 6078 11902 6130
rect 11954 6078 12292 6130
rect 11900 6076 12292 6078
rect 11900 6066 11956 6076
rect 11788 6020 11844 6030
rect 11676 6018 11844 6020
rect 11676 5966 11790 6018
rect 11842 5966 11844 6018
rect 11676 5964 11844 5966
rect 11788 5954 11844 5964
rect 12572 6018 12628 6412
rect 13244 6132 13300 7420
rect 13804 7364 13860 8204
rect 13916 8484 13972 8494
rect 13916 7588 13972 8428
rect 14364 8484 14420 8988
rect 15036 9044 15092 9054
rect 15036 8950 15092 8988
rect 15148 8820 15204 9212
rect 15260 9044 15316 9548
rect 15708 9826 15764 10556
rect 16044 10546 16100 10556
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9156 15764 9774
rect 16156 10386 16212 11230
rect 16716 10724 16772 10734
rect 16828 10724 16884 11340
rect 16940 11302 16996 11340
rect 17500 11396 17556 11406
rect 17612 11396 17668 11564
rect 17556 11340 17668 11396
rect 17500 11264 17556 11340
rect 17172 11004 17436 11014
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17172 10938 17436 10948
rect 16716 10722 16884 10724
rect 16716 10670 16718 10722
rect 16770 10670 16884 10722
rect 16716 10668 16884 10670
rect 17724 10722 17780 11564
rect 18172 11396 18228 12236
rect 18396 12198 18452 12236
rect 18956 12292 19012 13134
rect 19180 13188 19236 13198
rect 19180 12852 19236 13132
rect 19628 12964 19684 13468
rect 19832 13356 20096 13366
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 19832 13290 20096 13300
rect 19628 12908 19908 12964
rect 19516 12852 19572 12862
rect 19180 12850 19684 12852
rect 19180 12798 19518 12850
rect 19570 12798 19684 12850
rect 19180 12796 19684 12798
rect 19180 12402 19236 12796
rect 19516 12786 19572 12796
rect 19180 12350 19182 12402
rect 19234 12350 19236 12402
rect 19068 12292 19124 12302
rect 19012 12290 19124 12292
rect 19012 12238 19070 12290
rect 19122 12238 19124 12290
rect 19012 12236 19124 12238
rect 18508 11954 18564 11966
rect 18508 11902 18510 11954
rect 18562 11902 18564 11954
rect 18508 11732 18564 11902
rect 18172 11394 18452 11396
rect 18172 11342 18174 11394
rect 18226 11342 18452 11394
rect 18172 11340 18452 11342
rect 18172 11330 18228 11340
rect 17724 10670 17726 10722
rect 17778 10670 17780 10722
rect 16716 10658 16772 10668
rect 16156 10334 16158 10386
rect 16210 10334 16212 10386
rect 15260 8978 15316 8988
rect 15596 9154 15764 9156
rect 15596 9102 15710 9154
rect 15762 9102 15764 9154
rect 15596 9100 15764 9102
rect 15036 8764 15204 8820
rect 14512 8652 14776 8662
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14512 8586 14776 8596
rect 14364 8258 14420 8428
rect 14364 8206 14366 8258
rect 14418 8206 14420 8258
rect 14364 7700 14420 8206
rect 14476 8260 14532 8270
rect 14476 8166 14532 8204
rect 15036 8260 15092 8764
rect 15148 8484 15204 8522
rect 15148 8372 15316 8428
rect 15036 8166 15092 8204
rect 14700 7700 14756 7710
rect 14364 7698 14980 7700
rect 14364 7646 14702 7698
rect 14754 7646 14980 7698
rect 14364 7644 14980 7646
rect 14700 7634 14756 7644
rect 13916 7586 14196 7588
rect 13916 7534 13918 7586
rect 13970 7534 14196 7586
rect 13916 7532 14196 7534
rect 13916 7522 13972 7532
rect 14028 7364 14084 7374
rect 13804 7362 14084 7364
rect 13804 7310 14030 7362
rect 14082 7310 14084 7362
rect 13804 7308 14084 7310
rect 14028 6916 14084 7308
rect 14028 6850 14084 6860
rect 14140 6690 14196 7532
rect 14588 7476 14644 7486
rect 14364 7474 14644 7476
rect 14364 7422 14590 7474
rect 14642 7422 14644 7474
rect 14364 7420 14644 7422
rect 14252 6916 14308 6926
rect 14364 6916 14420 7420
rect 14588 7410 14644 7420
rect 14512 7084 14776 7094
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14512 7018 14776 7028
rect 14308 6860 14420 6916
rect 14588 6916 14644 6926
rect 14252 6822 14308 6860
rect 14140 6638 14142 6690
rect 14194 6638 14196 6690
rect 13356 6132 13412 6142
rect 13244 6130 13412 6132
rect 13244 6078 13358 6130
rect 13410 6078 13412 6130
rect 13244 6076 13412 6078
rect 13356 6066 13412 6076
rect 14028 6132 14084 6142
rect 14140 6132 14196 6638
rect 14028 6130 14196 6132
rect 14028 6078 14030 6130
rect 14082 6078 14196 6130
rect 14028 6076 14196 6078
rect 14028 6066 14084 6076
rect 12572 5966 12574 6018
rect 12626 5966 12628 6018
rect 10556 5294 10558 5346
rect 10610 5294 10612 5346
rect 10444 4452 10500 4462
rect 10556 4452 10612 5294
rect 11452 5124 11508 5134
rect 11564 5124 11620 5134
rect 11452 5122 11564 5124
rect 11452 5070 11454 5122
rect 11506 5070 11564 5122
rect 11452 5068 11564 5070
rect 11452 5058 11508 5068
rect 11564 5030 11620 5068
rect 12124 5124 12180 5134
rect 12124 5010 12180 5068
rect 12124 4958 12126 5010
rect 12178 4958 12180 5010
rect 12124 4900 12180 4958
rect 12572 5012 12628 5966
rect 13244 5906 13300 5918
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 12684 5682 12740 5694
rect 12684 5630 12686 5682
rect 12738 5630 12740 5682
rect 12684 5236 12740 5630
rect 13244 5236 13300 5854
rect 12684 5180 13300 5236
rect 13916 5906 13972 5918
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 12796 5012 12852 5022
rect 12572 5010 12852 5012
rect 12572 4958 12798 5010
rect 12850 4958 12852 5010
rect 12572 4956 12852 4958
rect 12236 4900 12292 4910
rect 12348 4900 12404 4910
rect 12124 4898 12348 4900
rect 12124 4846 12238 4898
rect 12290 4846 12348 4898
rect 12124 4844 12348 4846
rect 12236 4834 12292 4844
rect 11852 4732 12116 4742
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 11852 4666 12116 4676
rect 10444 4450 10612 4452
rect 10444 4398 10446 4450
rect 10498 4398 10612 4450
rect 10444 4396 10612 4398
rect 10444 4386 10500 4396
rect 11116 4340 11172 4350
rect 12348 4340 12404 4844
rect 12684 4340 12740 4956
rect 12796 4946 12852 4956
rect 12908 4900 12964 5180
rect 12908 4806 12964 4844
rect 13916 5012 13972 5854
rect 14140 5346 14196 6076
rect 14588 6692 14644 6860
rect 14924 6914 14980 7644
rect 15260 7586 15316 8372
rect 15596 8260 15652 9100
rect 15708 9090 15764 9100
rect 15820 9604 15876 9614
rect 16156 9604 16212 10334
rect 16828 10388 16884 10398
rect 15820 9602 16212 9604
rect 15820 9550 15822 9602
rect 15874 9550 16212 9602
rect 15820 9548 16212 9550
rect 16380 9714 16436 9726
rect 16380 9662 16382 9714
rect 16434 9662 16436 9714
rect 15820 8820 15876 9548
rect 16380 9044 16436 9662
rect 16828 9716 16884 10332
rect 17724 9828 17780 10670
rect 18284 11172 18340 11182
rect 17836 10388 17892 10398
rect 17836 10294 17892 10332
rect 18284 10388 18340 11116
rect 18284 10322 18340 10332
rect 18396 10722 18452 11340
rect 18508 11172 18564 11676
rect 18844 11396 18900 11406
rect 18956 11396 19012 12236
rect 19068 12226 19124 12236
rect 18844 11394 18956 11396
rect 18844 11342 18846 11394
rect 18898 11342 18956 11394
rect 18844 11340 18956 11342
rect 19012 11340 19124 11396
rect 18844 11330 18900 11340
rect 18956 11330 19012 11340
rect 18508 11106 18564 11116
rect 18956 11172 19012 11182
rect 18956 11078 19012 11116
rect 18396 10670 18398 10722
rect 18450 10670 18452 10722
rect 18396 10052 18452 10670
rect 19068 10722 19124 11340
rect 19068 10670 19070 10722
rect 19122 10670 19124 10722
rect 19068 10658 19124 10670
rect 19180 10834 19236 12350
rect 19628 12738 19684 12796
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19628 12292 19684 12686
rect 19852 12402 19908 12908
rect 22492 12572 22756 12582
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22492 12506 22756 12516
rect 19852 12350 19854 12402
rect 19906 12350 19908 12402
rect 19852 12338 19908 12350
rect 19740 12292 19796 12302
rect 19628 12236 19740 12292
rect 19628 11618 19684 12236
rect 19740 12160 19796 12236
rect 20412 12292 20468 12302
rect 20524 12292 20580 12302
rect 20468 12290 20580 12292
rect 20468 12238 20526 12290
rect 20578 12238 20580 12290
rect 20468 12236 20580 12238
rect 20412 12198 20468 12236
rect 20524 12226 20580 12236
rect 21084 12292 21140 12302
rect 19832 11788 20096 11798
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 19832 11722 20096 11732
rect 19628 11566 19630 11618
rect 19682 11566 19684 11618
rect 19516 11396 19572 11406
rect 19516 11302 19572 11340
rect 19180 10782 19182 10834
rect 19234 10782 19236 10834
rect 18508 10388 18564 10398
rect 18508 10294 18564 10332
rect 18508 10052 18564 10062
rect 18396 10050 18564 10052
rect 18396 9998 18510 10050
rect 18562 9998 18564 10050
rect 18396 9996 18564 9998
rect 18508 9986 18564 9996
rect 17836 9828 17892 9838
rect 17724 9826 17892 9828
rect 17724 9774 17838 9826
rect 17890 9774 17892 9826
rect 17724 9772 17892 9774
rect 17836 9762 17892 9772
rect 19068 9828 19124 9838
rect 19180 9828 19236 10782
rect 19068 9826 19236 9828
rect 19068 9774 19070 9826
rect 19122 9774 19236 9826
rect 19068 9772 19236 9774
rect 19628 10724 19684 11566
rect 19852 11396 19908 11406
rect 19852 10834 19908 11340
rect 19852 10782 19854 10834
rect 19906 10782 19908 10834
rect 19740 10724 19796 10734
rect 19628 10722 19796 10724
rect 19628 10670 19742 10722
rect 19794 10670 19796 10722
rect 19628 10668 19796 10670
rect 19628 9828 19684 10668
rect 19740 10658 19796 10668
rect 19852 10724 19908 10782
rect 19852 10658 19908 10668
rect 20188 11282 20244 11294
rect 20188 11230 20190 11282
rect 20242 11230 20244 11282
rect 20188 10724 20244 11230
rect 20300 11170 20356 11182
rect 20300 11118 20302 11170
rect 20354 11118 20356 11170
rect 20300 10724 20356 11118
rect 20412 10724 20468 10734
rect 20300 10722 20468 10724
rect 20300 10670 20414 10722
rect 20466 10670 20468 10722
rect 20300 10668 20468 10670
rect 20188 10658 20244 10668
rect 19832 10220 20096 10230
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 19832 10154 20096 10164
rect 19852 10052 19908 10062
rect 19740 9828 19796 9838
rect 19628 9826 19796 9828
rect 19628 9774 19742 9826
rect 19794 9774 19796 9826
rect 19628 9772 19796 9774
rect 17052 9716 17108 9726
rect 16828 9714 17108 9716
rect 16828 9662 17054 9714
rect 17106 9662 17108 9714
rect 16828 9660 17108 9662
rect 15596 8194 15652 8204
rect 15708 8818 15876 8820
rect 15708 8766 15822 8818
rect 15874 8766 15876 8818
rect 15708 8764 15876 8766
rect 15708 8484 15764 8764
rect 15820 8754 15876 8764
rect 16268 9042 16436 9044
rect 16268 8990 16382 9042
rect 16434 8990 16436 9042
rect 16268 8988 16436 8990
rect 15260 7534 15262 7586
rect 15314 7534 15316 7586
rect 15260 7522 15316 7534
rect 15708 8146 15764 8428
rect 15708 8094 15710 8146
rect 15762 8094 15764 8146
rect 15372 7252 15428 7262
rect 14924 6862 14926 6914
rect 14978 6862 14980 6914
rect 14812 6692 14868 6702
rect 14588 6690 14868 6692
rect 14588 6638 14814 6690
rect 14866 6638 14868 6690
rect 14588 6636 14868 6638
rect 14588 6132 14644 6636
rect 14812 6626 14868 6636
rect 14700 6132 14756 6142
rect 14588 6130 14756 6132
rect 14588 6078 14702 6130
rect 14754 6078 14756 6130
rect 14588 6076 14756 6078
rect 14588 6020 14644 6076
rect 14700 6066 14756 6076
rect 14140 5294 14142 5346
rect 14194 5294 14196 5346
rect 14140 5282 14196 5294
rect 14364 6018 14644 6020
rect 14364 5966 14590 6018
rect 14642 5966 14644 6018
rect 14364 5964 14644 5966
rect 14028 5012 14084 5022
rect 13916 5010 14084 5012
rect 13916 4958 14030 5010
rect 14082 4958 14084 5010
rect 13916 4956 14084 4958
rect 13020 4340 13076 4350
rect 13692 4340 13748 4350
rect 11116 4338 11284 4340
rect 11116 4286 11118 4338
rect 11170 4286 11284 4338
rect 11116 4284 11284 4286
rect 11116 4274 11172 4284
rect 10556 4116 10612 4126
rect 10444 4114 10612 4116
rect 10444 4062 10558 4114
rect 10610 4062 10612 4114
rect 10444 4060 10612 4062
rect 10332 3556 10388 3566
rect 10444 3556 10500 4060
rect 10556 4050 10612 4060
rect 11228 4114 11284 4284
rect 12348 4338 12516 4340
rect 12348 4286 12350 4338
rect 12402 4286 12516 4338
rect 12348 4284 12516 4286
rect 12684 4338 13748 4340
rect 12684 4286 13022 4338
rect 13074 4286 13694 4338
rect 13746 4286 13748 4338
rect 12684 4284 13748 4286
rect 12348 4274 12404 4284
rect 11228 4062 11230 4114
rect 11282 4062 11284 4114
rect 10388 3554 10500 3556
rect 10388 3502 10446 3554
rect 10498 3502 10500 3554
rect 10388 3500 10500 3502
rect 10332 3462 10388 3500
rect 10444 3490 10500 3500
rect 11116 3556 11172 3566
rect 11228 3556 11284 4062
rect 12460 4116 12516 4284
rect 13020 4274 13076 4284
rect 12460 4022 12516 4060
rect 13132 4116 13188 4126
rect 13132 4022 13188 4060
rect 11172 3500 11284 3556
rect 11676 3556 11732 3566
rect 11116 3462 11172 3500
rect 11676 3462 11732 3500
rect 11004 3444 11060 3454
rect 11004 3350 11060 3388
rect 11788 3444 11844 3454
rect 11788 3350 11844 3388
rect 11852 3164 12116 3174
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 11852 3098 12116 3108
rect 13692 2996 13748 4284
rect 13804 4116 13860 4126
rect 13916 4116 13972 4956
rect 14028 4946 14084 4956
rect 13860 4060 13972 4116
rect 13804 3984 13860 4060
rect 13916 3444 13972 4060
rect 14364 4450 14420 5964
rect 14588 5954 14644 5964
rect 14512 5516 14776 5526
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14512 5450 14776 5460
rect 14812 5348 14868 5358
rect 14924 5348 14980 6862
rect 15260 7250 15428 7252
rect 15260 7198 15374 7250
rect 15426 7198 15428 7250
rect 15260 7196 15428 7198
rect 15260 6916 15316 7196
rect 15372 7186 15428 7196
rect 15260 6692 15316 6860
rect 15596 6916 15652 6926
rect 15708 6916 15764 8094
rect 15820 8260 15876 8270
rect 15820 7588 15876 8204
rect 16268 8260 16324 8988
rect 16380 8978 16436 8988
rect 16492 9604 16548 9614
rect 16492 8820 16548 9548
rect 16268 8194 16324 8204
rect 16380 8818 16548 8820
rect 16380 8766 16494 8818
rect 16546 8766 16548 8818
rect 16380 8764 16548 8766
rect 16380 8484 16436 8764
rect 16492 8754 16548 8764
rect 16380 8146 16436 8428
rect 16492 8260 16548 8270
rect 16492 8166 16548 8204
rect 17052 8260 17108 9660
rect 18396 9714 18452 9726
rect 18396 9662 18398 9714
rect 18450 9662 18452 9714
rect 17164 9604 17220 9642
rect 17164 9538 17220 9548
rect 17724 9602 17780 9614
rect 17724 9550 17726 9602
rect 17778 9550 17780 9602
rect 17172 9436 17436 9446
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17172 9370 17436 9380
rect 17724 9154 17780 9550
rect 17724 9102 17726 9154
rect 17778 9102 17780 9154
rect 17164 8484 17220 8522
rect 17724 8428 17780 9102
rect 18396 9042 18452 9662
rect 18396 8990 18398 9042
rect 18450 8990 18452 9042
rect 17164 8418 17220 8428
rect 17052 8166 17108 8204
rect 17612 8372 17780 8428
rect 17836 8818 17892 8830
rect 17836 8766 17838 8818
rect 17890 8766 17892 8818
rect 17836 8484 17892 8766
rect 17836 8418 17892 8428
rect 18396 8372 18452 8990
rect 19068 9154 19124 9772
rect 19068 9102 19070 9154
rect 19122 9102 19124 9154
rect 18508 8818 18564 8830
rect 18508 8766 18510 8818
rect 18562 8766 18564 8818
rect 18508 8484 18564 8766
rect 18508 8418 18564 8428
rect 18956 8820 19012 8830
rect 18956 8484 19012 8764
rect 19068 8484 19124 9102
rect 19180 9604 19236 9614
rect 19180 8820 19236 9548
rect 19740 9268 19796 9772
rect 19852 9604 19908 9996
rect 19852 9510 19908 9548
rect 20412 9826 20468 10668
rect 21084 10724 21140 12236
rect 21084 10592 21140 10668
rect 21756 11172 21812 11182
rect 21756 10722 21812 11116
rect 22492 11004 22756 11014
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22492 10938 22756 10948
rect 21756 10670 21758 10722
rect 21810 10670 21812 10722
rect 21756 10658 21812 10670
rect 21868 10724 21924 10734
rect 20524 10388 20580 10398
rect 21196 10388 21252 10398
rect 20524 10386 21252 10388
rect 20524 10334 20526 10386
rect 20578 10334 21198 10386
rect 21250 10334 21252 10386
rect 20524 10332 21252 10334
rect 20524 10052 20580 10332
rect 21196 10322 21252 10332
rect 21868 10276 21924 10668
rect 20524 9920 20580 9996
rect 21756 10220 21924 10276
rect 21756 10050 21812 10220
rect 21756 9998 21758 10050
rect 21810 9998 21812 10050
rect 20412 9774 20414 9826
rect 20466 9774 20468 9826
rect 19852 9268 19908 9278
rect 20412 9268 20468 9774
rect 21644 9828 21700 9838
rect 21756 9828 21812 9998
rect 21644 9826 21812 9828
rect 21644 9774 21646 9826
rect 21698 9774 21812 9826
rect 21644 9772 21812 9774
rect 21644 9762 21700 9772
rect 20524 9268 20580 9278
rect 19740 9266 20580 9268
rect 19740 9214 19854 9266
rect 19906 9214 20526 9266
rect 20578 9214 20580 9266
rect 19740 9212 20580 9214
rect 19852 9202 19908 9212
rect 20412 9154 20468 9212
rect 20524 9202 20580 9212
rect 20412 9102 20414 9154
rect 20466 9102 20468 9154
rect 20412 9090 20468 9102
rect 19740 9044 19796 9054
rect 19180 8726 19236 8764
rect 19628 9042 19796 9044
rect 19628 8990 19742 9042
rect 19794 8990 19796 9042
rect 19628 8988 19796 8990
rect 19180 8484 19236 8494
rect 19068 8482 19236 8484
rect 19068 8430 19182 8482
rect 19234 8430 19236 8482
rect 19068 8428 19236 8430
rect 17612 8260 17668 8372
rect 17612 8194 17668 8204
rect 18396 8258 18452 8316
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 16380 8094 16382 8146
rect 16434 8094 16436 8146
rect 16380 7700 16436 8094
rect 17724 8148 17780 8158
rect 17724 8146 17892 8148
rect 17724 8094 17726 8146
rect 17778 8094 17892 8146
rect 17724 8092 17892 8094
rect 17724 8082 17780 8092
rect 17172 7868 17436 7878
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17172 7802 17436 7812
rect 16716 7700 16772 7710
rect 17836 7700 17892 8092
rect 16380 7698 16772 7700
rect 16380 7646 16718 7698
rect 16770 7646 16772 7698
rect 16380 7644 16772 7646
rect 16716 7634 16772 7644
rect 17612 7644 17836 7700
rect 15932 7588 15988 7598
rect 15820 7586 15988 7588
rect 15820 7534 15934 7586
rect 15986 7534 15988 7586
rect 15820 7532 15988 7534
rect 15932 7522 15988 7532
rect 16604 7476 16660 7486
rect 16604 7382 16660 7420
rect 17612 7476 17668 7644
rect 17836 7606 17892 7644
rect 18396 7700 18452 8206
rect 18508 7700 18564 7710
rect 18452 7698 18564 7700
rect 18452 7646 18510 7698
rect 18562 7646 18564 7698
rect 18452 7644 18564 7646
rect 18396 7634 18452 7644
rect 18508 7634 18564 7644
rect 16044 7250 16100 7262
rect 16044 7198 16046 7250
rect 16098 7198 16100 7250
rect 16044 6916 16100 7198
rect 15596 6914 16100 6916
rect 15596 6862 15598 6914
rect 15650 6862 16100 6914
rect 15596 6860 16100 6862
rect 17612 6914 17668 7420
rect 17612 6862 17614 6914
rect 17666 6862 17668 6914
rect 15596 6850 15652 6860
rect 17612 6850 17668 6862
rect 17724 7474 17780 7486
rect 17724 7422 17726 7474
rect 17778 7422 17780 7474
rect 17724 7364 17780 7422
rect 15484 6692 15540 6702
rect 15260 6690 15540 6692
rect 15260 6638 15486 6690
rect 15538 6638 15540 6690
rect 15260 6636 15540 6638
rect 15260 6132 15316 6636
rect 15484 6626 15540 6636
rect 16156 6580 16212 6590
rect 16268 6580 16324 6590
rect 16828 6580 16884 6590
rect 16940 6580 16996 6590
rect 16044 6578 16940 6580
rect 16044 6526 16158 6578
rect 16210 6526 16270 6578
rect 16322 6526 16830 6578
rect 16882 6526 16940 6578
rect 16044 6524 16940 6526
rect 15372 6132 15428 6142
rect 16044 6132 16100 6524
rect 16156 6514 16212 6524
rect 16268 6514 16324 6524
rect 15260 6130 16100 6132
rect 15260 6078 15374 6130
rect 15426 6078 16046 6130
rect 16098 6078 16100 6130
rect 15260 6076 16100 6078
rect 15260 6018 15316 6076
rect 15372 6066 15428 6076
rect 15260 5966 15262 6018
rect 15314 5966 15316 6018
rect 15260 5954 15316 5966
rect 14812 5346 15204 5348
rect 14812 5294 14814 5346
rect 14866 5294 15204 5346
rect 14812 5292 15204 5294
rect 14812 5282 14868 5292
rect 14364 4398 14366 4450
rect 14418 4398 14420 4450
rect 14364 3780 14420 4398
rect 14700 5012 14756 5022
rect 14476 4340 14532 4350
rect 14476 4246 14532 4284
rect 14700 4340 14756 4956
rect 15148 4564 15204 5292
rect 15484 5346 15540 6076
rect 15932 6018 15988 6076
rect 16044 6066 16100 6076
rect 16604 6132 16660 6524
rect 16828 6514 16884 6524
rect 16940 6448 16996 6524
rect 17500 6580 17556 6590
rect 17724 6580 17780 7308
rect 18396 7474 18452 7486
rect 18396 7422 18398 7474
rect 18450 7422 18452 7474
rect 18396 7364 18452 7422
rect 18956 7476 19012 8428
rect 19180 8372 19236 8428
rect 19180 8306 19236 8316
rect 19068 8260 19124 8270
rect 19068 8166 19124 8204
rect 19628 8260 19684 8988
rect 19740 8978 19796 8988
rect 19832 8652 20096 8662
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 19832 8586 20096 8596
rect 21756 8428 21812 9772
rect 22492 9436 22756 9446
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22492 9370 22756 9380
rect 21756 8372 22036 8428
rect 19740 8260 19796 8270
rect 19852 8260 19908 8270
rect 19684 8258 19908 8260
rect 19684 8206 19742 8258
rect 19794 8206 19854 8258
rect 19906 8206 19908 8258
rect 19684 8204 19908 8206
rect 19628 8194 19684 8204
rect 19740 8194 19796 8204
rect 19852 8194 19908 8204
rect 20524 8146 20580 8158
rect 20524 8094 20526 8146
rect 20578 8094 20580 8146
rect 20412 8036 20468 8046
rect 20524 8036 20580 8094
rect 20412 8034 20580 8036
rect 20412 7982 20414 8034
rect 20466 7982 20580 8034
rect 20412 7980 20580 7982
rect 20412 7970 20468 7980
rect 19068 7476 19124 7486
rect 19740 7476 19796 7486
rect 20412 7476 20468 7486
rect 18956 7474 19124 7476
rect 18956 7422 19070 7474
rect 19122 7422 19124 7474
rect 18956 7420 19124 7422
rect 18396 7298 18452 7308
rect 18956 6692 19012 6702
rect 18956 6598 19012 6636
rect 17556 6524 17780 6580
rect 18172 6578 18228 6590
rect 18172 6526 18174 6578
rect 18226 6526 18228 6578
rect 17500 6486 17556 6524
rect 17172 6300 17436 6310
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17172 6234 17436 6244
rect 16716 6132 16772 6142
rect 16604 6130 16772 6132
rect 16604 6078 16718 6130
rect 16770 6078 16772 6130
rect 16604 6076 16772 6078
rect 15932 5966 15934 6018
rect 15986 5966 15988 6018
rect 15932 5954 15988 5966
rect 16604 6018 16660 6076
rect 16716 6066 16772 6076
rect 16604 5966 16606 6018
rect 16658 5966 16660 6018
rect 16604 5954 16660 5966
rect 15484 5294 15486 5346
rect 15538 5294 15540 5346
rect 15372 5124 15428 5134
rect 15484 5124 15540 5294
rect 15372 5122 15540 5124
rect 15372 5070 15374 5122
rect 15426 5070 15540 5122
rect 15372 5068 15540 5070
rect 16156 5124 16212 5134
rect 15372 5058 15428 5068
rect 16044 5012 16100 5022
rect 16044 4918 16100 4956
rect 16156 4898 16212 5068
rect 16828 5124 16884 5134
rect 16828 5030 16884 5068
rect 17388 5124 17444 5134
rect 17388 5030 17444 5068
rect 17612 5124 17668 6524
rect 18172 6132 18228 6526
rect 18844 6578 18900 6590
rect 18844 6526 18846 6578
rect 18898 6526 18900 6578
rect 18284 6468 18340 6478
rect 18844 6468 18900 6526
rect 18284 6466 18900 6468
rect 18284 6414 18286 6466
rect 18338 6414 18900 6466
rect 18284 6412 18900 6414
rect 18284 6402 18340 6412
rect 16716 5012 16772 5022
rect 16716 4918 16772 4956
rect 16156 4846 16158 4898
rect 16210 4846 16212 4898
rect 15820 4564 15876 4574
rect 16156 4564 16212 4846
rect 17500 4898 17556 4910
rect 17500 4846 17502 4898
rect 17554 4846 17556 4898
rect 17172 4732 17436 4742
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17172 4666 17436 4676
rect 15148 4562 16436 4564
rect 15148 4510 15150 4562
rect 15202 4510 15822 4562
rect 15874 4510 16436 4562
rect 15148 4508 16436 4510
rect 15148 4498 15204 4508
rect 15820 4498 15876 4508
rect 16380 4450 16436 4508
rect 16380 4398 16382 4450
rect 16434 4398 16436 4450
rect 16380 4386 16436 4398
rect 16492 4452 16548 4462
rect 16492 4358 16548 4396
rect 17500 4452 17556 4846
rect 17612 4788 17668 5068
rect 17724 6076 18228 6132
rect 17724 5906 17780 6076
rect 17724 5854 17726 5906
rect 17778 5854 17780 5906
rect 17724 5012 17780 5854
rect 17836 5908 17892 5918
rect 17836 5682 17892 5852
rect 18396 5908 18452 6412
rect 18844 6020 18900 6412
rect 19068 6020 19124 7420
rect 19516 7474 20468 7476
rect 19516 7422 19742 7474
rect 19794 7422 20414 7474
rect 20466 7422 20468 7474
rect 19516 7420 20468 7422
rect 19180 7250 19236 7262
rect 19180 7198 19182 7250
rect 19234 7198 19236 7250
rect 19180 6692 19236 7198
rect 19180 6626 19236 6636
rect 19516 6578 19572 7420
rect 19740 7410 19796 7420
rect 20412 7410 20468 7420
rect 19852 7252 19908 7262
rect 19516 6526 19518 6578
rect 19570 6526 19572 6578
rect 19516 6020 19572 6526
rect 18844 6018 19572 6020
rect 18844 5966 19070 6018
rect 19122 5966 19572 6018
rect 18844 5964 19572 5966
rect 19628 7250 19908 7252
rect 19628 7198 19854 7250
rect 19906 7198 19908 7250
rect 19628 7196 19908 7198
rect 19628 6914 19684 7196
rect 19852 7186 19908 7196
rect 20524 7250 20580 7980
rect 20524 7198 20526 7250
rect 20578 7198 20580 7250
rect 19832 7084 20096 7094
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 19832 7018 20096 7028
rect 19628 6862 19630 6914
rect 19682 6862 19684 6914
rect 19628 6692 19684 6862
rect 19628 6020 19684 6636
rect 20300 6578 20356 6590
rect 20300 6526 20302 6578
rect 20354 6526 20356 6578
rect 20188 6466 20244 6478
rect 20188 6414 20190 6466
rect 20242 6414 20244 6466
rect 19740 6020 19796 6030
rect 19628 6018 19796 6020
rect 19628 5966 19742 6018
rect 19794 5966 19796 6018
rect 19628 5964 19796 5966
rect 19068 5954 19124 5964
rect 19628 5908 19684 5964
rect 19740 5954 19796 5964
rect 18396 5814 18452 5852
rect 19180 5852 19684 5908
rect 17836 5630 17838 5682
rect 17890 5630 17892 5682
rect 17836 5124 17892 5630
rect 18172 5796 18228 5806
rect 18172 5348 18228 5740
rect 18508 5796 18564 5806
rect 18508 5702 18564 5740
rect 18732 5796 18788 5806
rect 18172 5346 18452 5348
rect 18172 5294 18174 5346
rect 18226 5294 18452 5346
rect 18172 5292 18452 5294
rect 18172 5282 18228 5292
rect 18060 5124 18116 5134
rect 17836 5122 18116 5124
rect 17836 5070 18062 5122
rect 18114 5070 18116 5122
rect 17836 5068 18116 5070
rect 18060 5058 18116 5068
rect 17724 4946 17780 4956
rect 17612 4732 17892 4788
rect 17836 4562 17892 4732
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17724 4452 17780 4462
rect 17500 4396 17724 4452
rect 14700 4274 14756 4284
rect 15036 4340 15092 4350
rect 15036 4246 15092 4284
rect 15708 4340 15764 4350
rect 14512 3948 14776 3958
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14512 3882 14776 3892
rect 14364 3724 14644 3780
rect 14588 3668 14644 3724
rect 14588 3612 15652 3668
rect 14588 3554 14644 3612
rect 14588 3502 14590 3554
rect 14642 3502 14644 3554
rect 14588 3490 14644 3502
rect 15260 3554 15316 3612
rect 15260 3502 15262 3554
rect 15314 3502 15316 3554
rect 15260 3490 15316 3502
rect 15596 3554 15652 3612
rect 15596 3502 15598 3554
rect 15650 3502 15652 3554
rect 15596 3490 15652 3502
rect 14028 3444 14084 3454
rect 13916 3442 14028 3444
rect 13916 3390 13918 3442
rect 13970 3390 14028 3442
rect 13916 3388 14028 3390
rect 13916 3378 13972 3388
rect 14028 3350 14084 3388
rect 14700 3444 14756 3454
rect 14700 3350 14756 3388
rect 15372 3444 15428 3454
rect 15372 3350 15428 3388
rect 15708 3444 15764 4284
rect 15932 3612 16660 3668
rect 15820 3556 15876 3566
rect 15932 3556 15988 3612
rect 15820 3554 15988 3556
rect 15820 3502 15822 3554
rect 15874 3502 15988 3554
rect 15820 3500 15988 3502
rect 15820 3490 15876 3500
rect 15708 3378 15764 3388
rect 15932 3442 15988 3500
rect 16604 3554 16660 3612
rect 16604 3502 16606 3554
rect 16658 3502 16660 3554
rect 16604 3490 16660 3502
rect 17500 3554 17556 4396
rect 17724 4358 17780 4396
rect 17836 4228 17892 4510
rect 17612 4172 17892 4228
rect 18172 4452 18228 4462
rect 17612 3778 17668 4172
rect 17612 3726 17614 3778
rect 17666 3726 17668 3778
rect 17612 3714 17668 3726
rect 17500 3502 17502 3554
rect 17554 3502 17556 3554
rect 17500 3490 17556 3502
rect 18172 3554 18228 4396
rect 18396 4452 18452 5292
rect 18508 5124 18564 5134
rect 18508 4562 18564 5068
rect 18732 5122 18788 5740
rect 19180 5796 19236 5852
rect 19180 5664 19236 5740
rect 18732 5070 18734 5122
rect 18786 5070 18788 5122
rect 18732 5058 18788 5070
rect 18844 5124 18900 5134
rect 18844 5030 18900 5068
rect 19068 5124 19124 5134
rect 18508 4510 18510 4562
rect 18562 4510 18564 4562
rect 18508 4498 18564 4510
rect 19068 4452 19124 5068
rect 19404 5124 19460 5852
rect 19852 5684 19908 5760
rect 19628 5628 19852 5684
rect 19516 5236 19572 5246
rect 19628 5236 19684 5628
rect 19852 5618 19908 5628
rect 19832 5516 20096 5526
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 19832 5450 20096 5460
rect 19572 5180 19684 5236
rect 20188 5346 20244 6414
rect 20300 5684 20356 6526
rect 20300 5618 20356 5628
rect 20412 5908 20468 5918
rect 20524 5908 20580 7198
rect 20412 5906 20580 5908
rect 20412 5854 20414 5906
rect 20466 5854 20580 5906
rect 20412 5852 20580 5854
rect 21084 7474 21140 7486
rect 21084 7422 21086 7474
rect 21138 7422 21140 7474
rect 21084 5906 21140 7422
rect 21084 5854 21086 5906
rect 21138 5854 21140 5906
rect 20188 5294 20190 5346
rect 20242 5294 20244 5346
rect 19516 5142 19572 5180
rect 19404 4992 19460 5068
rect 19852 5124 19908 5134
rect 19852 4564 19908 5068
rect 18396 4320 18452 4396
rect 18844 4450 19124 4452
rect 18844 4398 19070 4450
rect 19122 4398 19124 4450
rect 18844 4396 19124 4398
rect 18172 3502 18174 3554
rect 18226 3502 18228 3554
rect 18172 3490 18228 3502
rect 18844 3554 18900 4396
rect 19068 4386 19124 4396
rect 19628 4562 19908 4564
rect 19628 4510 19854 4562
rect 19906 4510 19908 4562
rect 19628 4508 19908 4510
rect 20076 5124 20132 5134
rect 20076 4564 20132 5068
rect 20188 5012 20244 5294
rect 20412 5348 20468 5852
rect 20524 5684 20580 5694
rect 20524 5590 20580 5628
rect 20412 5292 20580 5348
rect 20188 4946 20244 4956
rect 20412 5012 20468 5022
rect 20076 4508 20356 4564
rect 18844 3502 18846 3554
rect 18898 3502 18900 3554
rect 18844 3490 18900 3502
rect 19180 4340 19236 4350
rect 19180 4114 19236 4284
rect 19180 4062 19182 4114
rect 19234 4062 19236 4114
rect 15932 3390 15934 3442
rect 15986 3390 15988 3442
rect 15932 3378 15988 3390
rect 16044 3444 16100 3454
rect 16044 3350 16100 3388
rect 16716 3444 16772 3454
rect 16716 3350 16772 3388
rect 17836 3444 17892 3454
rect 17172 3164 17436 3174
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17172 3098 17436 3108
rect 13692 2940 13972 2996
rect 13916 800 13972 2940
rect 17836 800 17892 3388
rect 18284 3444 18340 3454
rect 18284 3350 18340 3388
rect 18956 3444 19012 3454
rect 18956 3350 19012 3388
rect 19180 3444 19236 4062
rect 19628 3778 19684 4508
rect 19852 4498 19908 4508
rect 19740 4340 19796 4350
rect 19740 4246 19796 4284
rect 20300 4116 20356 4508
rect 20412 4450 20468 4956
rect 20412 4398 20414 4450
rect 20466 4398 20468 4450
rect 20412 4340 20468 4398
rect 20412 4274 20468 4284
rect 20524 4564 20580 5292
rect 20748 5012 20804 5022
rect 20748 4918 20804 4956
rect 20860 4898 20916 4910
rect 20860 4846 20862 4898
rect 20914 4846 20916 4898
rect 20860 4564 20916 4846
rect 20524 4562 20916 4564
rect 20524 4510 20526 4562
rect 20578 4510 20916 4562
rect 20524 4508 20916 4510
rect 20524 4116 20580 4508
rect 20860 4452 20916 4508
rect 21084 4452 21140 5854
rect 21196 7250 21252 7262
rect 21196 7198 21198 7250
rect 21250 7198 21252 7250
rect 21196 5684 21252 7198
rect 21644 6692 21700 6702
rect 21644 6690 21924 6692
rect 21644 6638 21646 6690
rect 21698 6638 21924 6690
rect 21644 6636 21924 6638
rect 21644 6626 21700 6636
rect 21756 6466 21812 6478
rect 21756 6414 21758 6466
rect 21810 6414 21812 6466
rect 21756 6244 21812 6414
rect 21196 5590 21252 5628
rect 21644 6188 21812 6244
rect 21644 5684 21700 6188
rect 21868 5906 21924 6636
rect 21868 5854 21870 5906
rect 21922 5854 21924 5906
rect 21644 5618 21700 5628
rect 21756 5682 21812 5694
rect 21756 5630 21758 5682
rect 21810 5630 21812 5682
rect 21756 5124 21812 5630
rect 21644 5068 21812 5124
rect 21644 5012 21700 5068
rect 21644 4918 21700 4956
rect 21756 4900 21812 4910
rect 21868 4900 21924 5854
rect 21980 5012 22036 8372
rect 22492 7868 22756 7878
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22492 7802 22756 7812
rect 22492 6300 22756 6310
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22492 6234 22756 6244
rect 21980 4946 22036 4956
rect 21756 4898 21924 4900
rect 21756 4846 21758 4898
rect 21810 4846 21924 4898
rect 21756 4844 21924 4846
rect 21196 4564 21252 4574
rect 21756 4564 21812 4844
rect 22492 4732 22756 4742
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22492 4666 22756 4676
rect 21196 4562 21812 4564
rect 21196 4510 21198 4562
rect 21250 4510 21812 4562
rect 21196 4508 21812 4510
rect 21196 4452 21252 4508
rect 20860 4450 21252 4452
rect 20860 4398 21086 4450
rect 21138 4398 21252 4450
rect 20860 4396 21252 4398
rect 21084 4386 21140 4396
rect 20300 4060 20580 4116
rect 21756 4340 21812 4508
rect 21868 4340 21924 4350
rect 21756 4338 21924 4340
rect 21756 4286 21870 4338
rect 21922 4286 21924 4338
rect 21756 4284 21924 4286
rect 21756 4114 21812 4284
rect 21868 4274 21924 4284
rect 21756 4062 21758 4114
rect 21810 4062 21812 4114
rect 19832 3948 20096 3958
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 19832 3882 20096 3892
rect 19628 3726 19630 3778
rect 19682 3726 19684 3778
rect 19628 3714 19684 3726
rect 20300 3778 20356 4060
rect 20300 3726 20302 3778
rect 20354 3726 20356 3778
rect 20188 3556 20244 3566
rect 20300 3556 20356 3726
rect 20188 3554 20356 3556
rect 20188 3502 20190 3554
rect 20242 3502 20356 3554
rect 20188 3500 20356 3502
rect 20188 3490 20244 3500
rect 19180 3378 19236 3388
rect 19516 3444 19572 3454
rect 19516 3350 19572 3388
rect 21756 800 21812 4062
rect 22492 3164 22756 3174
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22492 3098 22756 3108
rect 2128 0 2240 800
rect 6048 0 6160 800
rect 9968 0 10080 800
rect 13888 0 14000 800
rect 17808 0 17920 800
rect 21728 0 21840 800
<< via2 >>
rect 3872 16490 3928 16492
rect 3872 16438 3874 16490
rect 3874 16438 3926 16490
rect 3926 16438 3928 16490
rect 3872 16436 3928 16438
rect 3976 16490 4032 16492
rect 3976 16438 3978 16490
rect 3978 16438 4030 16490
rect 4030 16438 4032 16490
rect 3976 16436 4032 16438
rect 4080 16490 4136 16492
rect 4080 16438 4082 16490
rect 4082 16438 4134 16490
rect 4134 16438 4136 16490
rect 4080 16436 4136 16438
rect 9192 16490 9248 16492
rect 9192 16438 9194 16490
rect 9194 16438 9246 16490
rect 9246 16438 9248 16490
rect 9192 16436 9248 16438
rect 9296 16490 9352 16492
rect 9296 16438 9298 16490
rect 9298 16438 9350 16490
rect 9350 16438 9352 16490
rect 9296 16436 9352 16438
rect 9400 16490 9456 16492
rect 9400 16438 9402 16490
rect 9402 16438 9454 16490
rect 9454 16438 9456 16490
rect 9400 16436 9456 16438
rect 14512 16490 14568 16492
rect 14512 16438 14514 16490
rect 14514 16438 14566 16490
rect 14566 16438 14568 16490
rect 14512 16436 14568 16438
rect 14616 16490 14672 16492
rect 14616 16438 14618 16490
rect 14618 16438 14670 16490
rect 14670 16438 14672 16490
rect 14616 16436 14672 16438
rect 14720 16490 14776 16492
rect 14720 16438 14722 16490
rect 14722 16438 14774 16490
rect 14774 16438 14776 16490
rect 14720 16436 14776 16438
rect 19832 16490 19888 16492
rect 19832 16438 19834 16490
rect 19834 16438 19886 16490
rect 19886 16438 19888 16490
rect 19832 16436 19888 16438
rect 19936 16490 19992 16492
rect 19936 16438 19938 16490
rect 19938 16438 19990 16490
rect 19990 16438 19992 16490
rect 19936 16436 19992 16438
rect 20040 16490 20096 16492
rect 20040 16438 20042 16490
rect 20042 16438 20094 16490
rect 20094 16438 20096 16490
rect 20040 16436 20096 16438
rect 6532 15706 6588 15708
rect 6532 15654 6534 15706
rect 6534 15654 6586 15706
rect 6586 15654 6588 15706
rect 6532 15652 6588 15654
rect 6636 15706 6692 15708
rect 6636 15654 6638 15706
rect 6638 15654 6690 15706
rect 6690 15654 6692 15706
rect 6636 15652 6692 15654
rect 6740 15706 6796 15708
rect 6740 15654 6742 15706
rect 6742 15654 6794 15706
rect 6794 15654 6796 15706
rect 6740 15652 6796 15654
rect 11852 15706 11908 15708
rect 11852 15654 11854 15706
rect 11854 15654 11906 15706
rect 11906 15654 11908 15706
rect 11852 15652 11908 15654
rect 11956 15706 12012 15708
rect 11956 15654 11958 15706
rect 11958 15654 12010 15706
rect 12010 15654 12012 15706
rect 11956 15652 12012 15654
rect 12060 15706 12116 15708
rect 12060 15654 12062 15706
rect 12062 15654 12114 15706
rect 12114 15654 12116 15706
rect 12060 15652 12116 15654
rect 17172 15706 17228 15708
rect 17172 15654 17174 15706
rect 17174 15654 17226 15706
rect 17226 15654 17228 15706
rect 17172 15652 17228 15654
rect 17276 15706 17332 15708
rect 17276 15654 17278 15706
rect 17278 15654 17330 15706
rect 17330 15654 17332 15706
rect 17276 15652 17332 15654
rect 17380 15706 17436 15708
rect 17380 15654 17382 15706
rect 17382 15654 17434 15706
rect 17434 15654 17436 15706
rect 17380 15652 17436 15654
rect 22492 15706 22548 15708
rect 22492 15654 22494 15706
rect 22494 15654 22546 15706
rect 22546 15654 22548 15706
rect 22492 15652 22548 15654
rect 22596 15706 22652 15708
rect 22596 15654 22598 15706
rect 22598 15654 22650 15706
rect 22650 15654 22652 15706
rect 22596 15652 22652 15654
rect 22700 15706 22756 15708
rect 22700 15654 22702 15706
rect 22702 15654 22754 15706
rect 22754 15654 22756 15706
rect 22700 15652 22756 15654
rect 3612 14924 3668 14980
rect 3500 9154 3556 9156
rect 3500 9102 3502 9154
rect 3502 9102 3554 9154
rect 3554 9102 3556 9154
rect 3500 9100 3556 9102
rect 3872 14922 3928 14924
rect 3872 14870 3874 14922
rect 3874 14870 3926 14922
rect 3926 14870 3928 14922
rect 3872 14868 3928 14870
rect 3976 14922 4032 14924
rect 3976 14870 3978 14922
rect 3978 14870 4030 14922
rect 4030 14870 4032 14922
rect 3976 14868 4032 14870
rect 4080 14922 4136 14924
rect 4080 14870 4082 14922
rect 4082 14870 4134 14922
rect 4134 14870 4136 14922
rect 4080 14868 4136 14870
rect 9192 14922 9248 14924
rect 9192 14870 9194 14922
rect 9194 14870 9246 14922
rect 9246 14870 9248 14922
rect 9192 14868 9248 14870
rect 9296 14922 9352 14924
rect 9296 14870 9298 14922
rect 9298 14870 9350 14922
rect 9350 14870 9352 14922
rect 9296 14868 9352 14870
rect 9400 14922 9456 14924
rect 9400 14870 9402 14922
rect 9402 14870 9454 14922
rect 9454 14870 9456 14922
rect 9400 14868 9456 14870
rect 14512 14922 14568 14924
rect 14512 14870 14514 14922
rect 14514 14870 14566 14922
rect 14566 14870 14568 14922
rect 14512 14868 14568 14870
rect 14616 14922 14672 14924
rect 14616 14870 14618 14922
rect 14618 14870 14670 14922
rect 14670 14870 14672 14922
rect 14616 14868 14672 14870
rect 14720 14922 14776 14924
rect 14720 14870 14722 14922
rect 14722 14870 14774 14922
rect 14774 14870 14776 14922
rect 14720 14868 14776 14870
rect 19832 14922 19888 14924
rect 19832 14870 19834 14922
rect 19834 14870 19886 14922
rect 19886 14870 19888 14922
rect 19832 14868 19888 14870
rect 19936 14922 19992 14924
rect 19936 14870 19938 14922
rect 19938 14870 19990 14922
rect 19990 14870 19992 14922
rect 19936 14868 19992 14870
rect 20040 14922 20096 14924
rect 20040 14870 20042 14922
rect 20042 14870 20094 14922
rect 20094 14870 20096 14922
rect 20040 14868 20096 14870
rect 19628 14700 19684 14756
rect 6532 14138 6588 14140
rect 6532 14086 6534 14138
rect 6534 14086 6586 14138
rect 6586 14086 6588 14138
rect 6532 14084 6588 14086
rect 6636 14138 6692 14140
rect 6636 14086 6638 14138
rect 6638 14086 6690 14138
rect 6690 14086 6692 14138
rect 6636 14084 6692 14086
rect 6740 14138 6796 14140
rect 6740 14086 6742 14138
rect 6742 14086 6794 14138
rect 6794 14086 6796 14138
rect 6740 14084 6796 14086
rect 11852 14138 11908 14140
rect 11852 14086 11854 14138
rect 11854 14086 11906 14138
rect 11906 14086 11908 14138
rect 11852 14084 11908 14086
rect 11956 14138 12012 14140
rect 11956 14086 11958 14138
rect 11958 14086 12010 14138
rect 12010 14086 12012 14138
rect 11956 14084 12012 14086
rect 12060 14138 12116 14140
rect 12060 14086 12062 14138
rect 12062 14086 12114 14138
rect 12114 14086 12116 14138
rect 12060 14084 12116 14086
rect 3872 13354 3928 13356
rect 3872 13302 3874 13354
rect 3874 13302 3926 13354
rect 3926 13302 3928 13354
rect 3872 13300 3928 13302
rect 3976 13354 4032 13356
rect 3976 13302 3978 13354
rect 3978 13302 4030 13354
rect 4030 13302 4032 13354
rect 3976 13300 4032 13302
rect 4080 13354 4136 13356
rect 4080 13302 4082 13354
rect 4082 13302 4134 13354
rect 4134 13302 4136 13354
rect 4080 13300 4136 13302
rect 9192 13354 9248 13356
rect 9192 13302 9194 13354
rect 9194 13302 9246 13354
rect 9246 13302 9248 13354
rect 9192 13300 9248 13302
rect 9296 13354 9352 13356
rect 9296 13302 9298 13354
rect 9298 13302 9350 13354
rect 9350 13302 9352 13354
rect 9296 13300 9352 13302
rect 9400 13354 9456 13356
rect 9400 13302 9402 13354
rect 9402 13302 9454 13354
rect 9454 13302 9456 13354
rect 9400 13300 9456 13302
rect 14512 13354 14568 13356
rect 14512 13302 14514 13354
rect 14514 13302 14566 13354
rect 14566 13302 14568 13354
rect 14512 13300 14568 13302
rect 14616 13354 14672 13356
rect 14616 13302 14618 13354
rect 14618 13302 14670 13354
rect 14670 13302 14672 13354
rect 14616 13300 14672 13302
rect 14720 13354 14776 13356
rect 14720 13302 14722 13354
rect 14722 13302 14774 13354
rect 14774 13302 14776 13354
rect 14720 13300 14776 13302
rect 14924 13186 14980 13188
rect 14924 13134 14926 13186
rect 14926 13134 14978 13186
rect 14978 13134 14980 13186
rect 14924 13132 14980 13134
rect 16268 13522 16324 13524
rect 16268 13470 16270 13522
rect 16270 13470 16322 13522
rect 16322 13470 16324 13522
rect 16268 13468 16324 13470
rect 6532 12570 6588 12572
rect 6532 12518 6534 12570
rect 6534 12518 6586 12570
rect 6586 12518 6588 12570
rect 6532 12516 6588 12518
rect 6636 12570 6692 12572
rect 6636 12518 6638 12570
rect 6638 12518 6690 12570
rect 6690 12518 6692 12570
rect 6636 12516 6692 12518
rect 6740 12570 6796 12572
rect 6740 12518 6742 12570
rect 6742 12518 6794 12570
rect 6794 12518 6796 12570
rect 6740 12516 6796 12518
rect 11852 12570 11908 12572
rect 11852 12518 11854 12570
rect 11854 12518 11906 12570
rect 11906 12518 11908 12570
rect 11852 12516 11908 12518
rect 11956 12570 12012 12572
rect 11956 12518 11958 12570
rect 11958 12518 12010 12570
rect 12010 12518 12012 12570
rect 11956 12516 12012 12518
rect 12060 12570 12116 12572
rect 12060 12518 12062 12570
rect 12062 12518 12114 12570
rect 12114 12518 12116 12570
rect 12060 12516 12116 12518
rect 3872 11786 3928 11788
rect 3872 11734 3874 11786
rect 3874 11734 3926 11786
rect 3926 11734 3928 11786
rect 3872 11732 3928 11734
rect 3976 11786 4032 11788
rect 3976 11734 3978 11786
rect 3978 11734 4030 11786
rect 4030 11734 4032 11786
rect 3976 11732 4032 11734
rect 4080 11786 4136 11788
rect 4080 11734 4082 11786
rect 4082 11734 4134 11786
rect 4134 11734 4136 11786
rect 4080 11732 4136 11734
rect 9192 11786 9248 11788
rect 9192 11734 9194 11786
rect 9194 11734 9246 11786
rect 9246 11734 9248 11786
rect 9192 11732 9248 11734
rect 9296 11786 9352 11788
rect 9296 11734 9298 11786
rect 9298 11734 9350 11786
rect 9350 11734 9352 11786
rect 9296 11732 9352 11734
rect 9400 11786 9456 11788
rect 9400 11734 9402 11786
rect 9402 11734 9454 11786
rect 9454 11734 9456 11786
rect 9400 11732 9456 11734
rect 6188 11282 6244 11284
rect 6188 11230 6190 11282
rect 6190 11230 6242 11282
rect 6242 11230 6244 11282
rect 6188 11228 6244 11230
rect 5516 10722 5572 10724
rect 5516 10670 5518 10722
rect 5518 10670 5570 10722
rect 5570 10670 5572 10722
rect 5516 10668 5572 10670
rect 3872 10218 3928 10220
rect 3872 10166 3874 10218
rect 3874 10166 3926 10218
rect 3926 10166 3928 10218
rect 3872 10164 3928 10166
rect 3976 10218 4032 10220
rect 3976 10166 3978 10218
rect 3978 10166 4030 10218
rect 4030 10166 4032 10218
rect 3976 10164 4032 10166
rect 4080 10218 4136 10220
rect 4080 10166 4082 10218
rect 4082 10166 4134 10218
rect 4134 10166 4136 10218
rect 4080 10164 4136 10166
rect 4284 9826 4340 9828
rect 4284 9774 4286 9826
rect 4286 9774 4338 9826
rect 4338 9774 4340 9826
rect 4284 9772 4340 9774
rect 4844 9826 4900 9828
rect 4844 9774 4846 9826
rect 4846 9774 4898 9826
rect 4898 9774 4900 9826
rect 4844 9772 4900 9774
rect 6972 11282 7028 11284
rect 6972 11230 6974 11282
rect 6974 11230 7026 11282
rect 7026 11230 7028 11282
rect 6972 11228 7028 11230
rect 6532 11002 6588 11004
rect 6532 10950 6534 11002
rect 6534 10950 6586 11002
rect 6586 10950 6588 11002
rect 6532 10948 6588 10950
rect 6636 11002 6692 11004
rect 6636 10950 6638 11002
rect 6638 10950 6690 11002
rect 6690 10950 6692 11002
rect 6636 10948 6692 10950
rect 6740 11002 6796 11004
rect 6740 10950 6742 11002
rect 6742 10950 6794 11002
rect 6794 10950 6796 11002
rect 6740 10948 6796 10950
rect 6076 10722 6132 10724
rect 6076 10670 6078 10722
rect 6078 10670 6130 10722
rect 6130 10670 6132 10722
rect 6076 10668 6132 10670
rect 5404 9772 5460 9828
rect 5852 9714 5908 9716
rect 5852 9662 5854 9714
rect 5854 9662 5906 9714
rect 5906 9662 5908 9714
rect 5852 9660 5908 9662
rect 4060 9154 4116 9156
rect 4060 9102 4062 9154
rect 4062 9102 4114 9154
rect 4114 9102 4116 9154
rect 4060 9100 4116 9102
rect 3872 8650 3928 8652
rect 3872 8598 3874 8650
rect 3874 8598 3926 8650
rect 3926 8598 3928 8650
rect 3872 8596 3928 8598
rect 3976 8650 4032 8652
rect 3976 8598 3978 8650
rect 3978 8598 4030 8650
rect 4030 8598 4032 8650
rect 3976 8596 4032 8598
rect 4080 8650 4136 8652
rect 4080 8598 4082 8650
rect 4082 8598 4134 8650
rect 4134 8598 4136 8650
rect 4080 8596 4136 8598
rect 3612 8428 3668 8484
rect 4172 8428 4228 8484
rect 2156 7474 2212 7476
rect 2156 7422 2158 7474
rect 2158 7422 2210 7474
rect 2210 7422 2212 7474
rect 2156 7420 2212 7422
rect 2716 7474 2772 7476
rect 2716 7422 2718 7474
rect 2718 7422 2770 7474
rect 2770 7422 2772 7474
rect 2716 7420 2772 7422
rect 2156 6578 2212 6580
rect 2156 6526 2158 6578
rect 2158 6526 2210 6578
rect 2210 6526 2212 6578
rect 2156 6524 2212 6526
rect 2828 6748 2884 6804
rect 2828 6578 2884 6580
rect 2828 6526 2830 6578
rect 2830 6526 2882 6578
rect 2882 6526 2884 6578
rect 2828 6524 2884 6526
rect 3612 7196 3668 7252
rect 3388 6524 3444 6580
rect 2716 5068 2772 5124
rect 4284 8034 4340 8036
rect 4284 7982 4286 8034
rect 4286 7982 4338 8034
rect 4338 7982 4340 8034
rect 4284 7980 4340 7982
rect 4732 8428 4788 8484
rect 4172 7250 4228 7252
rect 4172 7198 4174 7250
rect 4174 7198 4226 7250
rect 4226 7198 4228 7250
rect 4172 7196 4228 7198
rect 3872 7082 3928 7084
rect 3872 7030 3874 7082
rect 3874 7030 3926 7082
rect 3926 7030 3928 7082
rect 3872 7028 3928 7030
rect 3976 7082 4032 7084
rect 3976 7030 3978 7082
rect 3978 7030 4030 7082
rect 4030 7030 4032 7082
rect 3976 7028 4032 7030
rect 4080 7082 4136 7084
rect 4080 7030 4082 7082
rect 4082 7030 4134 7082
rect 4134 7030 4136 7082
rect 4080 7028 4136 7030
rect 6524 9714 6580 9716
rect 6524 9662 6526 9714
rect 6526 9662 6578 9714
rect 6578 9662 6580 9714
rect 6524 9660 6580 9662
rect 9192 10218 9248 10220
rect 9192 10166 9194 10218
rect 9194 10166 9246 10218
rect 9246 10166 9248 10218
rect 9192 10164 9248 10166
rect 9296 10218 9352 10220
rect 9296 10166 9298 10218
rect 9298 10166 9350 10218
rect 9350 10166 9352 10218
rect 9296 10164 9352 10166
rect 9400 10218 9456 10220
rect 9400 10166 9402 10218
rect 9402 10166 9454 10218
rect 9454 10166 9456 10218
rect 9400 10164 9456 10166
rect 8988 9996 9044 10052
rect 9996 10108 10052 10164
rect 7196 9714 7252 9716
rect 7196 9662 7198 9714
rect 7198 9662 7250 9714
rect 7250 9662 7252 9714
rect 7196 9660 7252 9662
rect 4956 8482 5012 8484
rect 4956 8430 4958 8482
rect 4958 8430 5010 8482
rect 5010 8430 5012 8482
rect 4956 8428 5012 8430
rect 5404 8428 5460 8484
rect 4844 7980 4900 8036
rect 6532 9434 6588 9436
rect 6532 9382 6534 9434
rect 6534 9382 6586 9434
rect 6586 9382 6588 9434
rect 6532 9380 6588 9382
rect 6636 9434 6692 9436
rect 6636 9382 6638 9434
rect 6638 9382 6690 9434
rect 6690 9382 6692 9434
rect 6636 9380 6692 9382
rect 6740 9434 6796 9436
rect 6740 9382 6742 9434
rect 6742 9382 6794 9434
rect 6794 9382 6796 9434
rect 6740 9380 6796 9382
rect 5964 8482 6020 8484
rect 5964 8430 5966 8482
rect 5966 8430 6018 8482
rect 6018 8430 6020 8482
rect 5964 8428 6020 8430
rect 4844 7474 4900 7476
rect 4844 7422 4846 7474
rect 4846 7422 4898 7474
rect 4898 7422 4900 7474
rect 4844 7420 4900 7422
rect 6524 8428 6580 8484
rect 6532 7866 6588 7868
rect 6532 7814 6534 7866
rect 6534 7814 6586 7866
rect 6586 7814 6588 7866
rect 6532 7812 6588 7814
rect 6636 7866 6692 7868
rect 6636 7814 6638 7866
rect 6638 7814 6690 7866
rect 6690 7814 6692 7866
rect 6636 7812 6692 7814
rect 6740 7866 6796 7868
rect 6740 7814 6742 7866
rect 6742 7814 6794 7866
rect 6794 7814 6796 7866
rect 6740 7812 6796 7814
rect 5404 7474 5460 7476
rect 5404 7422 5406 7474
rect 5406 7422 5458 7474
rect 5458 7422 5460 7474
rect 5404 7420 5460 7422
rect 6076 7474 6132 7476
rect 6076 7422 6078 7474
rect 6078 7422 6130 7474
rect 6130 7422 6132 7474
rect 6076 7420 6132 7422
rect 3724 6748 3780 6804
rect 4620 6748 4676 6804
rect 3388 5068 3444 5124
rect 4060 5906 4116 5908
rect 4060 5854 4062 5906
rect 4062 5854 4114 5906
rect 4114 5854 4116 5906
rect 4060 5852 4116 5854
rect 2380 4450 2436 4452
rect 2380 4398 2382 4450
rect 2382 4398 2434 4450
rect 2434 4398 2436 4450
rect 2380 4396 2436 4398
rect 3052 4396 3108 4452
rect 2492 4338 2548 4340
rect 2492 4286 2494 4338
rect 2494 4286 2546 4338
rect 2546 4286 2548 4338
rect 2492 4284 2548 4286
rect 2828 4284 2884 4340
rect 2156 3500 2212 3556
rect 3164 4338 3220 4340
rect 3164 4286 3166 4338
rect 3166 4286 3218 4338
rect 3218 4286 3220 4338
rect 3164 4284 3220 4286
rect 5516 6748 5572 6804
rect 5740 6748 5796 6804
rect 4732 5906 4788 5908
rect 4732 5854 4734 5906
rect 4734 5854 4786 5906
rect 4786 5854 4788 5906
rect 4732 5852 4788 5854
rect 7196 8428 7252 8484
rect 8652 9602 8708 9604
rect 8652 9550 8654 9602
rect 8654 9550 8706 9602
rect 8706 9550 8708 9602
rect 8652 9548 8708 9550
rect 7980 8428 8036 8484
rect 7308 8034 7364 8036
rect 7308 7982 7310 8034
rect 7310 7982 7362 8034
rect 7362 7982 7364 8034
rect 7308 7980 7364 7982
rect 6748 7474 6804 7476
rect 6748 7422 6750 7474
rect 6750 7422 6802 7474
rect 6802 7422 6804 7474
rect 6748 7420 6804 7422
rect 6412 6748 6468 6804
rect 7308 7420 7364 7476
rect 7980 8034 8036 8036
rect 7980 7982 7982 8034
rect 7982 7982 8034 8034
rect 8034 7982 8036 8034
rect 7980 7980 8036 7982
rect 9324 9602 9380 9604
rect 9324 9550 9326 9602
rect 9326 9550 9378 9602
rect 9378 9550 9380 9602
rect 9324 9548 9380 9550
rect 8540 8428 8596 8484
rect 9192 8650 9248 8652
rect 9192 8598 9194 8650
rect 9194 8598 9246 8650
rect 9246 8598 9248 8650
rect 9192 8596 9248 8598
rect 9296 8650 9352 8652
rect 9296 8598 9298 8650
rect 9298 8598 9350 8650
rect 9350 8598 9352 8650
rect 9296 8596 9352 8598
rect 9400 8650 9456 8652
rect 9400 8598 9402 8650
rect 9402 8598 9454 8650
rect 9454 8598 9456 8650
rect 9400 8596 9456 8598
rect 9324 8482 9380 8484
rect 9324 8430 9326 8482
rect 9326 8430 9378 8482
rect 9378 8430 9380 8482
rect 9324 8428 9380 8430
rect 8316 7980 8372 8036
rect 8988 8316 9044 8372
rect 7532 6860 7588 6916
rect 6532 6298 6588 6300
rect 6532 6246 6534 6298
rect 6534 6246 6586 6298
rect 6586 6246 6588 6298
rect 6532 6244 6588 6246
rect 6636 6298 6692 6300
rect 6636 6246 6638 6298
rect 6638 6246 6690 6298
rect 6690 6246 6692 6298
rect 6636 6244 6692 6246
rect 6740 6298 6796 6300
rect 6740 6246 6742 6298
rect 6742 6246 6794 6298
rect 6794 6246 6796 6298
rect 6740 6244 6796 6246
rect 3872 5514 3928 5516
rect 3872 5462 3874 5514
rect 3874 5462 3926 5514
rect 3926 5462 3928 5514
rect 3872 5460 3928 5462
rect 3976 5514 4032 5516
rect 3976 5462 3978 5514
rect 3978 5462 4030 5514
rect 4030 5462 4032 5514
rect 3976 5460 4032 5462
rect 4080 5514 4136 5516
rect 4080 5462 4082 5514
rect 4082 5462 4134 5514
rect 4134 5462 4136 5514
rect 4080 5460 4136 5462
rect 4172 5122 4228 5124
rect 4172 5070 4174 5122
rect 4174 5070 4226 5122
rect 4226 5070 4228 5122
rect 4172 5068 4228 5070
rect 3612 5010 3668 5012
rect 3612 4958 3614 5010
rect 3614 4958 3666 5010
rect 3666 4958 3668 5010
rect 3612 4956 3668 4958
rect 3836 4562 3892 4564
rect 3836 4510 3838 4562
rect 3838 4510 3890 4562
rect 3890 4510 3892 4562
rect 3836 4508 3892 4510
rect 3500 4284 3556 4340
rect 3724 4338 3780 4340
rect 3724 4286 3726 4338
rect 3726 4286 3778 4338
rect 3778 4286 3780 4338
rect 3724 4284 3780 4286
rect 2828 3554 2884 3556
rect 2828 3502 2830 3554
rect 2830 3502 2882 3554
rect 2882 3502 2884 3554
rect 2828 3500 2884 3502
rect 4732 4844 4788 4900
rect 4508 4562 4564 4564
rect 4508 4510 4510 4562
rect 4510 4510 4562 4562
rect 4562 4510 4564 4562
rect 4508 4508 4564 4510
rect 4956 5068 5012 5124
rect 4956 4898 5012 4900
rect 4956 4846 4958 4898
rect 4958 4846 5010 4898
rect 5010 4846 5012 4898
rect 4956 4844 5012 4846
rect 4844 4508 4900 4564
rect 4396 4338 4452 4340
rect 4396 4286 4398 4338
rect 4398 4286 4450 4338
rect 4450 4286 4452 4338
rect 4396 4284 4452 4286
rect 4284 4060 4340 4116
rect 3872 3946 3928 3948
rect 3872 3894 3874 3946
rect 3874 3894 3926 3946
rect 3926 3894 3928 3946
rect 3872 3892 3928 3894
rect 3976 3946 4032 3948
rect 3976 3894 3978 3946
rect 3978 3894 4030 3946
rect 4030 3894 4032 3946
rect 3976 3892 4032 3894
rect 4080 3946 4136 3948
rect 4080 3894 4082 3946
rect 4082 3894 4134 3946
rect 4134 3894 4136 3946
rect 4080 3892 4136 3894
rect 3052 3500 3108 3556
rect 3500 3554 3556 3556
rect 3500 3502 3502 3554
rect 3502 3502 3554 3554
rect 3554 3502 3556 3554
rect 3500 3500 3556 3502
rect 4172 3554 4228 3556
rect 4172 3502 4174 3554
rect 4174 3502 4226 3554
rect 4226 3502 4228 3554
rect 4172 3500 4228 3502
rect 5404 4844 5460 4900
rect 5852 4844 5908 4900
rect 5740 4508 5796 4564
rect 4396 3388 4452 3444
rect 4844 3442 4900 3444
rect 4844 3390 4846 3442
rect 4846 3390 4898 3442
rect 4898 3390 4900 3442
rect 4844 3388 4900 3390
rect 5852 4114 5908 4116
rect 5852 4062 5854 4114
rect 5854 4062 5906 4114
rect 5906 4062 5908 4114
rect 5852 4060 5908 4062
rect 7084 5964 7140 6020
rect 7420 6018 7476 6020
rect 7420 5966 7422 6018
rect 7422 5966 7474 6018
rect 7474 5966 7476 6018
rect 7420 5964 7476 5966
rect 7756 5964 7812 6020
rect 9884 8316 9940 8372
rect 9212 8258 9268 8260
rect 9212 8206 9214 8258
rect 9214 8206 9266 8258
rect 9266 8206 9268 8258
rect 9212 8204 9268 8206
rect 11852 11002 11908 11004
rect 11852 10950 11854 11002
rect 11854 10950 11906 11002
rect 11906 10950 11908 11002
rect 11852 10948 11908 10950
rect 11956 11002 12012 11004
rect 11956 10950 11958 11002
rect 11958 10950 12010 11002
rect 12010 10950 12012 11002
rect 11956 10948 12012 10950
rect 12060 11002 12116 11004
rect 12060 10950 12062 11002
rect 12062 10950 12114 11002
rect 12114 10950 12116 11002
rect 12060 10948 12116 10950
rect 14812 12178 14868 12180
rect 14812 12126 14814 12178
rect 14814 12126 14866 12178
rect 14866 12126 14868 12178
rect 14812 12124 14868 12126
rect 14252 11954 14308 11956
rect 14252 11902 14254 11954
rect 14254 11902 14306 11954
rect 14306 11902 14308 11954
rect 14252 11900 14308 11902
rect 14924 11954 14980 11956
rect 14924 11902 14926 11954
rect 14926 11902 14978 11954
rect 14978 11902 14980 11954
rect 14924 11900 14980 11902
rect 14512 11786 14568 11788
rect 14512 11734 14514 11786
rect 14514 11734 14566 11786
rect 14566 11734 14568 11786
rect 14512 11732 14568 11734
rect 14616 11786 14672 11788
rect 14616 11734 14618 11786
rect 14618 11734 14670 11786
rect 14670 11734 14672 11786
rect 14616 11732 14672 11734
rect 14720 11786 14776 11788
rect 14720 11734 14722 11786
rect 14722 11734 14774 11786
rect 14774 11734 14776 11786
rect 14720 11732 14776 11734
rect 14924 11394 14980 11396
rect 14924 11342 14926 11394
rect 14926 11342 14978 11394
rect 14978 11342 14980 11394
rect 14924 11340 14980 11342
rect 11340 9996 11396 10052
rect 14512 10218 14568 10220
rect 14512 10166 14514 10218
rect 14514 10166 14566 10218
rect 14566 10166 14568 10218
rect 14512 10164 14568 10166
rect 14616 10218 14672 10220
rect 14616 10166 14618 10218
rect 14618 10166 14670 10218
rect 14670 10166 14672 10218
rect 14616 10164 14672 10166
rect 14720 10218 14776 10220
rect 14720 10166 14722 10218
rect 14722 10166 14774 10218
rect 14774 10166 14776 10218
rect 14720 10164 14776 10166
rect 12012 9996 12068 10052
rect 15484 12178 15540 12180
rect 15484 12126 15486 12178
rect 15486 12126 15538 12178
rect 15538 12126 15540 12178
rect 15484 12124 15540 12126
rect 15596 11394 15652 11396
rect 15596 11342 15598 11394
rect 15598 11342 15650 11394
rect 15650 11342 15652 11394
rect 15596 11340 15652 11342
rect 16156 12178 16212 12180
rect 16156 12126 16158 12178
rect 16158 12126 16210 12178
rect 16210 12126 16212 12178
rect 16156 12124 16212 12126
rect 16940 13522 16996 13524
rect 16940 13470 16942 13522
rect 16942 13470 16994 13522
rect 16994 13470 16996 13522
rect 16940 13468 16996 13470
rect 17172 14138 17228 14140
rect 17172 14086 17174 14138
rect 17174 14086 17226 14138
rect 17226 14086 17228 14138
rect 17172 14084 17228 14086
rect 17276 14138 17332 14140
rect 17276 14086 17278 14138
rect 17278 14086 17330 14138
rect 17330 14086 17332 14138
rect 17276 14084 17332 14086
rect 17380 14138 17436 14140
rect 17380 14086 17382 14138
rect 17382 14086 17434 14138
rect 17434 14086 17436 14138
rect 17380 14084 17436 14086
rect 17052 13132 17108 13188
rect 17388 13468 17444 13524
rect 16828 12178 16884 12180
rect 16828 12126 16830 12178
rect 16830 12126 16882 12178
rect 16882 12126 16884 12178
rect 16828 12124 16884 12126
rect 17612 13468 17668 13524
rect 17724 13132 17780 13188
rect 18396 13468 18452 13524
rect 18508 13244 18564 13300
rect 18956 13468 19012 13524
rect 18284 13186 18340 13188
rect 18284 13134 18286 13186
rect 18286 13134 18338 13186
rect 18338 13134 18340 13186
rect 18284 13132 18340 13134
rect 18844 13132 18900 13188
rect 17172 12570 17228 12572
rect 17172 12518 17174 12570
rect 17174 12518 17226 12570
rect 17226 12518 17228 12570
rect 17172 12516 17228 12518
rect 17276 12570 17332 12572
rect 17276 12518 17278 12570
rect 17278 12518 17330 12570
rect 17330 12518 17332 12570
rect 17276 12516 17332 12518
rect 17380 12570 17436 12572
rect 17380 12518 17382 12570
rect 17382 12518 17434 12570
rect 17434 12518 17436 12570
rect 17380 12516 17436 12518
rect 16268 11394 16324 11396
rect 16268 11342 16270 11394
rect 16270 11342 16322 11394
rect 16322 11342 16324 11394
rect 16268 11340 16324 11342
rect 17612 11788 17668 11844
rect 22492 14138 22548 14140
rect 22492 14086 22494 14138
rect 22494 14086 22546 14138
rect 22546 14086 22548 14138
rect 22492 14084 22548 14086
rect 22596 14138 22652 14140
rect 22596 14086 22598 14138
rect 22598 14086 22650 14138
rect 22650 14086 22652 14138
rect 22596 14084 22652 14086
rect 22700 14138 22756 14140
rect 22700 14086 22702 14138
rect 22702 14086 22754 14138
rect 22754 14086 22756 14138
rect 22700 14084 22756 14086
rect 19628 13468 19684 13524
rect 18396 12290 18452 12292
rect 18396 12238 18398 12290
rect 18398 12238 18450 12290
rect 18450 12238 18452 12290
rect 18396 12236 18452 12238
rect 16940 11394 16996 11396
rect 16940 11342 16942 11394
rect 16942 11342 16994 11394
rect 16994 11342 16996 11394
rect 16940 11340 16996 11342
rect 9996 8540 10052 8596
rect 11852 9434 11908 9436
rect 11852 9382 11854 9434
rect 11854 9382 11906 9434
rect 11906 9382 11908 9434
rect 11852 9380 11908 9382
rect 11956 9434 12012 9436
rect 11956 9382 11958 9434
rect 11958 9382 12010 9434
rect 12010 9382 12012 9434
rect 11956 9380 12012 9382
rect 12060 9434 12116 9436
rect 12060 9382 12062 9434
rect 12062 9382 12114 9434
rect 12114 9382 12116 9434
rect 12060 9380 12116 9382
rect 10556 8540 10612 8596
rect 10332 8316 10388 8372
rect 9996 8204 10052 8260
rect 12460 8204 12516 8260
rect 12796 8428 12852 8484
rect 14364 9042 14420 9044
rect 14364 8990 14366 9042
rect 14366 8990 14418 9042
rect 14418 8990 14420 9042
rect 14364 8988 14420 8990
rect 13692 8428 13748 8484
rect 12908 8258 12964 8260
rect 12908 8206 12910 8258
rect 12910 8206 12962 8258
rect 12962 8206 12964 8258
rect 12908 8204 12964 8206
rect 13356 8204 13412 8260
rect 8428 6578 8484 6580
rect 8428 6526 8430 6578
rect 8430 6526 8482 6578
rect 8482 6526 8484 6578
rect 8428 6524 8484 6526
rect 8540 6690 8596 6692
rect 8540 6638 8542 6690
rect 8542 6638 8594 6690
rect 8594 6638 8596 6690
rect 8540 6636 8596 6638
rect 8092 6018 8148 6020
rect 8092 5966 8094 6018
rect 8094 5966 8146 6018
rect 8146 5966 8148 6018
rect 8092 5964 8148 5966
rect 6076 4844 6132 4900
rect 6300 4508 6356 4564
rect 6532 4730 6588 4732
rect 6532 4678 6534 4730
rect 6534 4678 6586 4730
rect 6586 4678 6588 4730
rect 6532 4676 6588 4678
rect 6636 4730 6692 4732
rect 6636 4678 6638 4730
rect 6638 4678 6690 4730
rect 6690 4678 6692 4730
rect 6636 4676 6692 4678
rect 6740 4730 6796 4732
rect 6740 4678 6742 4730
rect 6742 4678 6794 4730
rect 6794 4678 6796 4730
rect 6740 4676 6796 4678
rect 6076 4060 6132 4116
rect 5180 3388 5236 3444
rect 5740 3442 5796 3444
rect 5740 3390 5742 3442
rect 5742 3390 5794 3442
rect 5794 3390 5796 3442
rect 5740 3388 5796 3390
rect 7308 5068 7364 5124
rect 6524 4114 6580 4116
rect 6524 4062 6526 4114
rect 6526 4062 6578 4114
rect 6578 4062 6580 4114
rect 6524 4060 6580 4062
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 7084 4060 7140 4116
rect 7084 3500 7140 3556
rect 9192 7082 9248 7084
rect 9192 7030 9194 7082
rect 9194 7030 9246 7082
rect 9246 7030 9248 7082
rect 9192 7028 9248 7030
rect 9296 7082 9352 7084
rect 9296 7030 9298 7082
rect 9298 7030 9350 7082
rect 9350 7030 9352 7082
rect 9296 7028 9352 7030
rect 9400 7082 9456 7084
rect 9400 7030 9402 7082
rect 9402 7030 9454 7082
rect 9454 7030 9456 7082
rect 9400 7028 9456 7030
rect 8764 6636 8820 6692
rect 8876 6860 8932 6916
rect 9212 6690 9268 6692
rect 9212 6638 9214 6690
rect 9214 6638 9266 6690
rect 9266 6638 9268 6690
rect 9212 6636 9268 6638
rect 9884 6636 9940 6692
rect 9100 6578 9156 6580
rect 9100 6526 9102 6578
rect 9102 6526 9154 6578
rect 9154 6526 9156 6578
rect 9100 6524 9156 6526
rect 9996 6860 10052 6916
rect 9884 6466 9940 6468
rect 9884 6414 9886 6466
rect 9886 6414 9938 6466
rect 9938 6414 9940 6466
rect 9884 6412 9940 6414
rect 9100 5852 9156 5908
rect 9772 5906 9828 5908
rect 9772 5854 9774 5906
rect 9774 5854 9826 5906
rect 9826 5854 9828 5906
rect 9772 5852 9828 5854
rect 9192 5514 9248 5516
rect 9192 5462 9194 5514
rect 9194 5462 9246 5514
rect 9246 5462 9248 5514
rect 9192 5460 9248 5462
rect 9296 5514 9352 5516
rect 9296 5462 9298 5514
rect 9298 5462 9350 5514
rect 9350 5462 9352 5514
rect 9296 5460 9352 5462
rect 9400 5514 9456 5516
rect 9400 5462 9402 5514
rect 9402 5462 9454 5514
rect 9454 5462 9456 5514
rect 9400 5460 9456 5462
rect 7756 5122 7812 5124
rect 7756 5070 7758 5122
rect 7758 5070 7810 5122
rect 7810 5070 7812 5122
rect 7756 5068 7812 5070
rect 11852 7866 11908 7868
rect 11852 7814 11854 7866
rect 11854 7814 11906 7866
rect 11906 7814 11908 7866
rect 11852 7812 11908 7814
rect 11956 7866 12012 7868
rect 11956 7814 11958 7866
rect 11958 7814 12010 7866
rect 12010 7814 12012 7866
rect 11956 7812 12012 7814
rect 12060 7866 12116 7868
rect 12060 7814 12062 7866
rect 12062 7814 12114 7866
rect 12114 7814 12116 7866
rect 12060 7812 12116 7814
rect 10556 6914 10612 6916
rect 10556 6862 10558 6914
rect 10558 6862 10610 6914
rect 10610 6862 10612 6914
rect 10556 6860 10612 6862
rect 10444 6690 10500 6692
rect 10444 6638 10446 6690
rect 10446 6638 10498 6690
rect 10498 6638 10500 6690
rect 10444 6636 10500 6638
rect 11228 6914 11284 6916
rect 11228 6862 11230 6914
rect 11230 6862 11282 6914
rect 11282 6862 11284 6914
rect 11228 6860 11284 6862
rect 10556 6412 10612 6468
rect 11116 6690 11172 6692
rect 11116 6638 11118 6690
rect 11118 6638 11170 6690
rect 11170 6638 11172 6690
rect 11116 6636 11172 6638
rect 10444 5906 10500 5908
rect 10444 5854 10446 5906
rect 10446 5854 10498 5906
rect 10498 5854 10500 5906
rect 10444 5852 10500 5854
rect 8540 5068 8596 5124
rect 9100 5122 9156 5124
rect 9100 5070 9102 5122
rect 9102 5070 9154 5122
rect 9154 5070 9156 5122
rect 9100 5068 9156 5070
rect 9660 5068 9716 5124
rect 7756 4338 7812 4340
rect 7756 4286 7758 4338
rect 7758 4286 7810 4338
rect 7810 4286 7812 4338
rect 7756 4284 7812 4286
rect 7756 3554 7812 3556
rect 7756 3502 7758 3554
rect 7758 3502 7810 3554
rect 7810 3502 7812 3554
rect 7756 3500 7812 3502
rect 8428 3554 8484 3556
rect 8428 3502 8430 3554
rect 8430 3502 8482 3554
rect 8482 3502 8484 3554
rect 8428 3500 8484 3502
rect 9192 3946 9248 3948
rect 9192 3894 9194 3946
rect 9194 3894 9246 3946
rect 9246 3894 9248 3946
rect 9192 3892 9248 3894
rect 9296 3946 9352 3948
rect 9296 3894 9298 3946
rect 9298 3894 9350 3946
rect 9350 3894 9352 3946
rect 9296 3892 9352 3894
rect 9400 3946 9456 3948
rect 9400 3894 9402 3946
rect 9402 3894 9454 3946
rect 9454 3894 9456 3946
rect 9400 3892 9456 3894
rect 9660 3554 9716 3556
rect 9660 3502 9662 3554
rect 9662 3502 9714 3554
rect 9714 3502 9716 3554
rect 9660 3500 9716 3502
rect 9884 3500 9940 3556
rect 6636 3388 6692 3444
rect 6532 3162 6588 3164
rect 6532 3110 6534 3162
rect 6534 3110 6586 3162
rect 6586 3110 6588 3162
rect 6532 3108 6588 3110
rect 6636 3162 6692 3164
rect 6636 3110 6638 3162
rect 6638 3110 6690 3162
rect 6690 3110 6692 3162
rect 6636 3108 6692 3110
rect 6740 3162 6796 3164
rect 6740 3110 6742 3162
rect 6742 3110 6794 3162
rect 6794 3110 6796 3162
rect 6740 3108 6796 3110
rect 11900 6636 11956 6692
rect 12012 6860 12068 6916
rect 13804 8258 13860 8260
rect 13804 8206 13806 8258
rect 13806 8206 13858 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 12460 6690 12516 6692
rect 12460 6638 12462 6690
rect 12462 6638 12514 6690
rect 12514 6638 12516 6690
rect 12460 6636 12516 6638
rect 11852 6298 11908 6300
rect 11852 6246 11854 6298
rect 11854 6246 11906 6298
rect 11906 6246 11908 6298
rect 11852 6244 11908 6246
rect 11956 6298 12012 6300
rect 11956 6246 11958 6298
rect 11958 6246 12010 6298
rect 12010 6246 12012 6298
rect 11956 6244 12012 6246
rect 12060 6298 12116 6300
rect 12060 6246 12062 6298
rect 12062 6246 12114 6298
rect 12114 6246 12116 6298
rect 12060 6244 12116 6246
rect 13916 8428 13972 8484
rect 15036 9042 15092 9044
rect 15036 8990 15038 9042
rect 15038 8990 15090 9042
rect 15090 8990 15092 9042
rect 15036 8988 15092 8990
rect 17500 11394 17556 11396
rect 17500 11342 17502 11394
rect 17502 11342 17554 11394
rect 17554 11342 17556 11394
rect 17500 11340 17556 11342
rect 17172 11002 17228 11004
rect 17172 10950 17174 11002
rect 17174 10950 17226 11002
rect 17226 10950 17228 11002
rect 17172 10948 17228 10950
rect 17276 11002 17332 11004
rect 17276 10950 17278 11002
rect 17278 10950 17330 11002
rect 17330 10950 17332 11002
rect 17276 10948 17332 10950
rect 17380 11002 17436 11004
rect 17380 10950 17382 11002
rect 17382 10950 17434 11002
rect 17434 10950 17436 11002
rect 17380 10948 17436 10950
rect 19180 13132 19236 13188
rect 19832 13354 19888 13356
rect 19832 13302 19834 13354
rect 19834 13302 19886 13354
rect 19886 13302 19888 13354
rect 19832 13300 19888 13302
rect 19936 13354 19992 13356
rect 19936 13302 19938 13354
rect 19938 13302 19990 13354
rect 19990 13302 19992 13354
rect 19936 13300 19992 13302
rect 20040 13354 20096 13356
rect 20040 13302 20042 13354
rect 20042 13302 20094 13354
rect 20094 13302 20096 13354
rect 20040 13300 20096 13302
rect 18956 12236 19012 12292
rect 18508 11676 18564 11732
rect 15260 8988 15316 9044
rect 14512 8650 14568 8652
rect 14512 8598 14514 8650
rect 14514 8598 14566 8650
rect 14566 8598 14568 8650
rect 14512 8596 14568 8598
rect 14616 8650 14672 8652
rect 14616 8598 14618 8650
rect 14618 8598 14670 8650
rect 14670 8598 14672 8650
rect 14616 8596 14672 8598
rect 14720 8650 14776 8652
rect 14720 8598 14722 8650
rect 14722 8598 14774 8650
rect 14774 8598 14776 8650
rect 14720 8596 14776 8598
rect 14364 8428 14420 8484
rect 14476 8258 14532 8260
rect 14476 8206 14478 8258
rect 14478 8206 14530 8258
rect 14530 8206 14532 8258
rect 14476 8204 14532 8206
rect 15148 8482 15204 8484
rect 15148 8430 15150 8482
rect 15150 8430 15202 8482
rect 15202 8430 15204 8482
rect 15148 8428 15204 8430
rect 15036 8258 15092 8260
rect 15036 8206 15038 8258
rect 15038 8206 15090 8258
rect 15090 8206 15092 8258
rect 15036 8204 15092 8206
rect 14028 6860 14084 6916
rect 14512 7082 14568 7084
rect 14512 7030 14514 7082
rect 14514 7030 14566 7082
rect 14566 7030 14568 7082
rect 14512 7028 14568 7030
rect 14616 7082 14672 7084
rect 14616 7030 14618 7082
rect 14618 7030 14670 7082
rect 14670 7030 14672 7082
rect 14616 7028 14672 7030
rect 14720 7082 14776 7084
rect 14720 7030 14722 7082
rect 14722 7030 14774 7082
rect 14774 7030 14776 7082
rect 14720 7028 14776 7030
rect 14252 6914 14308 6916
rect 14252 6862 14254 6914
rect 14254 6862 14306 6914
rect 14306 6862 14308 6914
rect 14252 6860 14308 6862
rect 14588 6860 14644 6916
rect 11564 5122 11620 5124
rect 11564 5070 11566 5122
rect 11566 5070 11618 5122
rect 11618 5070 11620 5122
rect 11564 5068 11620 5070
rect 12124 5068 12180 5124
rect 12348 4844 12404 4900
rect 11852 4730 11908 4732
rect 11852 4678 11854 4730
rect 11854 4678 11906 4730
rect 11906 4678 11908 4730
rect 11852 4676 11908 4678
rect 11956 4730 12012 4732
rect 11956 4678 11958 4730
rect 11958 4678 12010 4730
rect 12010 4678 12012 4730
rect 11956 4676 12012 4678
rect 12060 4730 12116 4732
rect 12060 4678 12062 4730
rect 12062 4678 12114 4730
rect 12114 4678 12116 4730
rect 12060 4676 12116 4678
rect 12908 4898 12964 4900
rect 12908 4846 12910 4898
rect 12910 4846 12962 4898
rect 12962 4846 12964 4898
rect 12908 4844 12964 4846
rect 16828 10386 16884 10388
rect 16828 10334 16830 10386
rect 16830 10334 16882 10386
rect 16882 10334 16884 10386
rect 16828 10332 16884 10334
rect 18284 11170 18340 11172
rect 18284 11118 18286 11170
rect 18286 11118 18338 11170
rect 18338 11118 18340 11170
rect 18284 11116 18340 11118
rect 17836 10386 17892 10388
rect 17836 10334 17838 10386
rect 17838 10334 17890 10386
rect 17890 10334 17892 10386
rect 17836 10332 17892 10334
rect 18284 10332 18340 10388
rect 18956 11340 19012 11396
rect 18508 11116 18564 11172
rect 18956 11170 19012 11172
rect 18956 11118 18958 11170
rect 18958 11118 19010 11170
rect 19010 11118 19012 11170
rect 18956 11116 19012 11118
rect 22492 12570 22548 12572
rect 22492 12518 22494 12570
rect 22494 12518 22546 12570
rect 22546 12518 22548 12570
rect 22492 12516 22548 12518
rect 22596 12570 22652 12572
rect 22596 12518 22598 12570
rect 22598 12518 22650 12570
rect 22650 12518 22652 12570
rect 22596 12516 22652 12518
rect 22700 12570 22756 12572
rect 22700 12518 22702 12570
rect 22702 12518 22754 12570
rect 22754 12518 22756 12570
rect 22700 12516 22756 12518
rect 19740 12290 19796 12292
rect 19740 12238 19742 12290
rect 19742 12238 19794 12290
rect 19794 12238 19796 12290
rect 19740 12236 19796 12238
rect 20412 12290 20468 12292
rect 20412 12238 20414 12290
rect 20414 12238 20466 12290
rect 20466 12238 20468 12290
rect 20412 12236 20468 12238
rect 21084 12236 21140 12292
rect 19832 11786 19888 11788
rect 19832 11734 19834 11786
rect 19834 11734 19886 11786
rect 19886 11734 19888 11786
rect 19832 11732 19888 11734
rect 19936 11786 19992 11788
rect 19936 11734 19938 11786
rect 19938 11734 19990 11786
rect 19990 11734 19992 11786
rect 19936 11732 19992 11734
rect 20040 11786 20096 11788
rect 20040 11734 20042 11786
rect 20042 11734 20094 11786
rect 20094 11734 20096 11786
rect 20040 11732 20096 11734
rect 19516 11394 19572 11396
rect 19516 11342 19518 11394
rect 19518 11342 19570 11394
rect 19570 11342 19572 11394
rect 19516 11340 19572 11342
rect 18508 10386 18564 10388
rect 18508 10334 18510 10386
rect 18510 10334 18562 10386
rect 18562 10334 18564 10386
rect 18508 10332 18564 10334
rect 19852 11340 19908 11396
rect 19852 10668 19908 10724
rect 20188 10668 20244 10724
rect 19832 10218 19888 10220
rect 19832 10166 19834 10218
rect 19834 10166 19886 10218
rect 19886 10166 19888 10218
rect 19832 10164 19888 10166
rect 19936 10218 19992 10220
rect 19936 10166 19938 10218
rect 19938 10166 19990 10218
rect 19990 10166 19992 10218
rect 19936 10164 19992 10166
rect 20040 10218 20096 10220
rect 20040 10166 20042 10218
rect 20042 10166 20094 10218
rect 20094 10166 20096 10218
rect 20040 10164 20096 10166
rect 19852 9996 19908 10052
rect 15596 8204 15652 8260
rect 15708 8428 15764 8484
rect 10332 3554 10388 3556
rect 10332 3502 10334 3554
rect 10334 3502 10386 3554
rect 10386 3502 10388 3554
rect 10332 3500 10388 3502
rect 12460 4114 12516 4116
rect 12460 4062 12462 4114
rect 12462 4062 12514 4114
rect 12514 4062 12516 4114
rect 12460 4060 12516 4062
rect 13132 4114 13188 4116
rect 13132 4062 13134 4114
rect 13134 4062 13186 4114
rect 13186 4062 13188 4114
rect 13132 4060 13188 4062
rect 11116 3554 11172 3556
rect 11116 3502 11118 3554
rect 11118 3502 11170 3554
rect 11170 3502 11172 3554
rect 11116 3500 11172 3502
rect 11676 3554 11732 3556
rect 11676 3502 11678 3554
rect 11678 3502 11730 3554
rect 11730 3502 11732 3554
rect 11676 3500 11732 3502
rect 11004 3442 11060 3444
rect 11004 3390 11006 3442
rect 11006 3390 11058 3442
rect 11058 3390 11060 3442
rect 11004 3388 11060 3390
rect 11788 3442 11844 3444
rect 11788 3390 11790 3442
rect 11790 3390 11842 3442
rect 11842 3390 11844 3442
rect 11788 3388 11844 3390
rect 11852 3162 11908 3164
rect 11852 3110 11854 3162
rect 11854 3110 11906 3162
rect 11906 3110 11908 3162
rect 11852 3108 11908 3110
rect 11956 3162 12012 3164
rect 11956 3110 11958 3162
rect 11958 3110 12010 3162
rect 12010 3110 12012 3162
rect 11956 3108 12012 3110
rect 12060 3162 12116 3164
rect 12060 3110 12062 3162
rect 12062 3110 12114 3162
rect 12114 3110 12116 3162
rect 12060 3108 12116 3110
rect 13804 4114 13860 4116
rect 13804 4062 13806 4114
rect 13806 4062 13858 4114
rect 13858 4062 13860 4114
rect 13804 4060 13860 4062
rect 14512 5514 14568 5516
rect 14512 5462 14514 5514
rect 14514 5462 14566 5514
rect 14566 5462 14568 5514
rect 14512 5460 14568 5462
rect 14616 5514 14672 5516
rect 14616 5462 14618 5514
rect 14618 5462 14670 5514
rect 14670 5462 14672 5514
rect 14616 5460 14672 5462
rect 14720 5514 14776 5516
rect 14720 5462 14722 5514
rect 14722 5462 14774 5514
rect 14774 5462 14776 5514
rect 14720 5460 14776 5462
rect 15260 6860 15316 6916
rect 15820 8258 15876 8260
rect 15820 8206 15822 8258
rect 15822 8206 15874 8258
rect 15874 8206 15876 8258
rect 15820 8204 15876 8206
rect 16492 9602 16548 9604
rect 16492 9550 16494 9602
rect 16494 9550 16546 9602
rect 16546 9550 16548 9602
rect 16492 9548 16548 9550
rect 16268 8204 16324 8260
rect 16380 8428 16436 8484
rect 16492 8258 16548 8260
rect 16492 8206 16494 8258
rect 16494 8206 16546 8258
rect 16546 8206 16548 8258
rect 16492 8204 16548 8206
rect 17164 9602 17220 9604
rect 17164 9550 17166 9602
rect 17166 9550 17218 9602
rect 17218 9550 17220 9602
rect 17164 9548 17220 9550
rect 17172 9434 17228 9436
rect 17172 9382 17174 9434
rect 17174 9382 17226 9434
rect 17226 9382 17228 9434
rect 17172 9380 17228 9382
rect 17276 9434 17332 9436
rect 17276 9382 17278 9434
rect 17278 9382 17330 9434
rect 17330 9382 17332 9434
rect 17276 9380 17332 9382
rect 17380 9434 17436 9436
rect 17380 9382 17382 9434
rect 17382 9382 17434 9434
rect 17434 9382 17436 9434
rect 17380 9380 17436 9382
rect 17164 8482 17220 8484
rect 17164 8430 17166 8482
rect 17166 8430 17218 8482
rect 17218 8430 17220 8482
rect 17164 8428 17220 8430
rect 17052 8258 17108 8260
rect 17052 8206 17054 8258
rect 17054 8206 17106 8258
rect 17106 8206 17108 8258
rect 17052 8204 17108 8206
rect 17836 8482 17892 8484
rect 17836 8430 17838 8482
rect 17838 8430 17890 8482
rect 17890 8430 17892 8482
rect 17836 8428 17892 8430
rect 18508 8482 18564 8484
rect 18508 8430 18510 8482
rect 18510 8430 18562 8482
rect 18562 8430 18564 8482
rect 18508 8428 18564 8430
rect 18956 8764 19012 8820
rect 18956 8428 19012 8484
rect 19180 9602 19236 9604
rect 19180 9550 19182 9602
rect 19182 9550 19234 9602
rect 19234 9550 19236 9602
rect 19180 9548 19236 9550
rect 19852 9602 19908 9604
rect 19852 9550 19854 9602
rect 19854 9550 19906 9602
rect 19906 9550 19908 9602
rect 19852 9548 19908 9550
rect 21084 10722 21140 10724
rect 21084 10670 21086 10722
rect 21086 10670 21138 10722
rect 21138 10670 21140 10722
rect 21084 10668 21140 10670
rect 21756 11116 21812 11172
rect 22492 11002 22548 11004
rect 22492 10950 22494 11002
rect 22494 10950 22546 11002
rect 22546 10950 22548 11002
rect 22492 10948 22548 10950
rect 22596 11002 22652 11004
rect 22596 10950 22598 11002
rect 22598 10950 22650 11002
rect 22650 10950 22652 11002
rect 22596 10948 22652 10950
rect 22700 11002 22756 11004
rect 22700 10950 22702 11002
rect 22702 10950 22754 11002
rect 22754 10950 22756 11002
rect 22700 10948 22756 10950
rect 21868 10722 21924 10724
rect 21868 10670 21870 10722
rect 21870 10670 21922 10722
rect 21922 10670 21924 10722
rect 21868 10668 21924 10670
rect 20524 10050 20580 10052
rect 20524 9998 20526 10050
rect 20526 9998 20578 10050
rect 20578 9998 20580 10050
rect 20524 9996 20580 9998
rect 19180 8818 19236 8820
rect 19180 8766 19182 8818
rect 19182 8766 19234 8818
rect 19234 8766 19236 8818
rect 19180 8764 19236 8766
rect 17612 8204 17668 8260
rect 18396 8316 18452 8372
rect 17172 7866 17228 7868
rect 17172 7814 17174 7866
rect 17174 7814 17226 7866
rect 17226 7814 17228 7866
rect 17172 7812 17228 7814
rect 17276 7866 17332 7868
rect 17276 7814 17278 7866
rect 17278 7814 17330 7866
rect 17330 7814 17332 7866
rect 17276 7812 17332 7814
rect 17380 7866 17436 7868
rect 17380 7814 17382 7866
rect 17382 7814 17434 7866
rect 17434 7814 17436 7866
rect 17380 7812 17436 7814
rect 17836 7698 17892 7700
rect 17836 7646 17838 7698
rect 17838 7646 17890 7698
rect 17890 7646 17892 7698
rect 17836 7644 17892 7646
rect 16604 7474 16660 7476
rect 16604 7422 16606 7474
rect 16606 7422 16658 7474
rect 16658 7422 16660 7474
rect 16604 7420 16660 7422
rect 18396 7644 18452 7700
rect 17612 7420 17668 7476
rect 17724 7308 17780 7364
rect 16940 6578 16996 6580
rect 16940 6526 16942 6578
rect 16942 6526 16994 6578
rect 16994 6526 16996 6578
rect 16940 6524 16996 6526
rect 14700 5010 14756 5012
rect 14700 4958 14702 5010
rect 14702 4958 14754 5010
rect 14754 4958 14756 5010
rect 14700 4956 14756 4958
rect 14476 4338 14532 4340
rect 14476 4286 14478 4338
rect 14478 4286 14530 4338
rect 14530 4286 14532 4338
rect 14476 4284 14532 4286
rect 19180 8316 19236 8372
rect 19068 8258 19124 8260
rect 19068 8206 19070 8258
rect 19070 8206 19122 8258
rect 19122 8206 19124 8258
rect 19068 8204 19124 8206
rect 19832 8650 19888 8652
rect 19832 8598 19834 8650
rect 19834 8598 19886 8650
rect 19886 8598 19888 8650
rect 19832 8596 19888 8598
rect 19936 8650 19992 8652
rect 19936 8598 19938 8650
rect 19938 8598 19990 8650
rect 19990 8598 19992 8650
rect 19936 8596 19992 8598
rect 20040 8650 20096 8652
rect 20040 8598 20042 8650
rect 20042 8598 20094 8650
rect 20094 8598 20096 8650
rect 20040 8596 20096 8598
rect 22492 9434 22548 9436
rect 22492 9382 22494 9434
rect 22494 9382 22546 9434
rect 22546 9382 22548 9434
rect 22492 9380 22548 9382
rect 22596 9434 22652 9436
rect 22596 9382 22598 9434
rect 22598 9382 22650 9434
rect 22650 9382 22652 9434
rect 22596 9380 22652 9382
rect 22700 9434 22756 9436
rect 22700 9382 22702 9434
rect 22702 9382 22754 9434
rect 22754 9382 22756 9434
rect 22700 9380 22756 9382
rect 19628 8204 19684 8260
rect 18396 7308 18452 7364
rect 18956 6690 19012 6692
rect 18956 6638 18958 6690
rect 18958 6638 19010 6690
rect 19010 6638 19012 6690
rect 18956 6636 19012 6638
rect 17500 6578 17556 6580
rect 17500 6526 17502 6578
rect 17502 6526 17554 6578
rect 17554 6526 17556 6578
rect 17500 6524 17556 6526
rect 17172 6298 17228 6300
rect 17172 6246 17174 6298
rect 17174 6246 17226 6298
rect 17226 6246 17228 6298
rect 17172 6244 17228 6246
rect 17276 6298 17332 6300
rect 17276 6246 17278 6298
rect 17278 6246 17330 6298
rect 17330 6246 17332 6298
rect 17276 6244 17332 6246
rect 17380 6298 17436 6300
rect 17380 6246 17382 6298
rect 17382 6246 17434 6298
rect 17434 6246 17436 6298
rect 17380 6244 17436 6246
rect 16156 5068 16212 5124
rect 16044 5010 16100 5012
rect 16044 4958 16046 5010
rect 16046 4958 16098 5010
rect 16098 4958 16100 5010
rect 16044 4956 16100 4958
rect 16828 5122 16884 5124
rect 16828 5070 16830 5122
rect 16830 5070 16882 5122
rect 16882 5070 16884 5122
rect 16828 5068 16884 5070
rect 17388 5122 17444 5124
rect 17388 5070 17390 5122
rect 17390 5070 17442 5122
rect 17442 5070 17444 5122
rect 17388 5068 17444 5070
rect 17612 5068 17668 5124
rect 16716 5010 16772 5012
rect 16716 4958 16718 5010
rect 16718 4958 16770 5010
rect 16770 4958 16772 5010
rect 16716 4956 16772 4958
rect 17172 4730 17228 4732
rect 17172 4678 17174 4730
rect 17174 4678 17226 4730
rect 17226 4678 17228 4730
rect 17172 4676 17228 4678
rect 17276 4730 17332 4732
rect 17276 4678 17278 4730
rect 17278 4678 17330 4730
rect 17330 4678 17332 4730
rect 17276 4676 17332 4678
rect 17380 4730 17436 4732
rect 17380 4678 17382 4730
rect 17382 4678 17434 4730
rect 17434 4678 17436 4730
rect 17380 4676 17436 4678
rect 16492 4450 16548 4452
rect 16492 4398 16494 4450
rect 16494 4398 16546 4450
rect 16546 4398 16548 4450
rect 16492 4396 16548 4398
rect 17836 5852 17892 5908
rect 19180 6636 19236 6692
rect 19832 7082 19888 7084
rect 19832 7030 19834 7082
rect 19834 7030 19886 7082
rect 19886 7030 19888 7082
rect 19832 7028 19888 7030
rect 19936 7082 19992 7084
rect 19936 7030 19938 7082
rect 19938 7030 19990 7082
rect 19990 7030 19992 7082
rect 19936 7028 19992 7030
rect 20040 7082 20096 7084
rect 20040 7030 20042 7082
rect 20042 7030 20094 7082
rect 20094 7030 20096 7082
rect 20040 7028 20096 7030
rect 19628 6636 19684 6692
rect 18396 5906 18452 5908
rect 18396 5854 18398 5906
rect 18398 5854 18450 5906
rect 18450 5854 18452 5906
rect 18396 5852 18452 5854
rect 18172 5740 18228 5796
rect 18508 5794 18564 5796
rect 18508 5742 18510 5794
rect 18510 5742 18562 5794
rect 18562 5742 18564 5794
rect 18508 5740 18564 5742
rect 18732 5740 18788 5796
rect 17724 4956 17780 5012
rect 17724 4450 17780 4452
rect 17724 4398 17726 4450
rect 17726 4398 17778 4450
rect 17778 4398 17780 4450
rect 17724 4396 17780 4398
rect 14700 4284 14756 4340
rect 15036 4338 15092 4340
rect 15036 4286 15038 4338
rect 15038 4286 15090 4338
rect 15090 4286 15092 4338
rect 15036 4284 15092 4286
rect 15708 4338 15764 4340
rect 15708 4286 15710 4338
rect 15710 4286 15762 4338
rect 15762 4286 15764 4338
rect 15708 4284 15764 4286
rect 14512 3946 14568 3948
rect 14512 3894 14514 3946
rect 14514 3894 14566 3946
rect 14566 3894 14568 3946
rect 14512 3892 14568 3894
rect 14616 3946 14672 3948
rect 14616 3894 14618 3946
rect 14618 3894 14670 3946
rect 14670 3894 14672 3946
rect 14616 3892 14672 3894
rect 14720 3946 14776 3948
rect 14720 3894 14722 3946
rect 14722 3894 14774 3946
rect 14774 3894 14776 3946
rect 14720 3892 14776 3894
rect 14028 3442 14084 3444
rect 14028 3390 14030 3442
rect 14030 3390 14082 3442
rect 14082 3390 14084 3442
rect 14028 3388 14084 3390
rect 14700 3442 14756 3444
rect 14700 3390 14702 3442
rect 14702 3390 14754 3442
rect 14754 3390 14756 3442
rect 14700 3388 14756 3390
rect 15372 3442 15428 3444
rect 15372 3390 15374 3442
rect 15374 3390 15426 3442
rect 15426 3390 15428 3442
rect 15372 3388 15428 3390
rect 15708 3388 15764 3444
rect 18172 4396 18228 4452
rect 18508 5068 18564 5124
rect 19180 5794 19236 5796
rect 19180 5742 19182 5794
rect 19182 5742 19234 5794
rect 19234 5742 19236 5794
rect 19180 5740 19236 5742
rect 18844 5122 18900 5124
rect 18844 5070 18846 5122
rect 18846 5070 18898 5122
rect 18898 5070 18900 5122
rect 18844 5068 18900 5070
rect 19068 5068 19124 5124
rect 19852 5682 19908 5684
rect 19852 5630 19854 5682
rect 19854 5630 19906 5682
rect 19906 5630 19908 5682
rect 19852 5628 19908 5630
rect 19832 5514 19888 5516
rect 19832 5462 19834 5514
rect 19834 5462 19886 5514
rect 19886 5462 19888 5514
rect 19832 5460 19888 5462
rect 19936 5514 19992 5516
rect 19936 5462 19938 5514
rect 19938 5462 19990 5514
rect 19990 5462 19992 5514
rect 19936 5460 19992 5462
rect 20040 5514 20096 5516
rect 20040 5462 20042 5514
rect 20042 5462 20094 5514
rect 20094 5462 20096 5514
rect 20040 5460 20096 5462
rect 19516 5234 19572 5236
rect 19516 5182 19518 5234
rect 19518 5182 19570 5234
rect 19570 5182 19572 5234
rect 19516 5180 19572 5182
rect 20300 5628 20356 5684
rect 19404 5122 19460 5124
rect 19404 5070 19406 5122
rect 19406 5070 19458 5122
rect 19458 5070 19460 5122
rect 19404 5068 19460 5070
rect 19852 5068 19908 5124
rect 18396 4450 18452 4452
rect 18396 4398 18398 4450
rect 18398 4398 18450 4450
rect 18450 4398 18452 4450
rect 18396 4396 18452 4398
rect 20076 5122 20132 5124
rect 20076 5070 20078 5122
rect 20078 5070 20130 5122
rect 20130 5070 20132 5122
rect 20076 5068 20132 5070
rect 20524 5682 20580 5684
rect 20524 5630 20526 5682
rect 20526 5630 20578 5682
rect 20578 5630 20580 5682
rect 20524 5628 20580 5630
rect 20188 4956 20244 5012
rect 20412 4956 20468 5012
rect 19180 4284 19236 4340
rect 16044 3442 16100 3444
rect 16044 3390 16046 3442
rect 16046 3390 16098 3442
rect 16098 3390 16100 3442
rect 16044 3388 16100 3390
rect 16716 3442 16772 3444
rect 16716 3390 16718 3442
rect 16718 3390 16770 3442
rect 16770 3390 16772 3442
rect 16716 3388 16772 3390
rect 17836 3388 17892 3444
rect 17172 3162 17228 3164
rect 17172 3110 17174 3162
rect 17174 3110 17226 3162
rect 17226 3110 17228 3162
rect 17172 3108 17228 3110
rect 17276 3162 17332 3164
rect 17276 3110 17278 3162
rect 17278 3110 17330 3162
rect 17330 3110 17332 3162
rect 17276 3108 17332 3110
rect 17380 3162 17436 3164
rect 17380 3110 17382 3162
rect 17382 3110 17434 3162
rect 17434 3110 17436 3162
rect 17380 3108 17436 3110
rect 18284 3442 18340 3444
rect 18284 3390 18286 3442
rect 18286 3390 18338 3442
rect 18338 3390 18340 3442
rect 18284 3388 18340 3390
rect 18956 3442 19012 3444
rect 18956 3390 18958 3442
rect 18958 3390 19010 3442
rect 19010 3390 19012 3442
rect 18956 3388 19012 3390
rect 19740 4338 19796 4340
rect 19740 4286 19742 4338
rect 19742 4286 19794 4338
rect 19794 4286 19796 4338
rect 19740 4284 19796 4286
rect 20412 4284 20468 4340
rect 20748 5010 20804 5012
rect 20748 4958 20750 5010
rect 20750 4958 20802 5010
rect 20802 4958 20804 5010
rect 20748 4956 20804 4958
rect 21196 5682 21252 5684
rect 21196 5630 21198 5682
rect 21198 5630 21250 5682
rect 21250 5630 21252 5682
rect 21196 5628 21252 5630
rect 21644 5628 21700 5684
rect 21644 5010 21700 5012
rect 21644 4958 21646 5010
rect 21646 4958 21698 5010
rect 21698 4958 21700 5010
rect 21644 4956 21700 4958
rect 22492 7866 22548 7868
rect 22492 7814 22494 7866
rect 22494 7814 22546 7866
rect 22546 7814 22548 7866
rect 22492 7812 22548 7814
rect 22596 7866 22652 7868
rect 22596 7814 22598 7866
rect 22598 7814 22650 7866
rect 22650 7814 22652 7866
rect 22596 7812 22652 7814
rect 22700 7866 22756 7868
rect 22700 7814 22702 7866
rect 22702 7814 22754 7866
rect 22754 7814 22756 7866
rect 22700 7812 22756 7814
rect 22492 6298 22548 6300
rect 22492 6246 22494 6298
rect 22494 6246 22546 6298
rect 22546 6246 22548 6298
rect 22492 6244 22548 6246
rect 22596 6298 22652 6300
rect 22596 6246 22598 6298
rect 22598 6246 22650 6298
rect 22650 6246 22652 6298
rect 22596 6244 22652 6246
rect 22700 6298 22756 6300
rect 22700 6246 22702 6298
rect 22702 6246 22754 6298
rect 22754 6246 22756 6298
rect 22700 6244 22756 6246
rect 21980 4956 22036 5012
rect 22492 4730 22548 4732
rect 22492 4678 22494 4730
rect 22494 4678 22546 4730
rect 22546 4678 22548 4730
rect 22492 4676 22548 4678
rect 22596 4730 22652 4732
rect 22596 4678 22598 4730
rect 22598 4678 22650 4730
rect 22650 4678 22652 4730
rect 22596 4676 22652 4678
rect 22700 4730 22756 4732
rect 22700 4678 22702 4730
rect 22702 4678 22754 4730
rect 22754 4678 22756 4730
rect 22700 4676 22756 4678
rect 19832 3946 19888 3948
rect 19832 3894 19834 3946
rect 19834 3894 19886 3946
rect 19886 3894 19888 3946
rect 19832 3892 19888 3894
rect 19936 3946 19992 3948
rect 19936 3894 19938 3946
rect 19938 3894 19990 3946
rect 19990 3894 19992 3946
rect 19936 3892 19992 3894
rect 20040 3946 20096 3948
rect 20040 3894 20042 3946
rect 20042 3894 20094 3946
rect 20094 3894 20096 3946
rect 20040 3892 20096 3894
rect 19180 3388 19236 3444
rect 19516 3442 19572 3444
rect 19516 3390 19518 3442
rect 19518 3390 19570 3442
rect 19570 3390 19572 3442
rect 19516 3388 19572 3390
rect 22492 3162 22548 3164
rect 22492 3110 22494 3162
rect 22494 3110 22546 3162
rect 22546 3110 22548 3162
rect 22492 3108 22548 3110
rect 22596 3162 22652 3164
rect 22596 3110 22598 3162
rect 22598 3110 22650 3162
rect 22650 3110 22652 3162
rect 22596 3108 22652 3110
rect 22700 3162 22756 3164
rect 22700 3110 22702 3162
rect 22702 3110 22754 3162
rect 22754 3110 22756 3162
rect 22700 3108 22756 3110
<< metal3 >>
rect 3862 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4146 16492
rect 9182 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9466 16492
rect 14502 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14786 16492
rect 19822 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20106 16492
rect 6522 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6806 15708
rect 11842 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12126 15708
rect 17162 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17446 15708
rect 22482 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22766 15708
rect 0 14980 800 15008
rect 23200 14980 24000 15008
rect 0 14924 3612 14980
rect 3668 14924 3678 14980
rect 21644 14924 24000 14980
rect 0 14896 800 14924
rect 3862 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4146 14924
rect 9182 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9466 14924
rect 14502 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14786 14924
rect 19822 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20106 14924
rect 21644 14756 21700 14924
rect 23200 14896 24000 14924
rect 19618 14700 19628 14756
rect 19684 14700 21700 14756
rect 6522 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6806 14140
rect 11842 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12126 14140
rect 17162 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17446 14140
rect 22482 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22766 14140
rect 16258 13468 16268 13524
rect 16324 13468 16940 13524
rect 16996 13468 17388 13524
rect 17444 13468 17612 13524
rect 17668 13468 18396 13524
rect 18452 13468 18462 13524
rect 18946 13468 18956 13524
rect 19012 13468 19628 13524
rect 19684 13468 19694 13524
rect 3862 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4146 13356
rect 9182 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9466 13356
rect 14502 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14786 13356
rect 19822 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20106 13356
rect 18498 13244 18508 13300
rect 18564 13244 18574 13300
rect 18508 13188 18564 13244
rect 14914 13132 14924 13188
rect 14980 13132 17052 13188
rect 17108 13132 17724 13188
rect 17780 13132 18284 13188
rect 18340 13132 18844 13188
rect 18900 13132 19180 13188
rect 19236 13132 19246 13188
rect 6522 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6806 12572
rect 11842 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12126 12572
rect 17162 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17446 12572
rect 22482 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22766 12572
rect 18386 12236 18396 12292
rect 18452 12236 18956 12292
rect 19012 12236 19022 12292
rect 19730 12236 19740 12292
rect 19796 12236 20412 12292
rect 20468 12236 21084 12292
rect 21140 12236 21150 12292
rect 14802 12124 14812 12180
rect 14868 12124 15484 12180
rect 15540 12124 15550 12180
rect 16146 12124 16156 12180
rect 16212 12124 16828 12180
rect 16884 12124 16894 12180
rect 14242 11900 14252 11956
rect 14308 11900 14924 11956
rect 14980 11900 14990 11956
rect 17602 11788 17612 11844
rect 17668 11788 17678 11844
rect 3862 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4146 11788
rect 9182 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9466 11788
rect 14502 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14786 11788
rect 17612 11732 17668 11788
rect 19822 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20106 11788
rect 17612 11676 18508 11732
rect 18564 11676 18574 11732
rect 14914 11340 14924 11396
rect 14980 11340 15596 11396
rect 15652 11340 16268 11396
rect 16324 11340 16940 11396
rect 16996 11340 17500 11396
rect 17556 11340 17566 11396
rect 18946 11340 18956 11396
rect 19012 11340 19516 11396
rect 19572 11340 19852 11396
rect 19908 11340 19918 11396
rect 6178 11228 6188 11284
rect 6244 11228 6972 11284
rect 7028 11228 7038 11284
rect 18274 11116 18284 11172
rect 18340 11116 18508 11172
rect 18564 11116 18956 11172
rect 19012 11116 21756 11172
rect 21812 11116 21822 11172
rect 6522 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6806 11004
rect 11842 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12126 11004
rect 17162 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17446 11004
rect 22482 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22766 11004
rect 5506 10668 5516 10724
rect 5572 10668 6076 10724
rect 6132 10668 6142 10724
rect 19842 10668 19852 10724
rect 19908 10668 20188 10724
rect 20244 10668 20254 10724
rect 21074 10668 21084 10724
rect 21140 10668 21868 10724
rect 21924 10668 21934 10724
rect 16818 10332 16828 10388
rect 16884 10332 17836 10388
rect 17892 10332 18284 10388
rect 18340 10332 18508 10388
rect 18564 10332 18574 10388
rect 3862 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4146 10220
rect 9182 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9466 10220
rect 14502 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14786 10220
rect 19822 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20106 10220
rect 9986 10108 9996 10164
rect 10052 10108 10062 10164
rect 9996 10052 10052 10108
rect 8978 9996 8988 10052
rect 9044 9996 11340 10052
rect 11396 9996 12012 10052
rect 12068 9996 12078 10052
rect 19842 9996 19852 10052
rect 19908 9996 20524 10052
rect 20580 9996 20590 10052
rect 4274 9772 4284 9828
rect 4340 9772 4844 9828
rect 4900 9772 5404 9828
rect 5460 9772 5470 9828
rect 5842 9660 5852 9716
rect 5908 9660 6524 9716
rect 6580 9660 7196 9716
rect 7252 9660 7262 9716
rect 8988 9604 9044 9996
rect 8642 9548 8652 9604
rect 8708 9548 9324 9604
rect 9380 9548 9390 9604
rect 16482 9548 16492 9604
rect 16548 9548 17164 9604
rect 17220 9548 17230 9604
rect 19170 9548 19180 9604
rect 19236 9548 19852 9604
rect 19908 9548 19918 9604
rect 6522 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6806 9436
rect 11842 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12126 9436
rect 17162 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17446 9436
rect 22482 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22766 9436
rect 3490 9100 3500 9156
rect 3556 9100 4060 9156
rect 4116 9100 4126 9156
rect 14354 8988 14364 9044
rect 14420 8988 15036 9044
rect 15092 8988 15260 9044
rect 15316 8988 15326 9044
rect 18946 8764 18956 8820
rect 19012 8764 19180 8820
rect 19236 8764 19246 8820
rect 3862 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4146 8652
rect 9182 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9466 8652
rect 14502 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14786 8652
rect 19822 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20106 8652
rect 9986 8540 9996 8596
rect 10052 8540 10556 8596
rect 10612 8540 10622 8596
rect 3602 8428 3612 8484
rect 3668 8428 4172 8484
rect 4228 8428 4732 8484
rect 4788 8428 4956 8484
rect 5012 8428 5404 8484
rect 5460 8428 5964 8484
rect 6020 8428 6524 8484
rect 6580 8428 6590 8484
rect 7186 8428 7196 8484
rect 7252 8428 7980 8484
rect 8036 8428 8540 8484
rect 8596 8428 9324 8484
rect 9380 8428 9390 8484
rect 12786 8428 12796 8484
rect 12852 8428 13692 8484
rect 13748 8428 13916 8484
rect 13972 8428 14364 8484
rect 14420 8428 15148 8484
rect 15204 8428 15708 8484
rect 15764 8428 16380 8484
rect 16436 8428 17164 8484
rect 17220 8428 17836 8484
rect 17892 8428 18508 8484
rect 18564 8428 18956 8484
rect 19012 8428 19022 8484
rect 8978 8316 8988 8372
rect 9044 8316 9884 8372
rect 9940 8316 10332 8372
rect 10388 8316 10398 8372
rect 18386 8316 18396 8372
rect 18452 8316 19180 8372
rect 19236 8316 19246 8372
rect 9202 8204 9212 8260
rect 9268 8204 9996 8260
rect 10052 8204 10062 8260
rect 12450 8204 12460 8260
rect 12516 8204 12908 8260
rect 12964 8204 13356 8260
rect 13412 8204 13804 8260
rect 13860 8204 14476 8260
rect 14532 8204 15036 8260
rect 15092 8204 15596 8260
rect 15652 8204 15820 8260
rect 15876 8204 16268 8260
rect 16324 8204 16492 8260
rect 16548 8204 17052 8260
rect 17108 8204 17612 8260
rect 17668 8204 19068 8260
rect 19124 8204 19628 8260
rect 19684 8204 19694 8260
rect 4274 7980 4284 8036
rect 4340 7980 4844 8036
rect 4900 7980 4910 8036
rect 7298 7980 7308 8036
rect 7364 7980 7980 8036
rect 8036 7980 8316 8036
rect 8372 7980 8382 8036
rect 6522 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6806 7868
rect 11842 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12126 7868
rect 17162 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17446 7868
rect 22482 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22766 7868
rect 17826 7644 17836 7700
rect 17892 7644 18396 7700
rect 18452 7644 18462 7700
rect 2146 7420 2156 7476
rect 2212 7420 2716 7476
rect 2772 7420 2782 7476
rect 4834 7420 4844 7476
rect 4900 7420 5404 7476
rect 5460 7420 6076 7476
rect 6132 7420 6142 7476
rect 6738 7420 6748 7476
rect 6804 7420 7308 7476
rect 7364 7420 7374 7476
rect 16594 7420 16604 7476
rect 16660 7420 17612 7476
rect 17668 7420 17678 7476
rect 17714 7308 17724 7364
rect 17780 7308 18396 7364
rect 18452 7308 18462 7364
rect 3602 7196 3612 7252
rect 3668 7196 4172 7252
rect 4228 7196 4238 7252
rect 3862 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4146 7084
rect 9182 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9466 7084
rect 14502 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14786 7084
rect 19822 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20106 7084
rect 7522 6860 7532 6916
rect 7588 6860 8876 6916
rect 8932 6860 9996 6916
rect 10052 6860 10062 6916
rect 10546 6860 10556 6916
rect 10612 6860 11228 6916
rect 11284 6860 12012 6916
rect 12068 6860 12078 6916
rect 14018 6860 14028 6916
rect 14084 6860 14252 6916
rect 14308 6860 14588 6916
rect 14644 6860 15260 6916
rect 15316 6860 15326 6916
rect 2818 6748 2828 6804
rect 2884 6748 3724 6804
rect 3780 6748 4620 6804
rect 4676 6748 5516 6804
rect 5572 6748 5740 6804
rect 5796 6748 6412 6804
rect 6468 6748 6478 6804
rect 8530 6636 8540 6692
rect 8596 6636 8764 6692
rect 8820 6636 9212 6692
rect 9268 6636 9884 6692
rect 9940 6636 10444 6692
rect 10500 6636 11116 6692
rect 11172 6636 11900 6692
rect 11956 6636 12460 6692
rect 12516 6636 12526 6692
rect 18946 6636 18956 6692
rect 19012 6636 19180 6692
rect 19236 6636 19628 6692
rect 19684 6636 19694 6692
rect 2146 6524 2156 6580
rect 2212 6524 2828 6580
rect 2884 6524 3388 6580
rect 3444 6524 3454 6580
rect 8418 6524 8428 6580
rect 8484 6524 9100 6580
rect 9156 6524 9166 6580
rect 16930 6524 16940 6580
rect 16996 6524 17500 6580
rect 17556 6524 17566 6580
rect 9874 6412 9884 6468
rect 9940 6412 10556 6468
rect 10612 6412 10622 6468
rect 6522 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6806 6300
rect 11842 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12126 6300
rect 17162 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17446 6300
rect 22482 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22766 6300
rect 7074 5964 7084 6020
rect 7140 5964 7420 6020
rect 7476 5964 7756 6020
rect 7812 5964 8092 6020
rect 8148 5964 8158 6020
rect 4050 5852 4060 5908
rect 4116 5852 4732 5908
rect 4788 5852 4798 5908
rect 9090 5852 9100 5908
rect 9156 5852 9772 5908
rect 9828 5852 10444 5908
rect 10500 5852 10510 5908
rect 17826 5852 17836 5908
rect 17892 5852 18396 5908
rect 18452 5852 18462 5908
rect 18162 5740 18172 5796
rect 18228 5740 18508 5796
rect 18564 5740 18732 5796
rect 18788 5740 19180 5796
rect 19236 5740 19246 5796
rect 19842 5628 19852 5684
rect 19908 5628 20300 5684
rect 20356 5628 20524 5684
rect 20580 5628 21196 5684
rect 21252 5628 21644 5684
rect 21700 5628 21710 5684
rect 3862 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4146 5516
rect 9182 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9466 5516
rect 14502 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14786 5516
rect 19822 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20106 5516
rect 18844 5180 19516 5236
rect 19572 5180 19582 5236
rect 18844 5124 18900 5180
rect 2706 5068 2716 5124
rect 2772 5068 2782 5124
rect 3378 5068 3388 5124
rect 3444 5068 4172 5124
rect 4228 5068 4956 5124
rect 5012 5068 5022 5124
rect 7298 5068 7308 5124
rect 7364 5068 7756 5124
rect 7812 5068 8540 5124
rect 8596 5068 9100 5124
rect 9156 5068 9660 5124
rect 9716 5068 9726 5124
rect 11554 5068 11564 5124
rect 11620 5068 12124 5124
rect 12180 5068 12190 5124
rect 16146 5068 16156 5124
rect 16212 5068 16828 5124
rect 16884 5068 17388 5124
rect 17444 5068 17454 5124
rect 17602 5068 17612 5124
rect 17668 5068 18508 5124
rect 18564 5068 18844 5124
rect 18900 5068 18910 5124
rect 19058 5068 19068 5124
rect 19124 5068 19404 5124
rect 19460 5068 19852 5124
rect 19908 5068 20076 5124
rect 20132 5068 20142 5124
rect 0 5012 800 5040
rect 2716 5012 2772 5068
rect 23200 5012 24000 5040
rect 0 4956 3612 5012
rect 3668 4956 3678 5012
rect 14690 4956 14700 5012
rect 14756 4956 16044 5012
rect 16100 4956 16716 5012
rect 16772 4956 17724 5012
rect 17780 4956 17790 5012
rect 20178 4956 20188 5012
rect 20244 4956 20412 5012
rect 20468 4956 20748 5012
rect 20804 4956 21644 5012
rect 21700 4956 21710 5012
rect 21970 4956 21980 5012
rect 22036 4956 24000 5012
rect 0 4928 800 4956
rect 23200 4928 24000 4956
rect 4722 4844 4732 4900
rect 4788 4844 4956 4900
rect 5012 4844 5404 4900
rect 5460 4844 5852 4900
rect 5908 4844 6076 4900
rect 6132 4844 6142 4900
rect 12338 4844 12348 4900
rect 12404 4844 12908 4900
rect 12964 4844 12974 4900
rect 6522 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6806 4732
rect 11842 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12126 4732
rect 17162 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17446 4732
rect 22482 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22766 4732
rect 3826 4508 3836 4564
rect 3892 4508 4508 4564
rect 4564 4508 4844 4564
rect 4900 4508 5740 4564
rect 5796 4508 6300 4564
rect 6356 4508 6366 4564
rect 2370 4396 2380 4452
rect 2436 4396 3052 4452
rect 3108 4396 3118 4452
rect 16482 4396 16492 4452
rect 16548 4396 17724 4452
rect 17780 4396 18172 4452
rect 18228 4396 18396 4452
rect 18452 4396 18462 4452
rect 2482 4284 2492 4340
rect 2548 4284 2828 4340
rect 2884 4284 3164 4340
rect 3220 4284 3500 4340
rect 3556 4284 3724 4340
rect 3780 4284 4396 4340
rect 4452 4284 4462 4340
rect 7074 4284 7084 4340
rect 7140 4284 7756 4340
rect 7812 4284 7822 4340
rect 14466 4284 14476 4340
rect 14532 4284 14700 4340
rect 14756 4284 15036 4340
rect 15092 4284 15708 4340
rect 15764 4284 15774 4340
rect 19170 4284 19180 4340
rect 19236 4284 19740 4340
rect 19796 4284 20412 4340
rect 20468 4284 20478 4340
rect 4274 4060 4284 4116
rect 4340 4060 5852 4116
rect 5908 4060 6076 4116
rect 6132 4060 6524 4116
rect 6580 4060 7084 4116
rect 7140 4060 7150 4116
rect 12450 4060 12460 4116
rect 12516 4060 13132 4116
rect 13188 4060 13804 4116
rect 13860 4060 13870 4116
rect 3862 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4146 3948
rect 9182 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9466 3948
rect 14502 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14786 3948
rect 19822 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20106 3948
rect 2146 3500 2156 3556
rect 2212 3500 2828 3556
rect 2884 3500 2894 3556
rect 3042 3500 3052 3556
rect 3108 3500 3500 3556
rect 3556 3500 4172 3556
rect 4228 3500 4238 3556
rect 7074 3500 7084 3556
rect 7140 3500 7756 3556
rect 7812 3500 8428 3556
rect 8484 3500 9660 3556
rect 9716 3500 9884 3556
rect 9940 3500 10332 3556
rect 10388 3500 11116 3556
rect 11172 3500 11676 3556
rect 11732 3500 11742 3556
rect 4386 3388 4396 3444
rect 4452 3388 4844 3444
rect 4900 3388 5180 3444
rect 5236 3388 5740 3444
rect 5796 3388 6636 3444
rect 6692 3388 11004 3444
rect 11060 3388 11788 3444
rect 11844 3388 11854 3444
rect 14018 3388 14028 3444
rect 14084 3388 14700 3444
rect 14756 3388 15372 3444
rect 15428 3388 15708 3444
rect 15764 3388 16044 3444
rect 16100 3388 16716 3444
rect 16772 3388 17836 3444
rect 17892 3388 18284 3444
rect 18340 3388 18956 3444
rect 19012 3388 19180 3444
rect 19236 3388 19516 3444
rect 19572 3388 19582 3444
rect 6522 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6806 3164
rect 11842 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12126 3164
rect 17162 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17446 3164
rect 22482 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22766 3164
<< via3 >>
rect 3872 16436 3928 16492
rect 3976 16436 4032 16492
rect 4080 16436 4136 16492
rect 9192 16436 9248 16492
rect 9296 16436 9352 16492
rect 9400 16436 9456 16492
rect 14512 16436 14568 16492
rect 14616 16436 14672 16492
rect 14720 16436 14776 16492
rect 19832 16436 19888 16492
rect 19936 16436 19992 16492
rect 20040 16436 20096 16492
rect 6532 15652 6588 15708
rect 6636 15652 6692 15708
rect 6740 15652 6796 15708
rect 11852 15652 11908 15708
rect 11956 15652 12012 15708
rect 12060 15652 12116 15708
rect 17172 15652 17228 15708
rect 17276 15652 17332 15708
rect 17380 15652 17436 15708
rect 22492 15652 22548 15708
rect 22596 15652 22652 15708
rect 22700 15652 22756 15708
rect 3872 14868 3928 14924
rect 3976 14868 4032 14924
rect 4080 14868 4136 14924
rect 9192 14868 9248 14924
rect 9296 14868 9352 14924
rect 9400 14868 9456 14924
rect 14512 14868 14568 14924
rect 14616 14868 14672 14924
rect 14720 14868 14776 14924
rect 19832 14868 19888 14924
rect 19936 14868 19992 14924
rect 20040 14868 20096 14924
rect 6532 14084 6588 14140
rect 6636 14084 6692 14140
rect 6740 14084 6796 14140
rect 11852 14084 11908 14140
rect 11956 14084 12012 14140
rect 12060 14084 12116 14140
rect 17172 14084 17228 14140
rect 17276 14084 17332 14140
rect 17380 14084 17436 14140
rect 22492 14084 22548 14140
rect 22596 14084 22652 14140
rect 22700 14084 22756 14140
rect 3872 13300 3928 13356
rect 3976 13300 4032 13356
rect 4080 13300 4136 13356
rect 9192 13300 9248 13356
rect 9296 13300 9352 13356
rect 9400 13300 9456 13356
rect 14512 13300 14568 13356
rect 14616 13300 14672 13356
rect 14720 13300 14776 13356
rect 19832 13300 19888 13356
rect 19936 13300 19992 13356
rect 20040 13300 20096 13356
rect 6532 12516 6588 12572
rect 6636 12516 6692 12572
rect 6740 12516 6796 12572
rect 11852 12516 11908 12572
rect 11956 12516 12012 12572
rect 12060 12516 12116 12572
rect 17172 12516 17228 12572
rect 17276 12516 17332 12572
rect 17380 12516 17436 12572
rect 22492 12516 22548 12572
rect 22596 12516 22652 12572
rect 22700 12516 22756 12572
rect 3872 11732 3928 11788
rect 3976 11732 4032 11788
rect 4080 11732 4136 11788
rect 9192 11732 9248 11788
rect 9296 11732 9352 11788
rect 9400 11732 9456 11788
rect 14512 11732 14568 11788
rect 14616 11732 14672 11788
rect 14720 11732 14776 11788
rect 19832 11732 19888 11788
rect 19936 11732 19992 11788
rect 20040 11732 20096 11788
rect 6532 10948 6588 11004
rect 6636 10948 6692 11004
rect 6740 10948 6796 11004
rect 11852 10948 11908 11004
rect 11956 10948 12012 11004
rect 12060 10948 12116 11004
rect 17172 10948 17228 11004
rect 17276 10948 17332 11004
rect 17380 10948 17436 11004
rect 22492 10948 22548 11004
rect 22596 10948 22652 11004
rect 22700 10948 22756 11004
rect 3872 10164 3928 10220
rect 3976 10164 4032 10220
rect 4080 10164 4136 10220
rect 9192 10164 9248 10220
rect 9296 10164 9352 10220
rect 9400 10164 9456 10220
rect 14512 10164 14568 10220
rect 14616 10164 14672 10220
rect 14720 10164 14776 10220
rect 19832 10164 19888 10220
rect 19936 10164 19992 10220
rect 20040 10164 20096 10220
rect 6532 9380 6588 9436
rect 6636 9380 6692 9436
rect 6740 9380 6796 9436
rect 11852 9380 11908 9436
rect 11956 9380 12012 9436
rect 12060 9380 12116 9436
rect 17172 9380 17228 9436
rect 17276 9380 17332 9436
rect 17380 9380 17436 9436
rect 22492 9380 22548 9436
rect 22596 9380 22652 9436
rect 22700 9380 22756 9436
rect 3872 8596 3928 8652
rect 3976 8596 4032 8652
rect 4080 8596 4136 8652
rect 9192 8596 9248 8652
rect 9296 8596 9352 8652
rect 9400 8596 9456 8652
rect 14512 8596 14568 8652
rect 14616 8596 14672 8652
rect 14720 8596 14776 8652
rect 19832 8596 19888 8652
rect 19936 8596 19992 8652
rect 20040 8596 20096 8652
rect 6532 7812 6588 7868
rect 6636 7812 6692 7868
rect 6740 7812 6796 7868
rect 11852 7812 11908 7868
rect 11956 7812 12012 7868
rect 12060 7812 12116 7868
rect 17172 7812 17228 7868
rect 17276 7812 17332 7868
rect 17380 7812 17436 7868
rect 22492 7812 22548 7868
rect 22596 7812 22652 7868
rect 22700 7812 22756 7868
rect 3872 7028 3928 7084
rect 3976 7028 4032 7084
rect 4080 7028 4136 7084
rect 9192 7028 9248 7084
rect 9296 7028 9352 7084
rect 9400 7028 9456 7084
rect 14512 7028 14568 7084
rect 14616 7028 14672 7084
rect 14720 7028 14776 7084
rect 19832 7028 19888 7084
rect 19936 7028 19992 7084
rect 20040 7028 20096 7084
rect 6532 6244 6588 6300
rect 6636 6244 6692 6300
rect 6740 6244 6796 6300
rect 11852 6244 11908 6300
rect 11956 6244 12012 6300
rect 12060 6244 12116 6300
rect 17172 6244 17228 6300
rect 17276 6244 17332 6300
rect 17380 6244 17436 6300
rect 22492 6244 22548 6300
rect 22596 6244 22652 6300
rect 22700 6244 22756 6300
rect 3872 5460 3928 5516
rect 3976 5460 4032 5516
rect 4080 5460 4136 5516
rect 9192 5460 9248 5516
rect 9296 5460 9352 5516
rect 9400 5460 9456 5516
rect 14512 5460 14568 5516
rect 14616 5460 14672 5516
rect 14720 5460 14776 5516
rect 19832 5460 19888 5516
rect 19936 5460 19992 5516
rect 20040 5460 20096 5516
rect 6532 4676 6588 4732
rect 6636 4676 6692 4732
rect 6740 4676 6796 4732
rect 11852 4676 11908 4732
rect 11956 4676 12012 4732
rect 12060 4676 12116 4732
rect 17172 4676 17228 4732
rect 17276 4676 17332 4732
rect 17380 4676 17436 4732
rect 22492 4676 22548 4732
rect 22596 4676 22652 4732
rect 22700 4676 22756 4732
rect 3872 3892 3928 3948
rect 3976 3892 4032 3948
rect 4080 3892 4136 3948
rect 9192 3892 9248 3948
rect 9296 3892 9352 3948
rect 9400 3892 9456 3948
rect 14512 3892 14568 3948
rect 14616 3892 14672 3948
rect 14720 3892 14776 3948
rect 19832 3892 19888 3948
rect 19936 3892 19992 3948
rect 20040 3892 20096 3948
rect 6532 3108 6588 3164
rect 6636 3108 6692 3164
rect 6740 3108 6796 3164
rect 11852 3108 11908 3164
rect 11956 3108 12012 3164
rect 12060 3108 12116 3164
rect 17172 3108 17228 3164
rect 17276 3108 17332 3164
rect 17380 3108 17436 3164
rect 22492 3108 22548 3164
rect 22596 3108 22652 3164
rect 22700 3108 22756 3164
<< metal4 >>
rect 3844 16492 4164 16524
rect 3844 16436 3872 16492
rect 3928 16436 3976 16492
rect 4032 16436 4080 16492
rect 4136 16436 4164 16492
rect 3844 14924 4164 16436
rect 3844 14868 3872 14924
rect 3928 14868 3976 14924
rect 4032 14868 4080 14924
rect 4136 14868 4164 14924
rect 3844 13356 4164 14868
rect 3844 13300 3872 13356
rect 3928 13300 3976 13356
rect 4032 13300 4080 13356
rect 4136 13300 4164 13356
rect 3844 11788 4164 13300
rect 3844 11732 3872 11788
rect 3928 11732 3976 11788
rect 4032 11732 4080 11788
rect 4136 11732 4164 11788
rect 3844 10220 4164 11732
rect 3844 10164 3872 10220
rect 3928 10164 3976 10220
rect 4032 10164 4080 10220
rect 4136 10164 4164 10220
rect 3844 8652 4164 10164
rect 3844 8596 3872 8652
rect 3928 8596 3976 8652
rect 4032 8596 4080 8652
rect 4136 8596 4164 8652
rect 3844 7084 4164 8596
rect 3844 7028 3872 7084
rect 3928 7028 3976 7084
rect 4032 7028 4080 7084
rect 4136 7028 4164 7084
rect 3844 5516 4164 7028
rect 3844 5460 3872 5516
rect 3928 5460 3976 5516
rect 4032 5460 4080 5516
rect 4136 5460 4164 5516
rect 3844 3948 4164 5460
rect 3844 3892 3872 3948
rect 3928 3892 3976 3948
rect 4032 3892 4080 3948
rect 4136 3892 4164 3948
rect 3844 3076 4164 3892
rect 6504 15708 6824 16524
rect 6504 15652 6532 15708
rect 6588 15652 6636 15708
rect 6692 15652 6740 15708
rect 6796 15652 6824 15708
rect 6504 14140 6824 15652
rect 6504 14084 6532 14140
rect 6588 14084 6636 14140
rect 6692 14084 6740 14140
rect 6796 14084 6824 14140
rect 6504 12572 6824 14084
rect 6504 12516 6532 12572
rect 6588 12516 6636 12572
rect 6692 12516 6740 12572
rect 6796 12516 6824 12572
rect 6504 11004 6824 12516
rect 6504 10948 6532 11004
rect 6588 10948 6636 11004
rect 6692 10948 6740 11004
rect 6796 10948 6824 11004
rect 6504 9436 6824 10948
rect 6504 9380 6532 9436
rect 6588 9380 6636 9436
rect 6692 9380 6740 9436
rect 6796 9380 6824 9436
rect 6504 7868 6824 9380
rect 6504 7812 6532 7868
rect 6588 7812 6636 7868
rect 6692 7812 6740 7868
rect 6796 7812 6824 7868
rect 6504 6300 6824 7812
rect 6504 6244 6532 6300
rect 6588 6244 6636 6300
rect 6692 6244 6740 6300
rect 6796 6244 6824 6300
rect 6504 4732 6824 6244
rect 6504 4676 6532 4732
rect 6588 4676 6636 4732
rect 6692 4676 6740 4732
rect 6796 4676 6824 4732
rect 6504 3164 6824 4676
rect 6504 3108 6532 3164
rect 6588 3108 6636 3164
rect 6692 3108 6740 3164
rect 6796 3108 6824 3164
rect 6504 3076 6824 3108
rect 9164 16492 9484 16524
rect 9164 16436 9192 16492
rect 9248 16436 9296 16492
rect 9352 16436 9400 16492
rect 9456 16436 9484 16492
rect 9164 14924 9484 16436
rect 9164 14868 9192 14924
rect 9248 14868 9296 14924
rect 9352 14868 9400 14924
rect 9456 14868 9484 14924
rect 9164 13356 9484 14868
rect 9164 13300 9192 13356
rect 9248 13300 9296 13356
rect 9352 13300 9400 13356
rect 9456 13300 9484 13356
rect 9164 11788 9484 13300
rect 9164 11732 9192 11788
rect 9248 11732 9296 11788
rect 9352 11732 9400 11788
rect 9456 11732 9484 11788
rect 9164 10220 9484 11732
rect 9164 10164 9192 10220
rect 9248 10164 9296 10220
rect 9352 10164 9400 10220
rect 9456 10164 9484 10220
rect 9164 8652 9484 10164
rect 9164 8596 9192 8652
rect 9248 8596 9296 8652
rect 9352 8596 9400 8652
rect 9456 8596 9484 8652
rect 9164 7084 9484 8596
rect 9164 7028 9192 7084
rect 9248 7028 9296 7084
rect 9352 7028 9400 7084
rect 9456 7028 9484 7084
rect 9164 5516 9484 7028
rect 9164 5460 9192 5516
rect 9248 5460 9296 5516
rect 9352 5460 9400 5516
rect 9456 5460 9484 5516
rect 9164 3948 9484 5460
rect 9164 3892 9192 3948
rect 9248 3892 9296 3948
rect 9352 3892 9400 3948
rect 9456 3892 9484 3948
rect 9164 3076 9484 3892
rect 11824 15708 12144 16524
rect 11824 15652 11852 15708
rect 11908 15652 11956 15708
rect 12012 15652 12060 15708
rect 12116 15652 12144 15708
rect 11824 14140 12144 15652
rect 11824 14084 11852 14140
rect 11908 14084 11956 14140
rect 12012 14084 12060 14140
rect 12116 14084 12144 14140
rect 11824 12572 12144 14084
rect 11824 12516 11852 12572
rect 11908 12516 11956 12572
rect 12012 12516 12060 12572
rect 12116 12516 12144 12572
rect 11824 11004 12144 12516
rect 11824 10948 11852 11004
rect 11908 10948 11956 11004
rect 12012 10948 12060 11004
rect 12116 10948 12144 11004
rect 11824 9436 12144 10948
rect 11824 9380 11852 9436
rect 11908 9380 11956 9436
rect 12012 9380 12060 9436
rect 12116 9380 12144 9436
rect 11824 7868 12144 9380
rect 11824 7812 11852 7868
rect 11908 7812 11956 7868
rect 12012 7812 12060 7868
rect 12116 7812 12144 7868
rect 11824 6300 12144 7812
rect 11824 6244 11852 6300
rect 11908 6244 11956 6300
rect 12012 6244 12060 6300
rect 12116 6244 12144 6300
rect 11824 4732 12144 6244
rect 11824 4676 11852 4732
rect 11908 4676 11956 4732
rect 12012 4676 12060 4732
rect 12116 4676 12144 4732
rect 11824 3164 12144 4676
rect 11824 3108 11852 3164
rect 11908 3108 11956 3164
rect 12012 3108 12060 3164
rect 12116 3108 12144 3164
rect 11824 3076 12144 3108
rect 14484 16492 14804 16524
rect 14484 16436 14512 16492
rect 14568 16436 14616 16492
rect 14672 16436 14720 16492
rect 14776 16436 14804 16492
rect 14484 14924 14804 16436
rect 14484 14868 14512 14924
rect 14568 14868 14616 14924
rect 14672 14868 14720 14924
rect 14776 14868 14804 14924
rect 14484 13356 14804 14868
rect 14484 13300 14512 13356
rect 14568 13300 14616 13356
rect 14672 13300 14720 13356
rect 14776 13300 14804 13356
rect 14484 11788 14804 13300
rect 14484 11732 14512 11788
rect 14568 11732 14616 11788
rect 14672 11732 14720 11788
rect 14776 11732 14804 11788
rect 14484 10220 14804 11732
rect 14484 10164 14512 10220
rect 14568 10164 14616 10220
rect 14672 10164 14720 10220
rect 14776 10164 14804 10220
rect 14484 8652 14804 10164
rect 14484 8596 14512 8652
rect 14568 8596 14616 8652
rect 14672 8596 14720 8652
rect 14776 8596 14804 8652
rect 14484 7084 14804 8596
rect 14484 7028 14512 7084
rect 14568 7028 14616 7084
rect 14672 7028 14720 7084
rect 14776 7028 14804 7084
rect 14484 5516 14804 7028
rect 14484 5460 14512 5516
rect 14568 5460 14616 5516
rect 14672 5460 14720 5516
rect 14776 5460 14804 5516
rect 14484 3948 14804 5460
rect 14484 3892 14512 3948
rect 14568 3892 14616 3948
rect 14672 3892 14720 3948
rect 14776 3892 14804 3948
rect 14484 3076 14804 3892
rect 17144 15708 17464 16524
rect 17144 15652 17172 15708
rect 17228 15652 17276 15708
rect 17332 15652 17380 15708
rect 17436 15652 17464 15708
rect 17144 14140 17464 15652
rect 17144 14084 17172 14140
rect 17228 14084 17276 14140
rect 17332 14084 17380 14140
rect 17436 14084 17464 14140
rect 17144 12572 17464 14084
rect 17144 12516 17172 12572
rect 17228 12516 17276 12572
rect 17332 12516 17380 12572
rect 17436 12516 17464 12572
rect 17144 11004 17464 12516
rect 17144 10948 17172 11004
rect 17228 10948 17276 11004
rect 17332 10948 17380 11004
rect 17436 10948 17464 11004
rect 17144 9436 17464 10948
rect 17144 9380 17172 9436
rect 17228 9380 17276 9436
rect 17332 9380 17380 9436
rect 17436 9380 17464 9436
rect 17144 7868 17464 9380
rect 17144 7812 17172 7868
rect 17228 7812 17276 7868
rect 17332 7812 17380 7868
rect 17436 7812 17464 7868
rect 17144 6300 17464 7812
rect 17144 6244 17172 6300
rect 17228 6244 17276 6300
rect 17332 6244 17380 6300
rect 17436 6244 17464 6300
rect 17144 4732 17464 6244
rect 17144 4676 17172 4732
rect 17228 4676 17276 4732
rect 17332 4676 17380 4732
rect 17436 4676 17464 4732
rect 17144 3164 17464 4676
rect 17144 3108 17172 3164
rect 17228 3108 17276 3164
rect 17332 3108 17380 3164
rect 17436 3108 17464 3164
rect 17144 3076 17464 3108
rect 19804 16492 20124 16524
rect 19804 16436 19832 16492
rect 19888 16436 19936 16492
rect 19992 16436 20040 16492
rect 20096 16436 20124 16492
rect 19804 14924 20124 16436
rect 19804 14868 19832 14924
rect 19888 14868 19936 14924
rect 19992 14868 20040 14924
rect 20096 14868 20124 14924
rect 19804 13356 20124 14868
rect 19804 13300 19832 13356
rect 19888 13300 19936 13356
rect 19992 13300 20040 13356
rect 20096 13300 20124 13356
rect 19804 11788 20124 13300
rect 19804 11732 19832 11788
rect 19888 11732 19936 11788
rect 19992 11732 20040 11788
rect 20096 11732 20124 11788
rect 19804 10220 20124 11732
rect 19804 10164 19832 10220
rect 19888 10164 19936 10220
rect 19992 10164 20040 10220
rect 20096 10164 20124 10220
rect 19804 8652 20124 10164
rect 19804 8596 19832 8652
rect 19888 8596 19936 8652
rect 19992 8596 20040 8652
rect 20096 8596 20124 8652
rect 19804 7084 20124 8596
rect 19804 7028 19832 7084
rect 19888 7028 19936 7084
rect 19992 7028 20040 7084
rect 20096 7028 20124 7084
rect 19804 5516 20124 7028
rect 19804 5460 19832 5516
rect 19888 5460 19936 5516
rect 19992 5460 20040 5516
rect 20096 5460 20124 5516
rect 19804 3948 20124 5460
rect 19804 3892 19832 3948
rect 19888 3892 19936 3948
rect 19992 3892 20040 3948
rect 20096 3892 20124 3948
rect 19804 3076 20124 3892
rect 22464 15708 22784 16524
rect 22464 15652 22492 15708
rect 22548 15652 22596 15708
rect 22652 15652 22700 15708
rect 22756 15652 22784 15708
rect 22464 14140 22784 15652
rect 22464 14084 22492 14140
rect 22548 14084 22596 14140
rect 22652 14084 22700 14140
rect 22756 14084 22784 14140
rect 22464 12572 22784 14084
rect 22464 12516 22492 12572
rect 22548 12516 22596 12572
rect 22652 12516 22700 12572
rect 22756 12516 22784 12572
rect 22464 11004 22784 12516
rect 22464 10948 22492 11004
rect 22548 10948 22596 11004
rect 22652 10948 22700 11004
rect 22756 10948 22784 11004
rect 22464 9436 22784 10948
rect 22464 9380 22492 9436
rect 22548 9380 22596 9436
rect 22652 9380 22700 9436
rect 22756 9380 22784 9436
rect 22464 7868 22784 9380
rect 22464 7812 22492 7868
rect 22548 7812 22596 7868
rect 22652 7812 22700 7868
rect 22756 7812 22784 7868
rect 22464 6300 22784 7812
rect 22464 6244 22492 6300
rect 22548 6244 22596 6300
rect 22652 6244 22700 6300
rect 22756 6244 22784 6300
rect 22464 4732 22784 6244
rect 22464 4676 22492 4732
rect 22548 4676 22596 4732
rect 22652 4676 22700 4732
rect 22756 4676 22784 4732
rect 22464 3164 22784 4676
rect 22464 3108 22492 3164
rect 22548 3108 22596 3164
rect 22652 3108 22700 3164
rect 22756 3108 22784 3164
rect 22464 3076 22784 3108
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16
timestamp 1667941163
transform 1 0 3136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22
timestamp 1667941163
transform 1 0 3808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28
timestamp 1667941163
transform 1 0 4480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1667941163
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42
timestamp 1667941163
transform 1 0 6048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48
timestamp 1667941163
transform 1 0 6720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 7392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60
timestamp 1667941163
transform 1 0 8064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1667941163
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77
timestamp 1667941163
transform 1 0 9968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83
timestamp 1667941163
transform 1 0 10640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89
timestamp 1667941163
transform 1 0 11312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95
timestamp 1667941163
transform 1 0 11984 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103
timestamp 1667941163
transform 1 0 12880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107
timestamp 1667941163
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115
timestamp 1667941163
transform 1 0 14224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121
timestamp 1667941163
transform 1 0 14896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127
timestamp 1667941163
transform 1 0 15568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133
timestamp 1667941163
transform 1 0 16240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1667941163
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147
timestamp 1667941163
transform 1 0 17808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_153
timestamp 1667941163
transform 1 0 18480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159
timestamp 1667941163
transform 1 0 19152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_165
timestamp 1667941163
transform 1 0 19824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171
timestamp 1667941163
transform 1 0 20496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_177
timestamp 1667941163
transform 1 0 21168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185
timestamp 1667941163
transform 1 0 22064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_187
timestamp 1667941163
transform 1 0 22288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1667941163
transform 1 0 1568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_6
timestamp 1667941163
transform 1 0 2016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_12
timestamp 1667941163
transform 1 0 2688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_18
timestamp 1667941163
transform 1 0 3360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_24
timestamp 1667941163
transform 1 0 4032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_30
timestamp 1667941163
transform 1 0 4704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_36
timestamp 1667941163
transform 1 0 5376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1667941163
transform 1 0 6048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_48
timestamp 1667941163
transform 1 0 6720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 7392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_60
timestamp 1667941163
transform 1 0 8064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1667941163
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_78
timestamp 1667941163
transform 1 0 10080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_84
timestamp 1667941163
transform 1 0 10752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_90
timestamp 1667941163
transform 1 0 11424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_94
timestamp 1667941163
transform 1 0 11872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_96
timestamp 1667941163
transform 1 0 12096 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_101
timestamp 1667941163
transform 1 0 12656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_107
timestamp 1667941163
transform 1 0 13328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 14000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_119
timestamp 1667941163
transform 1 0 14672 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_125
timestamp 1667941163
transform 1 0 15344 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_131
timestamp 1667941163
transform 1 0 16016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1667941163
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_149
timestamp 1667941163
transform 1 0 18032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_155
timestamp 1667941163
transform 1 0 18704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_161
timestamp 1667941163
transform 1 0 19376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_167
timestamp 1667941163
transform 1 0 20048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_173
timestamp 1667941163
transform 1 0 20720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_179
timestamp 1667941163
transform 1 0 21392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_185
timestamp 1667941163
transform 1 0 22064 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_187
timestamp 1667941163
transform 1 0 22288 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1667941163
transform 1 0 1568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_10
timestamp 1667941163
transform 1 0 2464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_16
timestamp 1667941163
transform 1 0 3136 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_22
timestamp 1667941163
transform 1 0 3808 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_28
timestamp 1667941163
transform 1 0 4480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1667941163
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_42
timestamp 1667941163
transform 1 0 6048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_48
timestamp 1667941163
transform 1 0 6720 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_54
timestamp 1667941163
transform 1 0 7392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_60
timestamp 1667941163
transform 1 0 8064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_66
timestamp 1667941163
transform 1 0 8736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_72
timestamp 1667941163
transform 1 0 9408 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_78
timestamp 1667941163
transform 1 0 10080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_84
timestamp 1667941163
transform 1 0 10752 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_88
timestamp 1667941163
transform 1 0 11200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_93
timestamp 1667941163
transform 1 0 11760 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_99
timestamp 1667941163
transform 1 0 12432 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_108
timestamp 1667941163
transform 1 0 13440 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_116
timestamp 1667941163
transform 1 0 14336 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_122
timestamp 1667941163
transform 1 0 15008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_128
timestamp 1667941163
transform 1 0 15680 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_134
timestamp 1667941163
transform 1 0 16352 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_140
timestamp 1667941163
transform 1 0 17024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_146
timestamp 1667941163
transform 1 0 17696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_152
timestamp 1667941163
transform 1 0 18368 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_158
timestamp 1667941163
transform 1 0 19040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_164
timestamp 1667941163
transform 1 0 19712 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_170
timestamp 1667941163
transform 1 0 20384 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1667941163
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_184
timestamp 1667941163
transform 1 0 21952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_2
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_4
timestamp 1667941163
transform 1 0 1792 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_9
timestamp 1667941163
transform 1 0 2352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_15
timestamp 1667941163
transform 1 0 3024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_21
timestamp 1667941163
transform 1 0 3696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_27
timestamp 1667941163
transform 1 0 4368 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_33
timestamp 1667941163
transform 1 0 5040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_39
timestamp 1667941163
transform 1 0 5712 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_45
timestamp 1667941163
transform 1 0 6384 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_51
timestamp 1667941163
transform 1 0 7056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 7728 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_63
timestamp 1667941163
transform 1 0 8400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_69
timestamp 1667941163
transform 1 0 9072 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1667941163
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_78
timestamp 1667941163
transform 1 0 10080 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_84
timestamp 1667941163
transform 1 0 10752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_90
timestamp 1667941163
transform 1 0 11424 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_96
timestamp 1667941163
transform 1 0 12096 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_98
timestamp 1667941163
transform 1 0 12320 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_103
timestamp 1667941163
transform 1 0 12880 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_109
timestamp 1667941163
transform 1 0 13552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_115
timestamp 1667941163
transform 1 0 14224 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_121
timestamp 1667941163
transform 1 0 14896 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_127
timestamp 1667941163
transform 1 0 15568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_133
timestamp 1667941163
transform 1 0 16240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_139
timestamp 1667941163
transform 1 0 16912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1667941163
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_149
timestamp 1667941163
transform 1 0 18032 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_155
timestamp 1667941163
transform 1 0 18704 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_161
timestamp 1667941163
transform 1 0 19376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_167
timestamp 1667941163
transform 1 0 20048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_173
timestamp 1667941163
transform 1 0 20720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_179
timestamp 1667941163
transform 1 0 21392 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_185
timestamp 1667941163
transform 1 0 22064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_187
timestamp 1667941163
transform 1 0 22288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1667941163
transform 1 0 1568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_10
timestamp 1667941163
transform 1 0 2464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_16
timestamp 1667941163
transform 1 0 3136 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_22
timestamp 1667941163
transform 1 0 3808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_28
timestamp 1667941163
transform 1 0 4480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1667941163
transform 1 0 5488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_42
timestamp 1667941163
transform 1 0 6048 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_48
timestamp 1667941163
transform 1 0 6720 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_54
timestamp 1667941163
transform 1 0 7392 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_60
timestamp 1667941163
transform 1 0 8064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_66
timestamp 1667941163
transform 1 0 8736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_72
timestamp 1667941163
transform 1 0 9408 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_78
timestamp 1667941163
transform 1 0 10080 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_84
timestamp 1667941163
transform 1 0 10752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_90
timestamp 1667941163
transform 1 0 11424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_96
timestamp 1667941163
transform 1 0 12096 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_102
timestamp 1667941163
transform 1 0 12768 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_108
timestamp 1667941163
transform 1 0 13440 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_112
timestamp 1667941163
transform 1 0 13888 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_117
timestamp 1667941163
transform 1 0 14448 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_123
timestamp 1667941163
transform 1 0 15120 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_129
timestamp 1667941163
transform 1 0 15792 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_135
timestamp 1667941163
transform 1 0 16464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 17136 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_147
timestamp 1667941163
transform 1 0 17808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_153
timestamp 1667941163
transform 1 0 18480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_159
timestamp 1667941163
transform 1 0 19152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_165
timestamp 1667941163
transform 1 0 19824 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1667941163
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_175
timestamp 1667941163
transform 1 0 20944 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1667941163
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_184
timestamp 1667941163
transform 1 0 21952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_2
timestamp 1667941163
transform 1 0 1568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_4
timestamp 1667941163
transform 1 0 1792 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_9
timestamp 1667941163
transform 1 0 2352 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_15
timestamp 1667941163
transform 1 0 3024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_21
timestamp 1667941163
transform 1 0 3696 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_27
timestamp 1667941163
transform 1 0 4368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_33
timestamp 1667941163
transform 1 0 5040 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_39
timestamp 1667941163
transform 1 0 5712 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_45
timestamp 1667941163
transform 1 0 6384 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_51
timestamp 1667941163
transform 1 0 7056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 7728 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_59
timestamp 1667941163
transform 1 0 7952 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_64
timestamp 1667941163
transform 1 0 8512 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_73
timestamp 1667941163
transform 1 0 9520 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_79
timestamp 1667941163
transform 1 0 10192 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_85
timestamp 1667941163
transform 1 0 10864 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_91
timestamp 1667941163
transform 1 0 11536 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_97
timestamp 1667941163
transform 1 0 12208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_103
timestamp 1667941163
transform 1 0 12880 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_109
timestamp 1667941163
transform 1 0 13552 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_115
timestamp 1667941163
transform 1 0 14224 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_121
timestamp 1667941163
transform 1 0 14896 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_127
timestamp 1667941163
transform 1 0 15568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_133
timestamp 1667941163
transform 1 0 16240 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_139
timestamp 1667941163
transform 1 0 16912 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1667941163
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_149
timestamp 1667941163
transform 1 0 18032 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_155
timestamp 1667941163
transform 1 0 18704 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_161
timestamp 1667941163
transform 1 0 19376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_167
timestamp 1667941163
transform 1 0 20048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_173
timestamp 1667941163
transform 1 0 20720 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_179
timestamp 1667941163
transform 1 0 21392 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_187
timestamp 1667941163
transform 1 0 22288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_2
timestamp 1667941163
transform 1 0 1568 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_10
timestamp 1667941163
transform 1 0 2464 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_16
timestamp 1667941163
transform 1 0 3136 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_22
timestamp 1667941163
transform 1 0 3808 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_28
timestamp 1667941163
transform 1 0 4480 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_37
timestamp 1667941163
transform 1 0 5488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_43
timestamp 1667941163
transform 1 0 6160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_49
timestamp 1667941163
transform 1 0 6832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_55
timestamp 1667941163
transform 1 0 7504 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_61
timestamp 1667941163
transform 1 0 8176 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_67
timestamp 1667941163
transform 1 0 8848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_73
timestamp 1667941163
transform 1 0 9520 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_79
timestamp 1667941163
transform 1 0 10192 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 10864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_91
timestamp 1667941163
transform 1 0 11536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_99
timestamp 1667941163
transform 1 0 12432 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1667941163
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_113
timestamp 1667941163
transform 1 0 14000 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_119
timestamp 1667941163
transform 1 0 14672 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_125
timestamp 1667941163
transform 1 0 15344 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_131
timestamp 1667941163
transform 1 0 16016 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_137
timestamp 1667941163
transform 1 0 16688 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_143
timestamp 1667941163
transform 1 0 17360 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_149
timestamp 1667941163
transform 1 0 18032 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_155
timestamp 1667941163
transform 1 0 18704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_161
timestamp 1667941163
transform 1 0 19376 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_167
timestamp 1667941163
transform 1 0 20048 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_173
timestamp 1667941163
transform 1 0 20720 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_179
timestamp 1667941163
transform 1 0 21392 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_187
timestamp 1667941163
transform 1 0 22288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_2
timestamp 1667941163
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_10
timestamp 1667941163
transform 1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_14
timestamp 1667941163
transform 1 0 2912 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_16
timestamp 1667941163
transform 1 0 3136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_21
timestamp 1667941163
transform 1 0 3696 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_27
timestamp 1667941163
transform 1 0 4368 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_33
timestamp 1667941163
transform 1 0 5040 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_39
timestamp 1667941163
transform 1 0 5712 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_45
timestamp 1667941163
transform 1 0 6384 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_51
timestamp 1667941163
transform 1 0 7056 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 7728 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_59
timestamp 1667941163
transform 1 0 7952 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_64
timestamp 1667941163
transform 1 0 8512 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_73
timestamp 1667941163
transform 1 0 9520 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_77
timestamp 1667941163
transform 1 0 9968 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_83
timestamp 1667941163
transform 1 0 10640 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_89
timestamp 1667941163
transform 1 0 11312 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_95
timestamp 1667941163
transform 1 0 11984 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_101
timestamp 1667941163
transform 1 0 12656 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_107
timestamp 1667941163
transform 1 0 13328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 14000 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_119
timestamp 1667941163
transform 1 0 14672 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_125
timestamp 1667941163
transform 1 0 15344 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_131
timestamp 1667941163
transform 1 0 16016 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1667941163
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_149
timestamp 1667941163
transform 1 0 18032 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_155
timestamp 1667941163
transform 1 0 18704 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_161
timestamp 1667941163
transform 1 0 19376 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_167
timestamp 1667941163
transform 1 0 20048 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_173
timestamp 1667941163
transform 1 0 20720 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_181
timestamp 1667941163
transform 1 0 21616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_185
timestamp 1667941163
transform 1 0 22064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_187
timestamp 1667941163
transform 1 0 22288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_18
timestamp 1667941163
transform 1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_22
timestamp 1667941163
transform 1 0 3808 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_28
timestamp 1667941163
transform 1 0 4480 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_37
timestamp 1667941163
transform 1 0 5488 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_43
timestamp 1667941163
transform 1 0 6160 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_49
timestamp 1667941163
transform 1 0 6832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_55
timestamp 1667941163
transform 1 0 7504 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_61
timestamp 1667941163
transform 1 0 8176 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_67
timestamp 1667941163
transform 1 0 8848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_73
timestamp 1667941163
transform 1 0 9520 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_79
timestamp 1667941163
transform 1 0 10192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_85
timestamp 1667941163
transform 1 0 10864 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_93
timestamp 1667941163
transform 1 0 11760 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_99
timestamp 1667941163
transform 1 0 12432 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1667941163
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_113
timestamp 1667941163
transform 1 0 14000 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_119
timestamp 1667941163
transform 1 0 14672 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_125
timestamp 1667941163
transform 1 0 15344 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_131
timestamp 1667941163
transform 1 0 16016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_137
timestamp 1667941163
transform 1 0 16688 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_143
timestamp 1667941163
transform 1 0 17360 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_149
timestamp 1667941163
transform 1 0 18032 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_155
timestamp 1667941163
transform 1 0 18704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_161
timestamp 1667941163
transform 1 0 19376 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_167
timestamp 1667941163
transform 1 0 20048 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_173
timestamp 1667941163
transform 1 0 20720 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_179
timestamp 1667941163
transform 1 0 21392 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_184
timestamp 1667941163
transform 1 0 21952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_34
timestamp 1667941163
transform 1 0 5152 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_39
timestamp 1667941163
transform 1 0 5712 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_45
timestamp 1667941163
transform 1 0 6384 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_51
timestamp 1667941163
transform 1 0 7056 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 7728 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_63
timestamp 1667941163
transform 1 0 8400 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_65
timestamp 1667941163
transform 1 0 8624 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_73
timestamp 1667941163
transform 1 0 9520 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_79
timestamp 1667941163
transform 1 0 10192 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_85
timestamp 1667941163
transform 1 0 10864 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_91
timestamp 1667941163
transform 1 0 11536 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_93
timestamp 1667941163
transform 1 0 11760 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_98
timestamp 1667941163
transform 1 0 12320 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_104
timestamp 1667941163
transform 1 0 12992 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 13664 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_116
timestamp 1667941163
transform 1 0 14336 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_122
timestamp 1667941163
transform 1 0 15008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_128
timestamp 1667941163
transform 1 0 15680 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_134
timestamp 1667941163
transform 1 0 16352 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_140
timestamp 1667941163
transform 1 0 17024 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1667941163
transform 1 0 17472 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_149
timestamp 1667941163
transform 1 0 18032 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_155
timestamp 1667941163
transform 1 0 18704 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_161
timestamp 1667941163
transform 1 0 19376 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_167
timestamp 1667941163
transform 1 0 20048 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_173
timestamp 1667941163
transform 1 0 20720 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_179
timestamp 1667941163
transform 1 0 21392 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_185
timestamp 1667941163
transform 1 0 22064 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_187
timestamp 1667941163
transform 1 0 22288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1667941163
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_37
timestamp 1667941163
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_45
timestamp 1667941163
transform 1 0 6384 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_47
timestamp 1667941163
transform 1 0 6608 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_52
timestamp 1667941163
transform 1 0 7168 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_58
timestamp 1667941163
transform 1 0 7840 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_64
timestamp 1667941163
transform 1 0 8512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_68
timestamp 1667941163
transform 1 0 8960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_73
timestamp 1667941163
transform 1 0 9520 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_79
timestamp 1667941163
transform 1 0 10192 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_85
timestamp 1667941163
transform 1 0 10864 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_93
timestamp 1667941163
transform 1 0 11760 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_99
timestamp 1667941163
transform 1 0 12432 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1667941163
transform 1 0 13440 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_113
timestamp 1667941163
transform 1 0 14000 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_117
timestamp 1667941163
transform 1 0 14448 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_123
timestamp 1667941163
transform 1 0 15120 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_129
timestamp 1667941163
transform 1 0 15792 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_135
timestamp 1667941163
transform 1 0 16464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 17136 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_147
timestamp 1667941163
transform 1 0 17808 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_153
timestamp 1667941163
transform 1 0 18480 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_159
timestamp 1667941163
transform 1 0 19152 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_165
timestamp 1667941163
transform 1 0 19824 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1667941163
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_175
timestamp 1667941163
transform 1 0 20944 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_179
timestamp 1667941163
transform 1 0 21392 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_187
timestamp 1667941163
transform 1 0 22288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_73
timestamp 1667941163
transform 1 0 9520 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_105
timestamp 1667941163
transform 1 0 13104 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_117
timestamp 1667941163
transform 1 0 14448 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_123
timestamp 1667941163
transform 1 0 15120 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_129
timestamp 1667941163
transform 1 0 15792 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_135
timestamp 1667941163
transform 1 0 16464 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1667941163
transform 1 0 17472 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_149
timestamp 1667941163
transform 1 0 18032 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_155
timestamp 1667941163
transform 1 0 18704 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_161
timestamp 1667941163
transform 1 0 19376 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_167
timestamp 1667941163
transform 1 0 20048 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_173
timestamp 1667941163
transform 1 0 20720 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_181
timestamp 1667941163
transform 1 0 21616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_185
timestamp 1667941163
transform 1 0 22064 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_187
timestamp 1667941163
transform 1 0 22288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1667941163
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1667941163
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1667941163
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_108
timestamp 1667941163
transform 1 0 13440 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_116
timestamp 1667941163
transform 1 0 14336 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_118
timestamp 1667941163
transform 1 0 14560 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_123
timestamp 1667941163
transform 1 0 15120 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_129
timestamp 1667941163
transform 1 0 15792 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_135
timestamp 1667941163
transform 1 0 16464 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 17136 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_147
timestamp 1667941163
transform 1 0 17808 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_153
timestamp 1667941163
transform 1 0 18480 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_159
timestamp 1667941163
transform 1 0 19152 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_165
timestamp 1667941163
transform 1 0 19824 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_173
timestamp 1667941163
transform 1 0 20720 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_179
timestamp 1667941163
transform 1 0 21392 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_187
timestamp 1667941163
transform 1 0 22288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1667941163
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_73
timestamp 1667941163
transform 1 0 9520 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_105
timestamp 1667941163
transform 1 0 13104 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_121
timestamp 1667941163
transform 1 0 14896 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_129
timestamp 1667941163
transform 1 0 15792 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_135
timestamp 1667941163
transform 1 0 16464 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_144
timestamp 1667941163
transform 1 0 17472 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_149
timestamp 1667941163
transform 1 0 18032 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_155
timestamp 1667941163
transform 1 0 18704 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_187
timestamp 1667941163
transform 1 0 22288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1667941163
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1667941163
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1667941163
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_108
timestamp 1667941163
transform 1 0 13440 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_124
timestamp 1667941163
transform 1 0 15232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_132
timestamp 1667941163
transform 1 0 16128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_136
timestamp 1667941163
transform 1 0 16576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 17136 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_147
timestamp 1667941163
transform 1 0 17808 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_163
timestamp 1667941163
transform 1 0 19600 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_171
timestamp 1667941163
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_175
timestamp 1667941163
transform 1 0 20944 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_179
timestamp 1667941163
transform 1 0 21392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_187
timestamp 1667941163
transform 1 0 22288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1667941163
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1667941163
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_144
timestamp 1667941163
transform 1 0 17472 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_176
timestamp 1667941163
transform 1 0 21056 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_184
timestamp 1667941163
transform 1 0 21952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1667941163
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1667941163
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_37
timestamp 1667941163
transform 1 0 5488 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_69
timestamp 1667941163
transform 1 0 9072 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_72
timestamp 1667941163
transform 1 0 9408 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_104
timestamp 1667941163
transform 1 0 12992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_107
timestamp 1667941163
transform 1 0 13328 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 16912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_142
timestamp 1667941163
transform 1 0 17248 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_174
timestamp 1667941163
transform 1 0 20832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_177
timestamp 1667941163
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_185
timestamp 1667941163
transform 1 0 22064 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_187
timestamp 1667941163
transform 1 0 22288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 22624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 22624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 22624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 22624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 22624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 22624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 22624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 22624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 22624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 22624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 22624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 22624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1667941163
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1667941163
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1667941163
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1667941163
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1667941163
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1667941163
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1667941163
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1667941163
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1667941163
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1667941163
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1667941163
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1667941163
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1667941163
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1667941163
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1667941163
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1667941163
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1667941163
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1667941163
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1667941163
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1667941163
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1667941163
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1667941163
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1667941163
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1667941163
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1667941163
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1667941163
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1667941163
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1667941163
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1667941163
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1667941163
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1667941163
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1667941163
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1667941163
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1667941163
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1667941163
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1667941163
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1667941163
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1667941163
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1667941163
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1667941163
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1667941163
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1667941163
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1667941163
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1667941163
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1667941163
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1667941163
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[0\].fbn pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 11872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 16464 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 13552 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 15792 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 13216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 11984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 15120 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 19600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 10976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 18928 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 11648 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 18928 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 11760 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 20272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 9632 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 18256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 10976 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 20272 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 10304 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 16464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 9744 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 17584 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 11648 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 20944 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 12320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 14448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 12880 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 15344 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 13552 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 15792 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 15120 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 15568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 15568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 15904 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f1.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 13776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 16016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 13552 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 15232 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 14560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 19600 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 15232 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 14448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 11088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 18704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 9744 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 16016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 10416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 18032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 9072 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 17360 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 8400 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 9072 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 17584 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 9744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[7\].thrun
timestamp 1667941163
transform -1 0 18032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 9072 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 7728 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 17584 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 16240 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 14896 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 14000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 14672 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 14224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 14896 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 13104 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_f2.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 16912 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 5264 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 6384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 8960 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 7280 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 7616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 5936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 8288 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 6608 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 8064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 10416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 10304 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 10192 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 10304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 9744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 7056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 10416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 8960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[4\].thrup
timestamp 1667941163
transform -1 0 11536 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 9632 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[5\].thrup
timestamp 1667941163
transform -1 0 11536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 7728 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 10416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 8064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 9744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 8400 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 8288 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 10416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 4592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 5936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 5712 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 6608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 4592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 8624 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 6608 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 6944 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[4\].crossn
timestamp 1667941163
transform -1 0 8512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r1.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 5712 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 20272 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 17360 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 21504 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 16688 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 19376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 17584 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 20272 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 16688 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 14672 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 21616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 15344 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 17584 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 15344 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 19600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 15344 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[4\].thrun
timestamp 1667941163
transform -1 0 17136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 16016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 16016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 14672 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 16016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 17360 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[8\].thrun
timestamp 1667941163
transform -1 0 17808 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 14000 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 18928 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 14672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 20048 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 18256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 18032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 17584 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 19376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 18704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 18928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 19600 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 18928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_nauta_series_r2.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 19600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[0\].fbn
timestamp 1667941163
transform -1 0 20720 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 13776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 20048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 11312 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 20944 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 11984 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[3\].fbn
timestamp 1667941163
transform -1 0 22064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 12208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 19600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 12880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 17248 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 16464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 20272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 15120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 19376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 12432 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 17920 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[5\].thrup
timestamp 1667941163
transform -1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 18928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 15792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 18704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 14448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 16240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 13552 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 18928 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 14224 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 19600 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 18704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 20272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 18032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 18928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 21504 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 19936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 19376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_f.gen_X\[4\].crossp
timestamp 1667941163
transform -1 0 22064 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 12432 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 13888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 11536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 12544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 16688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 11984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 10864 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 11984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 17584 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 17584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 18592 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 13776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 19264 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 13888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 20272 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 15904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 21504 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 18032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 20944 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[5\].thrup
timestamp 1667941163
transform 1 0 13104 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 19600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 14560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 20944 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 15568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 17360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 14896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 18256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 16576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 14896 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 11312 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 13552 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 16240 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 12208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 16912 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 14224 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 15568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_seriesgy.u_nauta_r.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 16240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 10976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 3248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 4032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[1\].fbp
timestamp 1667941163
transform -1 0 6384 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 2688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 4032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 10192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 5264 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 3248 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[1\].thrun
timestamp 1667941163
transform -1 0 7392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 3248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[2\].thrun
timestamp 1667941163
transform -1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 4032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 5600 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[3\].thrup
timestamp 1667941163
transform -1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 6272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 2016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 4592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[5\].thrup
timestamp 1667941163
transform -1 0 6720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 3920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 3920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[7\].thrun
timestamp 1667941163
transform -1 0 9968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 2688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 9632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 4928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 10304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 3360 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 2688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 2912 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[1\].crossn
timestamp 1667941163
transform -1 0 3136 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 2016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[2\].crossn
timestamp 1667941163
transform -1 0 2352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 3360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 10864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 2240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[4\].crossn
timestamp 1667941163
transform -1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_f.gen_X\[4\].crossp
timestamp 1667941163
transform 1 0 1904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[0\].fbn
timestamp 1667941163
transform 1 0 7280 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[0\].fbp
timestamp 1667941163
transform 1 0 5600 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[1\].fbn
timestamp 1667941163
transform 1 0 6384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[1\].fbp
timestamp 1667941163
transform 1 0 8288 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[2\].fbn
timestamp 1667941163
transform 1 0 7056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[2\].fbp
timestamp 1667941163
transform 1 0 6608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[3\].fbn
timestamp 1667941163
transform 1 0 7280 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_FB\[3\].fbp
timestamp 1667941163
transform 1 0 6272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[0\].thrun
timestamp 1667941163
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[0\].thrup
timestamp 1667941163
transform 1 0 5936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[1\].thrun
timestamp 1667941163
transform 1 0 5936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[1\].thrup
timestamp 1667941163
transform 1 0 3360 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[2\].thrun
timestamp 1667941163
transform 1 0 5264 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[2\].thrup
timestamp 1667941163
transform 1 0 2576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[3\].thrun
timestamp 1667941163
transform 1 0 6944 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[3\].thrup
timestamp 1667941163
transform 1 0 3920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[4\].thrun
timestamp 1667941163
transform 1 0 7616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[4\].thrup
timestamp 1667941163
transform 1 0 2576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[5\].thrun
timestamp 1667941163
transform 1 0 5600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[5\].thrup
timestamp 1667941163
transform -1 0 7168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[6\].thrun
timestamp 1667941163
transform 1 0 4032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[6\].thrup
timestamp 1667941163
transform 1 0 4256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[7\].thrun
timestamp 1667941163
transform 1 0 9632 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[7\].thrup
timestamp 1667941163
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[8\].thrun
timestamp 1667941163
transform 1 0 7616 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[8\].thrup
timestamp 1667941163
transform 1 0 3584 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[9\].thrun
timestamp 1667941163
transform 1 0 6272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_T\[9\].thrup
timestamp 1667941163
transform 1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[0\].crossn
timestamp 1667941163
transform 1 0 7616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[0\].crossp
timestamp 1667941163
transform 1 0 3360 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[1\].crossn
timestamp 1667941163
transform 1 0 7952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[1\].crossp
timestamp 1667941163
transform 1 0 6944 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[2\].crossn
timestamp 1667941163
transform 1 0 7952 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[2\].crossp
timestamp 1667941163
transform 1 0 4032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[3\].crossn
timestamp 1667941163
transform 1 0 7280 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[3\].crossp
timestamp 1667941163
transform 1 0 5264 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[4\].crossn
timestamp 1667941163
transform 1 0 4704 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_shuntgy.u_nauta_r.gen_X\[4\].crossp
timestamp 1667941163
transform -1 0 7840 0 1 10976
box -86 -86 534 870
<< labels >>
flabel metal3 s 0 14896 800 15008 0 FreeSans 448 0 0 0 nbusin_nshunt
port 0 nsew signal bidirectional
flabel metal3 s 23200 14896 24000 15008 0 FreeSans 448 0 0 0 nbusout
port 1 nsew signal bidirectional
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 nseries_gy
port 2 nsew signal bidirectional
flabel metal2 s 21728 0 21840 800 0 FreeSans 448 90 0 0 nseries_gygy
port 3 nsew signal bidirectional
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 nshunt_gy
port 4 nsew signal bidirectional
flabel metal3 s 0 4928 800 5040 0 FreeSans 448 0 0 0 pbusin_pshunt
port 5 nsew signal bidirectional
flabel metal3 s 23200 4928 24000 5040 0 FreeSans 448 0 0 0 pbusout
port 6 nsew signal bidirectional
flabel metal2 s 9968 0 10080 800 0 FreeSans 448 90 0 0 pseries_gy
port 7 nsew signal bidirectional
flabel metal2 s 17808 0 17920 800 0 FreeSans 448 90 0 0 pseries_gygy
port 8 nsew signal bidirectional
flabel metal2 s 2128 0 2240 800 0 FreeSans 448 90 0 0 pshunt_gy
port 9 nsew signal bidirectional
flabel metal4 s 3844 3076 4164 16524 0 FreeSans 1280 90 0 0 vdd
port 10 nsew power bidirectional
flabel metal4 s 9164 3076 9484 16524 0 FreeSans 1280 90 0 0 vdd
port 10 nsew power bidirectional
flabel metal4 s 14484 3076 14804 16524 0 FreeSans 1280 90 0 0 vdd
port 10 nsew power bidirectional
flabel metal4 s 19804 3076 20124 16524 0 FreeSans 1280 90 0 0 vdd
port 10 nsew power bidirectional
flabel metal4 s 6504 3076 6824 16524 0 FreeSans 1280 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 11824 3076 12144 16524 0 FreeSans 1280 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 17144 3076 17464 16524 0 FreeSans 1280 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 22464 3076 22784 16524 0 FreeSans 1280 90 0 0 vss
port 11 nsew ground bidirectional
rlabel metal1 11984 16464 11984 16464 0 vdd
rlabel via1 12064 15680 12064 15680 0 vss
rlabel metal3 4592 5096 4592 5096 0 nbusin_nshunt
rlabel metal2 20216 10976 20216 10976 0 nbusout
rlabel metal3 20888 5656 20888 5656 0 nseries_gy
rlabel metal2 21784 2422 21784 2422 0 nseries_gygy
rlabel metal3 5992 4088 5992 4088 0 nshunt_gy
rlabel metal2 2856 5600 2856 5600 0 pbusin_pshunt
rlabel metal3 22610 4984 22610 4984 0 pbusout
rlabel metal2 7896 8316 7896 8316 0 pseries_gy
rlabel metal2 20216 5880 20216 5880 0 pseries_gygy
rlabel metal2 6552 3752 6552 3752 0 pshunt_gy
<< properties >>
string FIXED_BBOX 0 0 24000 20000
<< end >>
