magic
tech gf180mcuC
magscale 1 5
timestamp 1669860616
<< obsm1 >>
rect 672 1538 5400 4342
<< obsm2 >>
rect 910 625 5386 5367
<< metal3 >>
rect 5600 5320 6000 5376
rect 0 4424 400 4480
rect 5600 4144 6000 4200
rect 5600 2968 6000 3024
rect 5600 1792 6000 1848
rect 0 1456 400 1512
rect 5600 616 6000 672
<< obsm3 >>
rect 400 5290 5570 5362
rect 400 4510 5600 5290
rect 430 4394 5600 4510
rect 400 4230 5600 4394
rect 400 4114 5570 4230
rect 400 3054 5600 4114
rect 400 2938 5570 3054
rect 400 1878 5600 2938
rect 400 1762 5570 1878
rect 400 1542 5600 1762
rect 430 1426 5600 1542
rect 400 702 5600 1426
rect 400 630 5570 702
<< metal4 >>
rect 1173 1538 1333 4342
rect 1754 1538 1914 4342
rect 2335 1538 2495 4342
rect 2916 1538 3076 4342
rect 3497 1538 3657 4342
rect 4078 1538 4238 4342
rect 4659 1538 4819 4342
rect 5240 1538 5400 4342
<< labels >>
rlabel metal3 s 0 4424 400 4480 6 nbus
port 1 nsew signal bidirectional
rlabel metal3 s 5600 1792 6000 1848 6 outn
port 2 nsew signal bidirectional
rlabel metal3 s 5600 4144 6000 4200 6 outnn
port 3 nsew signal output
rlabel metal3 s 5600 616 6000 672 6 outp
port 4 nsew signal bidirectional
rlabel metal3 s 5600 2968 6000 3024 6 outpn
port 5 nsew signal output
rlabel metal3 s 5600 5320 6000 5376 6 outxor
port 6 nsew signal output
rlabel metal3 s 0 1456 400 1512 6 pbus
port 7 nsew signal bidirectional
rlabel metal4 s 1173 1538 1333 4342 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 2335 1538 2495 4342 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 3497 1538 3657 4342 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 4659 1538 4819 4342 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 1754 1538 1914 4342 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 2916 1538 3076 4342 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 4078 1538 4238 4342 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 5240 1538 5400 4342 6 vss
port 9 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 6000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 118374
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/active_load/runs/22_11_30_21_09/results/signoff/active_load.magic.gds
string GDS_START 32722
<< end >>

