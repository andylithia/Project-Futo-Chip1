magic
tech gf180mcuC
magscale 1 10
timestamp 1669830126
<< nwell >>
rect 1258 8217 18678 8710
rect 1258 8192 3030 8217
rect 3403 8192 7846 8217
rect 8219 8192 11941 8217
rect 12314 8192 15077 8217
rect 15450 8192 18678 8217
rect 1258 7463 3030 7488
rect 3403 7463 7846 7488
rect 8219 7463 12662 7488
rect 13035 7463 15189 7488
rect 15562 7463 18678 7488
rect 1258 6624 18678 7463
rect 1258 5081 18678 5920
rect 1258 5056 17205 5081
rect 17578 5056 18678 5081
rect 1258 4327 3254 4352
rect 3627 4327 7909 4352
rect 8282 4327 12837 4352
rect 13210 4327 18678 4352
rect 1258 3513 18678 4327
rect 1258 3488 3429 3513
rect 3802 3488 8021 3513
rect 8394 3488 11941 3513
rect 12314 3488 15861 3513
rect 16234 3488 18678 3513
<< pwell >>
rect 3030 8192 3403 8217
rect 7846 8192 8219 8217
rect 11941 8192 12314 8217
rect 15077 8192 15450 8217
rect 1258 7488 18678 8192
rect 3030 7463 3403 7488
rect 7846 7463 8219 7488
rect 12662 7463 13035 7488
rect 15189 7463 15562 7488
rect 1258 5920 18678 6624
rect 17205 5056 17578 5081
rect 1258 4352 18678 5056
rect 3254 4327 3627 4352
rect 7909 4327 8282 4352
rect 12837 4327 13210 4352
rect 3429 3488 3802 3513
rect 8021 3488 8394 3513
rect 11941 3488 12314 3513
rect 15861 3488 16234 3513
rect 1258 3050 18678 3488
<< mvnmos >>
rect 1804 7908 1924 8072
rect 2476 7933 2596 8005
rect 2700 7933 2820 8005
rect 2924 7933 3044 8005
rect 3389 7908 3509 8072
rect 3757 7933 3877 8005
rect 4012 7933 4132 8005
rect 4640 7908 4760 8072
rect 4908 8000 5028 8072
rect 5612 7908 5812 8072
rect 6060 7908 6260 8072
rect 6700 7908 6820 8072
rect 7292 7933 7412 8005
rect 7516 7933 7636 8005
rect 7740 7933 7860 8005
rect 8205 7908 8325 8072
rect 8573 7933 8693 8005
rect 8828 7933 8948 8005
rect 9868 7908 9988 8072
rect 10620 7908 10740 8072
rect 11212 7933 11332 8005
rect 11467 7933 11587 8005
rect 11835 7908 11955 8072
rect 12300 7933 12420 8005
rect 12524 7933 12644 8005
rect 12748 7933 12868 8005
rect 13644 7908 13764 8072
rect 14348 7933 14468 8005
rect 14603 7933 14723 8005
rect 14971 7908 15091 8072
rect 15436 7933 15556 8005
rect 15660 7933 15780 8005
rect 15884 7933 16004 8005
rect 16476 7908 16596 8072
rect 17484 7908 17604 8072
rect 17932 7908 18132 8072
rect 1804 7608 1924 7772
rect 2476 7675 2596 7747
rect 2700 7675 2820 7747
rect 2924 7675 3044 7747
rect 3389 7608 3509 7772
rect 3757 7675 3877 7747
rect 4012 7675 4132 7747
rect 4684 7608 4804 7772
rect 5052 7608 5252 7772
rect 5500 7608 5700 7772
rect 5948 7608 6148 7772
rect 6396 7608 6596 7772
rect 6844 7608 7044 7772
rect 7292 7675 7412 7747
rect 7516 7675 7636 7747
rect 7740 7675 7860 7747
rect 8205 7608 8325 7772
rect 8573 7675 8693 7747
rect 8828 7675 8948 7747
rect 9644 7608 9844 7772
rect 10092 7608 10212 7772
rect 10764 7608 10884 7772
rect 11436 7608 11556 7772
rect 12108 7675 12228 7747
rect 12332 7675 12452 7747
rect 12556 7675 12676 7747
rect 13021 7608 13141 7772
rect 13389 7675 13509 7747
rect 13644 7675 13764 7747
rect 14012 7608 14212 7772
rect 14460 7675 14580 7747
rect 14715 7675 14835 7747
rect 15083 7608 15203 7772
rect 15548 7675 15668 7747
rect 15772 7675 15892 7747
rect 15996 7675 16116 7747
rect 16588 7608 16708 7772
rect 17708 7608 17828 7772
rect 1692 6340 1892 6504
rect 2161 6340 2281 6504
rect 2433 6365 2553 6437
rect 2657 6365 2777 6437
rect 3296 6340 3416 6504
rect 3564 6432 3684 6504
rect 3932 6340 4132 6504
rect 4380 6340 4580 6504
rect 4828 6340 5028 6504
rect 5612 6340 5812 6504
rect 6060 6340 6260 6504
rect 6923 6340 7043 6504
rect 7516 6340 7636 6504
rect 8188 6340 8308 6504
rect 8860 6340 8980 6504
rect 9532 6340 9652 6504
rect 10204 6340 10324 6504
rect 10876 6340 10996 6504
rect 11548 6340 11668 6504
rect 12220 6340 12340 6504
rect 12668 6340 12868 6504
rect 13676 6340 13796 6504
rect 14348 6340 14468 6504
rect 15020 6340 15140 6504
rect 15692 6340 15812 6504
rect 16364 6340 16484 6504
rect 17036 6340 17156 6504
rect 17708 6340 17828 6504
rect 1804 6040 1924 6113
rect 1988 6040 2108 6113
rect 2256 6040 2376 6203
rect 2924 6040 3044 6204
rect 3372 6040 3572 6204
rect 3820 6040 4020 6204
rect 4268 6040 4468 6204
rect 4716 6040 4916 6204
rect 5501 6040 5621 6204
rect 6252 6040 6372 6204
rect 6924 6040 7044 6204
rect 7516 6040 7636 6204
rect 8189 6040 8309 6204
rect 8860 6040 8980 6204
rect 9644 6040 9844 6204
rect 10316 6040 10436 6204
rect 10988 6040 11108 6204
rect 11660 6040 11780 6204
rect 12332 6040 12452 6204
rect 13004 6040 13124 6204
rect 13676 6040 13796 6204
rect 14348 6040 14468 6204
rect 15020 6040 15140 6204
rect 15692 6040 15812 6204
rect 16365 6040 16485 6204
rect 16812 6040 17012 6204
rect 17787 6040 17907 6204
rect 1692 4772 1892 4936
rect 2140 4772 2340 4936
rect 2588 4772 2788 4936
rect 3036 4772 3236 4936
rect 3484 4772 3684 4936
rect 4157 4772 4277 4936
rect 4829 4772 4949 4936
rect 5612 4772 5812 4936
rect 6285 4772 6405 4936
rect 7035 4772 7155 4936
rect 7708 4772 7828 4936
rect 8301 4772 8421 4936
rect 8972 4772 9092 4936
rect 9644 4772 9764 4936
rect 10316 4772 10436 4936
rect 10988 4772 11108 4936
rect 11660 4772 11780 4936
rect 12332 4772 12452 4936
rect 12780 4772 12980 4936
rect 13676 4772 13796 4936
rect 14348 4772 14468 4936
rect 15100 4772 15220 4936
rect 15771 4772 15891 4936
rect 16476 4797 16596 4869
rect 16731 4797 16851 4869
rect 17099 4772 17219 4936
rect 17564 4797 17684 4869
rect 17788 4797 17908 4869
rect 18012 4797 18132 4869
rect 1692 4472 1892 4636
rect 2140 4472 2340 4636
rect 2700 4539 2820 4611
rect 2924 4539 3044 4611
rect 3148 4539 3268 4611
rect 3613 4472 3733 4636
rect 3981 4539 4101 4611
rect 4236 4539 4356 4611
rect 4604 4472 4804 4636
rect 5165 4472 5285 4636
rect 5837 4472 5957 4636
rect 6509 4472 6629 4636
rect 7180 4539 7300 4611
rect 7435 4539 7555 4611
rect 7803 4472 7923 4636
rect 8268 4539 8388 4611
rect 8492 4539 8612 4611
rect 8716 4539 8836 4611
rect 9644 4472 9844 4636
rect 10093 4472 10213 4636
rect 10844 4472 10964 4636
rect 11516 4472 11636 4636
rect 12108 4539 12228 4611
rect 12363 4539 12483 4611
rect 12731 4472 12851 4636
rect 13196 4539 13316 4611
rect 13420 4539 13540 4611
rect 13644 4539 13764 4611
rect 14237 4472 14357 4636
rect 14908 4472 15028 4636
rect 15580 4472 15700 4636
rect 16252 4472 16372 4636
rect 16700 4472 16900 4636
rect 17708 4472 17828 4636
rect 2029 3204 2149 3368
rect 2700 3229 2820 3301
rect 2955 3229 3075 3301
rect 3323 3204 3443 3368
rect 3788 3229 3908 3301
rect 4012 3229 4132 3301
rect 4236 3229 4356 3301
rect 4829 3204 4949 3368
rect 5949 3204 6069 3368
rect 6621 3204 6741 3368
rect 7292 3229 7412 3301
rect 7547 3229 7667 3301
rect 7915 3204 8035 3368
rect 8380 3229 8500 3301
rect 8604 3229 8724 3301
rect 8828 3229 8948 3301
rect 9869 3204 9989 3368
rect 10541 3204 10661 3368
rect 11212 3229 11332 3301
rect 11467 3229 11587 3301
rect 11835 3204 11955 3368
rect 12300 3229 12420 3301
rect 12524 3229 12644 3301
rect 12748 3229 12868 3301
rect 13644 3204 13764 3368
rect 14237 3204 14357 3368
rect 14684 3204 14884 3368
rect 15132 3229 15252 3301
rect 15387 3229 15507 3301
rect 15755 3204 15875 3368
rect 16220 3229 16340 3301
rect 16444 3229 16564 3301
rect 16668 3229 16788 3301
rect 17563 3204 17683 3368
rect 17932 3204 18132 3368
<< mvpmos >>
rect 1824 8312 1924 8556
rect 2476 8400 2576 8524
rect 2680 8400 2780 8524
rect 2884 8400 2984 8524
rect 3346 8337 3446 8556
rect 3777 8432 3877 8556
rect 4012 8432 4112 8556
rect 4660 8312 4760 8556
rect 4908 8443 5008 8556
rect 5612 8312 5812 8556
rect 6060 8312 6260 8556
rect 6700 8312 6800 8556
rect 7292 8400 7392 8524
rect 7496 8400 7596 8524
rect 7700 8400 7800 8524
rect 8162 8337 8262 8556
rect 8593 8432 8693 8556
rect 8828 8432 8928 8556
rect 9888 8312 9988 8556
rect 10620 8312 10720 8556
rect 11232 8432 11332 8556
rect 11467 8432 11567 8556
rect 11898 8337 11998 8556
rect 12360 8400 12460 8524
rect 12564 8400 12664 8524
rect 12768 8400 12868 8524
rect 13644 8312 13744 8556
rect 14368 8432 14468 8556
rect 14603 8432 14703 8556
rect 15034 8337 15134 8556
rect 15496 8400 15596 8524
rect 15700 8400 15800 8524
rect 15904 8400 16004 8524
rect 16496 8312 16596 8556
rect 17504 8312 17604 8556
rect 17932 8312 18132 8556
rect 1824 7124 1924 7368
rect 2476 7156 2576 7280
rect 2680 7156 2780 7280
rect 2884 7156 2984 7280
rect 3346 7124 3446 7343
rect 3777 7124 3877 7248
rect 4012 7124 4112 7248
rect 4684 7124 4784 7368
rect 5052 7124 5252 7368
rect 5500 7124 5700 7368
rect 5948 7124 6148 7368
rect 6396 7124 6596 7368
rect 6844 7124 7044 7368
rect 7292 7156 7392 7280
rect 7496 7156 7596 7280
rect 7700 7156 7800 7280
rect 8162 7124 8262 7343
rect 8593 7124 8693 7248
rect 8828 7124 8928 7248
rect 9644 7124 9844 7368
rect 10112 7124 10212 7368
rect 10784 7124 10884 7368
rect 11456 7124 11556 7368
rect 12108 7156 12208 7280
rect 12312 7156 12412 7280
rect 12516 7156 12616 7280
rect 12978 7124 13078 7343
rect 13409 7124 13509 7248
rect 13644 7124 13744 7248
rect 14012 7124 14212 7368
rect 14480 7124 14580 7248
rect 14715 7124 14815 7248
rect 15146 7124 15246 7343
rect 15608 7156 15708 7280
rect 15812 7156 15912 7280
rect 16016 7156 16116 7280
rect 16608 7124 16708 7368
rect 17728 7124 17828 7368
rect 1692 6744 1892 6988
rect 2181 6744 2281 6988
rect 2453 6875 2553 6988
rect 2657 6875 2757 6988
rect 3316 6744 3416 6988
rect 3564 6875 3664 6988
rect 3932 6744 4132 6988
rect 4380 6744 4580 6988
rect 4828 6744 5028 6988
rect 5612 6744 5812 6988
rect 6060 6744 6260 6988
rect 6943 6744 7043 6988
rect 7536 6744 7636 6988
rect 8208 6744 8308 6988
rect 8880 6744 8980 6988
rect 9552 6744 9652 6988
rect 10224 6744 10324 6988
rect 10896 6744 10996 6988
rect 11568 6744 11668 6988
rect 12240 6744 12340 6988
rect 12668 6744 12868 6988
rect 13696 6744 13796 6988
rect 14368 6744 14468 6988
rect 15040 6744 15140 6988
rect 15712 6744 15812 6988
rect 16384 6744 16484 6988
rect 17056 6744 17156 6988
rect 17728 6744 17828 6988
rect 1804 5557 1904 5677
rect 2008 5557 2108 5677
rect 2276 5557 2376 5800
rect 2944 5556 3044 5800
rect 3372 5556 3572 5800
rect 3820 5556 4020 5800
rect 4268 5556 4468 5800
rect 4716 5556 4916 5800
rect 5501 5556 5601 5800
rect 6252 5556 6352 5800
rect 6924 5556 7024 5800
rect 7536 5556 7636 5800
rect 8189 5556 8289 5800
rect 8880 5556 8980 5800
rect 9644 5556 9844 5800
rect 10336 5556 10436 5800
rect 11008 5556 11108 5800
rect 11680 5556 11780 5800
rect 12352 5556 12452 5800
rect 13024 5556 13124 5800
rect 13696 5556 13796 5800
rect 14368 5556 14468 5800
rect 15040 5556 15140 5800
rect 15712 5556 15812 5800
rect 16365 5556 16465 5800
rect 16812 5556 17012 5800
rect 17807 5556 17907 5800
rect 1692 5176 1892 5420
rect 2140 5176 2340 5420
rect 2588 5176 2788 5420
rect 3036 5176 3236 5420
rect 3484 5176 3684 5420
rect 4157 5176 4257 5420
rect 4829 5176 4929 5420
rect 5612 5176 5812 5420
rect 6285 5176 6385 5420
rect 7055 5176 7155 5420
rect 7708 5176 7808 5420
rect 8301 5176 8401 5420
rect 8992 5176 9092 5420
rect 9664 5176 9764 5420
rect 10336 5176 10436 5420
rect 11008 5176 11108 5420
rect 11680 5176 11780 5420
rect 12352 5176 12452 5420
rect 12780 5176 12980 5420
rect 13696 5176 13796 5420
rect 14368 5176 14468 5420
rect 15100 5176 15200 5420
rect 15791 5176 15891 5420
rect 16496 5296 16596 5420
rect 16731 5296 16831 5420
rect 17162 5201 17262 5420
rect 17624 5264 17724 5388
rect 17828 5264 17928 5388
rect 18032 5264 18132 5388
rect 1692 3988 1892 4232
rect 2140 3988 2340 4232
rect 2700 4020 2800 4144
rect 2904 4020 3004 4144
rect 3108 4020 3208 4144
rect 3570 3988 3670 4207
rect 4001 3988 4101 4112
rect 4236 3988 4336 4112
rect 4604 3988 4804 4232
rect 5165 3988 5265 4232
rect 5837 3988 5937 4232
rect 6509 3988 6609 4232
rect 7200 3988 7300 4112
rect 7435 3988 7535 4112
rect 7866 3988 7966 4207
rect 8328 4020 8428 4144
rect 8532 4020 8632 4144
rect 8736 4020 8836 4144
rect 9644 3988 9844 4232
rect 10093 3988 10193 4232
rect 10844 3988 10944 4232
rect 11516 3988 11616 4232
rect 12128 3988 12228 4112
rect 12363 3988 12463 4112
rect 12794 3988 12894 4207
rect 13256 4020 13356 4144
rect 13460 4020 13560 4144
rect 13664 4020 13764 4144
rect 14237 3988 14337 4232
rect 14928 3988 15028 4232
rect 15600 3988 15700 4232
rect 16272 3988 16372 4232
rect 16700 3988 16900 4232
rect 17728 3988 17828 4232
rect 2029 3608 2129 3852
rect 2720 3728 2820 3852
rect 2955 3728 3055 3852
rect 3386 3633 3486 3852
rect 3848 3696 3948 3820
rect 4052 3696 4152 3820
rect 4256 3696 4356 3820
rect 4829 3608 4929 3852
rect 5949 3608 6049 3852
rect 6621 3608 6721 3852
rect 7312 3728 7412 3852
rect 7547 3728 7647 3852
rect 7978 3633 8078 3852
rect 8440 3696 8540 3820
rect 8644 3696 8744 3820
rect 8848 3696 8948 3820
rect 9869 3608 9969 3852
rect 10541 3608 10641 3852
rect 11232 3728 11332 3852
rect 11467 3728 11567 3852
rect 11898 3633 11998 3852
rect 12360 3696 12460 3820
rect 12564 3696 12664 3820
rect 12768 3696 12868 3820
rect 13644 3608 13744 3852
rect 14237 3608 14337 3852
rect 14684 3608 14884 3852
rect 15152 3728 15252 3852
rect 15387 3728 15487 3852
rect 15818 3633 15918 3852
rect 16280 3696 16380 3820
rect 16484 3696 16584 3820
rect 16688 3696 16788 3820
rect 17583 3608 17683 3852
rect 17932 3608 18132 3852
<< mvndiff >>
rect 1716 8032 1804 8072
rect 1716 7986 1729 8032
rect 1775 7986 1804 8032
rect 1716 7908 1804 7986
rect 1924 8032 2012 8072
rect 1924 7986 1953 8032
rect 1999 7986 2012 8032
rect 3104 8084 3176 8097
rect 3104 8038 3117 8084
rect 3163 8038 3176 8084
rect 3104 8005 3176 8038
rect 1924 7908 2012 7986
rect 2388 7992 2476 8005
rect 2388 7946 2401 7992
rect 2447 7946 2476 7992
rect 2388 7933 2476 7946
rect 2596 7992 2700 8005
rect 2596 7946 2625 7992
rect 2671 7946 2700 7992
rect 2596 7933 2700 7946
rect 2820 7992 2924 8005
rect 2820 7946 2849 7992
rect 2895 7946 2924 7992
rect 2820 7933 2924 7946
rect 3044 7933 3176 8005
rect 3256 8084 3329 8097
rect 3256 8038 3269 8084
rect 3315 8072 3329 8084
rect 3315 8038 3389 8072
rect 3256 7908 3389 8038
rect 3509 7982 3597 8072
rect 4552 8016 4640 8072
rect 3509 7936 3538 7982
rect 3584 7936 3597 7982
rect 3509 7908 3597 7936
rect 3669 7992 3757 8005
rect 3669 7946 3682 7992
rect 3728 7946 3757 7992
rect 3669 7933 3757 7946
rect 3877 7992 4012 8005
rect 3877 7946 3906 7992
rect 3952 7946 4012 7992
rect 3877 7933 4012 7946
rect 4132 7992 4220 8005
rect 4132 7946 4161 7992
rect 4207 7946 4220 7992
rect 4132 7933 4220 7946
rect 4552 7970 4565 8016
rect 4611 7970 4640 8016
rect 4552 7908 4640 7970
rect 4760 8000 4908 8072
rect 5028 8059 5116 8072
rect 5028 8013 5057 8059
rect 5103 8013 5116 8059
rect 5028 8000 5116 8013
rect 4760 7954 4789 8000
rect 4835 7954 4848 8000
rect 4760 7908 4848 7954
rect 5524 8032 5612 8072
rect 5524 7986 5537 8032
rect 5583 7986 5612 8032
rect 5524 7908 5612 7986
rect 5812 8032 5900 8072
rect 5812 7986 5841 8032
rect 5887 7986 5900 8032
rect 5812 7908 5900 7986
rect 5972 8032 6060 8072
rect 5972 7986 5985 8032
rect 6031 7986 6060 8032
rect 5972 7908 6060 7986
rect 6260 8032 6348 8072
rect 6260 7986 6289 8032
rect 6335 7986 6348 8032
rect 6260 7908 6348 7986
rect 6612 8032 6700 8072
rect 6612 7986 6625 8032
rect 6671 7986 6700 8032
rect 6612 7908 6700 7986
rect 6820 8032 6908 8072
rect 6820 7986 6849 8032
rect 6895 7986 6908 8032
rect 7920 8084 7992 8097
rect 7920 8038 7933 8084
rect 7979 8038 7992 8084
rect 7920 8005 7992 8038
rect 6820 7908 6908 7986
rect 7204 7992 7292 8005
rect 7204 7946 7217 7992
rect 7263 7946 7292 7992
rect 7204 7933 7292 7946
rect 7412 7992 7516 8005
rect 7412 7946 7441 7992
rect 7487 7946 7516 7992
rect 7412 7933 7516 7946
rect 7636 7992 7740 8005
rect 7636 7946 7665 7992
rect 7711 7946 7740 7992
rect 7636 7933 7740 7946
rect 7860 7933 7992 8005
rect 8072 8084 8145 8097
rect 8072 8038 8085 8084
rect 8131 8072 8145 8084
rect 8131 8038 8205 8072
rect 8072 7908 8205 8038
rect 8325 7982 8413 8072
rect 8325 7936 8354 7982
rect 8400 7936 8413 7982
rect 8325 7908 8413 7936
rect 8485 7992 8573 8005
rect 8485 7946 8498 7992
rect 8544 7946 8573 7992
rect 8485 7933 8573 7946
rect 8693 7992 8828 8005
rect 8693 7946 8722 7992
rect 8768 7946 8828 7992
rect 8693 7933 8828 7946
rect 8948 7992 9036 8005
rect 8948 7946 8977 7992
rect 9023 7946 9036 7992
rect 8948 7933 9036 7946
rect 9780 8032 9868 8072
rect 9780 7986 9793 8032
rect 9839 7986 9868 8032
rect 9780 7908 9868 7986
rect 9988 8032 10076 8072
rect 9988 7986 10017 8032
rect 10063 7986 10076 8032
rect 9988 7908 10076 7986
rect 10532 8032 10620 8072
rect 10532 7986 10545 8032
rect 10591 7986 10620 8032
rect 10532 7908 10620 7986
rect 10740 8032 10828 8072
rect 10740 7986 10769 8032
rect 10815 7986 10828 8032
rect 12015 8084 12088 8097
rect 12015 8072 12029 8084
rect 10740 7908 10828 7986
rect 11124 7992 11212 8005
rect 11124 7946 11137 7992
rect 11183 7946 11212 7992
rect 11124 7933 11212 7946
rect 11332 7992 11467 8005
rect 11332 7946 11392 7992
rect 11438 7946 11467 7992
rect 11332 7933 11467 7946
rect 11587 7992 11675 8005
rect 11587 7946 11616 7992
rect 11662 7946 11675 7992
rect 11587 7933 11675 7946
rect 11747 7982 11835 8072
rect 11747 7936 11760 7982
rect 11806 7936 11835 7982
rect 11747 7908 11835 7936
rect 11955 8038 12029 8072
rect 12075 8038 12088 8084
rect 11955 7908 12088 8038
rect 12168 8084 12240 8097
rect 12168 8038 12181 8084
rect 12227 8038 12240 8084
rect 12168 8005 12240 8038
rect 12168 7933 12300 8005
rect 12420 7992 12524 8005
rect 12420 7946 12449 7992
rect 12495 7946 12524 7992
rect 12420 7933 12524 7946
rect 12644 7992 12748 8005
rect 12644 7946 12673 7992
rect 12719 7946 12748 7992
rect 12644 7933 12748 7946
rect 12868 7992 12956 8005
rect 12868 7946 12897 7992
rect 12943 7946 12956 7992
rect 12868 7933 12956 7946
rect 13556 8032 13644 8072
rect 13556 7986 13569 8032
rect 13615 7986 13644 8032
rect 13556 7908 13644 7986
rect 13764 8032 13852 8072
rect 13764 7986 13793 8032
rect 13839 7986 13852 8032
rect 15151 8084 15224 8097
rect 15151 8072 15165 8084
rect 13764 7908 13852 7986
rect 14260 7992 14348 8005
rect 14260 7946 14273 7992
rect 14319 7946 14348 7992
rect 14260 7933 14348 7946
rect 14468 7992 14603 8005
rect 14468 7946 14528 7992
rect 14574 7946 14603 7992
rect 14468 7933 14603 7946
rect 14723 7992 14811 8005
rect 14723 7946 14752 7992
rect 14798 7946 14811 7992
rect 14723 7933 14811 7946
rect 14883 7982 14971 8072
rect 14883 7936 14896 7982
rect 14942 7936 14971 7982
rect 14883 7908 14971 7936
rect 15091 8038 15165 8072
rect 15211 8038 15224 8084
rect 15091 7908 15224 8038
rect 15304 8084 15376 8097
rect 15304 8038 15317 8084
rect 15363 8038 15376 8084
rect 15304 8005 15376 8038
rect 16388 8032 16476 8072
rect 15304 7933 15436 8005
rect 15556 7992 15660 8005
rect 15556 7946 15585 7992
rect 15631 7946 15660 7992
rect 15556 7933 15660 7946
rect 15780 7992 15884 8005
rect 15780 7946 15809 7992
rect 15855 7946 15884 7992
rect 15780 7933 15884 7946
rect 16004 7992 16092 8005
rect 16004 7946 16033 7992
rect 16079 7946 16092 7992
rect 16004 7933 16092 7946
rect 16388 7986 16401 8032
rect 16447 7986 16476 8032
rect 16388 7908 16476 7986
rect 16596 8032 16684 8072
rect 16596 7986 16625 8032
rect 16671 7986 16684 8032
rect 16596 7908 16684 7986
rect 17396 8032 17484 8072
rect 17396 7986 17409 8032
rect 17455 7986 17484 8032
rect 17396 7908 17484 7986
rect 17604 8032 17692 8072
rect 17604 7986 17633 8032
rect 17679 7986 17692 8032
rect 17604 7908 17692 7986
rect 17844 8032 17932 8072
rect 17844 7986 17857 8032
rect 17903 7986 17932 8032
rect 17844 7908 17932 7986
rect 18132 8032 18220 8072
rect 18132 7986 18161 8032
rect 18207 7986 18220 8032
rect 18132 7908 18220 7986
rect 1716 7694 1804 7772
rect 1716 7648 1729 7694
rect 1775 7648 1804 7694
rect 1716 7608 1804 7648
rect 1924 7694 2012 7772
rect 1924 7648 1953 7694
rect 1999 7648 2012 7694
rect 2388 7734 2476 7747
rect 2388 7688 2401 7734
rect 2447 7688 2476 7734
rect 2388 7675 2476 7688
rect 2596 7734 2700 7747
rect 2596 7688 2625 7734
rect 2671 7688 2700 7734
rect 2596 7675 2700 7688
rect 2820 7734 2924 7747
rect 2820 7688 2849 7734
rect 2895 7688 2924 7734
rect 2820 7675 2924 7688
rect 3044 7675 3176 7747
rect 1924 7608 2012 7648
rect 3104 7642 3176 7675
rect 3104 7596 3117 7642
rect 3163 7596 3176 7642
rect 3104 7583 3176 7596
rect 3256 7642 3389 7772
rect 3256 7596 3269 7642
rect 3315 7608 3389 7642
rect 3509 7744 3597 7772
rect 3509 7698 3538 7744
rect 3584 7698 3597 7744
rect 3509 7608 3597 7698
rect 3669 7734 3757 7747
rect 3669 7688 3682 7734
rect 3728 7688 3757 7734
rect 3669 7675 3757 7688
rect 3877 7734 4012 7747
rect 3877 7688 3906 7734
rect 3952 7688 4012 7734
rect 3877 7675 4012 7688
rect 4132 7734 4220 7747
rect 4132 7688 4161 7734
rect 4207 7688 4220 7734
rect 4132 7675 4220 7688
rect 4596 7694 4684 7772
rect 3315 7596 3329 7608
rect 3256 7583 3329 7596
rect 4596 7648 4609 7694
rect 4655 7648 4684 7694
rect 4596 7608 4684 7648
rect 4804 7694 4892 7772
rect 4804 7648 4833 7694
rect 4879 7648 4892 7694
rect 4804 7608 4892 7648
rect 4964 7694 5052 7772
rect 4964 7648 4977 7694
rect 5023 7648 5052 7694
rect 4964 7608 5052 7648
rect 5252 7694 5340 7772
rect 5252 7648 5281 7694
rect 5327 7648 5340 7694
rect 5252 7608 5340 7648
rect 5412 7694 5500 7772
rect 5412 7648 5425 7694
rect 5471 7648 5500 7694
rect 5412 7608 5500 7648
rect 5700 7694 5788 7772
rect 5700 7648 5729 7694
rect 5775 7648 5788 7694
rect 5700 7608 5788 7648
rect 5860 7694 5948 7772
rect 5860 7648 5873 7694
rect 5919 7648 5948 7694
rect 5860 7608 5948 7648
rect 6148 7694 6236 7772
rect 6148 7648 6177 7694
rect 6223 7648 6236 7694
rect 6148 7608 6236 7648
rect 6308 7694 6396 7772
rect 6308 7648 6321 7694
rect 6367 7648 6396 7694
rect 6308 7608 6396 7648
rect 6596 7694 6684 7772
rect 6596 7648 6625 7694
rect 6671 7648 6684 7694
rect 6596 7608 6684 7648
rect 6756 7694 6844 7772
rect 6756 7648 6769 7694
rect 6815 7648 6844 7694
rect 6756 7608 6844 7648
rect 7044 7694 7132 7772
rect 7044 7648 7073 7694
rect 7119 7648 7132 7694
rect 7204 7734 7292 7747
rect 7204 7688 7217 7734
rect 7263 7688 7292 7734
rect 7204 7675 7292 7688
rect 7412 7734 7516 7747
rect 7412 7688 7441 7734
rect 7487 7688 7516 7734
rect 7412 7675 7516 7688
rect 7636 7734 7740 7747
rect 7636 7688 7665 7734
rect 7711 7688 7740 7734
rect 7636 7675 7740 7688
rect 7860 7675 7992 7747
rect 7044 7608 7132 7648
rect 7920 7642 7992 7675
rect 7920 7596 7933 7642
rect 7979 7596 7992 7642
rect 7920 7583 7992 7596
rect 8072 7642 8205 7772
rect 8072 7596 8085 7642
rect 8131 7608 8205 7642
rect 8325 7744 8413 7772
rect 8325 7698 8354 7744
rect 8400 7698 8413 7744
rect 8325 7608 8413 7698
rect 8485 7734 8573 7747
rect 8485 7688 8498 7734
rect 8544 7688 8573 7734
rect 8485 7675 8573 7688
rect 8693 7734 8828 7747
rect 8693 7688 8722 7734
rect 8768 7688 8828 7734
rect 8693 7675 8828 7688
rect 8948 7734 9036 7747
rect 8948 7688 8977 7734
rect 9023 7688 9036 7734
rect 8948 7675 9036 7688
rect 8131 7596 8145 7608
rect 8072 7583 8145 7596
rect 9556 7694 9644 7772
rect 9556 7648 9569 7694
rect 9615 7648 9644 7694
rect 9556 7608 9644 7648
rect 9844 7694 9932 7772
rect 9844 7648 9873 7694
rect 9919 7648 9932 7694
rect 9844 7608 9932 7648
rect 10004 7694 10092 7772
rect 10004 7648 10017 7694
rect 10063 7648 10092 7694
rect 10004 7608 10092 7648
rect 10212 7694 10300 7772
rect 10212 7648 10241 7694
rect 10287 7648 10300 7694
rect 10212 7608 10300 7648
rect 10676 7694 10764 7772
rect 10676 7648 10689 7694
rect 10735 7648 10764 7694
rect 10676 7608 10764 7648
rect 10884 7694 10972 7772
rect 10884 7648 10913 7694
rect 10959 7648 10972 7694
rect 10884 7608 10972 7648
rect 11348 7694 11436 7772
rect 11348 7648 11361 7694
rect 11407 7648 11436 7694
rect 11348 7608 11436 7648
rect 11556 7694 11644 7772
rect 11556 7648 11585 7694
rect 11631 7648 11644 7694
rect 12020 7734 12108 7747
rect 12020 7688 12033 7734
rect 12079 7688 12108 7734
rect 12020 7675 12108 7688
rect 12228 7734 12332 7747
rect 12228 7688 12257 7734
rect 12303 7688 12332 7734
rect 12228 7675 12332 7688
rect 12452 7734 12556 7747
rect 12452 7688 12481 7734
rect 12527 7688 12556 7734
rect 12452 7675 12556 7688
rect 12676 7675 12808 7747
rect 11556 7608 11644 7648
rect 12736 7642 12808 7675
rect 12736 7596 12749 7642
rect 12795 7596 12808 7642
rect 12736 7583 12808 7596
rect 12888 7642 13021 7772
rect 12888 7596 12901 7642
rect 12947 7608 13021 7642
rect 13141 7744 13229 7772
rect 13141 7698 13170 7744
rect 13216 7698 13229 7744
rect 13141 7608 13229 7698
rect 13301 7734 13389 7747
rect 13301 7688 13314 7734
rect 13360 7688 13389 7734
rect 13301 7675 13389 7688
rect 13509 7734 13644 7747
rect 13509 7688 13538 7734
rect 13584 7688 13644 7734
rect 13509 7675 13644 7688
rect 13764 7734 13852 7747
rect 13764 7688 13793 7734
rect 13839 7688 13852 7734
rect 13764 7675 13852 7688
rect 13924 7694 14012 7772
rect 12947 7596 12961 7608
rect 12888 7583 12961 7596
rect 13924 7648 13937 7694
rect 13983 7648 14012 7694
rect 13924 7608 14012 7648
rect 14212 7694 14300 7772
rect 14212 7648 14241 7694
rect 14287 7648 14300 7694
rect 14372 7734 14460 7747
rect 14372 7688 14385 7734
rect 14431 7688 14460 7734
rect 14372 7675 14460 7688
rect 14580 7734 14715 7747
rect 14580 7688 14640 7734
rect 14686 7688 14715 7734
rect 14580 7675 14715 7688
rect 14835 7734 14923 7747
rect 14835 7688 14864 7734
rect 14910 7688 14923 7734
rect 14835 7675 14923 7688
rect 14995 7744 15083 7772
rect 14995 7698 15008 7744
rect 15054 7698 15083 7744
rect 14212 7608 14300 7648
rect 14995 7608 15083 7698
rect 15203 7642 15336 7772
rect 15203 7608 15277 7642
rect 15263 7596 15277 7608
rect 15323 7596 15336 7642
rect 15263 7583 15336 7596
rect 15416 7675 15548 7747
rect 15668 7734 15772 7747
rect 15668 7688 15697 7734
rect 15743 7688 15772 7734
rect 15668 7675 15772 7688
rect 15892 7734 15996 7747
rect 15892 7688 15921 7734
rect 15967 7688 15996 7734
rect 15892 7675 15996 7688
rect 16116 7734 16204 7747
rect 16116 7688 16145 7734
rect 16191 7688 16204 7734
rect 16116 7675 16204 7688
rect 16500 7694 16588 7772
rect 15416 7642 15488 7675
rect 15416 7596 15429 7642
rect 15475 7596 15488 7642
rect 15416 7583 15488 7596
rect 16500 7648 16513 7694
rect 16559 7648 16588 7694
rect 16500 7608 16588 7648
rect 16708 7694 16796 7772
rect 16708 7648 16737 7694
rect 16783 7648 16796 7694
rect 16708 7608 16796 7648
rect 17620 7694 17708 7772
rect 17620 7648 17633 7694
rect 17679 7648 17708 7694
rect 17620 7608 17708 7648
rect 17828 7694 17916 7772
rect 17828 7648 17857 7694
rect 17903 7648 17916 7694
rect 17828 7608 17916 7648
rect 1604 6464 1692 6504
rect 1604 6418 1617 6464
rect 1663 6418 1692 6464
rect 1604 6340 1692 6418
rect 1892 6464 1980 6504
rect 1892 6418 1921 6464
rect 1967 6418 1980 6464
rect 1892 6340 1980 6418
rect 2073 6464 2161 6504
rect 2073 6418 2086 6464
rect 2132 6418 2161 6464
rect 2073 6340 2161 6418
rect 2281 6437 2361 6504
rect 3208 6448 3296 6504
rect 2281 6423 2433 6437
rect 2281 6377 2310 6423
rect 2356 6377 2433 6423
rect 2281 6365 2433 6377
rect 2553 6424 2657 6437
rect 2553 6378 2582 6424
rect 2628 6378 2657 6424
rect 2553 6365 2657 6378
rect 2777 6424 2865 6437
rect 2777 6378 2806 6424
rect 2852 6378 2865 6424
rect 2777 6365 2865 6378
rect 3208 6402 3221 6448
rect 3267 6402 3296 6448
rect 2281 6340 2361 6365
rect 3208 6340 3296 6402
rect 3416 6432 3564 6504
rect 3684 6491 3772 6504
rect 3684 6445 3713 6491
rect 3759 6445 3772 6491
rect 3684 6432 3772 6445
rect 3844 6464 3932 6504
rect 3416 6386 3445 6432
rect 3491 6386 3504 6432
rect 3844 6418 3857 6464
rect 3903 6418 3932 6464
rect 3416 6340 3504 6386
rect 3844 6340 3932 6418
rect 4132 6464 4220 6504
rect 4132 6418 4161 6464
rect 4207 6418 4220 6464
rect 4132 6340 4220 6418
rect 4292 6464 4380 6504
rect 4292 6418 4305 6464
rect 4351 6418 4380 6464
rect 4292 6340 4380 6418
rect 4580 6464 4668 6504
rect 4580 6418 4609 6464
rect 4655 6418 4668 6464
rect 4580 6340 4668 6418
rect 4740 6464 4828 6504
rect 4740 6418 4753 6464
rect 4799 6418 4828 6464
rect 4740 6340 4828 6418
rect 5028 6464 5116 6504
rect 5028 6418 5057 6464
rect 5103 6418 5116 6464
rect 5028 6340 5116 6418
rect 5524 6464 5612 6504
rect 5524 6418 5537 6464
rect 5583 6418 5612 6464
rect 5524 6340 5612 6418
rect 5812 6464 5900 6504
rect 5812 6418 5841 6464
rect 5887 6418 5900 6464
rect 5812 6340 5900 6418
rect 5972 6464 6060 6504
rect 5972 6418 5985 6464
rect 6031 6418 6060 6464
rect 5972 6340 6060 6418
rect 6260 6464 6348 6504
rect 6260 6418 6289 6464
rect 6335 6418 6348 6464
rect 6260 6340 6348 6418
rect 6835 6447 6923 6504
rect 6835 6401 6848 6447
rect 6894 6401 6923 6447
rect 6835 6340 6923 6401
rect 7043 6444 7131 6504
rect 7043 6398 7072 6444
rect 7118 6398 7131 6444
rect 7043 6340 7131 6398
rect 7428 6464 7516 6504
rect 7428 6418 7441 6464
rect 7487 6418 7516 6464
rect 7428 6340 7516 6418
rect 7636 6464 7724 6504
rect 7636 6418 7665 6464
rect 7711 6418 7724 6464
rect 7636 6340 7724 6418
rect 8100 6464 8188 6504
rect 8100 6418 8113 6464
rect 8159 6418 8188 6464
rect 8100 6340 8188 6418
rect 8308 6464 8396 6504
rect 8308 6418 8337 6464
rect 8383 6418 8396 6464
rect 8308 6340 8396 6418
rect 8772 6464 8860 6504
rect 8772 6418 8785 6464
rect 8831 6418 8860 6464
rect 8772 6340 8860 6418
rect 8980 6464 9068 6504
rect 8980 6418 9009 6464
rect 9055 6418 9068 6464
rect 8980 6340 9068 6418
rect 9444 6464 9532 6504
rect 9444 6418 9457 6464
rect 9503 6418 9532 6464
rect 9444 6340 9532 6418
rect 9652 6464 9740 6504
rect 9652 6418 9681 6464
rect 9727 6418 9740 6464
rect 9652 6340 9740 6418
rect 10116 6464 10204 6504
rect 10116 6418 10129 6464
rect 10175 6418 10204 6464
rect 10116 6340 10204 6418
rect 10324 6464 10412 6504
rect 10324 6418 10353 6464
rect 10399 6418 10412 6464
rect 10324 6340 10412 6418
rect 10788 6464 10876 6504
rect 10788 6418 10801 6464
rect 10847 6418 10876 6464
rect 10788 6340 10876 6418
rect 10996 6464 11084 6504
rect 10996 6418 11025 6464
rect 11071 6418 11084 6464
rect 10996 6340 11084 6418
rect 11460 6464 11548 6504
rect 11460 6418 11473 6464
rect 11519 6418 11548 6464
rect 11460 6340 11548 6418
rect 11668 6464 11756 6504
rect 11668 6418 11697 6464
rect 11743 6418 11756 6464
rect 11668 6340 11756 6418
rect 12132 6464 12220 6504
rect 12132 6418 12145 6464
rect 12191 6418 12220 6464
rect 12132 6340 12220 6418
rect 12340 6464 12428 6504
rect 12340 6418 12369 6464
rect 12415 6418 12428 6464
rect 12340 6340 12428 6418
rect 12580 6464 12668 6504
rect 12580 6418 12593 6464
rect 12639 6418 12668 6464
rect 12580 6340 12668 6418
rect 12868 6464 12956 6504
rect 12868 6418 12897 6464
rect 12943 6418 12956 6464
rect 12868 6340 12956 6418
rect 13588 6464 13676 6504
rect 13588 6418 13601 6464
rect 13647 6418 13676 6464
rect 13588 6340 13676 6418
rect 13796 6464 13884 6504
rect 13796 6418 13825 6464
rect 13871 6418 13884 6464
rect 13796 6340 13884 6418
rect 14260 6464 14348 6504
rect 14260 6418 14273 6464
rect 14319 6418 14348 6464
rect 14260 6340 14348 6418
rect 14468 6464 14556 6504
rect 14468 6418 14497 6464
rect 14543 6418 14556 6464
rect 14468 6340 14556 6418
rect 14932 6464 15020 6504
rect 14932 6418 14945 6464
rect 14991 6418 15020 6464
rect 14932 6340 15020 6418
rect 15140 6464 15228 6504
rect 15140 6418 15169 6464
rect 15215 6418 15228 6464
rect 15140 6340 15228 6418
rect 15604 6464 15692 6504
rect 15604 6418 15617 6464
rect 15663 6418 15692 6464
rect 15604 6340 15692 6418
rect 15812 6464 15900 6504
rect 15812 6418 15841 6464
rect 15887 6418 15900 6464
rect 15812 6340 15900 6418
rect 16276 6464 16364 6504
rect 16276 6418 16289 6464
rect 16335 6418 16364 6464
rect 16276 6340 16364 6418
rect 16484 6464 16572 6504
rect 16484 6418 16513 6464
rect 16559 6418 16572 6464
rect 16484 6340 16572 6418
rect 16948 6464 17036 6504
rect 16948 6418 16961 6464
rect 17007 6418 17036 6464
rect 16948 6340 17036 6418
rect 17156 6464 17244 6504
rect 17156 6418 17185 6464
rect 17231 6418 17244 6464
rect 17156 6340 17244 6418
rect 17620 6464 17708 6504
rect 17620 6418 17633 6464
rect 17679 6418 17708 6464
rect 17620 6340 17708 6418
rect 17828 6464 17916 6504
rect 17828 6418 17857 6464
rect 17903 6418 17916 6464
rect 17828 6340 17916 6418
rect 2168 6176 2256 6203
rect 2168 6130 2181 6176
rect 2227 6130 2256 6176
rect 2168 6113 2256 6130
rect 1716 6100 1804 6113
rect 1716 6054 1729 6100
rect 1775 6054 1804 6100
rect 1716 6040 1804 6054
rect 1924 6040 1988 6113
rect 2108 6040 2256 6113
rect 2376 6100 2464 6203
rect 2376 6054 2405 6100
rect 2451 6054 2464 6100
rect 2376 6040 2464 6054
rect 2836 6126 2924 6204
rect 2836 6080 2849 6126
rect 2895 6080 2924 6126
rect 2836 6040 2924 6080
rect 3044 6126 3132 6204
rect 3044 6080 3073 6126
rect 3119 6080 3132 6126
rect 3044 6040 3132 6080
rect 3284 6126 3372 6204
rect 3284 6080 3297 6126
rect 3343 6080 3372 6126
rect 3284 6040 3372 6080
rect 3572 6126 3660 6204
rect 3572 6080 3601 6126
rect 3647 6080 3660 6126
rect 3572 6040 3660 6080
rect 3732 6126 3820 6204
rect 3732 6080 3745 6126
rect 3791 6080 3820 6126
rect 3732 6040 3820 6080
rect 4020 6126 4108 6204
rect 4020 6080 4049 6126
rect 4095 6080 4108 6126
rect 4020 6040 4108 6080
rect 4180 6126 4268 6204
rect 4180 6080 4193 6126
rect 4239 6080 4268 6126
rect 4180 6040 4268 6080
rect 4468 6126 4556 6204
rect 4468 6080 4497 6126
rect 4543 6080 4556 6126
rect 4468 6040 4556 6080
rect 4628 6126 4716 6204
rect 4628 6080 4641 6126
rect 4687 6080 4716 6126
rect 4628 6040 4716 6080
rect 4916 6126 5004 6204
rect 4916 6080 4945 6126
rect 4991 6080 5004 6126
rect 4916 6040 5004 6080
rect 5413 6146 5501 6204
rect 5413 6100 5426 6146
rect 5472 6100 5501 6146
rect 5413 6040 5501 6100
rect 5621 6143 5709 6204
rect 5621 6097 5650 6143
rect 5696 6097 5709 6143
rect 5621 6040 5709 6097
rect 6164 6126 6252 6204
rect 6164 6080 6177 6126
rect 6223 6080 6252 6126
rect 6164 6040 6252 6080
rect 6372 6126 6460 6204
rect 6372 6080 6401 6126
rect 6447 6080 6460 6126
rect 6372 6040 6460 6080
rect 6836 6126 6924 6204
rect 6836 6080 6849 6126
rect 6895 6080 6924 6126
rect 6836 6040 6924 6080
rect 7044 6126 7132 6204
rect 7044 6080 7073 6126
rect 7119 6080 7132 6126
rect 7044 6040 7132 6080
rect 7428 6126 7516 6204
rect 7428 6080 7441 6126
rect 7487 6080 7516 6126
rect 7428 6040 7516 6080
rect 7636 6126 7724 6204
rect 7636 6080 7665 6126
rect 7711 6080 7724 6126
rect 7636 6040 7724 6080
rect 8101 6146 8189 6204
rect 8101 6100 8114 6146
rect 8160 6100 8189 6146
rect 8101 6040 8189 6100
rect 8309 6143 8397 6204
rect 8309 6097 8338 6143
rect 8384 6097 8397 6143
rect 8309 6040 8397 6097
rect 8772 6126 8860 6204
rect 8772 6080 8785 6126
rect 8831 6080 8860 6126
rect 8772 6040 8860 6080
rect 8980 6126 9068 6204
rect 8980 6080 9009 6126
rect 9055 6080 9068 6126
rect 8980 6040 9068 6080
rect 9556 6126 9644 6204
rect 9556 6080 9569 6126
rect 9615 6080 9644 6126
rect 9556 6040 9644 6080
rect 9844 6126 9932 6204
rect 9844 6080 9873 6126
rect 9919 6080 9932 6126
rect 9844 6040 9932 6080
rect 10228 6126 10316 6204
rect 10228 6080 10241 6126
rect 10287 6080 10316 6126
rect 10228 6040 10316 6080
rect 10436 6126 10524 6204
rect 10436 6080 10465 6126
rect 10511 6080 10524 6126
rect 10436 6040 10524 6080
rect 10900 6126 10988 6204
rect 10900 6080 10913 6126
rect 10959 6080 10988 6126
rect 10900 6040 10988 6080
rect 11108 6126 11196 6204
rect 11108 6080 11137 6126
rect 11183 6080 11196 6126
rect 11108 6040 11196 6080
rect 11572 6126 11660 6204
rect 11572 6080 11585 6126
rect 11631 6080 11660 6126
rect 11572 6040 11660 6080
rect 11780 6126 11868 6204
rect 11780 6080 11809 6126
rect 11855 6080 11868 6126
rect 11780 6040 11868 6080
rect 12244 6126 12332 6204
rect 12244 6080 12257 6126
rect 12303 6080 12332 6126
rect 12244 6040 12332 6080
rect 12452 6126 12540 6204
rect 12452 6080 12481 6126
rect 12527 6080 12540 6126
rect 12452 6040 12540 6080
rect 12916 6126 13004 6204
rect 12916 6080 12929 6126
rect 12975 6080 13004 6126
rect 12916 6040 13004 6080
rect 13124 6126 13212 6204
rect 13124 6080 13153 6126
rect 13199 6080 13212 6126
rect 13124 6040 13212 6080
rect 13588 6126 13676 6204
rect 13588 6080 13601 6126
rect 13647 6080 13676 6126
rect 13588 6040 13676 6080
rect 13796 6126 13884 6204
rect 13796 6080 13825 6126
rect 13871 6080 13884 6126
rect 13796 6040 13884 6080
rect 14260 6126 14348 6204
rect 14260 6080 14273 6126
rect 14319 6080 14348 6126
rect 14260 6040 14348 6080
rect 14468 6126 14556 6204
rect 14468 6080 14497 6126
rect 14543 6080 14556 6126
rect 14468 6040 14556 6080
rect 14932 6126 15020 6204
rect 14932 6080 14945 6126
rect 14991 6080 15020 6126
rect 14932 6040 15020 6080
rect 15140 6126 15228 6204
rect 15140 6080 15169 6126
rect 15215 6080 15228 6126
rect 15140 6040 15228 6080
rect 15604 6126 15692 6204
rect 15604 6080 15617 6126
rect 15663 6080 15692 6126
rect 15604 6040 15692 6080
rect 15812 6126 15900 6204
rect 15812 6080 15841 6126
rect 15887 6080 15900 6126
rect 15812 6040 15900 6080
rect 16277 6146 16365 6204
rect 16277 6100 16290 6146
rect 16336 6100 16365 6146
rect 16277 6040 16365 6100
rect 16485 6143 16573 6204
rect 16485 6097 16514 6143
rect 16560 6097 16573 6143
rect 16485 6040 16573 6097
rect 16724 6126 16812 6204
rect 16724 6080 16737 6126
rect 16783 6080 16812 6126
rect 16724 6040 16812 6080
rect 17012 6126 17100 6204
rect 17012 6080 17041 6126
rect 17087 6080 17100 6126
rect 17012 6040 17100 6080
rect 17699 6143 17787 6204
rect 17699 6097 17712 6143
rect 17758 6097 17787 6143
rect 17699 6040 17787 6097
rect 17907 6146 17995 6204
rect 17907 6100 17936 6146
rect 17982 6100 17995 6146
rect 17907 6040 17995 6100
rect 1604 4896 1692 4936
rect 1604 4850 1617 4896
rect 1663 4850 1692 4896
rect 1604 4772 1692 4850
rect 1892 4896 1980 4936
rect 1892 4850 1921 4896
rect 1967 4850 1980 4896
rect 1892 4772 1980 4850
rect 2052 4896 2140 4936
rect 2052 4850 2065 4896
rect 2111 4850 2140 4896
rect 2052 4772 2140 4850
rect 2340 4896 2428 4936
rect 2340 4850 2369 4896
rect 2415 4850 2428 4896
rect 2340 4772 2428 4850
rect 2500 4896 2588 4936
rect 2500 4850 2513 4896
rect 2559 4850 2588 4896
rect 2500 4772 2588 4850
rect 2788 4896 2876 4936
rect 2788 4850 2817 4896
rect 2863 4850 2876 4896
rect 2788 4772 2876 4850
rect 2948 4896 3036 4936
rect 2948 4850 2961 4896
rect 3007 4850 3036 4896
rect 2948 4772 3036 4850
rect 3236 4896 3324 4936
rect 3236 4850 3265 4896
rect 3311 4850 3324 4896
rect 3236 4772 3324 4850
rect 3396 4896 3484 4936
rect 3396 4850 3409 4896
rect 3455 4850 3484 4896
rect 3396 4772 3484 4850
rect 3684 4896 3772 4936
rect 3684 4850 3713 4896
rect 3759 4850 3772 4896
rect 3684 4772 3772 4850
rect 4069 4876 4157 4936
rect 4069 4830 4082 4876
rect 4128 4830 4157 4876
rect 4069 4772 4157 4830
rect 4277 4879 4365 4936
rect 4277 4833 4306 4879
rect 4352 4833 4365 4879
rect 4277 4772 4365 4833
rect 4741 4876 4829 4936
rect 4741 4830 4754 4876
rect 4800 4830 4829 4876
rect 4741 4772 4829 4830
rect 4949 4879 5037 4936
rect 4949 4833 4978 4879
rect 5024 4833 5037 4879
rect 4949 4772 5037 4833
rect 5524 4896 5612 4936
rect 5524 4850 5537 4896
rect 5583 4850 5612 4896
rect 5524 4772 5612 4850
rect 5812 4896 5900 4936
rect 5812 4850 5841 4896
rect 5887 4850 5900 4896
rect 5812 4772 5900 4850
rect 6197 4876 6285 4936
rect 6197 4830 6210 4876
rect 6256 4830 6285 4876
rect 6197 4772 6285 4830
rect 6405 4879 6493 4936
rect 6405 4833 6434 4879
rect 6480 4833 6493 4879
rect 6405 4772 6493 4833
rect 6947 4879 7035 4936
rect 6947 4833 6960 4879
rect 7006 4833 7035 4879
rect 6947 4772 7035 4833
rect 7155 4876 7243 4936
rect 7155 4830 7184 4876
rect 7230 4830 7243 4876
rect 7155 4772 7243 4830
rect 7620 4896 7708 4936
rect 7620 4850 7633 4896
rect 7679 4850 7708 4896
rect 7620 4772 7708 4850
rect 7828 4896 7916 4936
rect 7828 4850 7857 4896
rect 7903 4850 7916 4896
rect 7828 4772 7916 4850
rect 8213 4876 8301 4936
rect 8213 4830 8226 4876
rect 8272 4830 8301 4876
rect 8213 4772 8301 4830
rect 8421 4879 8509 4936
rect 8421 4833 8450 4879
rect 8496 4833 8509 4879
rect 8421 4772 8509 4833
rect 8884 4896 8972 4936
rect 8884 4850 8897 4896
rect 8943 4850 8972 4896
rect 8884 4772 8972 4850
rect 9092 4896 9180 4936
rect 9092 4850 9121 4896
rect 9167 4850 9180 4896
rect 9092 4772 9180 4850
rect 9556 4896 9644 4936
rect 9556 4850 9569 4896
rect 9615 4850 9644 4896
rect 9556 4772 9644 4850
rect 9764 4896 9852 4936
rect 9764 4850 9793 4896
rect 9839 4850 9852 4896
rect 9764 4772 9852 4850
rect 10228 4896 10316 4936
rect 10228 4850 10241 4896
rect 10287 4850 10316 4896
rect 10228 4772 10316 4850
rect 10436 4896 10524 4936
rect 10436 4850 10465 4896
rect 10511 4850 10524 4896
rect 10436 4772 10524 4850
rect 10900 4896 10988 4936
rect 10900 4850 10913 4896
rect 10959 4850 10988 4896
rect 10900 4772 10988 4850
rect 11108 4896 11196 4936
rect 11108 4850 11137 4896
rect 11183 4850 11196 4896
rect 11108 4772 11196 4850
rect 11572 4896 11660 4936
rect 11572 4850 11585 4896
rect 11631 4850 11660 4896
rect 11572 4772 11660 4850
rect 11780 4896 11868 4936
rect 11780 4850 11809 4896
rect 11855 4850 11868 4896
rect 11780 4772 11868 4850
rect 12244 4896 12332 4936
rect 12244 4850 12257 4896
rect 12303 4850 12332 4896
rect 12244 4772 12332 4850
rect 12452 4896 12540 4936
rect 12452 4850 12481 4896
rect 12527 4850 12540 4896
rect 12452 4772 12540 4850
rect 12692 4896 12780 4936
rect 12692 4850 12705 4896
rect 12751 4850 12780 4896
rect 12692 4772 12780 4850
rect 12980 4896 13068 4936
rect 12980 4850 13009 4896
rect 13055 4850 13068 4896
rect 12980 4772 13068 4850
rect 13588 4896 13676 4936
rect 13588 4850 13601 4896
rect 13647 4850 13676 4896
rect 13588 4772 13676 4850
rect 13796 4896 13884 4936
rect 13796 4850 13825 4896
rect 13871 4850 13884 4896
rect 13796 4772 13884 4850
rect 14260 4896 14348 4936
rect 14260 4850 14273 4896
rect 14319 4850 14348 4896
rect 14260 4772 14348 4850
rect 14468 4896 14556 4936
rect 14468 4850 14497 4896
rect 14543 4850 14556 4896
rect 14468 4772 14556 4850
rect 15012 4896 15100 4936
rect 15012 4850 15025 4896
rect 15071 4850 15100 4896
rect 15012 4772 15100 4850
rect 15220 4896 15308 4936
rect 15220 4850 15249 4896
rect 15295 4850 15308 4896
rect 15220 4772 15308 4850
rect 15683 4879 15771 4936
rect 15683 4833 15696 4879
rect 15742 4833 15771 4879
rect 15683 4772 15771 4833
rect 15891 4876 15979 4936
rect 15891 4830 15920 4876
rect 15966 4830 15979 4876
rect 17279 4948 17352 4961
rect 17279 4936 17293 4948
rect 15891 4772 15979 4830
rect 16388 4856 16476 4869
rect 16388 4810 16401 4856
rect 16447 4810 16476 4856
rect 16388 4797 16476 4810
rect 16596 4856 16731 4869
rect 16596 4810 16656 4856
rect 16702 4810 16731 4856
rect 16596 4797 16731 4810
rect 16851 4856 16939 4869
rect 16851 4810 16880 4856
rect 16926 4810 16939 4856
rect 16851 4797 16939 4810
rect 17011 4846 17099 4936
rect 17011 4800 17024 4846
rect 17070 4800 17099 4846
rect 17011 4772 17099 4800
rect 17219 4902 17293 4936
rect 17339 4902 17352 4948
rect 17219 4772 17352 4902
rect 17432 4948 17504 4961
rect 17432 4902 17445 4948
rect 17491 4902 17504 4948
rect 17432 4869 17504 4902
rect 17432 4797 17564 4869
rect 17684 4856 17788 4869
rect 17684 4810 17713 4856
rect 17759 4810 17788 4856
rect 17684 4797 17788 4810
rect 17908 4856 18012 4869
rect 17908 4810 17937 4856
rect 17983 4810 18012 4856
rect 17908 4797 18012 4810
rect 18132 4856 18220 4869
rect 18132 4810 18161 4856
rect 18207 4810 18220 4856
rect 18132 4797 18220 4810
rect 1604 4558 1692 4636
rect 1604 4512 1617 4558
rect 1663 4512 1692 4558
rect 1604 4472 1692 4512
rect 1892 4558 1980 4636
rect 1892 4512 1921 4558
rect 1967 4512 1980 4558
rect 1892 4472 1980 4512
rect 2052 4558 2140 4636
rect 2052 4512 2065 4558
rect 2111 4512 2140 4558
rect 2052 4472 2140 4512
rect 2340 4558 2428 4636
rect 2340 4512 2369 4558
rect 2415 4512 2428 4558
rect 2612 4598 2700 4611
rect 2612 4552 2625 4598
rect 2671 4552 2700 4598
rect 2612 4539 2700 4552
rect 2820 4598 2924 4611
rect 2820 4552 2849 4598
rect 2895 4552 2924 4598
rect 2820 4539 2924 4552
rect 3044 4598 3148 4611
rect 3044 4552 3073 4598
rect 3119 4552 3148 4598
rect 3044 4539 3148 4552
rect 3268 4539 3400 4611
rect 2340 4472 2428 4512
rect 3328 4506 3400 4539
rect 3328 4460 3341 4506
rect 3387 4460 3400 4506
rect 3328 4447 3400 4460
rect 3480 4506 3613 4636
rect 3480 4460 3493 4506
rect 3539 4472 3613 4506
rect 3733 4608 3821 4636
rect 3733 4562 3762 4608
rect 3808 4562 3821 4608
rect 3733 4472 3821 4562
rect 3893 4598 3981 4611
rect 3893 4552 3906 4598
rect 3952 4552 3981 4598
rect 3893 4539 3981 4552
rect 4101 4598 4236 4611
rect 4101 4552 4130 4598
rect 4176 4552 4236 4598
rect 4101 4539 4236 4552
rect 4356 4598 4444 4611
rect 4356 4552 4385 4598
rect 4431 4552 4444 4598
rect 4356 4539 4444 4552
rect 4516 4558 4604 4636
rect 3539 4460 3553 4472
rect 3480 4447 3553 4460
rect 4516 4512 4529 4558
rect 4575 4512 4604 4558
rect 4516 4472 4604 4512
rect 4804 4558 4892 4636
rect 4804 4512 4833 4558
rect 4879 4512 4892 4558
rect 4804 4472 4892 4512
rect 5077 4578 5165 4636
rect 5077 4532 5090 4578
rect 5136 4532 5165 4578
rect 5077 4472 5165 4532
rect 5285 4575 5373 4636
rect 5285 4529 5314 4575
rect 5360 4529 5373 4575
rect 5285 4472 5373 4529
rect 5749 4578 5837 4636
rect 5749 4532 5762 4578
rect 5808 4532 5837 4578
rect 5749 4472 5837 4532
rect 5957 4575 6045 4636
rect 5957 4529 5986 4575
rect 6032 4529 6045 4575
rect 5957 4472 6045 4529
rect 6421 4578 6509 4636
rect 6421 4532 6434 4578
rect 6480 4532 6509 4578
rect 6421 4472 6509 4532
rect 6629 4575 6717 4636
rect 6629 4529 6658 4575
rect 6704 4529 6717 4575
rect 7092 4598 7180 4611
rect 7092 4552 7105 4598
rect 7151 4552 7180 4598
rect 7092 4539 7180 4552
rect 7300 4598 7435 4611
rect 7300 4552 7360 4598
rect 7406 4552 7435 4598
rect 7300 4539 7435 4552
rect 7555 4598 7643 4611
rect 7555 4552 7584 4598
rect 7630 4552 7643 4598
rect 7555 4539 7643 4552
rect 7715 4608 7803 4636
rect 7715 4562 7728 4608
rect 7774 4562 7803 4608
rect 6629 4472 6717 4529
rect 7715 4472 7803 4562
rect 7923 4506 8056 4636
rect 7923 4472 7997 4506
rect 7983 4460 7997 4472
rect 8043 4460 8056 4506
rect 7983 4447 8056 4460
rect 8136 4539 8268 4611
rect 8388 4598 8492 4611
rect 8388 4552 8417 4598
rect 8463 4552 8492 4598
rect 8388 4539 8492 4552
rect 8612 4598 8716 4611
rect 8612 4552 8641 4598
rect 8687 4552 8716 4598
rect 8612 4539 8716 4552
rect 8836 4598 8924 4611
rect 8836 4552 8865 4598
rect 8911 4552 8924 4598
rect 8836 4539 8924 4552
rect 8136 4506 8208 4539
rect 8136 4460 8149 4506
rect 8195 4460 8208 4506
rect 8136 4447 8208 4460
rect 9556 4558 9644 4636
rect 9556 4512 9569 4558
rect 9615 4512 9644 4558
rect 9556 4472 9644 4512
rect 9844 4558 9932 4636
rect 9844 4512 9873 4558
rect 9919 4512 9932 4558
rect 9844 4472 9932 4512
rect 10005 4578 10093 4636
rect 10005 4532 10018 4578
rect 10064 4532 10093 4578
rect 10005 4472 10093 4532
rect 10213 4575 10301 4636
rect 10213 4529 10242 4575
rect 10288 4529 10301 4575
rect 10213 4472 10301 4529
rect 10756 4558 10844 4636
rect 10756 4512 10769 4558
rect 10815 4512 10844 4558
rect 10756 4472 10844 4512
rect 10964 4558 11052 4636
rect 10964 4512 10993 4558
rect 11039 4512 11052 4558
rect 10964 4472 11052 4512
rect 11428 4558 11516 4636
rect 11428 4512 11441 4558
rect 11487 4512 11516 4558
rect 11428 4472 11516 4512
rect 11636 4558 11724 4636
rect 11636 4512 11665 4558
rect 11711 4512 11724 4558
rect 12020 4598 12108 4611
rect 12020 4552 12033 4598
rect 12079 4552 12108 4598
rect 12020 4539 12108 4552
rect 12228 4598 12363 4611
rect 12228 4552 12288 4598
rect 12334 4552 12363 4598
rect 12228 4539 12363 4552
rect 12483 4598 12571 4611
rect 12483 4552 12512 4598
rect 12558 4552 12571 4598
rect 12483 4539 12571 4552
rect 12643 4608 12731 4636
rect 12643 4562 12656 4608
rect 12702 4562 12731 4608
rect 11636 4472 11724 4512
rect 12643 4472 12731 4562
rect 12851 4506 12984 4636
rect 12851 4472 12925 4506
rect 12911 4460 12925 4472
rect 12971 4460 12984 4506
rect 12911 4447 12984 4460
rect 13064 4539 13196 4611
rect 13316 4598 13420 4611
rect 13316 4552 13345 4598
rect 13391 4552 13420 4598
rect 13316 4539 13420 4552
rect 13540 4598 13644 4611
rect 13540 4552 13569 4598
rect 13615 4552 13644 4598
rect 13540 4539 13644 4552
rect 13764 4598 13852 4611
rect 13764 4552 13793 4598
rect 13839 4552 13852 4598
rect 13764 4539 13852 4552
rect 14149 4578 14237 4636
rect 13064 4506 13136 4539
rect 13064 4460 13077 4506
rect 13123 4460 13136 4506
rect 13064 4447 13136 4460
rect 14149 4532 14162 4578
rect 14208 4532 14237 4578
rect 14149 4472 14237 4532
rect 14357 4575 14445 4636
rect 14357 4529 14386 4575
rect 14432 4529 14445 4575
rect 14357 4472 14445 4529
rect 14820 4558 14908 4636
rect 14820 4512 14833 4558
rect 14879 4512 14908 4558
rect 14820 4472 14908 4512
rect 15028 4558 15116 4636
rect 15028 4512 15057 4558
rect 15103 4512 15116 4558
rect 15028 4472 15116 4512
rect 15492 4558 15580 4636
rect 15492 4512 15505 4558
rect 15551 4512 15580 4558
rect 15492 4472 15580 4512
rect 15700 4558 15788 4636
rect 15700 4512 15729 4558
rect 15775 4512 15788 4558
rect 15700 4472 15788 4512
rect 16164 4558 16252 4636
rect 16164 4512 16177 4558
rect 16223 4512 16252 4558
rect 16164 4472 16252 4512
rect 16372 4558 16460 4636
rect 16372 4512 16401 4558
rect 16447 4512 16460 4558
rect 16372 4472 16460 4512
rect 16612 4558 16700 4636
rect 16612 4512 16625 4558
rect 16671 4512 16700 4558
rect 16612 4472 16700 4512
rect 16900 4558 16988 4636
rect 16900 4512 16929 4558
rect 16975 4512 16988 4558
rect 16900 4472 16988 4512
rect 17620 4558 17708 4636
rect 17620 4512 17633 4558
rect 17679 4512 17708 4558
rect 17620 4472 17708 4512
rect 17828 4558 17916 4636
rect 17828 4512 17857 4558
rect 17903 4512 17916 4558
rect 17828 4472 17916 4512
rect 1941 3308 2029 3368
rect 1941 3262 1954 3308
rect 2000 3262 2029 3308
rect 1941 3204 2029 3262
rect 2149 3311 2237 3368
rect 2149 3265 2178 3311
rect 2224 3265 2237 3311
rect 3503 3380 3576 3393
rect 3503 3368 3517 3380
rect 2149 3204 2237 3265
rect 2612 3288 2700 3301
rect 2612 3242 2625 3288
rect 2671 3242 2700 3288
rect 2612 3229 2700 3242
rect 2820 3288 2955 3301
rect 2820 3242 2880 3288
rect 2926 3242 2955 3288
rect 2820 3229 2955 3242
rect 3075 3288 3163 3301
rect 3075 3242 3104 3288
rect 3150 3242 3163 3288
rect 3075 3229 3163 3242
rect 3235 3278 3323 3368
rect 3235 3232 3248 3278
rect 3294 3232 3323 3278
rect 3235 3204 3323 3232
rect 3443 3334 3517 3368
rect 3563 3334 3576 3380
rect 3443 3204 3576 3334
rect 3656 3380 3728 3393
rect 3656 3334 3669 3380
rect 3715 3334 3728 3380
rect 3656 3301 3728 3334
rect 4741 3308 4829 3368
rect 3656 3229 3788 3301
rect 3908 3288 4012 3301
rect 3908 3242 3937 3288
rect 3983 3242 4012 3288
rect 3908 3229 4012 3242
rect 4132 3288 4236 3301
rect 4132 3242 4161 3288
rect 4207 3242 4236 3288
rect 4132 3229 4236 3242
rect 4356 3288 4444 3301
rect 4356 3242 4385 3288
rect 4431 3242 4444 3288
rect 4356 3229 4444 3242
rect 4741 3262 4754 3308
rect 4800 3262 4829 3308
rect 4741 3204 4829 3262
rect 4949 3311 5037 3368
rect 4949 3265 4978 3311
rect 5024 3265 5037 3311
rect 4949 3204 5037 3265
rect 5861 3308 5949 3368
rect 5861 3262 5874 3308
rect 5920 3262 5949 3308
rect 5861 3204 5949 3262
rect 6069 3311 6157 3368
rect 6069 3265 6098 3311
rect 6144 3265 6157 3311
rect 6069 3204 6157 3265
rect 6533 3308 6621 3368
rect 6533 3262 6546 3308
rect 6592 3262 6621 3308
rect 6533 3204 6621 3262
rect 6741 3311 6829 3368
rect 6741 3265 6770 3311
rect 6816 3265 6829 3311
rect 8095 3380 8168 3393
rect 8095 3368 8109 3380
rect 6741 3204 6829 3265
rect 7204 3288 7292 3301
rect 7204 3242 7217 3288
rect 7263 3242 7292 3288
rect 7204 3229 7292 3242
rect 7412 3288 7547 3301
rect 7412 3242 7472 3288
rect 7518 3242 7547 3288
rect 7412 3229 7547 3242
rect 7667 3288 7755 3301
rect 7667 3242 7696 3288
rect 7742 3242 7755 3288
rect 7667 3229 7755 3242
rect 7827 3278 7915 3368
rect 7827 3232 7840 3278
rect 7886 3232 7915 3278
rect 7827 3204 7915 3232
rect 8035 3334 8109 3368
rect 8155 3334 8168 3380
rect 8035 3204 8168 3334
rect 8248 3380 8320 3393
rect 8248 3334 8261 3380
rect 8307 3334 8320 3380
rect 8248 3301 8320 3334
rect 8248 3229 8380 3301
rect 8500 3288 8604 3301
rect 8500 3242 8529 3288
rect 8575 3242 8604 3288
rect 8500 3229 8604 3242
rect 8724 3288 8828 3301
rect 8724 3242 8753 3288
rect 8799 3242 8828 3288
rect 8724 3229 8828 3242
rect 8948 3288 9036 3301
rect 8948 3242 8977 3288
rect 9023 3242 9036 3288
rect 8948 3229 9036 3242
rect 9781 3308 9869 3368
rect 9781 3262 9794 3308
rect 9840 3262 9869 3308
rect 9781 3204 9869 3262
rect 9989 3311 10077 3368
rect 9989 3265 10018 3311
rect 10064 3265 10077 3311
rect 9989 3204 10077 3265
rect 10453 3308 10541 3368
rect 10453 3262 10466 3308
rect 10512 3262 10541 3308
rect 10453 3204 10541 3262
rect 10661 3311 10749 3368
rect 10661 3265 10690 3311
rect 10736 3265 10749 3311
rect 12015 3380 12088 3393
rect 12015 3368 12029 3380
rect 10661 3204 10749 3265
rect 11124 3288 11212 3301
rect 11124 3242 11137 3288
rect 11183 3242 11212 3288
rect 11124 3229 11212 3242
rect 11332 3288 11467 3301
rect 11332 3242 11392 3288
rect 11438 3242 11467 3288
rect 11332 3229 11467 3242
rect 11587 3288 11675 3301
rect 11587 3242 11616 3288
rect 11662 3242 11675 3288
rect 11587 3229 11675 3242
rect 11747 3278 11835 3368
rect 11747 3232 11760 3278
rect 11806 3232 11835 3278
rect 11747 3204 11835 3232
rect 11955 3334 12029 3368
rect 12075 3334 12088 3380
rect 11955 3204 12088 3334
rect 12168 3380 12240 3393
rect 12168 3334 12181 3380
rect 12227 3334 12240 3380
rect 12168 3301 12240 3334
rect 12168 3229 12300 3301
rect 12420 3288 12524 3301
rect 12420 3242 12449 3288
rect 12495 3242 12524 3288
rect 12420 3229 12524 3242
rect 12644 3288 12748 3301
rect 12644 3242 12673 3288
rect 12719 3242 12748 3288
rect 12644 3229 12748 3242
rect 12868 3288 12956 3301
rect 12868 3242 12897 3288
rect 12943 3242 12956 3288
rect 12868 3229 12956 3242
rect 13556 3328 13644 3368
rect 13556 3282 13569 3328
rect 13615 3282 13644 3328
rect 13556 3204 13644 3282
rect 13764 3328 13852 3368
rect 13764 3282 13793 3328
rect 13839 3282 13852 3328
rect 13764 3204 13852 3282
rect 14149 3308 14237 3368
rect 14149 3262 14162 3308
rect 14208 3262 14237 3308
rect 14149 3204 14237 3262
rect 14357 3311 14445 3368
rect 14357 3265 14386 3311
rect 14432 3265 14445 3311
rect 14357 3204 14445 3265
rect 14596 3328 14684 3368
rect 14596 3282 14609 3328
rect 14655 3282 14684 3328
rect 14596 3204 14684 3282
rect 14884 3328 14972 3368
rect 14884 3282 14913 3328
rect 14959 3282 14972 3328
rect 15935 3380 16008 3393
rect 15935 3368 15949 3380
rect 14884 3204 14972 3282
rect 15044 3288 15132 3301
rect 15044 3242 15057 3288
rect 15103 3242 15132 3288
rect 15044 3229 15132 3242
rect 15252 3288 15387 3301
rect 15252 3242 15312 3288
rect 15358 3242 15387 3288
rect 15252 3229 15387 3242
rect 15507 3288 15595 3301
rect 15507 3242 15536 3288
rect 15582 3242 15595 3288
rect 15507 3229 15595 3242
rect 15667 3278 15755 3368
rect 15667 3232 15680 3278
rect 15726 3232 15755 3278
rect 15667 3204 15755 3232
rect 15875 3334 15949 3368
rect 15995 3334 16008 3380
rect 15875 3204 16008 3334
rect 16088 3380 16160 3393
rect 16088 3334 16101 3380
rect 16147 3334 16160 3380
rect 16088 3301 16160 3334
rect 16088 3229 16220 3301
rect 16340 3288 16444 3301
rect 16340 3242 16369 3288
rect 16415 3242 16444 3288
rect 16340 3229 16444 3242
rect 16564 3288 16668 3301
rect 16564 3242 16593 3288
rect 16639 3242 16668 3288
rect 16564 3229 16668 3242
rect 16788 3288 16876 3301
rect 16788 3242 16817 3288
rect 16863 3242 16876 3288
rect 16788 3229 16876 3242
rect 17475 3311 17563 3368
rect 17475 3265 17488 3311
rect 17534 3265 17563 3311
rect 17475 3204 17563 3265
rect 17683 3308 17771 3368
rect 17683 3262 17712 3308
rect 17758 3262 17771 3308
rect 17683 3204 17771 3262
rect 17844 3328 17932 3368
rect 17844 3282 17857 3328
rect 17903 3282 17932 3328
rect 17844 3204 17932 3282
rect 18132 3328 18220 3368
rect 18132 3282 18161 3328
rect 18207 3282 18220 3328
rect 18132 3204 18220 3282
<< mvpdiff >>
rect 1736 8505 1824 8556
rect 1736 8365 1749 8505
rect 1795 8365 1824 8505
rect 1736 8312 1824 8365
rect 1924 8505 2012 8556
rect 1924 8365 1953 8505
rect 1999 8365 2012 8505
rect 2388 8485 2476 8524
rect 2388 8439 2401 8485
rect 2447 8439 2476 8485
rect 2388 8400 2476 8439
rect 2576 8485 2680 8524
rect 2576 8439 2605 8485
rect 2651 8439 2680 8485
rect 2576 8400 2680 8439
rect 2780 8485 2884 8524
rect 2780 8439 2809 8485
rect 2855 8439 2884 8485
rect 2780 8400 2884 8439
rect 2984 8421 3116 8524
rect 2984 8400 3057 8421
rect 1924 8312 2012 8365
rect 3044 8375 3057 8400
rect 3103 8375 3116 8421
rect 3044 8362 3116 8375
rect 3258 8407 3346 8556
rect 3258 8361 3271 8407
rect 3317 8361 3346 8407
rect 3258 8337 3346 8361
rect 3446 8527 3534 8556
rect 3446 8481 3475 8527
rect 3521 8481 3534 8527
rect 3446 8337 3534 8481
rect 3689 8502 3777 8556
rect 3689 8456 3702 8502
rect 3748 8456 3777 8502
rect 3689 8432 3777 8456
rect 3877 8520 4012 8556
rect 3877 8474 3906 8520
rect 3952 8474 4012 8520
rect 3877 8432 4012 8474
rect 4112 8502 4200 8556
rect 4112 8456 4141 8502
rect 4187 8456 4200 8502
rect 4112 8432 4200 8456
rect 4572 8505 4660 8556
rect 4572 8365 4585 8505
rect 4631 8365 4660 8505
rect 4572 8312 4660 8365
rect 4760 8527 4908 8556
rect 4760 8481 4789 8527
rect 4835 8481 4908 8527
rect 4760 8443 4908 8481
rect 5008 8508 5096 8556
rect 5008 8462 5037 8508
rect 5083 8462 5096 8508
rect 5008 8443 5096 8462
rect 4760 8312 4848 8443
rect 5524 8497 5612 8556
rect 5524 8357 5537 8497
rect 5583 8357 5612 8497
rect 5524 8312 5612 8357
rect 5812 8497 5900 8556
rect 5812 8357 5841 8497
rect 5887 8357 5900 8497
rect 5812 8312 5900 8357
rect 5972 8497 6060 8556
rect 5972 8357 5985 8497
rect 6031 8357 6060 8497
rect 5972 8312 6060 8357
rect 6260 8497 6348 8556
rect 6260 8357 6289 8497
rect 6335 8357 6348 8497
rect 6260 8312 6348 8357
rect 6612 8505 6700 8556
rect 6612 8365 6625 8505
rect 6671 8365 6700 8505
rect 6612 8312 6700 8365
rect 6800 8505 6888 8556
rect 6800 8365 6829 8505
rect 6875 8365 6888 8505
rect 7204 8485 7292 8524
rect 7204 8439 7217 8485
rect 7263 8439 7292 8485
rect 7204 8400 7292 8439
rect 7392 8485 7496 8524
rect 7392 8439 7421 8485
rect 7467 8439 7496 8485
rect 7392 8400 7496 8439
rect 7596 8485 7700 8524
rect 7596 8439 7625 8485
rect 7671 8439 7700 8485
rect 7596 8400 7700 8439
rect 7800 8421 7932 8524
rect 7800 8400 7873 8421
rect 6800 8312 6888 8365
rect 7860 8375 7873 8400
rect 7919 8375 7932 8421
rect 7860 8362 7932 8375
rect 8074 8407 8162 8556
rect 8074 8361 8087 8407
rect 8133 8361 8162 8407
rect 8074 8337 8162 8361
rect 8262 8527 8350 8556
rect 8262 8481 8291 8527
rect 8337 8481 8350 8527
rect 8262 8337 8350 8481
rect 8505 8502 8593 8556
rect 8505 8456 8518 8502
rect 8564 8456 8593 8502
rect 8505 8432 8593 8456
rect 8693 8520 8828 8556
rect 8693 8474 8722 8520
rect 8768 8474 8828 8520
rect 8693 8432 8828 8474
rect 8928 8502 9016 8556
rect 8928 8456 8957 8502
rect 9003 8456 9016 8502
rect 8928 8432 9016 8456
rect 9800 8505 9888 8556
rect 9800 8365 9813 8505
rect 9859 8365 9888 8505
rect 9800 8312 9888 8365
rect 9988 8505 10076 8556
rect 9988 8365 10017 8505
rect 10063 8365 10076 8505
rect 9988 8312 10076 8365
rect 10532 8505 10620 8556
rect 10532 8365 10545 8505
rect 10591 8365 10620 8505
rect 10532 8312 10620 8365
rect 10720 8505 10808 8556
rect 10720 8365 10749 8505
rect 10795 8365 10808 8505
rect 11144 8502 11232 8556
rect 11144 8456 11157 8502
rect 11203 8456 11232 8502
rect 11144 8432 11232 8456
rect 11332 8520 11467 8556
rect 11332 8474 11392 8520
rect 11438 8474 11467 8520
rect 11332 8432 11467 8474
rect 11567 8502 11655 8556
rect 11567 8456 11596 8502
rect 11642 8456 11655 8502
rect 11567 8432 11655 8456
rect 11810 8527 11898 8556
rect 11810 8481 11823 8527
rect 11869 8481 11898 8527
rect 10720 8312 10808 8365
rect 11810 8337 11898 8481
rect 11998 8407 12086 8556
rect 11998 8361 12027 8407
rect 12073 8361 12086 8407
rect 12228 8421 12360 8524
rect 12228 8375 12241 8421
rect 12287 8400 12360 8421
rect 12460 8485 12564 8524
rect 12460 8439 12489 8485
rect 12535 8439 12564 8485
rect 12460 8400 12564 8439
rect 12664 8485 12768 8524
rect 12664 8439 12693 8485
rect 12739 8439 12768 8485
rect 12664 8400 12768 8439
rect 12868 8485 12956 8524
rect 12868 8439 12897 8485
rect 12943 8439 12956 8485
rect 12868 8400 12956 8439
rect 12287 8375 12300 8400
rect 12228 8362 12300 8375
rect 11998 8337 12086 8361
rect 13556 8505 13644 8556
rect 13556 8365 13569 8505
rect 13615 8365 13644 8505
rect 13556 8312 13644 8365
rect 13744 8505 13832 8556
rect 13744 8365 13773 8505
rect 13819 8365 13832 8505
rect 14280 8502 14368 8556
rect 14280 8456 14293 8502
rect 14339 8456 14368 8502
rect 14280 8432 14368 8456
rect 14468 8520 14603 8556
rect 14468 8474 14528 8520
rect 14574 8474 14603 8520
rect 14468 8432 14603 8474
rect 14703 8502 14791 8556
rect 14703 8456 14732 8502
rect 14778 8456 14791 8502
rect 14703 8432 14791 8456
rect 14946 8527 15034 8556
rect 14946 8481 14959 8527
rect 15005 8481 15034 8527
rect 13744 8312 13832 8365
rect 14946 8337 15034 8481
rect 15134 8407 15222 8556
rect 15134 8361 15163 8407
rect 15209 8361 15222 8407
rect 15364 8421 15496 8524
rect 15364 8375 15377 8421
rect 15423 8400 15496 8421
rect 15596 8485 15700 8524
rect 15596 8439 15625 8485
rect 15671 8439 15700 8485
rect 15596 8400 15700 8439
rect 15800 8485 15904 8524
rect 15800 8439 15829 8485
rect 15875 8439 15904 8485
rect 15800 8400 15904 8439
rect 16004 8485 16092 8524
rect 16004 8439 16033 8485
rect 16079 8439 16092 8485
rect 16004 8400 16092 8439
rect 16408 8505 16496 8556
rect 15423 8375 15436 8400
rect 15364 8362 15436 8375
rect 15134 8337 15222 8361
rect 16408 8365 16421 8505
rect 16467 8365 16496 8505
rect 16408 8312 16496 8365
rect 16596 8505 16684 8556
rect 16596 8365 16625 8505
rect 16671 8365 16684 8505
rect 16596 8312 16684 8365
rect 17416 8505 17504 8556
rect 17416 8365 17429 8505
rect 17475 8365 17504 8505
rect 17416 8312 17504 8365
rect 17604 8505 17692 8556
rect 17604 8365 17633 8505
rect 17679 8365 17692 8505
rect 17604 8312 17692 8365
rect 17844 8497 17932 8556
rect 17844 8357 17857 8497
rect 17903 8357 17932 8497
rect 17844 8312 17932 8357
rect 18132 8497 18220 8556
rect 18132 8357 18161 8497
rect 18207 8357 18220 8497
rect 18132 8312 18220 8357
rect 1736 7315 1824 7368
rect 1736 7175 1749 7315
rect 1795 7175 1824 7315
rect 1736 7124 1824 7175
rect 1924 7315 2012 7368
rect 1924 7175 1953 7315
rect 1999 7175 2012 7315
rect 3258 7319 3346 7343
rect 3044 7305 3116 7318
rect 3044 7280 3057 7305
rect 1924 7124 2012 7175
rect 2388 7241 2476 7280
rect 2388 7195 2401 7241
rect 2447 7195 2476 7241
rect 2388 7156 2476 7195
rect 2576 7241 2680 7280
rect 2576 7195 2605 7241
rect 2651 7195 2680 7241
rect 2576 7156 2680 7195
rect 2780 7241 2884 7280
rect 2780 7195 2809 7241
rect 2855 7195 2884 7241
rect 2780 7156 2884 7195
rect 2984 7259 3057 7280
rect 3103 7259 3116 7305
rect 2984 7156 3116 7259
rect 3258 7273 3271 7319
rect 3317 7273 3346 7319
rect 3258 7124 3346 7273
rect 3446 7199 3534 7343
rect 4596 7315 4684 7368
rect 3446 7153 3475 7199
rect 3521 7153 3534 7199
rect 3446 7124 3534 7153
rect 3689 7224 3777 7248
rect 3689 7178 3702 7224
rect 3748 7178 3777 7224
rect 3689 7124 3777 7178
rect 3877 7206 4012 7248
rect 3877 7160 3906 7206
rect 3952 7160 4012 7206
rect 3877 7124 4012 7160
rect 4112 7224 4200 7248
rect 4112 7178 4141 7224
rect 4187 7178 4200 7224
rect 4112 7124 4200 7178
rect 4596 7175 4609 7315
rect 4655 7175 4684 7315
rect 4596 7124 4684 7175
rect 4784 7315 4872 7368
rect 4784 7175 4813 7315
rect 4859 7175 4872 7315
rect 4784 7124 4872 7175
rect 4964 7323 5052 7368
rect 4964 7183 4977 7323
rect 5023 7183 5052 7323
rect 4964 7124 5052 7183
rect 5252 7323 5340 7368
rect 5252 7183 5281 7323
rect 5327 7183 5340 7323
rect 5252 7124 5340 7183
rect 5412 7323 5500 7368
rect 5412 7183 5425 7323
rect 5471 7183 5500 7323
rect 5412 7124 5500 7183
rect 5700 7323 5788 7368
rect 5700 7183 5729 7323
rect 5775 7183 5788 7323
rect 5700 7124 5788 7183
rect 5860 7323 5948 7368
rect 5860 7183 5873 7323
rect 5919 7183 5948 7323
rect 5860 7124 5948 7183
rect 6148 7323 6236 7368
rect 6148 7183 6177 7323
rect 6223 7183 6236 7323
rect 6148 7124 6236 7183
rect 6308 7323 6396 7368
rect 6308 7183 6321 7323
rect 6367 7183 6396 7323
rect 6308 7124 6396 7183
rect 6596 7323 6684 7368
rect 6596 7183 6625 7323
rect 6671 7183 6684 7323
rect 6596 7124 6684 7183
rect 6756 7323 6844 7368
rect 6756 7183 6769 7323
rect 6815 7183 6844 7323
rect 6756 7124 6844 7183
rect 7044 7323 7132 7368
rect 7044 7183 7073 7323
rect 7119 7183 7132 7323
rect 8074 7319 8162 7343
rect 7860 7305 7932 7318
rect 7860 7280 7873 7305
rect 7044 7124 7132 7183
rect 7204 7241 7292 7280
rect 7204 7195 7217 7241
rect 7263 7195 7292 7241
rect 7204 7156 7292 7195
rect 7392 7241 7496 7280
rect 7392 7195 7421 7241
rect 7467 7195 7496 7241
rect 7392 7156 7496 7195
rect 7596 7241 7700 7280
rect 7596 7195 7625 7241
rect 7671 7195 7700 7241
rect 7596 7156 7700 7195
rect 7800 7259 7873 7280
rect 7919 7259 7932 7305
rect 7800 7156 7932 7259
rect 8074 7273 8087 7319
rect 8133 7273 8162 7319
rect 8074 7124 8162 7273
rect 8262 7199 8350 7343
rect 8262 7153 8291 7199
rect 8337 7153 8350 7199
rect 8262 7124 8350 7153
rect 8505 7224 8593 7248
rect 8505 7178 8518 7224
rect 8564 7178 8593 7224
rect 8505 7124 8593 7178
rect 8693 7206 8828 7248
rect 8693 7160 8722 7206
rect 8768 7160 8828 7206
rect 8693 7124 8828 7160
rect 8928 7224 9016 7248
rect 8928 7178 8957 7224
rect 9003 7178 9016 7224
rect 8928 7124 9016 7178
rect 9556 7323 9644 7368
rect 9556 7183 9569 7323
rect 9615 7183 9644 7323
rect 9556 7124 9644 7183
rect 9844 7323 9932 7368
rect 9844 7183 9873 7323
rect 9919 7183 9932 7323
rect 9844 7124 9932 7183
rect 10024 7315 10112 7368
rect 10024 7175 10037 7315
rect 10083 7175 10112 7315
rect 10024 7124 10112 7175
rect 10212 7315 10300 7368
rect 10212 7175 10241 7315
rect 10287 7175 10300 7315
rect 10212 7124 10300 7175
rect 10696 7315 10784 7368
rect 10696 7175 10709 7315
rect 10755 7175 10784 7315
rect 10696 7124 10784 7175
rect 10884 7315 10972 7368
rect 10884 7175 10913 7315
rect 10959 7175 10972 7315
rect 10884 7124 10972 7175
rect 11368 7315 11456 7368
rect 11368 7175 11381 7315
rect 11427 7175 11456 7315
rect 11368 7124 11456 7175
rect 11556 7315 11644 7368
rect 11556 7175 11585 7315
rect 11631 7175 11644 7315
rect 12890 7319 12978 7343
rect 12676 7305 12748 7318
rect 12676 7280 12689 7305
rect 11556 7124 11644 7175
rect 12020 7241 12108 7280
rect 12020 7195 12033 7241
rect 12079 7195 12108 7241
rect 12020 7156 12108 7195
rect 12208 7241 12312 7280
rect 12208 7195 12237 7241
rect 12283 7195 12312 7241
rect 12208 7156 12312 7195
rect 12412 7241 12516 7280
rect 12412 7195 12441 7241
rect 12487 7195 12516 7241
rect 12412 7156 12516 7195
rect 12616 7259 12689 7280
rect 12735 7259 12748 7305
rect 12616 7156 12748 7259
rect 12890 7273 12903 7319
rect 12949 7273 12978 7319
rect 12890 7124 12978 7273
rect 13078 7199 13166 7343
rect 13924 7323 14012 7368
rect 13078 7153 13107 7199
rect 13153 7153 13166 7199
rect 13078 7124 13166 7153
rect 13321 7224 13409 7248
rect 13321 7178 13334 7224
rect 13380 7178 13409 7224
rect 13321 7124 13409 7178
rect 13509 7206 13644 7248
rect 13509 7160 13538 7206
rect 13584 7160 13644 7206
rect 13509 7124 13644 7160
rect 13744 7224 13832 7248
rect 13744 7178 13773 7224
rect 13819 7178 13832 7224
rect 13744 7124 13832 7178
rect 13924 7183 13937 7323
rect 13983 7183 14012 7323
rect 13924 7124 14012 7183
rect 14212 7323 14300 7368
rect 14212 7183 14241 7323
rect 14287 7183 14300 7323
rect 14212 7124 14300 7183
rect 14392 7224 14480 7248
rect 14392 7178 14405 7224
rect 14451 7178 14480 7224
rect 14392 7124 14480 7178
rect 14580 7206 14715 7248
rect 14580 7160 14640 7206
rect 14686 7160 14715 7206
rect 14580 7124 14715 7160
rect 14815 7224 14903 7248
rect 14815 7178 14844 7224
rect 14890 7178 14903 7224
rect 14815 7124 14903 7178
rect 15058 7199 15146 7343
rect 15058 7153 15071 7199
rect 15117 7153 15146 7199
rect 15058 7124 15146 7153
rect 15246 7319 15334 7343
rect 15246 7273 15275 7319
rect 15321 7273 15334 7319
rect 15246 7124 15334 7273
rect 15476 7305 15548 7318
rect 15476 7259 15489 7305
rect 15535 7280 15548 7305
rect 16520 7315 16608 7368
rect 15535 7259 15608 7280
rect 15476 7156 15608 7259
rect 15708 7241 15812 7280
rect 15708 7195 15737 7241
rect 15783 7195 15812 7241
rect 15708 7156 15812 7195
rect 15912 7241 16016 7280
rect 15912 7195 15941 7241
rect 15987 7195 16016 7241
rect 15912 7156 16016 7195
rect 16116 7241 16204 7280
rect 16116 7195 16145 7241
rect 16191 7195 16204 7241
rect 16116 7156 16204 7195
rect 16520 7175 16533 7315
rect 16579 7175 16608 7315
rect 16520 7124 16608 7175
rect 16708 7315 16796 7368
rect 16708 7175 16737 7315
rect 16783 7175 16796 7315
rect 16708 7124 16796 7175
rect 17640 7315 17728 7368
rect 17640 7175 17653 7315
rect 17699 7175 17728 7315
rect 17640 7124 17728 7175
rect 17828 7315 17916 7368
rect 17828 7175 17857 7315
rect 17903 7175 17916 7315
rect 17828 7124 17916 7175
rect 1604 6929 1692 6988
rect 1604 6789 1617 6929
rect 1663 6789 1692 6929
rect 1604 6744 1692 6789
rect 1892 6929 1980 6988
rect 1892 6789 1921 6929
rect 1967 6789 1980 6929
rect 1892 6744 1980 6789
rect 2093 6937 2181 6988
rect 2093 6797 2106 6937
rect 2152 6797 2181 6937
rect 2093 6744 2181 6797
rect 2281 6937 2453 6988
rect 2281 6797 2310 6937
rect 2356 6875 2453 6937
rect 2553 6875 2657 6988
rect 2757 6944 2845 6988
rect 2757 6898 2786 6944
rect 2832 6898 2845 6944
rect 2757 6875 2845 6898
rect 3228 6937 3316 6988
rect 2356 6797 2369 6875
rect 2281 6744 2369 6797
rect 3228 6797 3241 6937
rect 3287 6797 3316 6937
rect 3228 6744 3316 6797
rect 3416 6959 3564 6988
rect 3416 6913 3445 6959
rect 3491 6913 3564 6959
rect 3416 6875 3564 6913
rect 3664 6940 3752 6988
rect 3664 6894 3693 6940
rect 3739 6894 3752 6940
rect 3664 6875 3752 6894
rect 3844 6929 3932 6988
rect 3416 6744 3504 6875
rect 3844 6789 3857 6929
rect 3903 6789 3932 6929
rect 3844 6744 3932 6789
rect 4132 6929 4220 6988
rect 4132 6789 4161 6929
rect 4207 6789 4220 6929
rect 4132 6744 4220 6789
rect 4292 6929 4380 6988
rect 4292 6789 4305 6929
rect 4351 6789 4380 6929
rect 4292 6744 4380 6789
rect 4580 6929 4668 6988
rect 4580 6789 4609 6929
rect 4655 6789 4668 6929
rect 4580 6744 4668 6789
rect 4740 6929 4828 6988
rect 4740 6789 4753 6929
rect 4799 6789 4828 6929
rect 4740 6744 4828 6789
rect 5028 6929 5116 6988
rect 5028 6789 5057 6929
rect 5103 6789 5116 6929
rect 5028 6744 5116 6789
rect 5524 6929 5612 6988
rect 5524 6789 5537 6929
rect 5583 6789 5612 6929
rect 5524 6744 5612 6789
rect 5812 6929 5900 6988
rect 5812 6789 5841 6929
rect 5887 6789 5900 6929
rect 5812 6744 5900 6789
rect 5972 6929 6060 6988
rect 5972 6789 5985 6929
rect 6031 6789 6060 6929
rect 5972 6744 6060 6789
rect 6260 6929 6348 6988
rect 6260 6789 6289 6929
rect 6335 6789 6348 6929
rect 6260 6744 6348 6789
rect 6855 6921 6943 6988
rect 6855 6781 6868 6921
rect 6914 6781 6943 6921
rect 6855 6744 6943 6781
rect 7043 6921 7131 6988
rect 7043 6781 7072 6921
rect 7118 6781 7131 6921
rect 7043 6744 7131 6781
rect 7448 6937 7536 6988
rect 7448 6797 7461 6937
rect 7507 6797 7536 6937
rect 7448 6744 7536 6797
rect 7636 6937 7724 6988
rect 7636 6797 7665 6937
rect 7711 6797 7724 6937
rect 7636 6744 7724 6797
rect 8120 6937 8208 6988
rect 8120 6797 8133 6937
rect 8179 6797 8208 6937
rect 8120 6744 8208 6797
rect 8308 6937 8396 6988
rect 8308 6797 8337 6937
rect 8383 6797 8396 6937
rect 8308 6744 8396 6797
rect 8792 6937 8880 6988
rect 8792 6797 8805 6937
rect 8851 6797 8880 6937
rect 8792 6744 8880 6797
rect 8980 6937 9068 6988
rect 8980 6797 9009 6937
rect 9055 6797 9068 6937
rect 8980 6744 9068 6797
rect 9464 6937 9552 6988
rect 9464 6797 9477 6937
rect 9523 6797 9552 6937
rect 9464 6744 9552 6797
rect 9652 6937 9740 6988
rect 9652 6797 9681 6937
rect 9727 6797 9740 6937
rect 9652 6744 9740 6797
rect 10136 6937 10224 6988
rect 10136 6797 10149 6937
rect 10195 6797 10224 6937
rect 10136 6744 10224 6797
rect 10324 6937 10412 6988
rect 10324 6797 10353 6937
rect 10399 6797 10412 6937
rect 10324 6744 10412 6797
rect 10808 6937 10896 6988
rect 10808 6797 10821 6937
rect 10867 6797 10896 6937
rect 10808 6744 10896 6797
rect 10996 6937 11084 6988
rect 10996 6797 11025 6937
rect 11071 6797 11084 6937
rect 10996 6744 11084 6797
rect 11480 6937 11568 6988
rect 11480 6797 11493 6937
rect 11539 6797 11568 6937
rect 11480 6744 11568 6797
rect 11668 6937 11756 6988
rect 11668 6797 11697 6937
rect 11743 6797 11756 6937
rect 11668 6744 11756 6797
rect 12152 6937 12240 6988
rect 12152 6797 12165 6937
rect 12211 6797 12240 6937
rect 12152 6744 12240 6797
rect 12340 6937 12428 6988
rect 12340 6797 12369 6937
rect 12415 6797 12428 6937
rect 12340 6744 12428 6797
rect 12580 6929 12668 6988
rect 12580 6789 12593 6929
rect 12639 6789 12668 6929
rect 12580 6744 12668 6789
rect 12868 6929 12956 6988
rect 12868 6789 12897 6929
rect 12943 6789 12956 6929
rect 12868 6744 12956 6789
rect 13608 6937 13696 6988
rect 13608 6797 13621 6937
rect 13667 6797 13696 6937
rect 13608 6744 13696 6797
rect 13796 6937 13884 6988
rect 13796 6797 13825 6937
rect 13871 6797 13884 6937
rect 13796 6744 13884 6797
rect 14280 6937 14368 6988
rect 14280 6797 14293 6937
rect 14339 6797 14368 6937
rect 14280 6744 14368 6797
rect 14468 6937 14556 6988
rect 14468 6797 14497 6937
rect 14543 6797 14556 6937
rect 14468 6744 14556 6797
rect 14952 6937 15040 6988
rect 14952 6797 14965 6937
rect 15011 6797 15040 6937
rect 14952 6744 15040 6797
rect 15140 6937 15228 6988
rect 15140 6797 15169 6937
rect 15215 6797 15228 6937
rect 15140 6744 15228 6797
rect 15624 6937 15712 6988
rect 15624 6797 15637 6937
rect 15683 6797 15712 6937
rect 15624 6744 15712 6797
rect 15812 6937 15900 6988
rect 15812 6797 15841 6937
rect 15887 6797 15900 6937
rect 15812 6744 15900 6797
rect 16296 6937 16384 6988
rect 16296 6797 16309 6937
rect 16355 6797 16384 6937
rect 16296 6744 16384 6797
rect 16484 6937 16572 6988
rect 16484 6797 16513 6937
rect 16559 6797 16572 6937
rect 16484 6744 16572 6797
rect 16968 6937 17056 6988
rect 16968 6797 16981 6937
rect 17027 6797 17056 6937
rect 16968 6744 17056 6797
rect 17156 6937 17244 6988
rect 17156 6797 17185 6937
rect 17231 6797 17244 6937
rect 17156 6744 17244 6797
rect 17640 6937 17728 6988
rect 17640 6797 17653 6937
rect 17699 6797 17728 6937
rect 17640 6744 17728 6797
rect 17828 6937 17916 6988
rect 17828 6797 17857 6937
rect 17903 6797 17916 6937
rect 17828 6744 17916 6797
rect 2176 5747 2276 5800
rect 2176 5677 2201 5747
rect 1716 5616 1804 5677
rect 1716 5570 1729 5616
rect 1775 5570 1804 5616
rect 1716 5557 1804 5570
rect 1904 5664 2008 5677
rect 1904 5618 1933 5664
rect 1979 5618 2008 5664
rect 1904 5557 2008 5618
rect 2108 5607 2201 5677
rect 2247 5607 2276 5747
rect 2108 5557 2276 5607
rect 2376 5747 2464 5800
rect 2376 5607 2405 5747
rect 2451 5607 2464 5747
rect 2376 5557 2464 5607
rect 2856 5747 2944 5800
rect 2856 5607 2869 5747
rect 2915 5607 2944 5747
rect 2856 5556 2944 5607
rect 3044 5747 3132 5800
rect 3044 5607 3073 5747
rect 3119 5607 3132 5747
rect 3044 5556 3132 5607
rect 3284 5755 3372 5800
rect 3284 5615 3297 5755
rect 3343 5615 3372 5755
rect 3284 5556 3372 5615
rect 3572 5755 3660 5800
rect 3572 5615 3601 5755
rect 3647 5615 3660 5755
rect 3572 5556 3660 5615
rect 3732 5755 3820 5800
rect 3732 5615 3745 5755
rect 3791 5615 3820 5755
rect 3732 5556 3820 5615
rect 4020 5755 4108 5800
rect 4020 5615 4049 5755
rect 4095 5615 4108 5755
rect 4020 5556 4108 5615
rect 4180 5755 4268 5800
rect 4180 5615 4193 5755
rect 4239 5615 4268 5755
rect 4180 5556 4268 5615
rect 4468 5755 4556 5800
rect 4468 5615 4497 5755
rect 4543 5615 4556 5755
rect 4468 5556 4556 5615
rect 4628 5755 4716 5800
rect 4628 5615 4641 5755
rect 4687 5615 4716 5755
rect 4628 5556 4716 5615
rect 4916 5755 5004 5800
rect 4916 5615 4945 5755
rect 4991 5615 5004 5755
rect 4916 5556 5004 5615
rect 5413 5763 5501 5800
rect 5413 5623 5426 5763
rect 5472 5623 5501 5763
rect 5413 5556 5501 5623
rect 5601 5763 5689 5800
rect 5601 5623 5630 5763
rect 5676 5623 5689 5763
rect 5601 5556 5689 5623
rect 6164 5747 6252 5800
rect 6164 5607 6177 5747
rect 6223 5607 6252 5747
rect 6164 5556 6252 5607
rect 6352 5747 6440 5800
rect 6352 5607 6381 5747
rect 6427 5607 6440 5747
rect 6352 5556 6440 5607
rect 6836 5747 6924 5800
rect 6836 5607 6849 5747
rect 6895 5607 6924 5747
rect 6836 5556 6924 5607
rect 7024 5747 7112 5800
rect 7024 5607 7053 5747
rect 7099 5607 7112 5747
rect 7024 5556 7112 5607
rect 7448 5747 7536 5800
rect 7448 5607 7461 5747
rect 7507 5607 7536 5747
rect 7448 5556 7536 5607
rect 7636 5747 7724 5800
rect 7636 5607 7665 5747
rect 7711 5607 7724 5747
rect 7636 5556 7724 5607
rect 8101 5763 8189 5800
rect 8101 5623 8114 5763
rect 8160 5623 8189 5763
rect 8101 5556 8189 5623
rect 8289 5763 8377 5800
rect 8289 5623 8318 5763
rect 8364 5623 8377 5763
rect 8289 5556 8377 5623
rect 8792 5747 8880 5800
rect 8792 5607 8805 5747
rect 8851 5607 8880 5747
rect 8792 5556 8880 5607
rect 8980 5747 9068 5800
rect 8980 5607 9009 5747
rect 9055 5607 9068 5747
rect 8980 5556 9068 5607
rect 9556 5755 9644 5800
rect 9556 5615 9569 5755
rect 9615 5615 9644 5755
rect 9556 5556 9644 5615
rect 9844 5755 9932 5800
rect 9844 5615 9873 5755
rect 9919 5615 9932 5755
rect 9844 5556 9932 5615
rect 10248 5747 10336 5800
rect 10248 5607 10261 5747
rect 10307 5607 10336 5747
rect 10248 5556 10336 5607
rect 10436 5747 10524 5800
rect 10436 5607 10465 5747
rect 10511 5607 10524 5747
rect 10436 5556 10524 5607
rect 10920 5747 11008 5800
rect 10920 5607 10933 5747
rect 10979 5607 11008 5747
rect 10920 5556 11008 5607
rect 11108 5747 11196 5800
rect 11108 5607 11137 5747
rect 11183 5607 11196 5747
rect 11108 5556 11196 5607
rect 11592 5747 11680 5800
rect 11592 5607 11605 5747
rect 11651 5607 11680 5747
rect 11592 5556 11680 5607
rect 11780 5747 11868 5800
rect 11780 5607 11809 5747
rect 11855 5607 11868 5747
rect 11780 5556 11868 5607
rect 12264 5747 12352 5800
rect 12264 5607 12277 5747
rect 12323 5607 12352 5747
rect 12264 5556 12352 5607
rect 12452 5747 12540 5800
rect 12452 5607 12481 5747
rect 12527 5607 12540 5747
rect 12452 5556 12540 5607
rect 12936 5747 13024 5800
rect 12936 5607 12949 5747
rect 12995 5607 13024 5747
rect 12936 5556 13024 5607
rect 13124 5747 13212 5800
rect 13124 5607 13153 5747
rect 13199 5607 13212 5747
rect 13124 5556 13212 5607
rect 13608 5747 13696 5800
rect 13608 5607 13621 5747
rect 13667 5607 13696 5747
rect 13608 5556 13696 5607
rect 13796 5747 13884 5800
rect 13796 5607 13825 5747
rect 13871 5607 13884 5747
rect 13796 5556 13884 5607
rect 14280 5747 14368 5800
rect 14280 5607 14293 5747
rect 14339 5607 14368 5747
rect 14280 5556 14368 5607
rect 14468 5747 14556 5800
rect 14468 5607 14497 5747
rect 14543 5607 14556 5747
rect 14468 5556 14556 5607
rect 14952 5747 15040 5800
rect 14952 5607 14965 5747
rect 15011 5607 15040 5747
rect 14952 5556 15040 5607
rect 15140 5747 15228 5800
rect 15140 5607 15169 5747
rect 15215 5607 15228 5747
rect 15140 5556 15228 5607
rect 15624 5747 15712 5800
rect 15624 5607 15637 5747
rect 15683 5607 15712 5747
rect 15624 5556 15712 5607
rect 15812 5747 15900 5800
rect 15812 5607 15841 5747
rect 15887 5607 15900 5747
rect 15812 5556 15900 5607
rect 16277 5763 16365 5800
rect 16277 5623 16290 5763
rect 16336 5623 16365 5763
rect 16277 5556 16365 5623
rect 16465 5763 16553 5800
rect 16465 5623 16494 5763
rect 16540 5623 16553 5763
rect 16465 5556 16553 5623
rect 16724 5755 16812 5800
rect 16724 5615 16737 5755
rect 16783 5615 16812 5755
rect 16724 5556 16812 5615
rect 17012 5755 17100 5800
rect 17012 5615 17041 5755
rect 17087 5615 17100 5755
rect 17012 5556 17100 5615
rect 17719 5763 17807 5800
rect 17719 5623 17732 5763
rect 17778 5623 17807 5763
rect 17719 5556 17807 5623
rect 17907 5763 17995 5800
rect 17907 5623 17936 5763
rect 17982 5623 17995 5763
rect 17907 5556 17995 5623
rect 1604 5361 1692 5420
rect 1604 5221 1617 5361
rect 1663 5221 1692 5361
rect 1604 5176 1692 5221
rect 1892 5361 1980 5420
rect 1892 5221 1921 5361
rect 1967 5221 1980 5361
rect 1892 5176 1980 5221
rect 2052 5361 2140 5420
rect 2052 5221 2065 5361
rect 2111 5221 2140 5361
rect 2052 5176 2140 5221
rect 2340 5361 2428 5420
rect 2340 5221 2369 5361
rect 2415 5221 2428 5361
rect 2340 5176 2428 5221
rect 2500 5361 2588 5420
rect 2500 5221 2513 5361
rect 2559 5221 2588 5361
rect 2500 5176 2588 5221
rect 2788 5361 2876 5420
rect 2788 5221 2817 5361
rect 2863 5221 2876 5361
rect 2788 5176 2876 5221
rect 2948 5361 3036 5420
rect 2948 5221 2961 5361
rect 3007 5221 3036 5361
rect 2948 5176 3036 5221
rect 3236 5361 3324 5420
rect 3236 5221 3265 5361
rect 3311 5221 3324 5361
rect 3236 5176 3324 5221
rect 3396 5361 3484 5420
rect 3396 5221 3409 5361
rect 3455 5221 3484 5361
rect 3396 5176 3484 5221
rect 3684 5361 3772 5420
rect 3684 5221 3713 5361
rect 3759 5221 3772 5361
rect 3684 5176 3772 5221
rect 4069 5353 4157 5420
rect 4069 5213 4082 5353
rect 4128 5213 4157 5353
rect 4069 5176 4157 5213
rect 4257 5353 4345 5420
rect 4257 5213 4286 5353
rect 4332 5213 4345 5353
rect 4257 5176 4345 5213
rect 4741 5353 4829 5420
rect 4741 5213 4754 5353
rect 4800 5213 4829 5353
rect 4741 5176 4829 5213
rect 4929 5353 5017 5420
rect 4929 5213 4958 5353
rect 5004 5213 5017 5353
rect 4929 5176 5017 5213
rect 5524 5361 5612 5420
rect 5524 5221 5537 5361
rect 5583 5221 5612 5361
rect 5524 5176 5612 5221
rect 5812 5361 5900 5420
rect 5812 5221 5841 5361
rect 5887 5221 5900 5361
rect 5812 5176 5900 5221
rect 6197 5353 6285 5420
rect 6197 5213 6210 5353
rect 6256 5213 6285 5353
rect 6197 5176 6285 5213
rect 6385 5353 6473 5420
rect 6385 5213 6414 5353
rect 6460 5213 6473 5353
rect 6385 5176 6473 5213
rect 6967 5353 7055 5420
rect 6967 5213 6980 5353
rect 7026 5213 7055 5353
rect 6967 5176 7055 5213
rect 7155 5353 7243 5420
rect 7155 5213 7184 5353
rect 7230 5213 7243 5353
rect 7155 5176 7243 5213
rect 7620 5369 7708 5420
rect 7620 5229 7633 5369
rect 7679 5229 7708 5369
rect 7620 5176 7708 5229
rect 7808 5369 7896 5420
rect 7808 5229 7837 5369
rect 7883 5229 7896 5369
rect 7808 5176 7896 5229
rect 8213 5353 8301 5420
rect 8213 5213 8226 5353
rect 8272 5213 8301 5353
rect 8213 5176 8301 5213
rect 8401 5353 8489 5420
rect 8401 5213 8430 5353
rect 8476 5213 8489 5353
rect 8401 5176 8489 5213
rect 8904 5369 8992 5420
rect 8904 5229 8917 5369
rect 8963 5229 8992 5369
rect 8904 5176 8992 5229
rect 9092 5369 9180 5420
rect 9092 5229 9121 5369
rect 9167 5229 9180 5369
rect 9092 5176 9180 5229
rect 9576 5369 9664 5420
rect 9576 5229 9589 5369
rect 9635 5229 9664 5369
rect 9576 5176 9664 5229
rect 9764 5369 9852 5420
rect 9764 5229 9793 5369
rect 9839 5229 9852 5369
rect 9764 5176 9852 5229
rect 10248 5369 10336 5420
rect 10248 5229 10261 5369
rect 10307 5229 10336 5369
rect 10248 5176 10336 5229
rect 10436 5369 10524 5420
rect 10436 5229 10465 5369
rect 10511 5229 10524 5369
rect 10436 5176 10524 5229
rect 10920 5369 11008 5420
rect 10920 5229 10933 5369
rect 10979 5229 11008 5369
rect 10920 5176 11008 5229
rect 11108 5369 11196 5420
rect 11108 5229 11137 5369
rect 11183 5229 11196 5369
rect 11108 5176 11196 5229
rect 11592 5369 11680 5420
rect 11592 5229 11605 5369
rect 11651 5229 11680 5369
rect 11592 5176 11680 5229
rect 11780 5369 11868 5420
rect 11780 5229 11809 5369
rect 11855 5229 11868 5369
rect 11780 5176 11868 5229
rect 12264 5369 12352 5420
rect 12264 5229 12277 5369
rect 12323 5229 12352 5369
rect 12264 5176 12352 5229
rect 12452 5369 12540 5420
rect 12452 5229 12481 5369
rect 12527 5229 12540 5369
rect 12452 5176 12540 5229
rect 12692 5361 12780 5420
rect 12692 5221 12705 5361
rect 12751 5221 12780 5361
rect 12692 5176 12780 5221
rect 12980 5361 13068 5420
rect 12980 5221 13009 5361
rect 13055 5221 13068 5361
rect 12980 5176 13068 5221
rect 13608 5369 13696 5420
rect 13608 5229 13621 5369
rect 13667 5229 13696 5369
rect 13608 5176 13696 5229
rect 13796 5369 13884 5420
rect 13796 5229 13825 5369
rect 13871 5229 13884 5369
rect 13796 5176 13884 5229
rect 14280 5369 14368 5420
rect 14280 5229 14293 5369
rect 14339 5229 14368 5369
rect 14280 5176 14368 5229
rect 14468 5369 14556 5420
rect 14468 5229 14497 5369
rect 14543 5229 14556 5369
rect 14468 5176 14556 5229
rect 15012 5369 15100 5420
rect 15012 5229 15025 5369
rect 15071 5229 15100 5369
rect 15012 5176 15100 5229
rect 15200 5369 15288 5420
rect 15200 5229 15229 5369
rect 15275 5229 15288 5369
rect 15200 5176 15288 5229
rect 15703 5353 15791 5420
rect 15703 5213 15716 5353
rect 15762 5213 15791 5353
rect 15703 5176 15791 5213
rect 15891 5353 15979 5420
rect 15891 5213 15920 5353
rect 15966 5213 15979 5353
rect 16408 5366 16496 5420
rect 16408 5320 16421 5366
rect 16467 5320 16496 5366
rect 16408 5296 16496 5320
rect 16596 5384 16731 5420
rect 16596 5338 16656 5384
rect 16702 5338 16731 5384
rect 16596 5296 16731 5338
rect 16831 5366 16919 5420
rect 16831 5320 16860 5366
rect 16906 5320 16919 5366
rect 16831 5296 16919 5320
rect 17074 5391 17162 5420
rect 17074 5345 17087 5391
rect 17133 5345 17162 5391
rect 15891 5176 15979 5213
rect 17074 5201 17162 5345
rect 17262 5271 17350 5420
rect 17262 5225 17291 5271
rect 17337 5225 17350 5271
rect 17492 5285 17624 5388
rect 17492 5239 17505 5285
rect 17551 5264 17624 5285
rect 17724 5349 17828 5388
rect 17724 5303 17753 5349
rect 17799 5303 17828 5349
rect 17724 5264 17828 5303
rect 17928 5349 18032 5388
rect 17928 5303 17957 5349
rect 18003 5303 18032 5349
rect 17928 5264 18032 5303
rect 18132 5349 18220 5388
rect 18132 5303 18161 5349
rect 18207 5303 18220 5349
rect 18132 5264 18220 5303
rect 17551 5239 17564 5264
rect 17492 5226 17564 5239
rect 17262 5201 17350 5225
rect 1604 4187 1692 4232
rect 1604 4047 1617 4187
rect 1663 4047 1692 4187
rect 1604 3988 1692 4047
rect 1892 4187 1980 4232
rect 1892 4047 1921 4187
rect 1967 4047 1980 4187
rect 1892 3988 1980 4047
rect 2052 4187 2140 4232
rect 2052 4047 2065 4187
rect 2111 4047 2140 4187
rect 2052 3988 2140 4047
rect 2340 4187 2428 4232
rect 2340 4047 2369 4187
rect 2415 4047 2428 4187
rect 3482 4183 3570 4207
rect 3268 4169 3340 4182
rect 3268 4144 3281 4169
rect 2340 3988 2428 4047
rect 2612 4105 2700 4144
rect 2612 4059 2625 4105
rect 2671 4059 2700 4105
rect 2612 4020 2700 4059
rect 2800 4105 2904 4144
rect 2800 4059 2829 4105
rect 2875 4059 2904 4105
rect 2800 4020 2904 4059
rect 3004 4105 3108 4144
rect 3004 4059 3033 4105
rect 3079 4059 3108 4105
rect 3004 4020 3108 4059
rect 3208 4123 3281 4144
rect 3327 4123 3340 4169
rect 3208 4020 3340 4123
rect 3482 4137 3495 4183
rect 3541 4137 3570 4183
rect 3482 3988 3570 4137
rect 3670 4063 3758 4207
rect 4516 4187 4604 4232
rect 3670 4017 3699 4063
rect 3745 4017 3758 4063
rect 3670 3988 3758 4017
rect 3913 4088 4001 4112
rect 3913 4042 3926 4088
rect 3972 4042 4001 4088
rect 3913 3988 4001 4042
rect 4101 4070 4236 4112
rect 4101 4024 4130 4070
rect 4176 4024 4236 4070
rect 4101 3988 4236 4024
rect 4336 4088 4424 4112
rect 4336 4042 4365 4088
rect 4411 4042 4424 4088
rect 4336 3988 4424 4042
rect 4516 4047 4529 4187
rect 4575 4047 4604 4187
rect 4516 3988 4604 4047
rect 4804 4187 4892 4232
rect 4804 4047 4833 4187
rect 4879 4047 4892 4187
rect 4804 3988 4892 4047
rect 5077 4195 5165 4232
rect 5077 4055 5090 4195
rect 5136 4055 5165 4195
rect 5077 3988 5165 4055
rect 5265 4195 5353 4232
rect 5265 4055 5294 4195
rect 5340 4055 5353 4195
rect 5265 3988 5353 4055
rect 5749 4195 5837 4232
rect 5749 4055 5762 4195
rect 5808 4055 5837 4195
rect 5749 3988 5837 4055
rect 5937 4195 6025 4232
rect 5937 4055 5966 4195
rect 6012 4055 6025 4195
rect 5937 3988 6025 4055
rect 6421 4195 6509 4232
rect 6421 4055 6434 4195
rect 6480 4055 6509 4195
rect 6421 3988 6509 4055
rect 6609 4195 6697 4232
rect 6609 4055 6638 4195
rect 6684 4055 6697 4195
rect 6609 3988 6697 4055
rect 7112 4088 7200 4112
rect 7112 4042 7125 4088
rect 7171 4042 7200 4088
rect 7112 3988 7200 4042
rect 7300 4070 7435 4112
rect 7300 4024 7360 4070
rect 7406 4024 7435 4070
rect 7300 3988 7435 4024
rect 7535 4088 7623 4112
rect 7535 4042 7564 4088
rect 7610 4042 7623 4088
rect 7535 3988 7623 4042
rect 7778 4063 7866 4207
rect 7778 4017 7791 4063
rect 7837 4017 7866 4063
rect 7778 3988 7866 4017
rect 7966 4183 8054 4207
rect 7966 4137 7995 4183
rect 8041 4137 8054 4183
rect 7966 3988 8054 4137
rect 8196 4169 8268 4182
rect 8196 4123 8209 4169
rect 8255 4144 8268 4169
rect 8255 4123 8328 4144
rect 8196 4020 8328 4123
rect 8428 4105 8532 4144
rect 8428 4059 8457 4105
rect 8503 4059 8532 4105
rect 8428 4020 8532 4059
rect 8632 4105 8736 4144
rect 8632 4059 8661 4105
rect 8707 4059 8736 4105
rect 8632 4020 8736 4059
rect 8836 4105 8924 4144
rect 8836 4059 8865 4105
rect 8911 4059 8924 4105
rect 8836 4020 8924 4059
rect 9556 4187 9644 4232
rect 9556 4047 9569 4187
rect 9615 4047 9644 4187
rect 9556 3988 9644 4047
rect 9844 4187 9932 4232
rect 9844 4047 9873 4187
rect 9919 4047 9932 4187
rect 9844 3988 9932 4047
rect 10005 4195 10093 4232
rect 10005 4055 10018 4195
rect 10064 4055 10093 4195
rect 10005 3988 10093 4055
rect 10193 4195 10281 4232
rect 10193 4055 10222 4195
rect 10268 4055 10281 4195
rect 10193 3988 10281 4055
rect 10756 4179 10844 4232
rect 10756 4039 10769 4179
rect 10815 4039 10844 4179
rect 10756 3988 10844 4039
rect 10944 4179 11032 4232
rect 10944 4039 10973 4179
rect 11019 4039 11032 4179
rect 10944 3988 11032 4039
rect 11428 4179 11516 4232
rect 11428 4039 11441 4179
rect 11487 4039 11516 4179
rect 11428 3988 11516 4039
rect 11616 4179 11704 4232
rect 11616 4039 11645 4179
rect 11691 4039 11704 4179
rect 11616 3988 11704 4039
rect 12040 4088 12128 4112
rect 12040 4042 12053 4088
rect 12099 4042 12128 4088
rect 12040 3988 12128 4042
rect 12228 4070 12363 4112
rect 12228 4024 12288 4070
rect 12334 4024 12363 4070
rect 12228 3988 12363 4024
rect 12463 4088 12551 4112
rect 12463 4042 12492 4088
rect 12538 4042 12551 4088
rect 12463 3988 12551 4042
rect 12706 4063 12794 4207
rect 12706 4017 12719 4063
rect 12765 4017 12794 4063
rect 12706 3988 12794 4017
rect 12894 4183 12982 4207
rect 12894 4137 12923 4183
rect 12969 4137 12982 4183
rect 12894 3988 12982 4137
rect 13124 4169 13196 4182
rect 13124 4123 13137 4169
rect 13183 4144 13196 4169
rect 14149 4195 14237 4232
rect 13183 4123 13256 4144
rect 13124 4020 13256 4123
rect 13356 4105 13460 4144
rect 13356 4059 13385 4105
rect 13431 4059 13460 4105
rect 13356 4020 13460 4059
rect 13560 4105 13664 4144
rect 13560 4059 13589 4105
rect 13635 4059 13664 4105
rect 13560 4020 13664 4059
rect 13764 4105 13852 4144
rect 13764 4059 13793 4105
rect 13839 4059 13852 4105
rect 13764 4020 13852 4059
rect 14149 4055 14162 4195
rect 14208 4055 14237 4195
rect 14149 3988 14237 4055
rect 14337 4195 14425 4232
rect 14337 4055 14366 4195
rect 14412 4055 14425 4195
rect 14337 3988 14425 4055
rect 14840 4179 14928 4232
rect 14840 4039 14853 4179
rect 14899 4039 14928 4179
rect 14840 3988 14928 4039
rect 15028 4179 15116 4232
rect 15028 4039 15057 4179
rect 15103 4039 15116 4179
rect 15028 3988 15116 4039
rect 15512 4179 15600 4232
rect 15512 4039 15525 4179
rect 15571 4039 15600 4179
rect 15512 3988 15600 4039
rect 15700 4179 15788 4232
rect 15700 4039 15729 4179
rect 15775 4039 15788 4179
rect 15700 3988 15788 4039
rect 16184 4179 16272 4232
rect 16184 4039 16197 4179
rect 16243 4039 16272 4179
rect 16184 3988 16272 4039
rect 16372 4179 16460 4232
rect 16372 4039 16401 4179
rect 16447 4039 16460 4179
rect 16372 3988 16460 4039
rect 16612 4187 16700 4232
rect 16612 4047 16625 4187
rect 16671 4047 16700 4187
rect 16612 3988 16700 4047
rect 16900 4187 16988 4232
rect 16900 4047 16929 4187
rect 16975 4047 16988 4187
rect 16900 3988 16988 4047
rect 17640 4179 17728 4232
rect 17640 4039 17653 4179
rect 17699 4039 17728 4179
rect 17640 3988 17728 4039
rect 17828 4179 17916 4232
rect 17828 4039 17857 4179
rect 17903 4039 17916 4179
rect 17828 3988 17916 4039
rect 1941 3785 2029 3852
rect 1941 3645 1954 3785
rect 2000 3645 2029 3785
rect 1941 3608 2029 3645
rect 2129 3785 2217 3852
rect 2129 3645 2158 3785
rect 2204 3645 2217 3785
rect 2632 3798 2720 3852
rect 2632 3752 2645 3798
rect 2691 3752 2720 3798
rect 2632 3728 2720 3752
rect 2820 3816 2955 3852
rect 2820 3770 2880 3816
rect 2926 3770 2955 3816
rect 2820 3728 2955 3770
rect 3055 3798 3143 3852
rect 3055 3752 3084 3798
rect 3130 3752 3143 3798
rect 3055 3728 3143 3752
rect 3298 3823 3386 3852
rect 3298 3777 3311 3823
rect 3357 3777 3386 3823
rect 2129 3608 2217 3645
rect 3298 3633 3386 3777
rect 3486 3703 3574 3852
rect 3486 3657 3515 3703
rect 3561 3657 3574 3703
rect 3716 3717 3848 3820
rect 3716 3671 3729 3717
rect 3775 3696 3848 3717
rect 3948 3781 4052 3820
rect 3948 3735 3977 3781
rect 4023 3735 4052 3781
rect 3948 3696 4052 3735
rect 4152 3781 4256 3820
rect 4152 3735 4181 3781
rect 4227 3735 4256 3781
rect 4152 3696 4256 3735
rect 4356 3781 4444 3820
rect 4356 3735 4385 3781
rect 4431 3735 4444 3781
rect 4356 3696 4444 3735
rect 4741 3785 4829 3852
rect 3775 3671 3788 3696
rect 3716 3658 3788 3671
rect 3486 3633 3574 3657
rect 4741 3645 4754 3785
rect 4800 3645 4829 3785
rect 4741 3608 4829 3645
rect 4929 3785 5017 3852
rect 4929 3645 4958 3785
rect 5004 3645 5017 3785
rect 4929 3608 5017 3645
rect 5861 3785 5949 3852
rect 5861 3645 5874 3785
rect 5920 3645 5949 3785
rect 5861 3608 5949 3645
rect 6049 3785 6137 3852
rect 6049 3645 6078 3785
rect 6124 3645 6137 3785
rect 6049 3608 6137 3645
rect 6533 3785 6621 3852
rect 6533 3645 6546 3785
rect 6592 3645 6621 3785
rect 6533 3608 6621 3645
rect 6721 3785 6809 3852
rect 6721 3645 6750 3785
rect 6796 3645 6809 3785
rect 7224 3798 7312 3852
rect 7224 3752 7237 3798
rect 7283 3752 7312 3798
rect 7224 3728 7312 3752
rect 7412 3816 7547 3852
rect 7412 3770 7472 3816
rect 7518 3770 7547 3816
rect 7412 3728 7547 3770
rect 7647 3798 7735 3852
rect 7647 3752 7676 3798
rect 7722 3752 7735 3798
rect 7647 3728 7735 3752
rect 7890 3823 7978 3852
rect 7890 3777 7903 3823
rect 7949 3777 7978 3823
rect 6721 3608 6809 3645
rect 7890 3633 7978 3777
rect 8078 3703 8166 3852
rect 8078 3657 8107 3703
rect 8153 3657 8166 3703
rect 8308 3717 8440 3820
rect 8308 3671 8321 3717
rect 8367 3696 8440 3717
rect 8540 3781 8644 3820
rect 8540 3735 8569 3781
rect 8615 3735 8644 3781
rect 8540 3696 8644 3735
rect 8744 3781 8848 3820
rect 8744 3735 8773 3781
rect 8819 3735 8848 3781
rect 8744 3696 8848 3735
rect 8948 3781 9036 3820
rect 8948 3735 8977 3781
rect 9023 3735 9036 3781
rect 8948 3696 9036 3735
rect 8367 3671 8380 3696
rect 8308 3658 8380 3671
rect 8078 3633 8166 3657
rect 9781 3785 9869 3852
rect 9781 3645 9794 3785
rect 9840 3645 9869 3785
rect 9781 3608 9869 3645
rect 9969 3785 10057 3852
rect 9969 3645 9998 3785
rect 10044 3645 10057 3785
rect 9969 3608 10057 3645
rect 10453 3785 10541 3852
rect 10453 3645 10466 3785
rect 10512 3645 10541 3785
rect 10453 3608 10541 3645
rect 10641 3785 10729 3852
rect 10641 3645 10670 3785
rect 10716 3645 10729 3785
rect 11144 3798 11232 3852
rect 11144 3752 11157 3798
rect 11203 3752 11232 3798
rect 11144 3728 11232 3752
rect 11332 3816 11467 3852
rect 11332 3770 11392 3816
rect 11438 3770 11467 3816
rect 11332 3728 11467 3770
rect 11567 3798 11655 3852
rect 11567 3752 11596 3798
rect 11642 3752 11655 3798
rect 11567 3728 11655 3752
rect 11810 3823 11898 3852
rect 11810 3777 11823 3823
rect 11869 3777 11898 3823
rect 10641 3608 10729 3645
rect 11810 3633 11898 3777
rect 11998 3703 12086 3852
rect 11998 3657 12027 3703
rect 12073 3657 12086 3703
rect 12228 3717 12360 3820
rect 12228 3671 12241 3717
rect 12287 3696 12360 3717
rect 12460 3781 12564 3820
rect 12460 3735 12489 3781
rect 12535 3735 12564 3781
rect 12460 3696 12564 3735
rect 12664 3781 12768 3820
rect 12664 3735 12693 3781
rect 12739 3735 12768 3781
rect 12664 3696 12768 3735
rect 12868 3781 12956 3820
rect 12868 3735 12897 3781
rect 12943 3735 12956 3781
rect 12868 3696 12956 3735
rect 12287 3671 12300 3696
rect 12228 3658 12300 3671
rect 11998 3633 12086 3657
rect 13556 3801 13644 3852
rect 13556 3661 13569 3801
rect 13615 3661 13644 3801
rect 13556 3608 13644 3661
rect 13744 3801 13832 3852
rect 13744 3661 13773 3801
rect 13819 3661 13832 3801
rect 13744 3608 13832 3661
rect 14149 3785 14237 3852
rect 14149 3645 14162 3785
rect 14208 3645 14237 3785
rect 14149 3608 14237 3645
rect 14337 3785 14425 3852
rect 14337 3645 14366 3785
rect 14412 3645 14425 3785
rect 14337 3608 14425 3645
rect 14596 3793 14684 3852
rect 14596 3653 14609 3793
rect 14655 3653 14684 3793
rect 14596 3608 14684 3653
rect 14884 3793 14972 3852
rect 14884 3653 14913 3793
rect 14959 3653 14972 3793
rect 15064 3798 15152 3852
rect 15064 3752 15077 3798
rect 15123 3752 15152 3798
rect 15064 3728 15152 3752
rect 15252 3816 15387 3852
rect 15252 3770 15312 3816
rect 15358 3770 15387 3816
rect 15252 3728 15387 3770
rect 15487 3798 15575 3852
rect 15487 3752 15516 3798
rect 15562 3752 15575 3798
rect 15487 3728 15575 3752
rect 15730 3823 15818 3852
rect 15730 3777 15743 3823
rect 15789 3777 15818 3823
rect 14884 3608 14972 3653
rect 15730 3633 15818 3777
rect 15918 3703 16006 3852
rect 15918 3657 15947 3703
rect 15993 3657 16006 3703
rect 16148 3717 16280 3820
rect 16148 3671 16161 3717
rect 16207 3696 16280 3717
rect 16380 3781 16484 3820
rect 16380 3735 16409 3781
rect 16455 3735 16484 3781
rect 16380 3696 16484 3735
rect 16584 3781 16688 3820
rect 16584 3735 16613 3781
rect 16659 3735 16688 3781
rect 16584 3696 16688 3735
rect 16788 3781 16876 3820
rect 16788 3735 16817 3781
rect 16863 3735 16876 3781
rect 16788 3696 16876 3735
rect 16207 3671 16220 3696
rect 16148 3658 16220 3671
rect 15918 3633 16006 3657
rect 17495 3785 17583 3852
rect 17495 3645 17508 3785
rect 17554 3645 17583 3785
rect 17495 3608 17583 3645
rect 17683 3785 17771 3852
rect 17683 3645 17712 3785
rect 17758 3645 17771 3785
rect 17683 3608 17771 3645
rect 17844 3793 17932 3852
rect 17844 3653 17857 3793
rect 17903 3653 17932 3793
rect 17844 3608 17932 3653
rect 18132 3793 18220 3852
rect 18132 3653 18161 3793
rect 18207 3653 18220 3793
rect 18132 3608 18220 3653
<< mvndiffc >>
rect 1729 7986 1775 8032
rect 1953 7986 1999 8032
rect 3117 8038 3163 8084
rect 2401 7946 2447 7992
rect 2625 7946 2671 7992
rect 2849 7946 2895 7992
rect 3269 8038 3315 8084
rect 3538 7936 3584 7982
rect 3682 7946 3728 7992
rect 3906 7946 3952 7992
rect 4161 7946 4207 7992
rect 4565 7970 4611 8016
rect 5057 8013 5103 8059
rect 4789 7954 4835 8000
rect 5537 7986 5583 8032
rect 5841 7986 5887 8032
rect 5985 7986 6031 8032
rect 6289 7986 6335 8032
rect 6625 7986 6671 8032
rect 6849 7986 6895 8032
rect 7933 8038 7979 8084
rect 7217 7946 7263 7992
rect 7441 7946 7487 7992
rect 7665 7946 7711 7992
rect 8085 8038 8131 8084
rect 8354 7936 8400 7982
rect 8498 7946 8544 7992
rect 8722 7946 8768 7992
rect 8977 7946 9023 7992
rect 9793 7986 9839 8032
rect 10017 7986 10063 8032
rect 10545 7986 10591 8032
rect 10769 7986 10815 8032
rect 11137 7946 11183 7992
rect 11392 7946 11438 7992
rect 11616 7946 11662 7992
rect 11760 7936 11806 7982
rect 12029 8038 12075 8084
rect 12181 8038 12227 8084
rect 12449 7946 12495 7992
rect 12673 7946 12719 7992
rect 12897 7946 12943 7992
rect 13569 7986 13615 8032
rect 13793 7986 13839 8032
rect 14273 7946 14319 7992
rect 14528 7946 14574 7992
rect 14752 7946 14798 7992
rect 14896 7936 14942 7982
rect 15165 8038 15211 8084
rect 15317 8038 15363 8084
rect 15585 7946 15631 7992
rect 15809 7946 15855 7992
rect 16033 7946 16079 7992
rect 16401 7986 16447 8032
rect 16625 7986 16671 8032
rect 17409 7986 17455 8032
rect 17633 7986 17679 8032
rect 17857 7986 17903 8032
rect 18161 7986 18207 8032
rect 1729 7648 1775 7694
rect 1953 7648 1999 7694
rect 2401 7688 2447 7734
rect 2625 7688 2671 7734
rect 2849 7688 2895 7734
rect 3117 7596 3163 7642
rect 3269 7596 3315 7642
rect 3538 7698 3584 7744
rect 3682 7688 3728 7734
rect 3906 7688 3952 7734
rect 4161 7688 4207 7734
rect 4609 7648 4655 7694
rect 4833 7648 4879 7694
rect 4977 7648 5023 7694
rect 5281 7648 5327 7694
rect 5425 7648 5471 7694
rect 5729 7648 5775 7694
rect 5873 7648 5919 7694
rect 6177 7648 6223 7694
rect 6321 7648 6367 7694
rect 6625 7648 6671 7694
rect 6769 7648 6815 7694
rect 7073 7648 7119 7694
rect 7217 7688 7263 7734
rect 7441 7688 7487 7734
rect 7665 7688 7711 7734
rect 7933 7596 7979 7642
rect 8085 7596 8131 7642
rect 8354 7698 8400 7744
rect 8498 7688 8544 7734
rect 8722 7688 8768 7734
rect 8977 7688 9023 7734
rect 9569 7648 9615 7694
rect 9873 7648 9919 7694
rect 10017 7648 10063 7694
rect 10241 7648 10287 7694
rect 10689 7648 10735 7694
rect 10913 7648 10959 7694
rect 11361 7648 11407 7694
rect 11585 7648 11631 7694
rect 12033 7688 12079 7734
rect 12257 7688 12303 7734
rect 12481 7688 12527 7734
rect 12749 7596 12795 7642
rect 12901 7596 12947 7642
rect 13170 7698 13216 7744
rect 13314 7688 13360 7734
rect 13538 7688 13584 7734
rect 13793 7688 13839 7734
rect 13937 7648 13983 7694
rect 14241 7648 14287 7694
rect 14385 7688 14431 7734
rect 14640 7688 14686 7734
rect 14864 7688 14910 7734
rect 15008 7698 15054 7744
rect 15277 7596 15323 7642
rect 15697 7688 15743 7734
rect 15921 7688 15967 7734
rect 16145 7688 16191 7734
rect 15429 7596 15475 7642
rect 16513 7648 16559 7694
rect 16737 7648 16783 7694
rect 17633 7648 17679 7694
rect 17857 7648 17903 7694
rect 1617 6418 1663 6464
rect 1921 6418 1967 6464
rect 2086 6418 2132 6464
rect 2310 6377 2356 6423
rect 2582 6378 2628 6424
rect 2806 6378 2852 6424
rect 3221 6402 3267 6448
rect 3713 6445 3759 6491
rect 3445 6386 3491 6432
rect 3857 6418 3903 6464
rect 4161 6418 4207 6464
rect 4305 6418 4351 6464
rect 4609 6418 4655 6464
rect 4753 6418 4799 6464
rect 5057 6418 5103 6464
rect 5537 6418 5583 6464
rect 5841 6418 5887 6464
rect 5985 6418 6031 6464
rect 6289 6418 6335 6464
rect 6848 6401 6894 6447
rect 7072 6398 7118 6444
rect 7441 6418 7487 6464
rect 7665 6418 7711 6464
rect 8113 6418 8159 6464
rect 8337 6418 8383 6464
rect 8785 6418 8831 6464
rect 9009 6418 9055 6464
rect 9457 6418 9503 6464
rect 9681 6418 9727 6464
rect 10129 6418 10175 6464
rect 10353 6418 10399 6464
rect 10801 6418 10847 6464
rect 11025 6418 11071 6464
rect 11473 6418 11519 6464
rect 11697 6418 11743 6464
rect 12145 6418 12191 6464
rect 12369 6418 12415 6464
rect 12593 6418 12639 6464
rect 12897 6418 12943 6464
rect 13601 6418 13647 6464
rect 13825 6418 13871 6464
rect 14273 6418 14319 6464
rect 14497 6418 14543 6464
rect 14945 6418 14991 6464
rect 15169 6418 15215 6464
rect 15617 6418 15663 6464
rect 15841 6418 15887 6464
rect 16289 6418 16335 6464
rect 16513 6418 16559 6464
rect 16961 6418 17007 6464
rect 17185 6418 17231 6464
rect 17633 6418 17679 6464
rect 17857 6418 17903 6464
rect 2181 6130 2227 6176
rect 1729 6054 1775 6100
rect 2405 6054 2451 6100
rect 2849 6080 2895 6126
rect 3073 6080 3119 6126
rect 3297 6080 3343 6126
rect 3601 6080 3647 6126
rect 3745 6080 3791 6126
rect 4049 6080 4095 6126
rect 4193 6080 4239 6126
rect 4497 6080 4543 6126
rect 4641 6080 4687 6126
rect 4945 6080 4991 6126
rect 5426 6100 5472 6146
rect 5650 6097 5696 6143
rect 6177 6080 6223 6126
rect 6401 6080 6447 6126
rect 6849 6080 6895 6126
rect 7073 6080 7119 6126
rect 7441 6080 7487 6126
rect 7665 6080 7711 6126
rect 8114 6100 8160 6146
rect 8338 6097 8384 6143
rect 8785 6080 8831 6126
rect 9009 6080 9055 6126
rect 9569 6080 9615 6126
rect 9873 6080 9919 6126
rect 10241 6080 10287 6126
rect 10465 6080 10511 6126
rect 10913 6080 10959 6126
rect 11137 6080 11183 6126
rect 11585 6080 11631 6126
rect 11809 6080 11855 6126
rect 12257 6080 12303 6126
rect 12481 6080 12527 6126
rect 12929 6080 12975 6126
rect 13153 6080 13199 6126
rect 13601 6080 13647 6126
rect 13825 6080 13871 6126
rect 14273 6080 14319 6126
rect 14497 6080 14543 6126
rect 14945 6080 14991 6126
rect 15169 6080 15215 6126
rect 15617 6080 15663 6126
rect 15841 6080 15887 6126
rect 16290 6100 16336 6146
rect 16514 6097 16560 6143
rect 16737 6080 16783 6126
rect 17041 6080 17087 6126
rect 17712 6097 17758 6143
rect 17936 6100 17982 6146
rect 1617 4850 1663 4896
rect 1921 4850 1967 4896
rect 2065 4850 2111 4896
rect 2369 4850 2415 4896
rect 2513 4850 2559 4896
rect 2817 4850 2863 4896
rect 2961 4850 3007 4896
rect 3265 4850 3311 4896
rect 3409 4850 3455 4896
rect 3713 4850 3759 4896
rect 4082 4830 4128 4876
rect 4306 4833 4352 4879
rect 4754 4830 4800 4876
rect 4978 4833 5024 4879
rect 5537 4850 5583 4896
rect 5841 4850 5887 4896
rect 6210 4830 6256 4876
rect 6434 4833 6480 4879
rect 6960 4833 7006 4879
rect 7184 4830 7230 4876
rect 7633 4850 7679 4896
rect 7857 4850 7903 4896
rect 8226 4830 8272 4876
rect 8450 4833 8496 4879
rect 8897 4850 8943 4896
rect 9121 4850 9167 4896
rect 9569 4850 9615 4896
rect 9793 4850 9839 4896
rect 10241 4850 10287 4896
rect 10465 4850 10511 4896
rect 10913 4850 10959 4896
rect 11137 4850 11183 4896
rect 11585 4850 11631 4896
rect 11809 4850 11855 4896
rect 12257 4850 12303 4896
rect 12481 4850 12527 4896
rect 12705 4850 12751 4896
rect 13009 4850 13055 4896
rect 13601 4850 13647 4896
rect 13825 4850 13871 4896
rect 14273 4850 14319 4896
rect 14497 4850 14543 4896
rect 15025 4850 15071 4896
rect 15249 4850 15295 4896
rect 15696 4833 15742 4879
rect 15920 4830 15966 4876
rect 16401 4810 16447 4856
rect 16656 4810 16702 4856
rect 16880 4810 16926 4856
rect 17024 4800 17070 4846
rect 17293 4902 17339 4948
rect 17445 4902 17491 4948
rect 17713 4810 17759 4856
rect 17937 4810 17983 4856
rect 18161 4810 18207 4856
rect 1617 4512 1663 4558
rect 1921 4512 1967 4558
rect 2065 4512 2111 4558
rect 2369 4512 2415 4558
rect 2625 4552 2671 4598
rect 2849 4552 2895 4598
rect 3073 4552 3119 4598
rect 3341 4460 3387 4506
rect 3493 4460 3539 4506
rect 3762 4562 3808 4608
rect 3906 4552 3952 4598
rect 4130 4552 4176 4598
rect 4385 4552 4431 4598
rect 4529 4512 4575 4558
rect 4833 4512 4879 4558
rect 5090 4532 5136 4578
rect 5314 4529 5360 4575
rect 5762 4532 5808 4578
rect 5986 4529 6032 4575
rect 6434 4532 6480 4578
rect 6658 4529 6704 4575
rect 7105 4552 7151 4598
rect 7360 4552 7406 4598
rect 7584 4552 7630 4598
rect 7728 4562 7774 4608
rect 7997 4460 8043 4506
rect 8417 4552 8463 4598
rect 8641 4552 8687 4598
rect 8865 4552 8911 4598
rect 8149 4460 8195 4506
rect 9569 4512 9615 4558
rect 9873 4512 9919 4558
rect 10018 4532 10064 4578
rect 10242 4529 10288 4575
rect 10769 4512 10815 4558
rect 10993 4512 11039 4558
rect 11441 4512 11487 4558
rect 11665 4512 11711 4558
rect 12033 4552 12079 4598
rect 12288 4552 12334 4598
rect 12512 4552 12558 4598
rect 12656 4562 12702 4608
rect 12925 4460 12971 4506
rect 13345 4552 13391 4598
rect 13569 4552 13615 4598
rect 13793 4552 13839 4598
rect 13077 4460 13123 4506
rect 14162 4532 14208 4578
rect 14386 4529 14432 4575
rect 14833 4512 14879 4558
rect 15057 4512 15103 4558
rect 15505 4512 15551 4558
rect 15729 4512 15775 4558
rect 16177 4512 16223 4558
rect 16401 4512 16447 4558
rect 16625 4512 16671 4558
rect 16929 4512 16975 4558
rect 17633 4512 17679 4558
rect 17857 4512 17903 4558
rect 1954 3262 2000 3308
rect 2178 3265 2224 3311
rect 2625 3242 2671 3288
rect 2880 3242 2926 3288
rect 3104 3242 3150 3288
rect 3248 3232 3294 3278
rect 3517 3334 3563 3380
rect 3669 3334 3715 3380
rect 3937 3242 3983 3288
rect 4161 3242 4207 3288
rect 4385 3242 4431 3288
rect 4754 3262 4800 3308
rect 4978 3265 5024 3311
rect 5874 3262 5920 3308
rect 6098 3265 6144 3311
rect 6546 3262 6592 3308
rect 6770 3265 6816 3311
rect 7217 3242 7263 3288
rect 7472 3242 7518 3288
rect 7696 3242 7742 3288
rect 7840 3232 7886 3278
rect 8109 3334 8155 3380
rect 8261 3334 8307 3380
rect 8529 3242 8575 3288
rect 8753 3242 8799 3288
rect 8977 3242 9023 3288
rect 9794 3262 9840 3308
rect 10018 3265 10064 3311
rect 10466 3262 10512 3308
rect 10690 3265 10736 3311
rect 11137 3242 11183 3288
rect 11392 3242 11438 3288
rect 11616 3242 11662 3288
rect 11760 3232 11806 3278
rect 12029 3334 12075 3380
rect 12181 3334 12227 3380
rect 12449 3242 12495 3288
rect 12673 3242 12719 3288
rect 12897 3242 12943 3288
rect 13569 3282 13615 3328
rect 13793 3282 13839 3328
rect 14162 3262 14208 3308
rect 14386 3265 14432 3311
rect 14609 3282 14655 3328
rect 14913 3282 14959 3328
rect 15057 3242 15103 3288
rect 15312 3242 15358 3288
rect 15536 3242 15582 3288
rect 15680 3232 15726 3278
rect 15949 3334 15995 3380
rect 16101 3334 16147 3380
rect 16369 3242 16415 3288
rect 16593 3242 16639 3288
rect 16817 3242 16863 3288
rect 17488 3265 17534 3311
rect 17712 3262 17758 3308
rect 17857 3282 17903 3328
rect 18161 3282 18207 3328
<< mvpdiffc >>
rect 1749 8365 1795 8505
rect 1953 8365 1999 8505
rect 2401 8439 2447 8485
rect 2605 8439 2651 8485
rect 2809 8439 2855 8485
rect 3057 8375 3103 8421
rect 3271 8361 3317 8407
rect 3475 8481 3521 8527
rect 3702 8456 3748 8502
rect 3906 8474 3952 8520
rect 4141 8456 4187 8502
rect 4585 8365 4631 8505
rect 4789 8481 4835 8527
rect 5037 8462 5083 8508
rect 5537 8357 5583 8497
rect 5841 8357 5887 8497
rect 5985 8357 6031 8497
rect 6289 8357 6335 8497
rect 6625 8365 6671 8505
rect 6829 8365 6875 8505
rect 7217 8439 7263 8485
rect 7421 8439 7467 8485
rect 7625 8439 7671 8485
rect 7873 8375 7919 8421
rect 8087 8361 8133 8407
rect 8291 8481 8337 8527
rect 8518 8456 8564 8502
rect 8722 8474 8768 8520
rect 8957 8456 9003 8502
rect 9813 8365 9859 8505
rect 10017 8365 10063 8505
rect 10545 8365 10591 8505
rect 10749 8365 10795 8505
rect 11157 8456 11203 8502
rect 11392 8474 11438 8520
rect 11596 8456 11642 8502
rect 11823 8481 11869 8527
rect 12027 8361 12073 8407
rect 12241 8375 12287 8421
rect 12489 8439 12535 8485
rect 12693 8439 12739 8485
rect 12897 8439 12943 8485
rect 13569 8365 13615 8505
rect 13773 8365 13819 8505
rect 14293 8456 14339 8502
rect 14528 8474 14574 8520
rect 14732 8456 14778 8502
rect 14959 8481 15005 8527
rect 15163 8361 15209 8407
rect 15377 8375 15423 8421
rect 15625 8439 15671 8485
rect 15829 8439 15875 8485
rect 16033 8439 16079 8485
rect 16421 8365 16467 8505
rect 16625 8365 16671 8505
rect 17429 8365 17475 8505
rect 17633 8365 17679 8505
rect 17857 8357 17903 8497
rect 18161 8357 18207 8497
rect 1749 7175 1795 7315
rect 1953 7175 1999 7315
rect 2401 7195 2447 7241
rect 2605 7195 2651 7241
rect 2809 7195 2855 7241
rect 3057 7259 3103 7305
rect 3271 7273 3317 7319
rect 3475 7153 3521 7199
rect 3702 7178 3748 7224
rect 3906 7160 3952 7206
rect 4141 7178 4187 7224
rect 4609 7175 4655 7315
rect 4813 7175 4859 7315
rect 4977 7183 5023 7323
rect 5281 7183 5327 7323
rect 5425 7183 5471 7323
rect 5729 7183 5775 7323
rect 5873 7183 5919 7323
rect 6177 7183 6223 7323
rect 6321 7183 6367 7323
rect 6625 7183 6671 7323
rect 6769 7183 6815 7323
rect 7073 7183 7119 7323
rect 7217 7195 7263 7241
rect 7421 7195 7467 7241
rect 7625 7195 7671 7241
rect 7873 7259 7919 7305
rect 8087 7273 8133 7319
rect 8291 7153 8337 7199
rect 8518 7178 8564 7224
rect 8722 7160 8768 7206
rect 8957 7178 9003 7224
rect 9569 7183 9615 7323
rect 9873 7183 9919 7323
rect 10037 7175 10083 7315
rect 10241 7175 10287 7315
rect 10709 7175 10755 7315
rect 10913 7175 10959 7315
rect 11381 7175 11427 7315
rect 11585 7175 11631 7315
rect 12033 7195 12079 7241
rect 12237 7195 12283 7241
rect 12441 7195 12487 7241
rect 12689 7259 12735 7305
rect 12903 7273 12949 7319
rect 13107 7153 13153 7199
rect 13334 7178 13380 7224
rect 13538 7160 13584 7206
rect 13773 7178 13819 7224
rect 13937 7183 13983 7323
rect 14241 7183 14287 7323
rect 14405 7178 14451 7224
rect 14640 7160 14686 7206
rect 14844 7178 14890 7224
rect 15071 7153 15117 7199
rect 15275 7273 15321 7319
rect 15489 7259 15535 7305
rect 15737 7195 15783 7241
rect 15941 7195 15987 7241
rect 16145 7195 16191 7241
rect 16533 7175 16579 7315
rect 16737 7175 16783 7315
rect 17653 7175 17699 7315
rect 17857 7175 17903 7315
rect 1617 6789 1663 6929
rect 1921 6789 1967 6929
rect 2106 6797 2152 6937
rect 2310 6797 2356 6937
rect 2786 6898 2832 6944
rect 3241 6797 3287 6937
rect 3445 6913 3491 6959
rect 3693 6894 3739 6940
rect 3857 6789 3903 6929
rect 4161 6789 4207 6929
rect 4305 6789 4351 6929
rect 4609 6789 4655 6929
rect 4753 6789 4799 6929
rect 5057 6789 5103 6929
rect 5537 6789 5583 6929
rect 5841 6789 5887 6929
rect 5985 6789 6031 6929
rect 6289 6789 6335 6929
rect 6868 6781 6914 6921
rect 7072 6781 7118 6921
rect 7461 6797 7507 6937
rect 7665 6797 7711 6937
rect 8133 6797 8179 6937
rect 8337 6797 8383 6937
rect 8805 6797 8851 6937
rect 9009 6797 9055 6937
rect 9477 6797 9523 6937
rect 9681 6797 9727 6937
rect 10149 6797 10195 6937
rect 10353 6797 10399 6937
rect 10821 6797 10867 6937
rect 11025 6797 11071 6937
rect 11493 6797 11539 6937
rect 11697 6797 11743 6937
rect 12165 6797 12211 6937
rect 12369 6797 12415 6937
rect 12593 6789 12639 6929
rect 12897 6789 12943 6929
rect 13621 6797 13667 6937
rect 13825 6797 13871 6937
rect 14293 6797 14339 6937
rect 14497 6797 14543 6937
rect 14965 6797 15011 6937
rect 15169 6797 15215 6937
rect 15637 6797 15683 6937
rect 15841 6797 15887 6937
rect 16309 6797 16355 6937
rect 16513 6797 16559 6937
rect 16981 6797 17027 6937
rect 17185 6797 17231 6937
rect 17653 6797 17699 6937
rect 17857 6797 17903 6937
rect 1729 5570 1775 5616
rect 1933 5618 1979 5664
rect 2201 5607 2247 5747
rect 2405 5607 2451 5747
rect 2869 5607 2915 5747
rect 3073 5607 3119 5747
rect 3297 5615 3343 5755
rect 3601 5615 3647 5755
rect 3745 5615 3791 5755
rect 4049 5615 4095 5755
rect 4193 5615 4239 5755
rect 4497 5615 4543 5755
rect 4641 5615 4687 5755
rect 4945 5615 4991 5755
rect 5426 5623 5472 5763
rect 5630 5623 5676 5763
rect 6177 5607 6223 5747
rect 6381 5607 6427 5747
rect 6849 5607 6895 5747
rect 7053 5607 7099 5747
rect 7461 5607 7507 5747
rect 7665 5607 7711 5747
rect 8114 5623 8160 5763
rect 8318 5623 8364 5763
rect 8805 5607 8851 5747
rect 9009 5607 9055 5747
rect 9569 5615 9615 5755
rect 9873 5615 9919 5755
rect 10261 5607 10307 5747
rect 10465 5607 10511 5747
rect 10933 5607 10979 5747
rect 11137 5607 11183 5747
rect 11605 5607 11651 5747
rect 11809 5607 11855 5747
rect 12277 5607 12323 5747
rect 12481 5607 12527 5747
rect 12949 5607 12995 5747
rect 13153 5607 13199 5747
rect 13621 5607 13667 5747
rect 13825 5607 13871 5747
rect 14293 5607 14339 5747
rect 14497 5607 14543 5747
rect 14965 5607 15011 5747
rect 15169 5607 15215 5747
rect 15637 5607 15683 5747
rect 15841 5607 15887 5747
rect 16290 5623 16336 5763
rect 16494 5623 16540 5763
rect 16737 5615 16783 5755
rect 17041 5615 17087 5755
rect 17732 5623 17778 5763
rect 17936 5623 17982 5763
rect 1617 5221 1663 5361
rect 1921 5221 1967 5361
rect 2065 5221 2111 5361
rect 2369 5221 2415 5361
rect 2513 5221 2559 5361
rect 2817 5221 2863 5361
rect 2961 5221 3007 5361
rect 3265 5221 3311 5361
rect 3409 5221 3455 5361
rect 3713 5221 3759 5361
rect 4082 5213 4128 5353
rect 4286 5213 4332 5353
rect 4754 5213 4800 5353
rect 4958 5213 5004 5353
rect 5537 5221 5583 5361
rect 5841 5221 5887 5361
rect 6210 5213 6256 5353
rect 6414 5213 6460 5353
rect 6980 5213 7026 5353
rect 7184 5213 7230 5353
rect 7633 5229 7679 5369
rect 7837 5229 7883 5369
rect 8226 5213 8272 5353
rect 8430 5213 8476 5353
rect 8917 5229 8963 5369
rect 9121 5229 9167 5369
rect 9589 5229 9635 5369
rect 9793 5229 9839 5369
rect 10261 5229 10307 5369
rect 10465 5229 10511 5369
rect 10933 5229 10979 5369
rect 11137 5229 11183 5369
rect 11605 5229 11651 5369
rect 11809 5229 11855 5369
rect 12277 5229 12323 5369
rect 12481 5229 12527 5369
rect 12705 5221 12751 5361
rect 13009 5221 13055 5361
rect 13621 5229 13667 5369
rect 13825 5229 13871 5369
rect 14293 5229 14339 5369
rect 14497 5229 14543 5369
rect 15025 5229 15071 5369
rect 15229 5229 15275 5369
rect 15716 5213 15762 5353
rect 15920 5213 15966 5353
rect 16421 5320 16467 5366
rect 16656 5338 16702 5384
rect 16860 5320 16906 5366
rect 17087 5345 17133 5391
rect 17291 5225 17337 5271
rect 17505 5239 17551 5285
rect 17753 5303 17799 5349
rect 17957 5303 18003 5349
rect 18161 5303 18207 5349
rect 1617 4047 1663 4187
rect 1921 4047 1967 4187
rect 2065 4047 2111 4187
rect 2369 4047 2415 4187
rect 2625 4059 2671 4105
rect 2829 4059 2875 4105
rect 3033 4059 3079 4105
rect 3281 4123 3327 4169
rect 3495 4137 3541 4183
rect 3699 4017 3745 4063
rect 3926 4042 3972 4088
rect 4130 4024 4176 4070
rect 4365 4042 4411 4088
rect 4529 4047 4575 4187
rect 4833 4047 4879 4187
rect 5090 4055 5136 4195
rect 5294 4055 5340 4195
rect 5762 4055 5808 4195
rect 5966 4055 6012 4195
rect 6434 4055 6480 4195
rect 6638 4055 6684 4195
rect 7125 4042 7171 4088
rect 7360 4024 7406 4070
rect 7564 4042 7610 4088
rect 7791 4017 7837 4063
rect 7995 4137 8041 4183
rect 8209 4123 8255 4169
rect 8457 4059 8503 4105
rect 8661 4059 8707 4105
rect 8865 4059 8911 4105
rect 9569 4047 9615 4187
rect 9873 4047 9919 4187
rect 10018 4055 10064 4195
rect 10222 4055 10268 4195
rect 10769 4039 10815 4179
rect 10973 4039 11019 4179
rect 11441 4039 11487 4179
rect 11645 4039 11691 4179
rect 12053 4042 12099 4088
rect 12288 4024 12334 4070
rect 12492 4042 12538 4088
rect 12719 4017 12765 4063
rect 12923 4137 12969 4183
rect 13137 4123 13183 4169
rect 13385 4059 13431 4105
rect 13589 4059 13635 4105
rect 13793 4059 13839 4105
rect 14162 4055 14208 4195
rect 14366 4055 14412 4195
rect 14853 4039 14899 4179
rect 15057 4039 15103 4179
rect 15525 4039 15571 4179
rect 15729 4039 15775 4179
rect 16197 4039 16243 4179
rect 16401 4039 16447 4179
rect 16625 4047 16671 4187
rect 16929 4047 16975 4187
rect 17653 4039 17699 4179
rect 17857 4039 17903 4179
rect 1954 3645 2000 3785
rect 2158 3645 2204 3785
rect 2645 3752 2691 3798
rect 2880 3770 2926 3816
rect 3084 3752 3130 3798
rect 3311 3777 3357 3823
rect 3515 3657 3561 3703
rect 3729 3671 3775 3717
rect 3977 3735 4023 3781
rect 4181 3735 4227 3781
rect 4385 3735 4431 3781
rect 4754 3645 4800 3785
rect 4958 3645 5004 3785
rect 5874 3645 5920 3785
rect 6078 3645 6124 3785
rect 6546 3645 6592 3785
rect 6750 3645 6796 3785
rect 7237 3752 7283 3798
rect 7472 3770 7518 3816
rect 7676 3752 7722 3798
rect 7903 3777 7949 3823
rect 8107 3657 8153 3703
rect 8321 3671 8367 3717
rect 8569 3735 8615 3781
rect 8773 3735 8819 3781
rect 8977 3735 9023 3781
rect 9794 3645 9840 3785
rect 9998 3645 10044 3785
rect 10466 3645 10512 3785
rect 10670 3645 10716 3785
rect 11157 3752 11203 3798
rect 11392 3770 11438 3816
rect 11596 3752 11642 3798
rect 11823 3777 11869 3823
rect 12027 3657 12073 3703
rect 12241 3671 12287 3717
rect 12489 3735 12535 3781
rect 12693 3735 12739 3781
rect 12897 3735 12943 3781
rect 13569 3661 13615 3801
rect 13773 3661 13819 3801
rect 14162 3645 14208 3785
rect 14366 3645 14412 3785
rect 14609 3653 14655 3793
rect 14913 3653 14959 3793
rect 15077 3752 15123 3798
rect 15312 3770 15358 3816
rect 15516 3752 15562 3798
rect 15743 3777 15789 3823
rect 15947 3657 15993 3703
rect 16161 3671 16207 3717
rect 16409 3735 16455 3781
rect 16613 3735 16659 3781
rect 16817 3735 16863 3781
rect 17508 3645 17554 3785
rect 17712 3645 17758 3785
rect 17857 3653 17903 3793
rect 18161 3653 18207 3793
<< mvpsubdiff >>
rect 1400 8066 1504 8096
rect 1400 7919 1429 8066
rect 1475 7919 1504 8066
rect 1400 7896 1504 7919
rect 5320 8066 5432 8096
rect 5320 7919 5353 8066
rect 5399 7919 5432 8066
rect 5320 7896 5432 7919
rect 9240 8066 9352 8096
rect 9240 7919 9273 8066
rect 9319 7919 9352 8066
rect 9240 7896 9352 7919
rect 13160 8066 13272 8096
rect 13160 7919 13193 8066
rect 13239 7919 13272 8066
rect 13160 7896 13272 7919
rect 17080 8066 17192 8096
rect 17080 7919 17113 8066
rect 17159 7919 17192 8066
rect 17080 7896 17192 7919
rect 18432 8066 18536 8096
rect 18432 7919 18461 8066
rect 18507 7919 18536 8066
rect 18432 7896 18536 7919
rect 1400 7761 1504 7784
rect 1400 7614 1429 7761
rect 1475 7614 1504 7761
rect 1400 7584 1504 7614
rect 9352 7761 9464 7784
rect 9352 7614 9385 7761
rect 9431 7614 9464 7761
rect 9352 7584 9464 7614
rect 17304 7761 17416 7784
rect 17304 7614 17337 7761
rect 17383 7614 17416 7761
rect 17304 7584 17416 7614
rect 18432 7761 18536 7784
rect 18432 7614 18461 7761
rect 18507 7614 18536 7761
rect 18432 7584 18536 7614
rect 1400 6498 1504 6528
rect 1400 6351 1429 6498
rect 1475 6351 1504 6498
rect 1400 6328 1504 6351
rect 5320 6498 5432 6528
rect 5320 6351 5353 6498
rect 5399 6351 5432 6498
rect 5320 6328 5432 6351
rect 13272 6498 13384 6528
rect 13272 6351 13305 6498
rect 13351 6351 13384 6498
rect 13272 6328 13384 6351
rect 18432 6498 18536 6528
rect 18432 6351 18461 6498
rect 18507 6351 18536 6498
rect 18432 6328 18536 6351
rect 1400 6193 1504 6216
rect 1400 6046 1429 6193
rect 1475 6046 1504 6193
rect 1400 6016 1504 6046
rect 9352 6193 9464 6216
rect 9352 6046 9385 6193
rect 9431 6046 9464 6193
rect 9352 6016 9464 6046
rect 17304 6193 17416 6216
rect 17304 6046 17337 6193
rect 17383 6046 17416 6193
rect 17304 6016 17416 6046
rect 18432 6193 18536 6216
rect 18432 6046 18461 6193
rect 18507 6046 18536 6193
rect 18432 6016 18536 6046
rect 1400 4930 1504 4960
rect 1400 4783 1429 4930
rect 1475 4783 1504 4930
rect 1400 4760 1504 4783
rect 5320 4930 5432 4960
rect 5320 4783 5353 4930
rect 5399 4783 5432 4930
rect 5320 4760 5432 4783
rect 13272 4930 13384 4960
rect 13272 4783 13305 4930
rect 13351 4783 13384 4930
rect 13272 4760 13384 4783
rect 18432 4930 18536 4960
rect 18432 4783 18461 4930
rect 18507 4783 18536 4930
rect 18432 4760 18536 4783
rect 1400 4625 1504 4648
rect 1400 4478 1429 4625
rect 1475 4478 1504 4625
rect 1400 4448 1504 4478
rect 9352 4625 9464 4648
rect 9352 4478 9385 4625
rect 9431 4478 9464 4625
rect 9352 4448 9464 4478
rect 17304 4625 17416 4648
rect 17304 4478 17337 4625
rect 17383 4478 17416 4625
rect 17304 4448 17416 4478
rect 18432 4625 18536 4648
rect 18432 4478 18461 4625
rect 18507 4478 18536 4625
rect 18432 4448 18536 4478
rect 1400 3362 1504 3392
rect 1400 3215 1429 3362
rect 1475 3215 1504 3362
rect 1400 3192 1504 3215
rect 5320 3362 5432 3392
rect 5320 3215 5353 3362
rect 5399 3215 5432 3362
rect 5320 3192 5432 3215
rect 9240 3362 9352 3392
rect 9240 3215 9273 3362
rect 9319 3215 9352 3362
rect 9240 3192 9352 3215
rect 13160 3362 13272 3392
rect 13160 3215 13193 3362
rect 13239 3215 13272 3362
rect 13160 3192 13272 3215
rect 17080 3362 17192 3392
rect 17080 3215 17113 3362
rect 17159 3215 17192 3362
rect 17080 3192 17192 3215
rect 18432 3362 18536 3392
rect 18432 3215 18461 3362
rect 18507 3215 18536 3362
rect 18432 3192 18536 3215
<< mvnsubdiff >>
rect 1416 8539 1488 8552
rect 1416 8493 1429 8539
rect 1475 8493 1488 8539
rect 1416 8411 1488 8493
rect 1416 8365 1429 8411
rect 1475 8365 1488 8411
rect 1416 8283 1488 8365
rect 1416 8237 1429 8283
rect 1475 8237 1488 8283
rect 1416 8224 1488 8237
rect 5336 8539 5416 8552
rect 5336 8493 5353 8539
rect 5399 8493 5416 8539
rect 5336 8411 5416 8493
rect 5336 8365 5353 8411
rect 5399 8365 5416 8411
rect 5336 8283 5416 8365
rect 5336 8237 5353 8283
rect 5399 8237 5416 8283
rect 5336 8224 5416 8237
rect 9256 8539 9336 8552
rect 9256 8493 9273 8539
rect 9319 8493 9336 8539
rect 9256 8411 9336 8493
rect 9256 8365 9273 8411
rect 9319 8365 9336 8411
rect 9256 8283 9336 8365
rect 9256 8237 9273 8283
rect 9319 8237 9336 8283
rect 9256 8224 9336 8237
rect 13176 8539 13256 8552
rect 13176 8493 13193 8539
rect 13239 8493 13256 8539
rect 13176 8411 13256 8493
rect 13176 8365 13193 8411
rect 13239 8365 13256 8411
rect 13176 8283 13256 8365
rect 13176 8237 13193 8283
rect 13239 8237 13256 8283
rect 13176 8224 13256 8237
rect 17096 8539 17176 8552
rect 17096 8493 17113 8539
rect 17159 8493 17176 8539
rect 17096 8411 17176 8493
rect 17096 8365 17113 8411
rect 17159 8365 17176 8411
rect 17096 8283 17176 8365
rect 18448 8539 18520 8552
rect 18448 8493 18461 8539
rect 18507 8493 18520 8539
rect 18448 8411 18520 8493
rect 18448 8365 18461 8411
rect 18507 8365 18520 8411
rect 17096 8237 17113 8283
rect 17159 8237 17176 8283
rect 17096 8224 17176 8237
rect 18448 8283 18520 8365
rect 18448 8237 18461 8283
rect 18507 8237 18520 8283
rect 18448 8224 18520 8237
rect 1416 7443 1488 7456
rect 1416 7397 1429 7443
rect 1475 7397 1488 7443
rect 1416 7315 1488 7397
rect 1416 7269 1429 7315
rect 1475 7269 1488 7315
rect 1416 7187 1488 7269
rect 1416 7141 1429 7187
rect 1475 7141 1488 7187
rect 1416 7128 1488 7141
rect 9368 7443 9448 7456
rect 9368 7397 9385 7443
rect 9431 7397 9448 7443
rect 9368 7315 9448 7397
rect 9368 7269 9385 7315
rect 9431 7269 9448 7315
rect 9368 7187 9448 7269
rect 9368 7141 9385 7187
rect 9431 7141 9448 7187
rect 9368 7128 9448 7141
rect 17320 7443 17400 7456
rect 17320 7397 17337 7443
rect 17383 7397 17400 7443
rect 17320 7315 17400 7397
rect 18448 7443 18520 7456
rect 18448 7397 18461 7443
rect 18507 7397 18520 7443
rect 17320 7269 17337 7315
rect 17383 7269 17400 7315
rect 17320 7187 17400 7269
rect 17320 7141 17337 7187
rect 17383 7141 17400 7187
rect 17320 7128 17400 7141
rect 18448 7315 18520 7397
rect 18448 7269 18461 7315
rect 18507 7269 18520 7315
rect 18448 7187 18520 7269
rect 18448 7141 18461 7187
rect 18507 7141 18520 7187
rect 18448 7128 18520 7141
rect 1416 6971 1488 6984
rect 1416 6925 1429 6971
rect 1475 6925 1488 6971
rect 1416 6843 1488 6925
rect 1416 6797 1429 6843
rect 1475 6797 1488 6843
rect 1416 6715 1488 6797
rect 1416 6669 1429 6715
rect 1475 6669 1488 6715
rect 1416 6656 1488 6669
rect 5336 6971 5416 6984
rect 5336 6925 5353 6971
rect 5399 6925 5416 6971
rect 5336 6843 5416 6925
rect 5336 6797 5353 6843
rect 5399 6797 5416 6843
rect 5336 6715 5416 6797
rect 13288 6971 13368 6984
rect 13288 6925 13305 6971
rect 13351 6925 13368 6971
rect 13288 6843 13368 6925
rect 13288 6797 13305 6843
rect 13351 6797 13368 6843
rect 5336 6669 5353 6715
rect 5399 6669 5416 6715
rect 5336 6656 5416 6669
rect 13288 6715 13368 6797
rect 18448 6971 18520 6984
rect 18448 6925 18461 6971
rect 18507 6925 18520 6971
rect 18448 6843 18520 6925
rect 18448 6797 18461 6843
rect 18507 6797 18520 6843
rect 13288 6669 13305 6715
rect 13351 6669 13368 6715
rect 13288 6656 13368 6669
rect 18448 6715 18520 6797
rect 18448 6669 18461 6715
rect 18507 6669 18520 6715
rect 18448 6656 18520 6669
rect 1416 5875 1488 5888
rect 1416 5829 1429 5875
rect 1475 5829 1488 5875
rect 1416 5747 1488 5829
rect 1416 5701 1429 5747
rect 1475 5701 1488 5747
rect 1416 5619 1488 5701
rect 9368 5875 9448 5888
rect 9368 5829 9385 5875
rect 9431 5829 9448 5875
rect 1416 5573 1429 5619
rect 1475 5573 1488 5619
rect 1416 5560 1488 5573
rect 9368 5747 9448 5829
rect 17320 5875 17400 5888
rect 17320 5829 17337 5875
rect 17383 5829 17400 5875
rect 9368 5701 9385 5747
rect 9431 5701 9448 5747
rect 9368 5619 9448 5701
rect 9368 5573 9385 5619
rect 9431 5573 9448 5619
rect 9368 5560 9448 5573
rect 17320 5747 17400 5829
rect 18448 5875 18520 5888
rect 18448 5829 18461 5875
rect 18507 5829 18520 5875
rect 17320 5701 17337 5747
rect 17383 5701 17400 5747
rect 17320 5619 17400 5701
rect 17320 5573 17337 5619
rect 17383 5573 17400 5619
rect 17320 5560 17400 5573
rect 18448 5747 18520 5829
rect 18448 5701 18461 5747
rect 18507 5701 18520 5747
rect 18448 5619 18520 5701
rect 18448 5573 18461 5619
rect 18507 5573 18520 5619
rect 18448 5560 18520 5573
rect 1416 5403 1488 5416
rect 1416 5357 1429 5403
rect 1475 5357 1488 5403
rect 1416 5275 1488 5357
rect 1416 5229 1429 5275
rect 1475 5229 1488 5275
rect 1416 5147 1488 5229
rect 5336 5403 5416 5416
rect 5336 5357 5353 5403
rect 5399 5357 5416 5403
rect 5336 5275 5416 5357
rect 5336 5229 5353 5275
rect 5399 5229 5416 5275
rect 1416 5101 1429 5147
rect 1475 5101 1488 5147
rect 1416 5088 1488 5101
rect 5336 5147 5416 5229
rect 13288 5403 13368 5416
rect 13288 5357 13305 5403
rect 13351 5357 13368 5403
rect 13288 5275 13368 5357
rect 13288 5229 13305 5275
rect 13351 5229 13368 5275
rect 5336 5101 5353 5147
rect 5399 5101 5416 5147
rect 5336 5088 5416 5101
rect 13288 5147 13368 5229
rect 13288 5101 13305 5147
rect 13351 5101 13368 5147
rect 13288 5088 13368 5101
rect 18448 5403 18520 5416
rect 18448 5357 18461 5403
rect 18507 5357 18520 5403
rect 18448 5275 18520 5357
rect 18448 5229 18461 5275
rect 18507 5229 18520 5275
rect 18448 5147 18520 5229
rect 18448 5101 18461 5147
rect 18507 5101 18520 5147
rect 18448 5088 18520 5101
rect 1416 4307 1488 4320
rect 1416 4261 1429 4307
rect 1475 4261 1488 4307
rect 1416 4179 1488 4261
rect 1416 4133 1429 4179
rect 1475 4133 1488 4179
rect 1416 4051 1488 4133
rect 1416 4005 1429 4051
rect 1475 4005 1488 4051
rect 1416 3992 1488 4005
rect 9368 4307 9448 4320
rect 9368 4261 9385 4307
rect 9431 4261 9448 4307
rect 9368 4179 9448 4261
rect 9368 4133 9385 4179
rect 9431 4133 9448 4179
rect 9368 4051 9448 4133
rect 9368 4005 9385 4051
rect 9431 4005 9448 4051
rect 9368 3992 9448 4005
rect 17320 4307 17400 4320
rect 17320 4261 17337 4307
rect 17383 4261 17400 4307
rect 17320 4179 17400 4261
rect 18448 4307 18520 4320
rect 18448 4261 18461 4307
rect 18507 4261 18520 4307
rect 17320 4133 17337 4179
rect 17383 4133 17400 4179
rect 17320 4051 17400 4133
rect 17320 4005 17337 4051
rect 17383 4005 17400 4051
rect 17320 3992 17400 4005
rect 18448 4179 18520 4261
rect 18448 4133 18461 4179
rect 18507 4133 18520 4179
rect 18448 4051 18520 4133
rect 18448 4005 18461 4051
rect 18507 4005 18520 4051
rect 18448 3992 18520 4005
rect 1416 3835 1488 3848
rect 1416 3789 1429 3835
rect 1475 3789 1488 3835
rect 1416 3707 1488 3789
rect 1416 3661 1429 3707
rect 1475 3661 1488 3707
rect 1416 3579 1488 3661
rect 1416 3533 1429 3579
rect 1475 3533 1488 3579
rect 1416 3520 1488 3533
rect 5336 3835 5416 3848
rect 5336 3789 5353 3835
rect 5399 3789 5416 3835
rect 5336 3707 5416 3789
rect 5336 3661 5353 3707
rect 5399 3661 5416 3707
rect 5336 3579 5416 3661
rect 5336 3533 5353 3579
rect 5399 3533 5416 3579
rect 5336 3520 5416 3533
rect 9256 3835 9336 3848
rect 9256 3789 9273 3835
rect 9319 3789 9336 3835
rect 9256 3707 9336 3789
rect 9256 3661 9273 3707
rect 9319 3661 9336 3707
rect 9256 3579 9336 3661
rect 9256 3533 9273 3579
rect 9319 3533 9336 3579
rect 9256 3520 9336 3533
rect 13176 3835 13256 3848
rect 13176 3789 13193 3835
rect 13239 3789 13256 3835
rect 13176 3707 13256 3789
rect 13176 3661 13193 3707
rect 13239 3661 13256 3707
rect 13176 3579 13256 3661
rect 13176 3533 13193 3579
rect 13239 3533 13256 3579
rect 13176 3520 13256 3533
rect 17096 3835 17176 3848
rect 17096 3789 17113 3835
rect 17159 3789 17176 3835
rect 17096 3707 17176 3789
rect 17096 3661 17113 3707
rect 17159 3661 17176 3707
rect 17096 3579 17176 3661
rect 18448 3835 18520 3848
rect 18448 3789 18461 3835
rect 18507 3789 18520 3835
rect 18448 3707 18520 3789
rect 18448 3661 18461 3707
rect 18507 3661 18520 3707
rect 17096 3533 17113 3579
rect 17159 3533 17176 3579
rect 17096 3520 17176 3533
rect 18448 3579 18520 3661
rect 18448 3533 18461 3579
rect 18507 3533 18520 3579
rect 18448 3520 18520 3533
<< mvpsubdiffcont >>
rect 1429 7919 1475 8066
rect 5353 7919 5399 8066
rect 9273 7919 9319 8066
rect 13193 7919 13239 8066
rect 17113 7919 17159 8066
rect 18461 7919 18507 8066
rect 1429 7614 1475 7761
rect 9385 7614 9431 7761
rect 17337 7614 17383 7761
rect 18461 7614 18507 7761
rect 1429 6351 1475 6498
rect 5353 6351 5399 6498
rect 13305 6351 13351 6498
rect 18461 6351 18507 6498
rect 1429 6046 1475 6193
rect 9385 6046 9431 6193
rect 17337 6046 17383 6193
rect 18461 6046 18507 6193
rect 1429 4783 1475 4930
rect 5353 4783 5399 4930
rect 13305 4783 13351 4930
rect 18461 4783 18507 4930
rect 1429 4478 1475 4625
rect 9385 4478 9431 4625
rect 17337 4478 17383 4625
rect 18461 4478 18507 4625
rect 1429 3215 1475 3362
rect 5353 3215 5399 3362
rect 9273 3215 9319 3362
rect 13193 3215 13239 3362
rect 17113 3215 17159 3362
rect 18461 3215 18507 3362
<< mvnsubdiffcont >>
rect 1429 8493 1475 8539
rect 1429 8365 1475 8411
rect 1429 8237 1475 8283
rect 5353 8493 5399 8539
rect 5353 8365 5399 8411
rect 5353 8237 5399 8283
rect 9273 8493 9319 8539
rect 9273 8365 9319 8411
rect 9273 8237 9319 8283
rect 13193 8493 13239 8539
rect 13193 8365 13239 8411
rect 13193 8237 13239 8283
rect 17113 8493 17159 8539
rect 17113 8365 17159 8411
rect 18461 8493 18507 8539
rect 18461 8365 18507 8411
rect 17113 8237 17159 8283
rect 18461 8237 18507 8283
rect 1429 7397 1475 7443
rect 1429 7269 1475 7315
rect 1429 7141 1475 7187
rect 9385 7397 9431 7443
rect 9385 7269 9431 7315
rect 9385 7141 9431 7187
rect 17337 7397 17383 7443
rect 18461 7397 18507 7443
rect 17337 7269 17383 7315
rect 17337 7141 17383 7187
rect 18461 7269 18507 7315
rect 18461 7141 18507 7187
rect 1429 6925 1475 6971
rect 1429 6797 1475 6843
rect 1429 6669 1475 6715
rect 5353 6925 5399 6971
rect 5353 6797 5399 6843
rect 13305 6925 13351 6971
rect 13305 6797 13351 6843
rect 5353 6669 5399 6715
rect 18461 6925 18507 6971
rect 18461 6797 18507 6843
rect 13305 6669 13351 6715
rect 18461 6669 18507 6715
rect 1429 5829 1475 5875
rect 1429 5701 1475 5747
rect 9385 5829 9431 5875
rect 1429 5573 1475 5619
rect 17337 5829 17383 5875
rect 9385 5701 9431 5747
rect 9385 5573 9431 5619
rect 18461 5829 18507 5875
rect 17337 5701 17383 5747
rect 17337 5573 17383 5619
rect 18461 5701 18507 5747
rect 18461 5573 18507 5619
rect 1429 5357 1475 5403
rect 1429 5229 1475 5275
rect 5353 5357 5399 5403
rect 5353 5229 5399 5275
rect 1429 5101 1475 5147
rect 13305 5357 13351 5403
rect 13305 5229 13351 5275
rect 5353 5101 5399 5147
rect 13305 5101 13351 5147
rect 18461 5357 18507 5403
rect 18461 5229 18507 5275
rect 18461 5101 18507 5147
rect 1429 4261 1475 4307
rect 1429 4133 1475 4179
rect 1429 4005 1475 4051
rect 9385 4261 9431 4307
rect 9385 4133 9431 4179
rect 9385 4005 9431 4051
rect 17337 4261 17383 4307
rect 18461 4261 18507 4307
rect 17337 4133 17383 4179
rect 17337 4005 17383 4051
rect 18461 4133 18507 4179
rect 18461 4005 18507 4051
rect 1429 3789 1475 3835
rect 1429 3661 1475 3707
rect 1429 3533 1475 3579
rect 5353 3789 5399 3835
rect 5353 3661 5399 3707
rect 5353 3533 5399 3579
rect 9273 3789 9319 3835
rect 9273 3661 9319 3707
rect 9273 3533 9319 3579
rect 13193 3789 13239 3835
rect 13193 3661 13239 3707
rect 13193 3533 13239 3579
rect 17113 3789 17159 3835
rect 17113 3661 17159 3707
rect 18461 3789 18507 3835
rect 18461 3661 18507 3707
rect 17113 3533 17159 3579
rect 18461 3533 18507 3579
<< polysilicon >>
rect 1824 8556 1924 8600
rect 2476 8524 2576 8568
rect 2680 8524 2780 8568
rect 2884 8524 2984 8568
rect 3346 8556 3446 8600
rect 3777 8556 3877 8600
rect 4012 8556 4112 8600
rect 4660 8556 4760 8600
rect 4908 8556 5008 8600
rect 5612 8556 5812 8600
rect 6060 8556 6260 8600
rect 6700 8556 6800 8600
rect 1824 8263 1924 8312
rect 1824 8226 1837 8263
rect 1804 8123 1837 8226
rect 1883 8123 1924 8263
rect 1804 8072 1924 8123
rect 2476 8252 2576 8400
rect 2680 8252 2780 8400
rect 2884 8367 2984 8400
rect 2884 8321 2897 8367
rect 2943 8321 2984 8367
rect 3777 8397 3877 8432
rect 2884 8308 2984 8321
rect 3346 8279 3446 8337
rect 2476 8239 3044 8252
rect 2476 8193 2489 8239
rect 2817 8193 3044 8239
rect 3346 8233 3382 8279
rect 3428 8233 3446 8279
rect 3346 8220 3446 8233
rect 2476 8180 3044 8193
rect 2476 8005 2596 8180
rect 2700 8085 2820 8098
rect 2700 8039 2737 8085
rect 2783 8039 2820 8085
rect 2700 8005 2820 8039
rect 2924 8005 3044 8180
rect 3389 8151 3509 8164
rect 3389 8105 3421 8151
rect 3467 8105 3509 8151
rect 3777 8127 3804 8397
rect 3389 8072 3509 8105
rect 1804 7864 1924 7908
rect 2476 7864 2596 7933
rect 2700 7864 2820 7933
rect 2924 7864 3044 7933
rect 3757 8069 3804 8127
rect 3850 8069 3877 8397
rect 3757 8005 3877 8069
rect 4012 8303 4112 8432
rect 4012 8163 4040 8303
rect 4086 8163 4112 8303
rect 4012 8127 4112 8163
rect 4660 8263 4760 8312
rect 4660 8217 4701 8263
rect 4747 8217 4760 8263
rect 4660 8128 4760 8217
rect 4012 8005 4132 8127
rect 4640 8072 4760 8128
rect 4908 8267 5008 8443
rect 7292 8524 7392 8568
rect 7496 8524 7596 8568
rect 7700 8524 7800 8568
rect 8162 8556 8262 8600
rect 8593 8556 8693 8600
rect 8828 8556 8928 8600
rect 9888 8556 9988 8600
rect 10620 8556 10720 8600
rect 11232 8556 11332 8600
rect 11467 8556 11567 8600
rect 11898 8556 11998 8600
rect 4908 8237 5028 8267
rect 4908 8191 4931 8237
rect 4977 8191 5028 8237
rect 5612 8278 5812 8312
rect 5612 8232 5648 8278
rect 5788 8232 5812 8278
rect 5612 8215 5812 8232
rect 6060 8278 6260 8312
rect 6060 8232 6096 8278
rect 6236 8232 6260 8278
rect 6060 8215 6260 8232
rect 6700 8263 6800 8312
rect 4908 8072 5028 8191
rect 5612 8151 5812 8164
rect 5612 8105 5640 8151
rect 5780 8105 5812 8151
rect 3389 7864 3509 7908
rect 3757 7889 3877 7933
rect 4012 7889 4132 7933
rect 5612 8072 5812 8105
rect 6060 8151 6260 8164
rect 6060 8105 6088 8151
rect 6228 8105 6260 8151
rect 6060 8072 6260 8105
rect 6700 8123 6741 8263
rect 6787 8226 6800 8263
rect 7292 8252 7392 8400
rect 7496 8252 7596 8400
rect 7700 8367 7800 8400
rect 7700 8321 7713 8367
rect 7759 8321 7800 8367
rect 8593 8397 8693 8432
rect 7700 8308 7800 8321
rect 8162 8279 8262 8337
rect 7292 8239 7860 8252
rect 6787 8123 6820 8226
rect 6700 8072 6820 8123
rect 7292 8193 7305 8239
rect 7633 8193 7860 8239
rect 8162 8233 8198 8279
rect 8244 8233 8262 8279
rect 8162 8220 8262 8233
rect 7292 8180 7860 8193
rect 4908 7956 5028 8000
rect 4640 7864 4760 7908
rect 7292 8005 7412 8180
rect 7516 8085 7636 8098
rect 7516 8039 7553 8085
rect 7599 8039 7636 8085
rect 7516 8005 7636 8039
rect 7740 8005 7860 8180
rect 8205 8151 8325 8164
rect 8205 8105 8237 8151
rect 8283 8105 8325 8151
rect 8593 8127 8620 8397
rect 8205 8072 8325 8105
rect 5612 7864 5812 7908
rect 6060 7864 6260 7908
rect 6700 7864 6820 7908
rect 7292 7864 7412 7933
rect 7516 7864 7636 7933
rect 7740 7864 7860 7933
rect 8573 8069 8620 8127
rect 8666 8069 8693 8397
rect 8573 8005 8693 8069
rect 8828 8303 8928 8432
rect 8828 8163 8856 8303
rect 8902 8163 8928 8303
rect 9888 8263 9988 8312
rect 9888 8226 9901 8263
rect 8828 8127 8928 8163
rect 8828 8005 8948 8127
rect 9868 8123 9901 8226
rect 9947 8123 9988 8263
rect 9868 8072 9988 8123
rect 10620 8263 10720 8312
rect 10620 8123 10661 8263
rect 10707 8226 10720 8263
rect 11232 8303 11332 8432
rect 10707 8123 10740 8226
rect 11232 8163 11258 8303
rect 11304 8163 11332 8303
rect 11232 8127 11332 8163
rect 10620 8072 10740 8123
rect 8205 7864 8325 7908
rect 8573 7889 8693 7933
rect 8828 7889 8948 7933
rect 11212 8005 11332 8127
rect 11467 8397 11567 8432
rect 11467 8069 11494 8397
rect 11540 8127 11567 8397
rect 12360 8524 12460 8568
rect 12564 8524 12664 8568
rect 12768 8524 12868 8568
rect 13644 8556 13744 8600
rect 14368 8556 14468 8600
rect 14603 8556 14703 8600
rect 15034 8556 15134 8600
rect 12360 8367 12460 8400
rect 11898 8279 11998 8337
rect 12360 8321 12401 8367
rect 12447 8321 12460 8367
rect 12360 8308 12460 8321
rect 11898 8233 11916 8279
rect 11962 8233 11998 8279
rect 12564 8252 12664 8400
rect 12768 8252 12868 8400
rect 11898 8220 11998 8233
rect 12300 8239 12868 8252
rect 12300 8193 12527 8239
rect 12855 8193 12868 8239
rect 13644 8263 13744 8312
rect 12300 8180 12868 8193
rect 11835 8151 11955 8164
rect 11540 8069 11587 8127
rect 11835 8105 11877 8151
rect 11923 8105 11955 8151
rect 11835 8072 11955 8105
rect 11467 8005 11587 8069
rect 9868 7864 9988 7908
rect 10620 7864 10740 7908
rect 11212 7889 11332 7933
rect 11467 7889 11587 7933
rect 12300 8005 12420 8180
rect 12524 8085 12644 8098
rect 12524 8039 12561 8085
rect 12607 8039 12644 8085
rect 12524 8005 12644 8039
rect 12748 8005 12868 8180
rect 13644 8123 13685 8263
rect 13731 8226 13744 8263
rect 14368 8303 14468 8432
rect 13731 8123 13764 8226
rect 14368 8163 14394 8303
rect 14440 8163 14468 8303
rect 14368 8127 14468 8163
rect 13644 8072 13764 8123
rect 11835 7864 11955 7908
rect 12300 7864 12420 7933
rect 12524 7864 12644 7933
rect 12748 7864 12868 7933
rect 14348 8005 14468 8127
rect 14603 8397 14703 8432
rect 14603 8069 14630 8397
rect 14676 8127 14703 8397
rect 15496 8524 15596 8568
rect 15700 8524 15800 8568
rect 15904 8524 16004 8568
rect 16496 8556 16596 8600
rect 17504 8556 17604 8600
rect 17932 8556 18132 8600
rect 15496 8367 15596 8400
rect 15034 8279 15134 8337
rect 15496 8321 15537 8367
rect 15583 8321 15596 8367
rect 15496 8308 15596 8321
rect 15034 8233 15052 8279
rect 15098 8233 15134 8279
rect 15700 8252 15800 8400
rect 15904 8252 16004 8400
rect 15034 8220 15134 8233
rect 15436 8239 16004 8252
rect 15436 8193 15663 8239
rect 15991 8193 16004 8239
rect 16496 8263 16596 8312
rect 16496 8226 16509 8263
rect 15436 8180 16004 8193
rect 14971 8151 15091 8164
rect 14676 8069 14723 8127
rect 14971 8105 15013 8151
rect 15059 8105 15091 8151
rect 14971 8072 15091 8105
rect 14603 8005 14723 8069
rect 13644 7864 13764 7908
rect 14348 7889 14468 7933
rect 14603 7889 14723 7933
rect 15436 8005 15556 8180
rect 15660 8085 15780 8098
rect 15660 8039 15697 8085
rect 15743 8039 15780 8085
rect 15660 8005 15780 8039
rect 15884 8005 16004 8180
rect 16476 8123 16509 8226
rect 16555 8123 16596 8263
rect 17504 8263 17604 8312
rect 17504 8226 17517 8263
rect 16476 8072 16596 8123
rect 17484 8123 17517 8226
rect 17563 8123 17604 8263
rect 17932 8278 18132 8312
rect 17932 8232 17968 8278
rect 18108 8232 18132 8278
rect 17932 8215 18132 8232
rect 14971 7864 15091 7908
rect 15436 7864 15556 7933
rect 15660 7864 15780 7933
rect 15884 7864 16004 7933
rect 17484 8072 17604 8123
rect 17932 8151 18132 8164
rect 17932 8105 17960 8151
rect 18100 8105 18132 8151
rect 17932 8072 18132 8105
rect 16476 7864 16596 7908
rect 17484 7864 17604 7908
rect 17932 7864 18132 7908
rect 1804 7772 1924 7816
rect 2476 7747 2596 7816
rect 2700 7747 2820 7816
rect 2924 7747 3044 7816
rect 3389 7772 3509 7816
rect 1804 7557 1924 7608
rect 1804 7454 1837 7557
rect 1824 7417 1837 7454
rect 1883 7417 1924 7557
rect 1824 7368 1924 7417
rect 2476 7500 2596 7675
rect 2700 7641 2820 7675
rect 2700 7595 2737 7641
rect 2783 7595 2820 7641
rect 2700 7582 2820 7595
rect 2924 7500 3044 7675
rect 3757 7747 3877 7791
rect 4012 7747 4132 7791
rect 4684 7772 4804 7816
rect 5052 7772 5252 7816
rect 5500 7772 5700 7816
rect 5948 7772 6148 7816
rect 6396 7772 6596 7816
rect 6844 7772 7044 7816
rect 3757 7611 3877 7675
rect 3389 7575 3509 7608
rect 3389 7529 3421 7575
rect 3467 7529 3509 7575
rect 3757 7553 3804 7611
rect 3389 7516 3509 7529
rect 2476 7487 3044 7500
rect 2476 7441 2489 7487
rect 2817 7441 3044 7487
rect 2476 7428 3044 7441
rect 3346 7447 3446 7460
rect 2476 7280 2576 7428
rect 2680 7280 2780 7428
rect 3346 7401 3382 7447
rect 3428 7401 3446 7447
rect 2884 7359 2984 7372
rect 2884 7313 2897 7359
rect 2943 7313 2984 7359
rect 3346 7343 3446 7401
rect 2884 7280 2984 7313
rect 1824 7080 1924 7124
rect 2476 7112 2576 7156
rect 2680 7112 2780 7156
rect 2884 7112 2984 7156
rect 3777 7283 3804 7553
rect 3850 7283 3877 7611
rect 3777 7248 3877 7283
rect 4012 7553 4132 7675
rect 7292 7747 7412 7816
rect 7516 7747 7636 7816
rect 7740 7747 7860 7816
rect 8205 7772 8325 7816
rect 4684 7557 4804 7608
rect 4012 7517 4112 7553
rect 4012 7377 4040 7517
rect 4086 7377 4112 7517
rect 4012 7248 4112 7377
rect 4684 7417 4725 7557
rect 4771 7454 4804 7557
rect 5052 7575 5252 7608
rect 5052 7529 5080 7575
rect 5220 7529 5252 7575
rect 5052 7516 5252 7529
rect 5500 7575 5700 7608
rect 5500 7529 5528 7575
rect 5668 7529 5700 7575
rect 5500 7516 5700 7529
rect 5948 7575 6148 7608
rect 5948 7529 5976 7575
rect 6116 7529 6148 7575
rect 5948 7516 6148 7529
rect 6396 7575 6596 7608
rect 6396 7529 6424 7575
rect 6564 7529 6596 7575
rect 6396 7516 6596 7529
rect 6844 7575 7044 7608
rect 6844 7529 6872 7575
rect 7012 7529 7044 7575
rect 6844 7516 7044 7529
rect 7292 7500 7412 7675
rect 7516 7641 7636 7675
rect 7516 7595 7553 7641
rect 7599 7595 7636 7641
rect 7516 7582 7636 7595
rect 7740 7500 7860 7675
rect 8573 7747 8693 7791
rect 8828 7747 8948 7791
rect 9644 7772 9844 7816
rect 10092 7772 10212 7816
rect 10764 7772 10884 7816
rect 11436 7772 11556 7816
rect 8573 7611 8693 7675
rect 8205 7575 8325 7608
rect 8205 7529 8237 7575
rect 8283 7529 8325 7575
rect 8573 7553 8620 7611
rect 8205 7516 8325 7529
rect 7292 7487 7860 7500
rect 4771 7417 4784 7454
rect 4684 7368 4784 7417
rect 5052 7448 5252 7465
rect 5052 7402 5088 7448
rect 5228 7402 5252 7448
rect 5052 7368 5252 7402
rect 5500 7448 5700 7465
rect 5500 7402 5536 7448
rect 5676 7402 5700 7448
rect 5500 7368 5700 7402
rect 5948 7448 6148 7465
rect 5948 7402 5984 7448
rect 6124 7402 6148 7448
rect 5948 7368 6148 7402
rect 6396 7448 6596 7465
rect 6396 7402 6432 7448
rect 6572 7402 6596 7448
rect 6396 7368 6596 7402
rect 6844 7448 7044 7465
rect 6844 7402 6880 7448
rect 7020 7402 7044 7448
rect 6844 7368 7044 7402
rect 7292 7441 7305 7487
rect 7633 7441 7860 7487
rect 7292 7428 7860 7441
rect 8162 7447 8262 7460
rect 7292 7280 7392 7428
rect 7496 7280 7596 7428
rect 8162 7401 8198 7447
rect 8244 7401 8262 7447
rect 7700 7359 7800 7372
rect 7700 7313 7713 7359
rect 7759 7313 7800 7359
rect 8162 7343 8262 7401
rect 7700 7280 7800 7313
rect 3346 7080 3446 7124
rect 3777 7080 3877 7124
rect 4012 7080 4112 7124
rect 4684 7080 4784 7124
rect 5052 7080 5252 7124
rect 5500 7080 5700 7124
rect 5948 7080 6148 7124
rect 6396 7080 6596 7124
rect 6844 7080 7044 7124
rect 7292 7112 7392 7156
rect 7496 7112 7596 7156
rect 7700 7112 7800 7156
rect 8593 7283 8620 7553
rect 8666 7283 8693 7611
rect 8593 7248 8693 7283
rect 8828 7553 8948 7675
rect 12108 7747 12228 7816
rect 12332 7747 12452 7816
rect 12556 7747 12676 7816
rect 13021 7772 13141 7816
rect 9644 7575 9844 7608
rect 8828 7517 8928 7553
rect 8828 7377 8856 7517
rect 8902 7377 8928 7517
rect 9644 7529 9672 7575
rect 9812 7529 9844 7575
rect 9644 7516 9844 7529
rect 10092 7557 10212 7608
rect 8828 7248 8928 7377
rect 9644 7448 9844 7465
rect 10092 7454 10125 7557
rect 9644 7402 9680 7448
rect 9820 7402 9844 7448
rect 9644 7368 9844 7402
rect 10112 7417 10125 7454
rect 10171 7417 10212 7557
rect 10764 7557 10884 7608
rect 10764 7454 10797 7557
rect 10112 7368 10212 7417
rect 10784 7417 10797 7454
rect 10843 7417 10884 7557
rect 11436 7557 11556 7608
rect 11436 7454 11469 7557
rect 10784 7368 10884 7417
rect 11456 7417 11469 7454
rect 11515 7417 11556 7557
rect 11456 7368 11556 7417
rect 12108 7500 12228 7675
rect 12332 7641 12452 7675
rect 12332 7595 12369 7641
rect 12415 7595 12452 7641
rect 12332 7582 12452 7595
rect 12556 7500 12676 7675
rect 13389 7747 13509 7791
rect 13644 7747 13764 7791
rect 14012 7772 14212 7816
rect 13389 7611 13509 7675
rect 13021 7575 13141 7608
rect 13021 7529 13053 7575
rect 13099 7529 13141 7575
rect 13389 7553 13436 7611
rect 13021 7516 13141 7529
rect 12108 7487 12676 7500
rect 12108 7441 12121 7487
rect 12449 7441 12676 7487
rect 12108 7428 12676 7441
rect 12978 7447 13078 7460
rect 12108 7280 12208 7428
rect 12312 7280 12412 7428
rect 12978 7401 13014 7447
rect 13060 7401 13078 7447
rect 12516 7359 12616 7372
rect 12516 7313 12529 7359
rect 12575 7313 12616 7359
rect 12978 7343 13078 7401
rect 12516 7280 12616 7313
rect 8162 7080 8262 7124
rect 8593 7080 8693 7124
rect 8828 7080 8928 7124
rect 9644 7080 9844 7124
rect 10112 7080 10212 7124
rect 10784 7080 10884 7124
rect 11456 7080 11556 7124
rect 12108 7112 12208 7156
rect 12312 7112 12412 7156
rect 12516 7112 12616 7156
rect 13409 7283 13436 7553
rect 13482 7283 13509 7611
rect 13409 7248 13509 7283
rect 13644 7553 13764 7675
rect 14460 7747 14580 7791
rect 14715 7747 14835 7791
rect 15083 7772 15203 7816
rect 14012 7575 14212 7608
rect 13644 7517 13744 7553
rect 13644 7377 13672 7517
rect 13718 7377 13744 7517
rect 14012 7529 14040 7575
rect 14180 7529 14212 7575
rect 14460 7553 14580 7675
rect 14012 7516 14212 7529
rect 14480 7517 14580 7553
rect 13644 7248 13744 7377
rect 14012 7448 14212 7465
rect 14012 7402 14048 7448
rect 14188 7402 14212 7448
rect 14012 7368 14212 7402
rect 14480 7377 14506 7517
rect 14552 7377 14580 7517
rect 14480 7248 14580 7377
rect 14715 7611 14835 7675
rect 14715 7283 14742 7611
rect 14788 7553 14835 7611
rect 15548 7747 15668 7816
rect 15772 7747 15892 7816
rect 15996 7747 16116 7816
rect 16588 7772 16708 7816
rect 15083 7575 15203 7608
rect 14788 7283 14815 7553
rect 15083 7529 15125 7575
rect 15171 7529 15203 7575
rect 15083 7516 15203 7529
rect 15548 7500 15668 7675
rect 15772 7641 15892 7675
rect 15772 7595 15809 7641
rect 15855 7595 15892 7641
rect 15772 7582 15892 7595
rect 15996 7500 16116 7675
rect 17708 7772 17828 7816
rect 15548 7487 16116 7500
rect 15146 7447 15246 7460
rect 15146 7401 15164 7447
rect 15210 7401 15246 7447
rect 15548 7441 15775 7487
rect 16103 7441 16116 7487
rect 16588 7557 16708 7608
rect 16588 7454 16621 7557
rect 15548 7428 16116 7441
rect 15146 7343 15246 7401
rect 15608 7359 15708 7372
rect 14715 7248 14815 7283
rect 15608 7313 15649 7359
rect 15695 7313 15708 7359
rect 15608 7280 15708 7313
rect 15812 7280 15912 7428
rect 16016 7280 16116 7428
rect 16608 7417 16621 7454
rect 16667 7417 16708 7557
rect 17708 7557 17828 7608
rect 16608 7368 16708 7417
rect 17708 7454 17741 7557
rect 12978 7080 13078 7124
rect 13409 7080 13509 7124
rect 13644 7080 13744 7124
rect 14012 7080 14212 7124
rect 14480 7080 14580 7124
rect 14715 7080 14815 7124
rect 15146 7080 15246 7124
rect 15608 7112 15708 7156
rect 15812 7112 15912 7156
rect 16016 7112 16116 7156
rect 17728 7417 17741 7454
rect 17787 7417 17828 7557
rect 17728 7368 17828 7417
rect 16608 7080 16708 7124
rect 17728 7080 17828 7124
rect 1692 6988 1892 7032
rect 2181 6988 2281 7032
rect 2453 6988 2553 7032
rect 2657 6988 2757 7032
rect 3316 6988 3416 7032
rect 3564 6988 3664 7032
rect 3932 6988 4132 7032
rect 4380 6988 4580 7032
rect 4828 6988 5028 7032
rect 5612 6988 5812 7032
rect 6060 6988 6260 7032
rect 6943 6988 7043 7032
rect 7536 6988 7636 7032
rect 8208 6988 8308 7032
rect 8880 6988 8980 7032
rect 9552 6988 9652 7032
rect 10224 6988 10324 7032
rect 10896 6988 10996 7032
rect 11568 6988 11668 7032
rect 12240 6988 12340 7032
rect 12668 6988 12868 7032
rect 13696 6988 13796 7032
rect 14368 6988 14468 7032
rect 15040 6988 15140 7032
rect 15712 6988 15812 7032
rect 16384 6988 16484 7032
rect 17056 6988 17156 7032
rect 17728 6988 17828 7032
rect 2453 6744 2553 6875
rect 1692 6710 1892 6744
rect 1692 6664 1728 6710
rect 1868 6664 1892 6710
rect 1692 6647 1892 6664
rect 1692 6583 1892 6596
rect 1692 6537 1720 6583
rect 1860 6537 1892 6583
rect 2181 6589 2281 6744
rect 2453 6698 2494 6744
rect 2540 6698 2553 6744
rect 2453 6641 2553 6698
rect 2181 6548 2216 6589
rect 1692 6504 1892 6537
rect 2161 6543 2216 6548
rect 2262 6543 2281 6589
rect 2161 6504 2281 6543
rect 2433 6437 2553 6641
rect 2657 6736 2757 6875
rect 2657 6690 2698 6736
rect 2744 6690 2757 6736
rect 2657 6641 2757 6690
rect 3316 6695 3416 6744
rect 3316 6649 3357 6695
rect 3403 6649 3416 6695
rect 2657 6437 2777 6641
rect 3316 6560 3416 6649
rect 3296 6504 3416 6560
rect 3564 6699 3664 6875
rect 3932 6710 4132 6744
rect 3564 6669 3684 6699
rect 3564 6623 3587 6669
rect 3633 6623 3684 6669
rect 3932 6664 3968 6710
rect 4108 6664 4132 6710
rect 3932 6647 4132 6664
rect 4380 6710 4580 6744
rect 4380 6664 4416 6710
rect 4556 6664 4580 6710
rect 4380 6647 4580 6664
rect 4828 6710 5028 6744
rect 4828 6664 4864 6710
rect 5004 6664 5028 6710
rect 4828 6647 5028 6664
rect 5612 6710 5812 6744
rect 5612 6664 5648 6710
rect 5788 6664 5812 6710
rect 5612 6647 5812 6664
rect 6060 6710 6260 6744
rect 6060 6664 6096 6710
rect 6236 6664 6260 6710
rect 6060 6647 6260 6664
rect 3564 6504 3684 6623
rect 6943 6599 7043 6744
rect 7536 6695 7636 6744
rect 7536 6658 7549 6695
rect 3932 6583 4132 6596
rect 3932 6537 3960 6583
rect 4100 6537 4132 6583
rect 3932 6504 4132 6537
rect 4380 6583 4580 6596
rect 4380 6537 4408 6583
rect 4548 6537 4580 6583
rect 4380 6504 4580 6537
rect 4828 6583 5028 6596
rect 4828 6537 4856 6583
rect 4996 6537 5028 6583
rect 4828 6504 5028 6537
rect 5612 6583 5812 6596
rect 5612 6537 5640 6583
rect 5780 6537 5812 6583
rect 1692 6296 1892 6340
rect 2161 6296 2281 6340
rect 2433 6320 2553 6365
rect 2657 6320 2777 6365
rect 3564 6388 3684 6432
rect 5612 6504 5812 6537
rect 6060 6583 6260 6596
rect 6060 6537 6088 6583
rect 6228 6537 6260 6583
rect 6060 6504 6260 6537
rect 6923 6586 7043 6599
rect 6923 6540 6936 6586
rect 6982 6540 7043 6586
rect 6923 6504 7043 6540
rect 7516 6555 7549 6658
rect 7595 6555 7636 6695
rect 8208 6695 8308 6744
rect 8208 6658 8221 6695
rect 7516 6504 7636 6555
rect 8188 6555 8221 6658
rect 8267 6555 8308 6695
rect 8880 6695 8980 6744
rect 8880 6658 8893 6695
rect 8188 6504 8308 6555
rect 8860 6555 8893 6658
rect 8939 6555 8980 6695
rect 9552 6695 9652 6744
rect 9552 6658 9565 6695
rect 8860 6504 8980 6555
rect 9532 6555 9565 6658
rect 9611 6555 9652 6695
rect 10224 6695 10324 6744
rect 10224 6658 10237 6695
rect 9532 6504 9652 6555
rect 10204 6555 10237 6658
rect 10283 6555 10324 6695
rect 10896 6695 10996 6744
rect 10896 6658 10909 6695
rect 10204 6504 10324 6555
rect 10876 6555 10909 6658
rect 10955 6555 10996 6695
rect 11568 6695 11668 6744
rect 11568 6658 11581 6695
rect 10876 6504 10996 6555
rect 11548 6555 11581 6658
rect 11627 6555 11668 6695
rect 12240 6695 12340 6744
rect 12240 6658 12253 6695
rect 11548 6504 11668 6555
rect 12220 6555 12253 6658
rect 12299 6555 12340 6695
rect 12668 6710 12868 6744
rect 12668 6664 12704 6710
rect 12844 6664 12868 6710
rect 12668 6647 12868 6664
rect 13696 6695 13796 6744
rect 13696 6658 13709 6695
rect 12220 6504 12340 6555
rect 12668 6583 12868 6596
rect 12668 6537 12696 6583
rect 12836 6537 12868 6583
rect 12668 6504 12868 6537
rect 13676 6555 13709 6658
rect 13755 6555 13796 6695
rect 14368 6695 14468 6744
rect 14368 6658 14381 6695
rect 3296 6296 3416 6340
rect 3932 6296 4132 6340
rect 4380 6296 4580 6340
rect 4828 6296 5028 6340
rect 13676 6504 13796 6555
rect 14348 6555 14381 6658
rect 14427 6555 14468 6695
rect 15040 6695 15140 6744
rect 15040 6658 15053 6695
rect 14348 6504 14468 6555
rect 15020 6555 15053 6658
rect 15099 6555 15140 6695
rect 15712 6695 15812 6744
rect 15712 6658 15725 6695
rect 15020 6504 15140 6555
rect 15692 6555 15725 6658
rect 15771 6555 15812 6695
rect 16384 6695 16484 6744
rect 16384 6658 16397 6695
rect 15692 6504 15812 6555
rect 16364 6555 16397 6658
rect 16443 6555 16484 6695
rect 17056 6695 17156 6744
rect 17056 6658 17069 6695
rect 16364 6504 16484 6555
rect 17036 6555 17069 6658
rect 17115 6555 17156 6695
rect 17728 6695 17828 6744
rect 17728 6658 17741 6695
rect 17036 6504 17156 6555
rect 17708 6555 17741 6658
rect 17787 6555 17828 6695
rect 17708 6504 17828 6555
rect 5612 6296 5812 6340
rect 6060 6296 6260 6340
rect 6923 6296 7043 6340
rect 7516 6296 7636 6340
rect 8188 6296 8308 6340
rect 8860 6296 8980 6340
rect 9532 6296 9652 6340
rect 10204 6296 10324 6340
rect 10876 6296 10996 6340
rect 11548 6296 11668 6340
rect 12220 6296 12340 6340
rect 12668 6296 12868 6340
rect 13676 6296 13796 6340
rect 14348 6296 14468 6340
rect 15020 6296 15140 6340
rect 15692 6296 15812 6340
rect 16364 6296 16484 6340
rect 17036 6296 17156 6340
rect 17708 6296 17828 6340
rect 2256 6203 2376 6248
rect 2924 6204 3044 6248
rect 3372 6204 3572 6248
rect 3820 6204 4020 6248
rect 4268 6204 4468 6248
rect 4716 6204 4916 6248
rect 5501 6204 5621 6248
rect 6252 6204 6372 6248
rect 6924 6204 7044 6248
rect 7516 6204 7636 6248
rect 8189 6204 8309 6248
rect 8860 6204 8980 6248
rect 1804 6113 1924 6157
rect 1988 6113 2108 6157
rect 9644 6204 9844 6248
rect 10316 6204 10436 6248
rect 10988 6204 11108 6248
rect 11660 6204 11780 6248
rect 12332 6204 12452 6248
rect 13004 6204 13124 6248
rect 13676 6204 13796 6248
rect 14348 6204 14468 6248
rect 15020 6204 15140 6248
rect 15692 6204 15812 6248
rect 16365 6204 16485 6248
rect 16812 6204 17012 6248
rect 1804 5996 1924 6040
rect 1988 5996 2108 6040
rect 1804 5903 1904 5996
rect 1804 5857 1825 5903
rect 1871 5857 1904 5903
rect 1804 5677 1904 5857
rect 2008 5903 2108 5996
rect 2008 5857 2049 5903
rect 2095 5857 2108 5903
rect 2256 5956 2376 6040
rect 2256 5910 2269 5956
rect 2315 5910 2376 5956
rect 2256 5883 2376 5910
rect 2924 5989 3044 6040
rect 2924 5886 2957 5989
rect 2008 5677 2108 5857
rect 2276 5800 2376 5883
rect 2944 5849 2957 5886
rect 3003 5849 3044 5989
rect 3372 6007 3572 6040
rect 3372 5961 3400 6007
rect 3540 5961 3572 6007
rect 3372 5948 3572 5961
rect 3820 6007 4020 6040
rect 3820 5961 3848 6007
rect 3988 5961 4020 6007
rect 3820 5948 4020 5961
rect 4268 6007 4468 6040
rect 4268 5961 4296 6007
rect 4436 5961 4468 6007
rect 4268 5948 4468 5961
rect 4716 6007 4916 6040
rect 4716 5961 4744 6007
rect 4884 5961 4916 6007
rect 4716 5948 4916 5961
rect 5501 6004 5621 6040
rect 5501 5958 5562 6004
rect 5608 5958 5621 6004
rect 5501 5945 5621 5958
rect 6252 5989 6372 6040
rect 2944 5800 3044 5849
rect 3372 5880 3572 5897
rect 3372 5834 3408 5880
rect 3548 5834 3572 5880
rect 3372 5800 3572 5834
rect 3820 5880 4020 5897
rect 3820 5834 3856 5880
rect 3996 5834 4020 5880
rect 3820 5800 4020 5834
rect 4268 5880 4468 5897
rect 4268 5834 4304 5880
rect 4444 5834 4468 5880
rect 4268 5800 4468 5834
rect 4716 5880 4916 5897
rect 4716 5834 4752 5880
rect 4892 5834 4916 5880
rect 4716 5800 4916 5834
rect 5501 5800 5601 5945
rect 6252 5849 6293 5989
rect 6339 5886 6372 5989
rect 6924 5989 7044 6040
rect 6339 5849 6352 5886
rect 6252 5800 6352 5849
rect 6924 5849 6965 5989
rect 7011 5886 7044 5989
rect 7516 5989 7636 6040
rect 7516 5886 7549 5989
rect 7011 5849 7024 5886
rect 6924 5800 7024 5849
rect 7536 5849 7549 5886
rect 7595 5849 7636 5989
rect 7536 5800 7636 5849
rect 8189 6004 8309 6040
rect 8189 5958 8250 6004
rect 8296 5958 8309 6004
rect 8189 5945 8309 5958
rect 8860 5989 8980 6040
rect 17787 6204 17907 6248
rect 8189 5800 8289 5945
rect 8860 5886 8893 5989
rect 8880 5849 8893 5886
rect 8939 5849 8980 5989
rect 9644 6007 9844 6040
rect 9644 5961 9672 6007
rect 9812 5961 9844 6007
rect 9644 5948 9844 5961
rect 10316 5989 10436 6040
rect 8880 5800 8980 5849
rect 1804 5512 1904 5557
rect 2008 5512 2108 5557
rect 2276 5512 2376 5557
rect 9644 5880 9844 5897
rect 10316 5886 10349 5989
rect 9644 5834 9680 5880
rect 9820 5834 9844 5880
rect 9644 5800 9844 5834
rect 10336 5849 10349 5886
rect 10395 5849 10436 5989
rect 10988 5989 11108 6040
rect 10988 5886 11021 5989
rect 10336 5800 10436 5849
rect 11008 5849 11021 5886
rect 11067 5849 11108 5989
rect 11660 5989 11780 6040
rect 11660 5886 11693 5989
rect 11008 5800 11108 5849
rect 11680 5849 11693 5886
rect 11739 5849 11780 5989
rect 12332 5989 12452 6040
rect 12332 5886 12365 5989
rect 11680 5800 11780 5849
rect 12352 5849 12365 5886
rect 12411 5849 12452 5989
rect 13004 5989 13124 6040
rect 13004 5886 13037 5989
rect 12352 5800 12452 5849
rect 13024 5849 13037 5886
rect 13083 5849 13124 5989
rect 13676 5989 13796 6040
rect 13676 5886 13709 5989
rect 13024 5800 13124 5849
rect 13696 5849 13709 5886
rect 13755 5849 13796 5989
rect 14348 5989 14468 6040
rect 14348 5886 14381 5989
rect 13696 5800 13796 5849
rect 14368 5849 14381 5886
rect 14427 5849 14468 5989
rect 15020 5989 15140 6040
rect 15020 5886 15053 5989
rect 14368 5800 14468 5849
rect 15040 5849 15053 5886
rect 15099 5849 15140 5989
rect 15692 5989 15812 6040
rect 15692 5886 15725 5989
rect 15040 5800 15140 5849
rect 15712 5849 15725 5886
rect 15771 5849 15812 5989
rect 15712 5800 15812 5849
rect 16365 6004 16485 6040
rect 16365 5958 16426 6004
rect 16472 5958 16485 6004
rect 16365 5945 16485 5958
rect 16812 6007 17012 6040
rect 16812 5961 16840 6007
rect 16980 5961 17012 6007
rect 16812 5948 17012 5961
rect 17787 6004 17907 6040
rect 17787 5958 17800 6004
rect 17846 5958 17907 6004
rect 17787 5945 17907 5958
rect 16365 5800 16465 5945
rect 16812 5880 17012 5897
rect 16812 5834 16848 5880
rect 16988 5834 17012 5880
rect 16812 5800 17012 5834
rect 17807 5800 17907 5945
rect 2944 5512 3044 5556
rect 3372 5512 3572 5556
rect 3820 5512 4020 5556
rect 4268 5512 4468 5556
rect 4716 5512 4916 5556
rect 5501 5512 5601 5556
rect 6252 5512 6352 5556
rect 6924 5512 7024 5556
rect 7536 5512 7636 5556
rect 8189 5512 8289 5556
rect 8880 5512 8980 5556
rect 9644 5512 9844 5556
rect 10336 5512 10436 5556
rect 11008 5512 11108 5556
rect 11680 5512 11780 5556
rect 12352 5512 12452 5556
rect 13024 5512 13124 5556
rect 13696 5512 13796 5556
rect 14368 5512 14468 5556
rect 15040 5512 15140 5556
rect 15712 5512 15812 5556
rect 16365 5512 16465 5556
rect 16812 5512 17012 5556
rect 17807 5512 17907 5556
rect 1692 5420 1892 5464
rect 2140 5420 2340 5464
rect 2588 5420 2788 5464
rect 3036 5420 3236 5464
rect 3484 5420 3684 5464
rect 4157 5420 4257 5464
rect 4829 5420 4929 5464
rect 5612 5420 5812 5464
rect 6285 5420 6385 5464
rect 7055 5420 7155 5464
rect 7708 5420 7808 5464
rect 8301 5420 8401 5464
rect 8992 5420 9092 5464
rect 9664 5420 9764 5464
rect 10336 5420 10436 5464
rect 11008 5420 11108 5464
rect 11680 5420 11780 5464
rect 12352 5420 12452 5464
rect 12780 5420 12980 5464
rect 13696 5420 13796 5464
rect 14368 5420 14468 5464
rect 15100 5420 15200 5464
rect 15791 5420 15891 5464
rect 16496 5420 16596 5464
rect 16731 5420 16831 5464
rect 17162 5420 17262 5464
rect 1692 5142 1892 5176
rect 1692 5096 1728 5142
rect 1868 5096 1892 5142
rect 1692 5079 1892 5096
rect 2140 5142 2340 5176
rect 2140 5096 2176 5142
rect 2316 5096 2340 5142
rect 2140 5079 2340 5096
rect 2588 5142 2788 5176
rect 2588 5096 2624 5142
rect 2764 5096 2788 5142
rect 2588 5079 2788 5096
rect 3036 5142 3236 5176
rect 3036 5096 3072 5142
rect 3212 5096 3236 5142
rect 3036 5079 3236 5096
rect 3484 5142 3684 5176
rect 3484 5096 3520 5142
rect 3660 5096 3684 5142
rect 3484 5079 3684 5096
rect 4157 5031 4257 5176
rect 4829 5031 4929 5176
rect 5612 5142 5812 5176
rect 5612 5096 5648 5142
rect 5788 5096 5812 5142
rect 5612 5079 5812 5096
rect 6285 5031 6385 5176
rect 7055 5031 7155 5176
rect 1692 5015 1892 5028
rect 1692 4969 1720 5015
rect 1860 4969 1892 5015
rect 1692 4936 1892 4969
rect 2140 5015 2340 5028
rect 2140 4969 2168 5015
rect 2308 4969 2340 5015
rect 2140 4936 2340 4969
rect 2588 5015 2788 5028
rect 2588 4969 2616 5015
rect 2756 4969 2788 5015
rect 2588 4936 2788 4969
rect 3036 5015 3236 5028
rect 3036 4969 3064 5015
rect 3204 4969 3236 5015
rect 3036 4936 3236 4969
rect 3484 5015 3684 5028
rect 3484 4969 3512 5015
rect 3652 4969 3684 5015
rect 3484 4936 3684 4969
rect 4157 5018 4277 5031
rect 4157 4972 4218 5018
rect 4264 4972 4277 5018
rect 4157 4936 4277 4972
rect 4829 5018 4949 5031
rect 4829 4972 4890 5018
rect 4936 4972 4949 5018
rect 4829 4936 4949 4972
rect 5612 5015 5812 5028
rect 5612 4969 5640 5015
rect 5780 4969 5812 5015
rect 5612 4936 5812 4969
rect 6285 5018 6405 5031
rect 6285 4972 6346 5018
rect 6392 4972 6405 5018
rect 6285 4936 6405 4972
rect 7035 5018 7155 5031
rect 7035 4972 7048 5018
rect 7094 4972 7155 5018
rect 7035 4936 7155 4972
rect 7708 5127 7808 5176
rect 7708 4987 7749 5127
rect 7795 5090 7808 5127
rect 7795 4987 7828 5090
rect 7708 4936 7828 4987
rect 8301 5031 8401 5176
rect 8992 5127 9092 5176
rect 8992 5090 9005 5127
rect 8301 5018 8421 5031
rect 8301 4972 8362 5018
rect 8408 4972 8421 5018
rect 8301 4936 8421 4972
rect 8972 4987 9005 5090
rect 9051 4987 9092 5127
rect 9664 5127 9764 5176
rect 9664 5090 9677 5127
rect 8972 4936 9092 4987
rect 9644 4987 9677 5090
rect 9723 4987 9764 5127
rect 10336 5127 10436 5176
rect 10336 5090 10349 5127
rect 9644 4936 9764 4987
rect 10316 4987 10349 5090
rect 10395 4987 10436 5127
rect 11008 5127 11108 5176
rect 11008 5090 11021 5127
rect 10316 4936 10436 4987
rect 10988 4987 11021 5090
rect 11067 4987 11108 5127
rect 11680 5127 11780 5176
rect 11680 5090 11693 5127
rect 10988 4936 11108 4987
rect 11660 4987 11693 5090
rect 11739 4987 11780 5127
rect 12352 5127 12452 5176
rect 12352 5090 12365 5127
rect 11660 4936 11780 4987
rect 12332 4987 12365 5090
rect 12411 4987 12452 5127
rect 12780 5142 12980 5176
rect 12780 5096 12816 5142
rect 12956 5096 12980 5142
rect 12780 5079 12980 5096
rect 13696 5127 13796 5176
rect 13696 5090 13709 5127
rect 12332 4936 12452 4987
rect 12780 5015 12980 5028
rect 12780 4969 12808 5015
rect 12948 4969 12980 5015
rect 12780 4936 12980 4969
rect 13676 4987 13709 5090
rect 13755 4987 13796 5127
rect 14368 5127 14468 5176
rect 14368 5090 14381 5127
rect 1692 4728 1892 4772
rect 2140 4728 2340 4772
rect 2588 4728 2788 4772
rect 3036 4728 3236 4772
rect 3484 4728 3684 4772
rect 4157 4728 4277 4772
rect 4829 4728 4949 4772
rect 13676 4936 13796 4987
rect 14348 4987 14381 5090
rect 14427 4987 14468 5127
rect 14348 4936 14468 4987
rect 15100 5127 15200 5176
rect 15100 4987 15141 5127
rect 15187 5090 15200 5127
rect 15187 4987 15220 5090
rect 15791 5031 15891 5176
rect 15100 4936 15220 4987
rect 15771 5018 15891 5031
rect 15771 4972 15784 5018
rect 15830 4972 15891 5018
rect 16496 5167 16596 5296
rect 16496 5027 16522 5167
rect 16568 5027 16596 5167
rect 16496 4991 16596 5027
rect 15771 4936 15891 4972
rect 5612 4728 5812 4772
rect 6285 4728 6405 4772
rect 7035 4728 7155 4772
rect 7708 4728 7828 4772
rect 8301 4728 8421 4772
rect 8972 4728 9092 4772
rect 9644 4728 9764 4772
rect 10316 4728 10436 4772
rect 10988 4728 11108 4772
rect 11660 4728 11780 4772
rect 12332 4728 12452 4772
rect 12780 4728 12980 4772
rect 16476 4869 16596 4991
rect 16731 5261 16831 5296
rect 16731 4933 16758 5261
rect 16804 4991 16831 5261
rect 17624 5388 17724 5432
rect 17828 5388 17928 5432
rect 18032 5388 18132 5432
rect 17624 5231 17724 5264
rect 17162 5143 17262 5201
rect 17624 5185 17665 5231
rect 17711 5185 17724 5231
rect 17624 5172 17724 5185
rect 17162 5097 17180 5143
rect 17226 5097 17262 5143
rect 17828 5116 17928 5264
rect 18032 5116 18132 5264
rect 17162 5084 17262 5097
rect 17564 5103 18132 5116
rect 17564 5057 17791 5103
rect 18119 5057 18132 5103
rect 17564 5044 18132 5057
rect 17099 5015 17219 5028
rect 16804 4933 16851 4991
rect 17099 4969 17141 5015
rect 17187 4969 17219 5015
rect 17099 4936 17219 4969
rect 16731 4869 16851 4933
rect 13676 4728 13796 4772
rect 14348 4728 14468 4772
rect 15100 4728 15220 4772
rect 15771 4728 15891 4772
rect 16476 4753 16596 4797
rect 16731 4753 16851 4797
rect 17564 4869 17684 5044
rect 17788 4949 17908 4962
rect 17788 4903 17825 4949
rect 17871 4903 17908 4949
rect 17788 4869 17908 4903
rect 18012 4869 18132 5044
rect 17099 4728 17219 4772
rect 17564 4728 17684 4797
rect 17788 4728 17908 4797
rect 18012 4728 18132 4797
rect 1692 4636 1892 4680
rect 2140 4636 2340 4680
rect 2700 4611 2820 4680
rect 2924 4611 3044 4680
rect 3148 4611 3268 4680
rect 3613 4636 3733 4680
rect 1692 4439 1892 4472
rect 1692 4393 1720 4439
rect 1860 4393 1892 4439
rect 1692 4380 1892 4393
rect 2140 4439 2340 4472
rect 2140 4393 2168 4439
rect 2308 4393 2340 4439
rect 2140 4380 2340 4393
rect 2700 4364 2820 4539
rect 2924 4505 3044 4539
rect 2924 4459 2961 4505
rect 3007 4459 3044 4505
rect 2924 4446 3044 4459
rect 3148 4364 3268 4539
rect 3981 4611 4101 4655
rect 4236 4611 4356 4655
rect 4604 4636 4804 4680
rect 5165 4636 5285 4680
rect 5837 4636 5957 4680
rect 6509 4636 6629 4680
rect 3981 4475 4101 4539
rect 3613 4439 3733 4472
rect 3613 4393 3645 4439
rect 3691 4393 3733 4439
rect 3981 4417 4028 4475
rect 3613 4380 3733 4393
rect 2700 4351 3268 4364
rect 1692 4312 1892 4329
rect 1692 4266 1728 4312
rect 1868 4266 1892 4312
rect 1692 4232 1892 4266
rect 2140 4312 2340 4329
rect 2140 4266 2176 4312
rect 2316 4266 2340 4312
rect 2140 4232 2340 4266
rect 2700 4305 2713 4351
rect 3041 4305 3268 4351
rect 2700 4292 3268 4305
rect 3570 4311 3670 4324
rect 2700 4144 2800 4292
rect 2904 4144 3004 4292
rect 3570 4265 3606 4311
rect 3652 4265 3670 4311
rect 3108 4223 3208 4236
rect 3108 4177 3121 4223
rect 3167 4177 3208 4223
rect 3570 4207 3670 4265
rect 3108 4144 3208 4177
rect 1692 3944 1892 3988
rect 2140 3944 2340 3988
rect 2700 3976 2800 4020
rect 2904 3976 3004 4020
rect 3108 3976 3208 4020
rect 4001 4147 4028 4417
rect 4074 4147 4101 4475
rect 4001 4112 4101 4147
rect 4236 4417 4356 4539
rect 7180 4611 7300 4655
rect 7435 4611 7555 4655
rect 7803 4636 7923 4680
rect 4604 4439 4804 4472
rect 4236 4381 4336 4417
rect 4236 4241 4264 4381
rect 4310 4241 4336 4381
rect 4604 4393 4632 4439
rect 4772 4393 4804 4439
rect 4604 4380 4804 4393
rect 5165 4436 5285 4472
rect 5165 4390 5226 4436
rect 5272 4390 5285 4436
rect 5165 4377 5285 4390
rect 5837 4436 5957 4472
rect 5837 4390 5898 4436
rect 5944 4390 5957 4436
rect 5837 4377 5957 4390
rect 6509 4436 6629 4472
rect 6509 4390 6570 4436
rect 6616 4390 6629 4436
rect 7180 4417 7300 4539
rect 6509 4377 6629 4390
rect 7200 4381 7300 4417
rect 4236 4112 4336 4241
rect 4604 4312 4804 4329
rect 4604 4266 4640 4312
rect 4780 4266 4804 4312
rect 4604 4232 4804 4266
rect 5165 4232 5265 4377
rect 5837 4232 5937 4377
rect 6509 4232 6609 4377
rect 7200 4241 7226 4381
rect 7272 4241 7300 4381
rect 7200 4112 7300 4241
rect 7435 4475 7555 4539
rect 7435 4147 7462 4475
rect 7508 4417 7555 4475
rect 8268 4611 8388 4680
rect 8492 4611 8612 4680
rect 8716 4611 8836 4680
rect 9644 4636 9844 4680
rect 10093 4636 10213 4680
rect 10844 4636 10964 4680
rect 11516 4636 11636 4680
rect 7803 4439 7923 4472
rect 7508 4147 7535 4417
rect 7803 4393 7845 4439
rect 7891 4393 7923 4439
rect 7803 4380 7923 4393
rect 8268 4364 8388 4539
rect 8492 4505 8612 4539
rect 8492 4459 8529 4505
rect 8575 4459 8612 4505
rect 8492 4446 8612 4459
rect 8716 4364 8836 4539
rect 12108 4611 12228 4655
rect 12363 4611 12483 4655
rect 12731 4636 12851 4680
rect 9644 4439 9844 4472
rect 9644 4393 9672 4439
rect 9812 4393 9844 4439
rect 9644 4380 9844 4393
rect 10093 4436 10213 4472
rect 10093 4390 10154 4436
rect 10200 4390 10213 4436
rect 8268 4351 8836 4364
rect 7866 4311 7966 4324
rect 7866 4265 7884 4311
rect 7930 4265 7966 4311
rect 8268 4305 8495 4351
rect 8823 4305 8836 4351
rect 10093 4377 10213 4390
rect 10844 4421 10964 4472
rect 8268 4292 8836 4305
rect 7866 4207 7966 4265
rect 8328 4223 8428 4236
rect 7435 4112 7535 4147
rect 8328 4177 8369 4223
rect 8415 4177 8428 4223
rect 8328 4144 8428 4177
rect 8532 4144 8632 4292
rect 8736 4144 8836 4292
rect 9644 4312 9844 4329
rect 9644 4266 9680 4312
rect 9820 4266 9844 4312
rect 9644 4232 9844 4266
rect 10093 4232 10193 4377
rect 10844 4281 10885 4421
rect 10931 4318 10964 4421
rect 11516 4421 11636 4472
rect 10931 4281 10944 4318
rect 10844 4232 10944 4281
rect 11516 4281 11557 4421
rect 11603 4318 11636 4421
rect 12108 4417 12228 4539
rect 12128 4381 12228 4417
rect 11603 4281 11616 4318
rect 11516 4232 11616 4281
rect 12128 4241 12154 4381
rect 12200 4241 12228 4381
rect 3570 3944 3670 3988
rect 4001 3944 4101 3988
rect 4236 3944 4336 3988
rect 4604 3944 4804 3988
rect 5165 3944 5265 3988
rect 5837 3944 5937 3988
rect 6509 3944 6609 3988
rect 7200 3944 7300 3988
rect 7435 3944 7535 3988
rect 7866 3944 7966 3988
rect 8328 3976 8428 4020
rect 8532 3976 8632 4020
rect 8736 3976 8836 4020
rect 12128 4112 12228 4241
rect 12363 4475 12483 4539
rect 12363 4147 12390 4475
rect 12436 4417 12483 4475
rect 13196 4611 13316 4680
rect 13420 4611 13540 4680
rect 13644 4611 13764 4680
rect 14237 4636 14357 4680
rect 14908 4636 15028 4680
rect 15580 4636 15700 4680
rect 16252 4636 16372 4680
rect 16700 4636 16900 4680
rect 12731 4439 12851 4472
rect 12436 4147 12463 4417
rect 12731 4393 12773 4439
rect 12819 4393 12851 4439
rect 12731 4380 12851 4393
rect 13196 4364 13316 4539
rect 13420 4505 13540 4539
rect 13420 4459 13457 4505
rect 13503 4459 13540 4505
rect 13420 4446 13540 4459
rect 13644 4364 13764 4539
rect 17708 4636 17828 4680
rect 13196 4351 13764 4364
rect 12794 4311 12894 4324
rect 12794 4265 12812 4311
rect 12858 4265 12894 4311
rect 13196 4305 13423 4351
rect 13751 4305 13764 4351
rect 13196 4292 13764 4305
rect 12794 4207 12894 4265
rect 13256 4223 13356 4236
rect 12363 4112 12463 4147
rect 13256 4177 13297 4223
rect 13343 4177 13356 4223
rect 13256 4144 13356 4177
rect 13460 4144 13560 4292
rect 13664 4144 13764 4292
rect 14237 4436 14357 4472
rect 14237 4390 14298 4436
rect 14344 4390 14357 4436
rect 14237 4377 14357 4390
rect 14908 4421 15028 4472
rect 14237 4232 14337 4377
rect 14908 4318 14941 4421
rect 14928 4281 14941 4318
rect 14987 4281 15028 4421
rect 15580 4421 15700 4472
rect 15580 4318 15613 4421
rect 14928 4232 15028 4281
rect 15600 4281 15613 4318
rect 15659 4281 15700 4421
rect 16252 4421 16372 4472
rect 16252 4318 16285 4421
rect 15600 4232 15700 4281
rect 16272 4281 16285 4318
rect 16331 4281 16372 4421
rect 16700 4439 16900 4472
rect 16700 4393 16728 4439
rect 16868 4393 16900 4439
rect 16700 4380 16900 4393
rect 17708 4421 17828 4472
rect 16272 4232 16372 4281
rect 16700 4312 16900 4329
rect 16700 4266 16736 4312
rect 16876 4266 16900 4312
rect 16700 4232 16900 4266
rect 17708 4318 17741 4421
rect 9644 3944 9844 3988
rect 10093 3944 10193 3988
rect 10844 3944 10944 3988
rect 11516 3944 11616 3988
rect 12128 3944 12228 3988
rect 12363 3944 12463 3988
rect 12794 3944 12894 3988
rect 13256 3976 13356 4020
rect 13460 3976 13560 4020
rect 13664 3976 13764 4020
rect 17728 4281 17741 4318
rect 17787 4281 17828 4421
rect 17728 4232 17828 4281
rect 14237 3944 14337 3988
rect 14928 3944 15028 3988
rect 15600 3944 15700 3988
rect 16272 3944 16372 3988
rect 16700 3944 16900 3988
rect 17728 3944 17828 3988
rect 2029 3852 2129 3896
rect 2720 3852 2820 3896
rect 2955 3852 3055 3896
rect 3386 3852 3486 3896
rect 2029 3463 2129 3608
rect 2720 3599 2820 3728
rect 2029 3450 2149 3463
rect 2029 3404 2090 3450
rect 2136 3404 2149 3450
rect 2720 3459 2746 3599
rect 2792 3459 2820 3599
rect 2720 3423 2820 3459
rect 2029 3368 2149 3404
rect 2700 3301 2820 3423
rect 2955 3693 3055 3728
rect 2955 3365 2982 3693
rect 3028 3423 3055 3693
rect 3848 3820 3948 3864
rect 4052 3820 4152 3864
rect 4256 3820 4356 3864
rect 4829 3852 4929 3896
rect 5949 3852 6049 3896
rect 6621 3852 6721 3896
rect 7312 3852 7412 3896
rect 7547 3852 7647 3896
rect 7978 3852 8078 3896
rect 3848 3663 3948 3696
rect 3386 3575 3486 3633
rect 3848 3617 3889 3663
rect 3935 3617 3948 3663
rect 3848 3604 3948 3617
rect 3386 3529 3404 3575
rect 3450 3529 3486 3575
rect 4052 3548 4152 3696
rect 4256 3548 4356 3696
rect 3386 3516 3486 3529
rect 3788 3535 4356 3548
rect 3788 3489 4015 3535
rect 4343 3489 4356 3535
rect 3788 3476 4356 3489
rect 3323 3447 3443 3460
rect 3028 3365 3075 3423
rect 3323 3401 3365 3447
rect 3411 3401 3443 3447
rect 3323 3368 3443 3401
rect 2955 3301 3075 3365
rect 2029 3160 2149 3204
rect 2700 3185 2820 3229
rect 2955 3185 3075 3229
rect 3788 3301 3908 3476
rect 4012 3381 4132 3394
rect 4012 3335 4049 3381
rect 4095 3335 4132 3381
rect 4012 3301 4132 3335
rect 4236 3301 4356 3476
rect 4829 3463 4929 3608
rect 5949 3463 6049 3608
rect 6621 3463 6721 3608
rect 7312 3599 7412 3728
rect 4829 3450 4949 3463
rect 4829 3404 4890 3450
rect 4936 3404 4949 3450
rect 4829 3368 4949 3404
rect 5949 3450 6069 3463
rect 5949 3404 6010 3450
rect 6056 3404 6069 3450
rect 3323 3160 3443 3204
rect 3788 3160 3908 3229
rect 4012 3160 4132 3229
rect 4236 3160 4356 3229
rect 5949 3368 6069 3404
rect 6621 3450 6741 3463
rect 6621 3404 6682 3450
rect 6728 3404 6741 3450
rect 7312 3459 7338 3599
rect 7384 3459 7412 3599
rect 7312 3423 7412 3459
rect 6621 3368 6741 3404
rect 4829 3160 4949 3204
rect 7292 3301 7412 3423
rect 7547 3693 7647 3728
rect 7547 3365 7574 3693
rect 7620 3423 7647 3693
rect 8440 3820 8540 3864
rect 8644 3820 8744 3864
rect 8848 3820 8948 3864
rect 9869 3852 9969 3896
rect 10541 3852 10641 3896
rect 11232 3852 11332 3896
rect 11467 3852 11567 3896
rect 11898 3852 11998 3896
rect 8440 3663 8540 3696
rect 7978 3575 8078 3633
rect 8440 3617 8481 3663
rect 8527 3617 8540 3663
rect 8440 3604 8540 3617
rect 7978 3529 7996 3575
rect 8042 3529 8078 3575
rect 8644 3548 8744 3696
rect 8848 3548 8948 3696
rect 7978 3516 8078 3529
rect 8380 3535 8948 3548
rect 8380 3489 8607 3535
rect 8935 3489 8948 3535
rect 8380 3476 8948 3489
rect 7915 3447 8035 3460
rect 7620 3365 7667 3423
rect 7915 3401 7957 3447
rect 8003 3401 8035 3447
rect 7915 3368 8035 3401
rect 7547 3301 7667 3365
rect 5949 3160 6069 3204
rect 6621 3160 6741 3204
rect 7292 3185 7412 3229
rect 7547 3185 7667 3229
rect 8380 3301 8500 3476
rect 8604 3381 8724 3394
rect 8604 3335 8641 3381
rect 8687 3335 8724 3381
rect 8604 3301 8724 3335
rect 8828 3301 8948 3476
rect 9869 3463 9969 3608
rect 10541 3463 10641 3608
rect 11232 3599 11332 3728
rect 9869 3450 9989 3463
rect 9869 3404 9930 3450
rect 9976 3404 9989 3450
rect 9869 3368 9989 3404
rect 10541 3450 10661 3463
rect 10541 3404 10602 3450
rect 10648 3404 10661 3450
rect 11232 3459 11258 3599
rect 11304 3459 11332 3599
rect 11232 3423 11332 3459
rect 10541 3368 10661 3404
rect 7915 3160 8035 3204
rect 8380 3160 8500 3229
rect 8604 3160 8724 3229
rect 8828 3160 8948 3229
rect 11212 3301 11332 3423
rect 11467 3693 11567 3728
rect 11467 3365 11494 3693
rect 11540 3423 11567 3693
rect 12360 3820 12460 3864
rect 12564 3820 12664 3864
rect 12768 3820 12868 3864
rect 13644 3852 13744 3896
rect 14237 3852 14337 3896
rect 14684 3852 14884 3896
rect 15152 3852 15252 3896
rect 15387 3852 15487 3896
rect 15818 3852 15918 3896
rect 12360 3663 12460 3696
rect 11898 3575 11998 3633
rect 12360 3617 12401 3663
rect 12447 3617 12460 3663
rect 12360 3604 12460 3617
rect 11898 3529 11916 3575
rect 11962 3529 11998 3575
rect 12564 3548 12664 3696
rect 12768 3548 12868 3696
rect 11898 3516 11998 3529
rect 12300 3535 12868 3548
rect 12300 3489 12527 3535
rect 12855 3489 12868 3535
rect 13644 3559 13744 3608
rect 12300 3476 12868 3489
rect 11835 3447 11955 3460
rect 11540 3365 11587 3423
rect 11835 3401 11877 3447
rect 11923 3401 11955 3447
rect 11835 3368 11955 3401
rect 11467 3301 11587 3365
rect 9869 3160 9989 3204
rect 10541 3160 10661 3204
rect 11212 3185 11332 3229
rect 11467 3185 11587 3229
rect 12300 3301 12420 3476
rect 12524 3381 12644 3394
rect 12524 3335 12561 3381
rect 12607 3335 12644 3381
rect 12524 3301 12644 3335
rect 12748 3301 12868 3476
rect 13644 3419 13685 3559
rect 13731 3522 13744 3559
rect 13731 3419 13764 3522
rect 13644 3368 13764 3419
rect 14237 3463 14337 3608
rect 14684 3574 14884 3608
rect 14684 3528 14720 3574
rect 14860 3528 14884 3574
rect 14684 3511 14884 3528
rect 15152 3599 15252 3728
rect 14237 3450 14357 3463
rect 14237 3404 14298 3450
rect 14344 3404 14357 3450
rect 14237 3368 14357 3404
rect 14684 3447 14884 3460
rect 14684 3401 14712 3447
rect 14852 3401 14884 3447
rect 15152 3459 15178 3599
rect 15224 3459 15252 3599
rect 15152 3423 15252 3459
rect 14684 3368 14884 3401
rect 11835 3160 11955 3204
rect 12300 3160 12420 3229
rect 12524 3160 12644 3229
rect 12748 3160 12868 3229
rect 15132 3301 15252 3423
rect 15387 3693 15487 3728
rect 15387 3365 15414 3693
rect 15460 3423 15487 3693
rect 16280 3820 16380 3864
rect 16484 3820 16584 3864
rect 16688 3820 16788 3864
rect 17583 3852 17683 3896
rect 17932 3852 18132 3896
rect 16280 3663 16380 3696
rect 15818 3575 15918 3633
rect 16280 3617 16321 3663
rect 16367 3617 16380 3663
rect 16280 3604 16380 3617
rect 15818 3529 15836 3575
rect 15882 3529 15918 3575
rect 16484 3548 16584 3696
rect 16688 3548 16788 3696
rect 15818 3516 15918 3529
rect 16220 3535 16788 3548
rect 16220 3489 16447 3535
rect 16775 3489 16788 3535
rect 16220 3476 16788 3489
rect 15755 3447 15875 3460
rect 15460 3365 15507 3423
rect 15755 3401 15797 3447
rect 15843 3401 15875 3447
rect 15755 3368 15875 3401
rect 15387 3301 15507 3365
rect 13644 3160 13764 3204
rect 14237 3160 14357 3204
rect 14684 3160 14884 3204
rect 15132 3185 15252 3229
rect 15387 3185 15507 3229
rect 16220 3301 16340 3476
rect 16444 3381 16564 3394
rect 16444 3335 16481 3381
rect 16527 3335 16564 3381
rect 16444 3301 16564 3335
rect 16668 3301 16788 3476
rect 17583 3463 17683 3608
rect 17932 3574 18132 3608
rect 17932 3528 17968 3574
rect 18108 3528 18132 3574
rect 17932 3511 18132 3528
rect 17563 3450 17683 3463
rect 17563 3404 17576 3450
rect 17622 3404 17683 3450
rect 17563 3368 17683 3404
rect 17932 3447 18132 3460
rect 17932 3401 17960 3447
rect 18100 3401 18132 3447
rect 17932 3368 18132 3401
rect 15755 3160 15875 3204
rect 16220 3160 16340 3229
rect 16444 3160 16564 3229
rect 16668 3160 16788 3229
rect 17563 3160 17683 3204
rect 17932 3160 18132 3204
<< polycontact >>
rect 1837 8123 1883 8263
rect 2897 8321 2943 8367
rect 2489 8193 2817 8239
rect 3382 8233 3428 8279
rect 2737 8039 2783 8085
rect 3421 8105 3467 8151
rect 3804 8069 3850 8397
rect 4040 8163 4086 8303
rect 4701 8217 4747 8263
rect 4931 8191 4977 8237
rect 5648 8232 5788 8278
rect 6096 8232 6236 8278
rect 5640 8105 5780 8151
rect 6088 8105 6228 8151
rect 6741 8123 6787 8263
rect 7713 8321 7759 8367
rect 7305 8193 7633 8239
rect 8198 8233 8244 8279
rect 7553 8039 7599 8085
rect 8237 8105 8283 8151
rect 8620 8069 8666 8397
rect 8856 8163 8902 8303
rect 9901 8123 9947 8263
rect 10661 8123 10707 8263
rect 11258 8163 11304 8303
rect 11494 8069 11540 8397
rect 12401 8321 12447 8367
rect 11916 8233 11962 8279
rect 12527 8193 12855 8239
rect 11877 8105 11923 8151
rect 12561 8039 12607 8085
rect 13685 8123 13731 8263
rect 14394 8163 14440 8303
rect 14630 8069 14676 8397
rect 15537 8321 15583 8367
rect 15052 8233 15098 8279
rect 15663 8193 15991 8239
rect 15013 8105 15059 8151
rect 15697 8039 15743 8085
rect 16509 8123 16555 8263
rect 17517 8123 17563 8263
rect 17968 8232 18108 8278
rect 17960 8105 18100 8151
rect 1837 7417 1883 7557
rect 2737 7595 2783 7641
rect 3421 7529 3467 7575
rect 2489 7441 2817 7487
rect 3382 7401 3428 7447
rect 2897 7313 2943 7359
rect 3804 7283 3850 7611
rect 4040 7377 4086 7517
rect 4725 7417 4771 7557
rect 5080 7529 5220 7575
rect 5528 7529 5668 7575
rect 5976 7529 6116 7575
rect 6424 7529 6564 7575
rect 6872 7529 7012 7575
rect 7553 7595 7599 7641
rect 8237 7529 8283 7575
rect 5088 7402 5228 7448
rect 5536 7402 5676 7448
rect 5984 7402 6124 7448
rect 6432 7402 6572 7448
rect 6880 7402 7020 7448
rect 7305 7441 7633 7487
rect 8198 7401 8244 7447
rect 7713 7313 7759 7359
rect 8620 7283 8666 7611
rect 8856 7377 8902 7517
rect 9672 7529 9812 7575
rect 9680 7402 9820 7448
rect 10125 7417 10171 7557
rect 10797 7417 10843 7557
rect 11469 7417 11515 7557
rect 12369 7595 12415 7641
rect 13053 7529 13099 7575
rect 12121 7441 12449 7487
rect 13014 7401 13060 7447
rect 12529 7313 12575 7359
rect 13436 7283 13482 7611
rect 13672 7377 13718 7517
rect 14040 7529 14180 7575
rect 14048 7402 14188 7448
rect 14506 7377 14552 7517
rect 14742 7283 14788 7611
rect 15125 7529 15171 7575
rect 15809 7595 15855 7641
rect 15164 7401 15210 7447
rect 15775 7441 16103 7487
rect 15649 7313 15695 7359
rect 16621 7417 16667 7557
rect 17741 7417 17787 7557
rect 1728 6664 1868 6710
rect 1720 6537 1860 6583
rect 2494 6698 2540 6744
rect 2216 6543 2262 6589
rect 2698 6690 2744 6736
rect 3357 6649 3403 6695
rect 3587 6623 3633 6669
rect 3968 6664 4108 6710
rect 4416 6664 4556 6710
rect 4864 6664 5004 6710
rect 5648 6664 5788 6710
rect 6096 6664 6236 6710
rect 3960 6537 4100 6583
rect 4408 6537 4548 6583
rect 4856 6537 4996 6583
rect 5640 6537 5780 6583
rect 6088 6537 6228 6583
rect 6936 6540 6982 6586
rect 7549 6555 7595 6695
rect 8221 6555 8267 6695
rect 8893 6555 8939 6695
rect 9565 6555 9611 6695
rect 10237 6555 10283 6695
rect 10909 6555 10955 6695
rect 11581 6555 11627 6695
rect 12253 6555 12299 6695
rect 12704 6664 12844 6710
rect 12696 6537 12836 6583
rect 13709 6555 13755 6695
rect 14381 6555 14427 6695
rect 15053 6555 15099 6695
rect 15725 6555 15771 6695
rect 16397 6555 16443 6695
rect 17069 6555 17115 6695
rect 17741 6555 17787 6695
rect 1825 5857 1871 5903
rect 2049 5857 2095 5903
rect 2269 5910 2315 5956
rect 2957 5849 3003 5989
rect 3400 5961 3540 6007
rect 3848 5961 3988 6007
rect 4296 5961 4436 6007
rect 4744 5961 4884 6007
rect 5562 5958 5608 6004
rect 3408 5834 3548 5880
rect 3856 5834 3996 5880
rect 4304 5834 4444 5880
rect 4752 5834 4892 5880
rect 6293 5849 6339 5989
rect 6965 5849 7011 5989
rect 7549 5849 7595 5989
rect 8250 5958 8296 6004
rect 8893 5849 8939 5989
rect 9672 5961 9812 6007
rect 9680 5834 9820 5880
rect 10349 5849 10395 5989
rect 11021 5849 11067 5989
rect 11693 5849 11739 5989
rect 12365 5849 12411 5989
rect 13037 5849 13083 5989
rect 13709 5849 13755 5989
rect 14381 5849 14427 5989
rect 15053 5849 15099 5989
rect 15725 5849 15771 5989
rect 16426 5958 16472 6004
rect 16840 5961 16980 6007
rect 17800 5958 17846 6004
rect 16848 5834 16988 5880
rect 1728 5096 1868 5142
rect 2176 5096 2316 5142
rect 2624 5096 2764 5142
rect 3072 5096 3212 5142
rect 3520 5096 3660 5142
rect 5648 5096 5788 5142
rect 1720 4969 1860 5015
rect 2168 4969 2308 5015
rect 2616 4969 2756 5015
rect 3064 4969 3204 5015
rect 3512 4969 3652 5015
rect 4218 4972 4264 5018
rect 4890 4972 4936 5018
rect 5640 4969 5780 5015
rect 6346 4972 6392 5018
rect 7048 4972 7094 5018
rect 7749 4987 7795 5127
rect 8362 4972 8408 5018
rect 9005 4987 9051 5127
rect 9677 4987 9723 5127
rect 10349 4987 10395 5127
rect 11021 4987 11067 5127
rect 11693 4987 11739 5127
rect 12365 4987 12411 5127
rect 12816 5096 12956 5142
rect 12808 4969 12948 5015
rect 13709 4987 13755 5127
rect 14381 4987 14427 5127
rect 15141 4987 15187 5127
rect 15784 4972 15830 5018
rect 16522 5027 16568 5167
rect 16758 4933 16804 5261
rect 17665 5185 17711 5231
rect 17180 5097 17226 5143
rect 17791 5057 18119 5103
rect 17141 4969 17187 5015
rect 17825 4903 17871 4949
rect 1720 4393 1860 4439
rect 2168 4393 2308 4439
rect 2961 4459 3007 4505
rect 3645 4393 3691 4439
rect 1728 4266 1868 4312
rect 2176 4266 2316 4312
rect 2713 4305 3041 4351
rect 3606 4265 3652 4311
rect 3121 4177 3167 4223
rect 4028 4147 4074 4475
rect 4264 4241 4310 4381
rect 4632 4393 4772 4439
rect 5226 4390 5272 4436
rect 5898 4390 5944 4436
rect 6570 4390 6616 4436
rect 4640 4266 4780 4312
rect 7226 4241 7272 4381
rect 7462 4147 7508 4475
rect 7845 4393 7891 4439
rect 8529 4459 8575 4505
rect 9672 4393 9812 4439
rect 10154 4390 10200 4436
rect 7884 4265 7930 4311
rect 8495 4305 8823 4351
rect 8369 4177 8415 4223
rect 9680 4266 9820 4312
rect 10885 4281 10931 4421
rect 11557 4281 11603 4421
rect 12154 4241 12200 4381
rect 12390 4147 12436 4475
rect 12773 4393 12819 4439
rect 13457 4459 13503 4505
rect 12812 4265 12858 4311
rect 13423 4305 13751 4351
rect 13297 4177 13343 4223
rect 14298 4390 14344 4436
rect 14941 4281 14987 4421
rect 15613 4281 15659 4421
rect 16285 4281 16331 4421
rect 16728 4393 16868 4439
rect 16736 4266 16876 4312
rect 17741 4281 17787 4421
rect 2090 3404 2136 3450
rect 2746 3459 2792 3599
rect 2982 3365 3028 3693
rect 3889 3617 3935 3663
rect 3404 3529 3450 3575
rect 4015 3489 4343 3535
rect 3365 3401 3411 3447
rect 4049 3335 4095 3381
rect 4890 3404 4936 3450
rect 6010 3404 6056 3450
rect 6682 3404 6728 3450
rect 7338 3459 7384 3599
rect 7574 3365 7620 3693
rect 8481 3617 8527 3663
rect 7996 3529 8042 3575
rect 8607 3489 8935 3535
rect 7957 3401 8003 3447
rect 8641 3335 8687 3381
rect 9930 3404 9976 3450
rect 10602 3404 10648 3450
rect 11258 3459 11304 3599
rect 11494 3365 11540 3693
rect 12401 3617 12447 3663
rect 11916 3529 11962 3575
rect 12527 3489 12855 3535
rect 11877 3401 11923 3447
rect 12561 3335 12607 3381
rect 13685 3419 13731 3559
rect 14720 3528 14860 3574
rect 14298 3404 14344 3450
rect 14712 3401 14852 3447
rect 15178 3459 15224 3599
rect 15414 3365 15460 3693
rect 16321 3617 16367 3663
rect 15836 3529 15882 3575
rect 16447 3489 16775 3535
rect 15797 3401 15843 3447
rect 16481 3335 16527 3381
rect 17968 3528 18108 3574
rect 17576 3404 17622 3450
rect 17960 3401 18100 3447
<< metal1 >>
rect 1344 8650 18592 8684
rect 1344 8598 3370 8650
rect 3630 8598 7682 8650
rect 7942 8598 11994 8650
rect 12254 8598 16306 8650
rect 16566 8598 18592 8650
rect 1344 8564 18592 8598
rect 1418 8539 1486 8564
rect 1418 8493 1429 8539
rect 1475 8493 1486 8539
rect 1418 8411 1486 8493
rect 1418 8365 1429 8411
rect 1475 8365 1486 8411
rect 1418 8283 1486 8365
rect 1749 8505 1795 8564
rect 1749 8346 1795 8365
rect 1933 8505 1999 8518
rect 1933 8365 1953 8505
rect 1418 8237 1429 8283
rect 1475 8237 1486 8283
rect 1418 8224 1486 8237
rect 1822 8263 1887 8280
rect 1822 8146 1837 8263
rect 1883 8123 1887 8263
rect 1874 8094 1887 8123
rect 1822 8080 1887 8094
rect 1418 8066 1486 8078
rect 1418 7919 1429 8066
rect 1475 7919 1486 8066
rect 1418 7900 1486 7919
rect 1729 8032 1775 8072
rect 1729 7900 1775 7986
rect 1933 8034 1999 8365
rect 2401 8485 2447 8518
rect 2401 8367 2447 8439
rect 2605 8485 2651 8564
rect 3475 8527 3521 8564
rect 2605 8413 2651 8439
rect 2809 8485 3429 8518
rect 2855 8472 3429 8485
rect 2809 8413 2855 8439
rect 3000 8421 3116 8422
rect 3000 8375 3057 8421
rect 3103 8375 3116 8421
rect 2401 8321 2897 8367
rect 2943 8321 2954 8367
rect 2434 8258 2837 8264
rect 2434 8239 2494 8258
rect 2546 8239 2837 8258
rect 2434 8193 2489 8239
rect 2817 8193 2837 8239
rect 2434 8180 2837 8193
rect 2894 8085 2954 8321
rect 1933 7982 1934 8034
rect 1986 8032 1999 8034
rect 1986 7982 1999 7986
rect 1933 7946 1999 7982
rect 2388 8039 2737 8085
rect 2783 8039 2954 8085
rect 3000 8362 3116 8375
rect 2388 7992 2460 8039
rect 3000 7992 3046 8362
rect 3162 8316 3208 8472
rect 3106 8270 3208 8316
rect 3258 8407 3336 8426
rect 3258 8361 3271 8407
rect 3317 8361 3336 8407
rect 3106 8084 3174 8270
rect 3106 8038 3117 8084
rect 3163 8038 3174 8084
rect 3258 8146 3336 8361
rect 3382 8394 3429 8472
rect 3906 8520 3952 8564
rect 3475 8440 3521 8481
rect 3702 8502 3748 8515
rect 4778 8527 4846 8564
rect 3906 8463 3952 8474
rect 4141 8502 4187 8515
rect 3702 8394 3748 8456
rect 4141 8417 4187 8456
rect 3382 8347 3748 8394
rect 3804 8397 4187 8417
rect 3382 8279 3428 8347
rect 3382 8220 3428 8233
rect 3258 8094 3278 8146
rect 3330 8094 3336 8146
rect 3258 8084 3336 8094
rect 3258 8038 3269 8084
rect 3315 8038 3336 8084
rect 3421 8151 3467 8164
rect 3467 8105 3739 8113
rect 3421 8067 3739 8105
rect 3421 7992 3467 8067
rect 2388 7946 2401 7992
rect 2447 7946 2460 7992
rect 2614 7946 2625 7992
rect 2671 7946 2682 7992
rect 2832 7946 2849 7992
rect 2895 7946 3467 7992
rect 3538 7982 3584 8021
rect 2614 7900 2682 7946
rect 3669 7992 3739 8067
rect 3850 8370 4187 8397
rect 4561 8505 4655 8516
rect 4561 8365 4585 8505
rect 4631 8365 4655 8505
rect 4778 8481 4789 8527
rect 4835 8481 4846 8527
rect 5342 8539 5410 8564
rect 4778 8466 4846 8481
rect 5026 8508 5103 8518
rect 5026 8462 5037 8508
rect 5083 8462 5103 8508
rect 5026 8403 5103 8462
rect 3900 8303 4232 8315
rect 3900 8163 4040 8303
rect 4086 8258 4232 8303
rect 4086 8206 4174 8258
rect 4226 8206 4232 8258
rect 4086 8163 4232 8206
rect 3900 8152 4232 8163
rect 4561 8160 4655 8365
rect 4701 8356 5103 8403
rect 4701 8263 4758 8356
rect 4747 8217 4758 8263
rect 4701 8206 4758 8217
rect 4834 8237 5011 8278
rect 4834 8191 4931 8237
rect 4977 8191 5011 8237
rect 4834 8166 5011 8191
rect 4561 8146 4686 8160
rect 3850 8069 4044 8095
rect 3804 8049 4044 8069
rect 3669 7946 3682 7992
rect 3728 7946 3739 7992
rect 3906 7992 3952 8003
rect 3998 7992 4044 8049
rect 4561 8094 4622 8146
rect 4674 8094 4686 8146
rect 4561 8016 4686 8094
rect 3998 7946 4161 7992
rect 4207 7946 4220 7992
rect 4561 7970 4565 8016
rect 4611 7970 4686 8016
rect 4908 8034 5011 8166
rect 4561 7955 4686 7970
rect 4789 8000 4835 8013
rect 4908 7982 4958 8034
rect 5010 7982 5011 8034
rect 5057 8059 5103 8356
rect 5342 8493 5353 8539
rect 5399 8493 5410 8539
rect 5342 8411 5410 8493
rect 5342 8365 5353 8411
rect 5399 8365 5410 8411
rect 5342 8283 5410 8365
rect 5342 8237 5353 8283
rect 5399 8237 5410 8283
rect 5342 8226 5410 8237
rect 5537 8497 5583 8518
rect 5537 8151 5583 8357
rect 5841 8497 5887 8564
rect 5841 8338 5887 8357
rect 5985 8497 6031 8518
rect 5634 8232 5648 8278
rect 5788 8232 5887 8278
rect 5537 8105 5640 8151
rect 5780 8105 5792 8151
rect 5057 8000 5103 8013
rect 5342 8066 5410 8077
rect 4908 7970 5011 7982
rect 3538 7900 3584 7936
rect 3906 7900 3952 7946
rect 4789 7900 4835 7954
rect 5342 7919 5353 8066
rect 5399 7919 5410 8066
rect 5342 7900 5410 7919
rect 5537 8032 5583 8057
rect 5537 7900 5583 7986
rect 5841 8032 5887 8232
rect 5985 8151 6031 8357
rect 6289 8497 6335 8564
rect 6289 8338 6335 8357
rect 6625 8505 6691 8518
rect 6671 8365 6691 8505
rect 6082 8232 6096 8278
rect 6236 8232 6335 8278
rect 5985 8105 6088 8151
rect 6228 8105 6240 8151
rect 5841 7946 5887 7986
rect 5985 8032 6031 8057
rect 5985 7900 6031 7986
rect 6289 8032 6335 8232
rect 6289 7946 6335 7986
rect 6625 8034 6691 8365
rect 6829 8505 6875 8564
rect 6829 8346 6875 8365
rect 7217 8485 7263 8518
rect 7217 8367 7263 8439
rect 7421 8485 7467 8564
rect 8291 8527 8337 8564
rect 7421 8413 7467 8439
rect 7625 8485 8245 8518
rect 7671 8472 8245 8485
rect 7625 8413 7671 8439
rect 7816 8421 7932 8422
rect 7816 8375 7873 8421
rect 7919 8375 7932 8421
rect 7217 8321 7713 8367
rect 7759 8321 7770 8367
rect 6737 8263 6802 8280
rect 6737 8123 6741 8263
rect 6787 8146 6802 8263
rect 7250 8258 7653 8264
rect 7250 8239 7310 8258
rect 7362 8239 7653 8258
rect 7250 8193 7305 8239
rect 7633 8193 7653 8239
rect 7250 8180 7653 8193
rect 6737 8094 6750 8123
rect 6737 8080 6802 8094
rect 7710 8085 7770 8321
rect 6625 8032 6638 8034
rect 6625 7982 6638 7986
rect 6690 7982 6691 8034
rect 6625 7946 6691 7982
rect 6849 8032 6895 8072
rect 6849 7900 6895 7986
rect 7204 8039 7553 8085
rect 7599 8039 7770 8085
rect 7816 8362 7932 8375
rect 7204 7992 7276 8039
rect 7816 7992 7862 8362
rect 7978 8316 8024 8472
rect 7922 8270 8024 8316
rect 8074 8407 8152 8426
rect 8074 8361 8087 8407
rect 8133 8361 8152 8407
rect 7922 8084 7990 8270
rect 7922 8038 7933 8084
rect 7979 8038 7990 8084
rect 8074 8146 8152 8361
rect 8198 8394 8245 8472
rect 8722 8520 8768 8564
rect 8291 8440 8337 8481
rect 8518 8502 8564 8515
rect 9262 8539 9330 8564
rect 8722 8463 8768 8474
rect 8957 8502 9003 8515
rect 8518 8394 8564 8456
rect 8957 8417 9003 8456
rect 8198 8347 8564 8394
rect 8620 8397 9003 8417
rect 8198 8279 8244 8347
rect 8198 8220 8244 8233
rect 8074 8094 8094 8146
rect 8146 8094 8152 8146
rect 8074 8084 8152 8094
rect 8074 8038 8085 8084
rect 8131 8038 8152 8084
rect 8237 8151 8283 8164
rect 8283 8105 8555 8113
rect 8237 8067 8555 8105
rect 8237 7992 8283 8067
rect 7204 7946 7217 7992
rect 7263 7946 7276 7992
rect 7430 7946 7441 7992
rect 7487 7946 7498 7992
rect 7648 7946 7665 7992
rect 7711 7946 8283 7992
rect 8354 7982 8400 8021
rect 7430 7900 7498 7946
rect 8485 7992 8555 8067
rect 8666 8370 9003 8397
rect 9262 8493 9273 8539
rect 9319 8493 9330 8539
rect 9262 8411 9330 8493
rect 9262 8365 9273 8411
rect 9319 8365 9330 8411
rect 8716 8303 9048 8315
rect 8716 8163 8856 8303
rect 8902 8258 9048 8303
rect 8930 8206 9048 8258
rect 9262 8283 9330 8365
rect 9813 8505 9859 8564
rect 9813 8346 9859 8365
rect 9997 8505 10063 8518
rect 9997 8365 10017 8505
rect 9262 8237 9273 8283
rect 9319 8237 9330 8283
rect 9262 8226 9330 8237
rect 9886 8263 9951 8280
rect 9886 8258 9901 8263
rect 8902 8163 9048 8206
rect 8716 8152 9048 8163
rect 9886 8123 9901 8206
rect 9947 8123 9951 8263
rect 8666 8069 8860 8095
rect 9886 8080 9951 8123
rect 8620 8049 8860 8069
rect 8485 7946 8498 7992
rect 8544 7946 8555 7992
rect 8722 7992 8768 8003
rect 8814 7992 8860 8049
rect 9262 8066 9330 8077
rect 8814 7946 8977 7992
rect 9023 7946 9036 7992
rect 8354 7900 8400 7936
rect 8722 7900 8768 7946
rect 9262 7919 9273 8066
rect 9319 7919 9330 8066
rect 9262 7900 9330 7919
rect 9793 8032 9839 8072
rect 9793 7900 9839 7986
rect 9997 8034 10063 8365
rect 9997 7982 9998 8034
rect 10050 8032 10063 8034
rect 10050 7982 10063 7986
rect 9997 7946 10063 7982
rect 10545 8505 10611 8518
rect 10591 8370 10611 8505
rect 10545 8318 10558 8365
rect 10610 8318 10611 8370
rect 10749 8505 10795 8564
rect 11392 8520 11438 8564
rect 11157 8502 11203 8515
rect 11823 8527 11869 8564
rect 11392 8463 11438 8474
rect 11596 8502 11642 8515
rect 11157 8417 11203 8456
rect 11157 8397 11540 8417
rect 11157 8370 11494 8397
rect 10749 8346 10795 8365
rect 10545 8032 10611 8318
rect 11112 8303 11444 8315
rect 10657 8263 10722 8280
rect 10657 8123 10661 8263
rect 10707 8146 10722 8263
rect 11112 8163 11258 8303
rect 11304 8258 11444 8303
rect 11304 8206 11342 8258
rect 11394 8206 11444 8258
rect 11304 8163 11444 8206
rect 11112 8152 11444 8163
rect 10657 8094 10670 8123
rect 10657 8080 10722 8094
rect 10591 7986 10611 8032
rect 10545 7946 10611 7986
rect 10769 8032 10815 8072
rect 11300 8069 11494 8095
rect 11596 8394 11642 8456
rect 11823 8440 11869 8481
rect 11915 8485 12535 8518
rect 11915 8472 12489 8485
rect 11915 8394 11962 8472
rect 11596 8347 11962 8394
rect 11916 8279 11962 8347
rect 11916 8220 11962 8233
rect 12008 8407 12086 8426
rect 12008 8361 12027 8407
rect 12073 8361 12086 8407
rect 11877 8151 11923 8164
rect 11300 8049 11540 8069
rect 11605 8105 11877 8113
rect 11605 8067 11923 8105
rect 11300 7992 11346 8049
rect 10769 7900 10815 7986
rect 11124 7946 11137 7992
rect 11183 7946 11346 7992
rect 11392 7992 11438 8003
rect 11605 7992 11675 8067
rect 11605 7946 11616 7992
rect 11662 7946 11675 7992
rect 11760 7982 11806 8021
rect 11392 7900 11438 7946
rect 11877 7992 11923 8067
rect 12008 8146 12086 8361
rect 12136 8316 12182 8472
rect 12228 8421 12344 8422
rect 12228 8375 12241 8421
rect 12287 8375 12344 8421
rect 12489 8413 12535 8439
rect 12693 8485 12739 8564
rect 13182 8539 13250 8564
rect 12693 8413 12739 8439
rect 12897 8485 12943 8518
rect 12228 8362 12344 8375
rect 12897 8367 12943 8439
rect 12136 8270 12238 8316
rect 12008 8094 12014 8146
rect 12066 8094 12086 8146
rect 12008 8084 12086 8094
rect 12008 8038 12029 8084
rect 12075 8038 12086 8084
rect 12170 8084 12238 8270
rect 12170 8038 12181 8084
rect 12227 8038 12238 8084
rect 12298 7992 12344 8362
rect 12390 8321 12401 8367
rect 12447 8321 12943 8367
rect 13182 8493 13193 8539
rect 13239 8493 13250 8539
rect 13182 8411 13250 8493
rect 13182 8365 13193 8411
rect 13239 8365 13250 8411
rect 12390 8085 12450 8321
rect 13182 8283 13250 8365
rect 12507 8258 12910 8264
rect 12507 8239 12574 8258
rect 12626 8239 12910 8258
rect 12507 8193 12527 8239
rect 12855 8193 12910 8239
rect 13182 8237 13193 8283
rect 13239 8237 13250 8283
rect 13182 8226 13250 8237
rect 13569 8505 13635 8518
rect 13615 8365 13635 8505
rect 12507 8180 12910 8193
rect 12390 8039 12561 8085
rect 12607 8039 12956 8085
rect 12884 7992 12956 8039
rect 11877 7946 12449 7992
rect 12495 7946 12512 7992
rect 12662 7946 12673 7992
rect 12719 7946 12730 7992
rect 12884 7946 12897 7992
rect 12943 7946 12956 7992
rect 13182 8066 13250 8077
rect 11760 7900 11806 7936
rect 12662 7900 12730 7946
rect 13182 7919 13193 8066
rect 13239 7919 13250 8066
rect 13569 8034 13635 8365
rect 13773 8505 13819 8564
rect 14528 8520 14574 8564
rect 14293 8502 14339 8515
rect 14959 8527 15005 8564
rect 14528 8463 14574 8474
rect 14732 8502 14778 8515
rect 14293 8417 14339 8456
rect 14293 8397 14676 8417
rect 14293 8370 14630 8397
rect 13773 8346 13819 8365
rect 14248 8303 14580 8315
rect 13681 8263 13746 8280
rect 13681 8123 13685 8263
rect 13731 8146 13746 8263
rect 14248 8163 14394 8303
rect 14440 8258 14580 8303
rect 14440 8206 14478 8258
rect 14530 8206 14580 8258
rect 14440 8163 14580 8206
rect 14248 8152 14580 8163
rect 13681 8094 13694 8123
rect 13681 8080 13746 8094
rect 13569 8032 13582 8034
rect 13569 7982 13582 7986
rect 13634 7982 13635 8034
rect 13569 7946 13635 7982
rect 13793 8032 13839 8072
rect 14436 8069 14630 8095
rect 14732 8394 14778 8456
rect 14959 8440 15005 8481
rect 15051 8485 15671 8518
rect 15051 8472 15625 8485
rect 15051 8394 15098 8472
rect 14732 8347 15098 8394
rect 15052 8279 15098 8347
rect 15052 8220 15098 8233
rect 15144 8407 15222 8426
rect 15144 8361 15163 8407
rect 15209 8361 15222 8407
rect 15013 8151 15059 8164
rect 14436 8049 14676 8069
rect 14741 8105 15013 8113
rect 14741 8067 15059 8105
rect 14436 7992 14482 8049
rect 13182 7900 13250 7919
rect 13793 7900 13839 7986
rect 14260 7946 14273 7992
rect 14319 7946 14482 7992
rect 14528 7992 14574 8003
rect 14741 7992 14811 8067
rect 14741 7946 14752 7992
rect 14798 7946 14811 7992
rect 14896 7982 14942 8021
rect 14528 7900 14574 7946
rect 15013 7992 15059 8067
rect 15144 8146 15222 8361
rect 15272 8316 15318 8472
rect 15364 8421 15480 8422
rect 15364 8375 15377 8421
rect 15423 8375 15480 8421
rect 15625 8413 15671 8439
rect 15829 8485 15875 8564
rect 15829 8413 15875 8439
rect 16033 8485 16079 8518
rect 15364 8362 15480 8375
rect 16033 8367 16079 8439
rect 15272 8270 15374 8316
rect 15144 8094 15150 8146
rect 15202 8094 15222 8146
rect 15144 8084 15222 8094
rect 15144 8038 15165 8084
rect 15211 8038 15222 8084
rect 15306 8084 15374 8270
rect 15306 8038 15317 8084
rect 15363 8038 15374 8084
rect 15434 7992 15480 8362
rect 15526 8321 15537 8367
rect 15583 8321 16079 8367
rect 16421 8505 16467 8564
rect 17102 8539 17170 8564
rect 16421 8346 16467 8365
rect 16605 8505 16671 8518
rect 16605 8370 16625 8505
rect 15526 8085 15586 8321
rect 16605 8318 16606 8370
rect 16658 8318 16671 8365
rect 15643 8258 16046 8264
rect 15643 8239 15822 8258
rect 15874 8239 16046 8258
rect 15643 8193 15663 8239
rect 15991 8193 16046 8239
rect 15643 8180 16046 8193
rect 16494 8263 16559 8280
rect 16494 8146 16509 8263
rect 16555 8123 16559 8263
rect 16546 8094 16559 8123
rect 15526 8039 15697 8085
rect 15743 8039 16092 8085
rect 16494 8080 16559 8094
rect 16020 7992 16092 8039
rect 15013 7946 15585 7992
rect 15631 7946 15648 7992
rect 15798 7946 15809 7992
rect 15855 7946 15866 7992
rect 16020 7946 16033 7992
rect 16079 7946 16092 7992
rect 16401 8032 16447 8072
rect 14896 7900 14942 7936
rect 15798 7900 15866 7946
rect 16401 7900 16447 7986
rect 16605 8032 16671 8318
rect 17102 8493 17113 8539
rect 17159 8493 17170 8539
rect 17102 8411 17170 8493
rect 17102 8365 17113 8411
rect 17159 8365 17170 8411
rect 17102 8283 17170 8365
rect 17429 8505 17475 8564
rect 17429 8346 17475 8365
rect 17613 8505 17679 8518
rect 17613 8365 17633 8505
rect 17102 8237 17113 8283
rect 17159 8237 17170 8283
rect 17102 8226 17170 8237
rect 17502 8263 17567 8280
rect 17502 8146 17517 8263
rect 17563 8123 17567 8263
rect 17554 8094 17567 8123
rect 17502 8080 17567 8094
rect 16605 7986 16625 8032
rect 16605 7946 16671 7986
rect 17102 8066 17170 8077
rect 17102 7919 17113 8066
rect 17159 7919 17170 8066
rect 17102 7900 17170 7919
rect 17409 8032 17455 8072
rect 17409 7900 17455 7986
rect 17613 8034 17679 8365
rect 17857 8497 17903 8518
rect 17857 8151 17903 8357
rect 18161 8497 18207 8564
rect 18161 8338 18207 8357
rect 18450 8539 18518 8564
rect 18450 8493 18461 8539
rect 18507 8493 18518 8539
rect 18450 8411 18518 8493
rect 18450 8365 18461 8411
rect 18507 8365 18518 8411
rect 18450 8283 18518 8365
rect 17954 8232 17968 8278
rect 18108 8232 18207 8278
rect 17857 8105 17960 8151
rect 18100 8105 18112 8151
rect 17613 7982 17614 8034
rect 17666 8032 17679 8034
rect 17666 7982 17679 7986
rect 17613 7946 17679 7982
rect 17857 8032 17903 8059
rect 17857 7900 17903 7986
rect 18161 8032 18207 8232
rect 18450 8237 18461 8283
rect 18507 8237 18518 8283
rect 18450 8224 18518 8237
rect 18161 7946 18207 7986
rect 18450 8066 18518 8078
rect 18450 7919 18461 8066
rect 18507 7919 18518 8066
rect 18450 7900 18518 7919
rect 1344 7866 18752 7900
rect 1344 7814 5526 7866
rect 5786 7814 9838 7866
rect 10098 7814 14150 7866
rect 14410 7814 18462 7866
rect 18722 7814 18752 7866
rect 1344 7780 18752 7814
rect 1418 7761 1486 7780
rect 1418 7614 1429 7761
rect 1475 7614 1486 7761
rect 1418 7602 1486 7614
rect 1729 7694 1775 7780
rect 2614 7734 2682 7780
rect 3538 7744 3584 7780
rect 1729 7608 1775 7648
rect 1933 7698 1999 7734
rect 1933 7646 1934 7698
rect 1986 7694 1999 7698
rect 1986 7646 1999 7648
rect 1822 7557 1887 7600
rect 1822 7474 1837 7557
rect 1418 7443 1486 7456
rect 1418 7397 1429 7443
rect 1475 7397 1486 7443
rect 1822 7417 1837 7422
rect 1883 7417 1887 7557
rect 1822 7400 1887 7417
rect 1418 7315 1486 7397
rect 1418 7269 1429 7315
rect 1475 7269 1486 7315
rect 1418 7187 1486 7269
rect 1418 7141 1429 7187
rect 1475 7141 1486 7187
rect 1418 7116 1486 7141
rect 1749 7315 1795 7334
rect 1749 7116 1795 7175
rect 1933 7315 1999 7646
rect 2388 7688 2401 7734
rect 2447 7688 2460 7734
rect 2614 7688 2625 7734
rect 2671 7688 2682 7734
rect 2832 7688 2849 7734
rect 2895 7688 3467 7734
rect 2388 7641 2460 7688
rect 2388 7595 2737 7641
rect 2783 7595 2954 7641
rect 2434 7487 2837 7500
rect 2434 7441 2489 7487
rect 2817 7441 2837 7487
rect 2434 7422 2494 7441
rect 2546 7422 2837 7441
rect 2434 7416 2837 7422
rect 2894 7359 2954 7595
rect 1933 7175 1953 7315
rect 1933 7162 1999 7175
rect 2401 7313 2897 7359
rect 2943 7313 2954 7359
rect 3000 7318 3046 7688
rect 3106 7596 3117 7642
rect 3163 7596 3174 7642
rect 3106 7410 3174 7596
rect 3258 7596 3269 7642
rect 3315 7596 3336 7642
rect 3258 7474 3336 7596
rect 3421 7613 3467 7688
rect 3906 7734 3952 7780
rect 3538 7659 3584 7698
rect 3669 7688 3682 7734
rect 3728 7688 3739 7734
rect 3669 7613 3739 7688
rect 3906 7677 3952 7688
rect 3998 7688 4161 7734
rect 4207 7688 4220 7734
rect 4609 7694 4675 7734
rect 3998 7631 4044 7688
rect 3421 7575 3739 7613
rect 3467 7567 3739 7575
rect 3804 7611 4044 7631
rect 3421 7516 3467 7529
rect 3258 7422 3278 7474
rect 3330 7422 3336 7474
rect 3106 7364 3208 7410
rect 2401 7241 2447 7313
rect 3000 7305 3116 7318
rect 2401 7162 2447 7195
rect 2605 7241 2651 7267
rect 2605 7116 2651 7195
rect 2809 7241 2855 7267
rect 3000 7259 3057 7305
rect 3103 7259 3116 7305
rect 3000 7258 3116 7259
rect 3162 7208 3208 7364
rect 3258 7319 3336 7422
rect 3258 7273 3271 7319
rect 3317 7273 3336 7319
rect 3258 7254 3336 7273
rect 3382 7447 3428 7460
rect 3382 7333 3428 7401
rect 3382 7286 3748 7333
rect 3382 7208 3429 7286
rect 2855 7195 3429 7208
rect 2809 7162 3429 7195
rect 3475 7199 3521 7240
rect 3702 7224 3748 7286
rect 3850 7585 4044 7611
rect 4655 7648 4675 7694
rect 3900 7517 4232 7528
rect 3900 7377 4040 7517
rect 4086 7474 4232 7517
rect 4086 7422 4174 7474
rect 4226 7422 4232 7474
rect 4086 7377 4232 7422
rect 3900 7365 4232 7377
rect 4609 7315 4675 7648
rect 4833 7694 4879 7780
rect 4833 7608 4879 7648
rect 4977 7694 5023 7780
rect 4977 7626 5023 7648
rect 5281 7694 5327 7734
rect 4721 7557 4786 7600
rect 4721 7417 4725 7557
rect 4771 7474 4786 7557
rect 4771 7417 4786 7422
rect 4721 7400 4786 7417
rect 4977 7529 5080 7575
rect 5220 7529 5232 7575
rect 3850 7283 4187 7310
rect 3804 7263 4187 7283
rect 4141 7224 4187 7263
rect 3702 7165 3748 7178
rect 3906 7206 3952 7217
rect 3475 7116 3521 7153
rect 4141 7165 4187 7178
rect 4655 7250 4675 7315
rect 4674 7198 4675 7250
rect 4655 7175 4675 7198
rect 4609 7162 4675 7175
rect 4813 7315 4859 7334
rect 3906 7116 3952 7160
rect 4813 7116 4859 7175
rect 4977 7323 5023 7529
rect 5281 7448 5327 7648
rect 5425 7694 5471 7780
rect 5425 7626 5471 7648
rect 5729 7694 5775 7734
rect 5074 7402 5088 7448
rect 5228 7402 5327 7448
rect 5425 7529 5528 7575
rect 5668 7529 5680 7575
rect 4977 7162 5023 7183
rect 5281 7323 5327 7342
rect 5281 7116 5327 7183
rect 5425 7323 5471 7529
rect 5729 7448 5775 7648
rect 5873 7694 5919 7780
rect 5873 7626 5919 7648
rect 6177 7694 6223 7734
rect 5522 7402 5536 7448
rect 5676 7402 5775 7448
rect 5873 7529 5976 7575
rect 6116 7529 6128 7575
rect 5425 7162 5471 7183
rect 5729 7323 5775 7342
rect 5729 7116 5775 7183
rect 5873 7323 5919 7529
rect 6177 7448 6223 7648
rect 6321 7694 6367 7780
rect 6321 7626 6367 7648
rect 6625 7694 6671 7734
rect 5970 7402 5984 7448
rect 6124 7402 6223 7448
rect 6321 7529 6424 7575
rect 6564 7529 6576 7575
rect 5873 7162 5919 7183
rect 6177 7323 6223 7342
rect 6177 7116 6223 7183
rect 6321 7323 6367 7529
rect 6625 7448 6671 7648
rect 6769 7694 6815 7780
rect 7430 7734 7498 7780
rect 8354 7744 8400 7780
rect 6769 7621 6815 7648
rect 7073 7694 7119 7734
rect 6418 7402 6432 7448
rect 6572 7402 6671 7448
rect 6769 7529 6872 7575
rect 7012 7529 7024 7575
rect 6321 7162 6367 7183
rect 6625 7323 6671 7342
rect 6625 7116 6671 7183
rect 6769 7323 6815 7529
rect 7073 7448 7119 7648
rect 7204 7688 7217 7734
rect 7263 7688 7276 7734
rect 7430 7688 7441 7734
rect 7487 7688 7498 7734
rect 7648 7688 7665 7734
rect 7711 7688 8283 7734
rect 7204 7641 7276 7688
rect 7204 7595 7553 7641
rect 7599 7595 7770 7641
rect 6866 7402 6880 7448
rect 7020 7402 7119 7448
rect 7250 7487 7653 7500
rect 7250 7441 7305 7487
rect 7633 7441 7653 7487
rect 7250 7422 7310 7441
rect 7362 7422 7653 7441
rect 7250 7416 7653 7422
rect 7710 7359 7770 7595
rect 6769 7162 6815 7183
rect 7073 7323 7119 7342
rect 7073 7116 7119 7183
rect 7217 7313 7713 7359
rect 7759 7313 7770 7359
rect 7816 7318 7862 7688
rect 7922 7596 7933 7642
rect 7979 7596 7990 7642
rect 7922 7410 7990 7596
rect 8074 7596 8085 7642
rect 8131 7596 8152 7642
rect 7922 7364 8024 7410
rect 7217 7241 7263 7313
rect 7816 7305 7932 7318
rect 7217 7162 7263 7195
rect 7421 7241 7467 7267
rect 7421 7116 7467 7195
rect 7625 7241 7671 7267
rect 7816 7259 7873 7305
rect 7919 7259 7932 7305
rect 7816 7258 7932 7259
rect 7978 7208 8024 7364
rect 8074 7362 8152 7596
rect 8237 7613 8283 7688
rect 8722 7734 8768 7780
rect 9374 7761 9442 7780
rect 8354 7659 8400 7698
rect 8485 7688 8498 7734
rect 8544 7688 8555 7734
rect 8485 7613 8555 7688
rect 8722 7677 8768 7688
rect 8814 7688 8977 7734
rect 9023 7688 9036 7734
rect 8814 7631 8860 7688
rect 8237 7575 8555 7613
rect 8283 7567 8555 7575
rect 8620 7611 8860 7631
rect 8237 7516 8283 7529
rect 8074 7319 8094 7362
rect 8074 7273 8087 7319
rect 8146 7310 8152 7362
rect 8133 7273 8152 7310
rect 8074 7254 8152 7273
rect 8198 7447 8244 7460
rect 8198 7333 8244 7401
rect 8198 7286 8564 7333
rect 8198 7208 8245 7286
rect 7671 7195 8245 7208
rect 7625 7162 8245 7195
rect 8291 7199 8337 7240
rect 8518 7224 8564 7286
rect 8666 7585 8860 7611
rect 9374 7614 9385 7761
rect 9431 7614 9442 7761
rect 9569 7694 9615 7780
rect 9569 7621 9615 7648
rect 9873 7694 9919 7734
rect 9374 7603 9442 7614
rect 9569 7529 9672 7575
rect 9812 7529 9824 7575
rect 8716 7517 9048 7528
rect 8716 7377 8856 7517
rect 8902 7474 9048 7517
rect 8930 7422 9048 7474
rect 8902 7377 9048 7422
rect 8716 7365 9048 7377
rect 9374 7443 9442 7454
rect 9374 7397 9385 7443
rect 9431 7397 9442 7443
rect 9374 7315 9442 7397
rect 8666 7283 9003 7310
rect 8620 7263 9003 7283
rect 8957 7224 9003 7263
rect 8518 7165 8564 7178
rect 8722 7206 8768 7217
rect 8291 7116 8337 7153
rect 8957 7165 9003 7178
rect 9374 7269 9385 7315
rect 9431 7269 9442 7315
rect 9374 7187 9442 7269
rect 8722 7116 8768 7160
rect 9374 7141 9385 7187
rect 9431 7141 9442 7187
rect 9569 7323 9615 7529
rect 9873 7448 9919 7648
rect 10017 7694 10063 7780
rect 10017 7608 10063 7648
rect 10221 7694 10287 7734
rect 10221 7648 10241 7694
rect 9666 7402 9680 7448
rect 9820 7402 9919 7448
rect 10110 7557 10175 7600
rect 10110 7474 10125 7557
rect 10110 7417 10125 7422
rect 10171 7417 10175 7557
rect 10110 7400 10175 7417
rect 9569 7162 9615 7183
rect 9873 7323 9919 7342
rect 9374 7116 9442 7141
rect 9873 7116 9919 7183
rect 10037 7315 10083 7334
rect 10037 7116 10083 7175
rect 10221 7315 10287 7648
rect 10689 7694 10735 7780
rect 10689 7608 10735 7648
rect 10893 7694 10959 7734
rect 10893 7648 10913 7694
rect 10782 7557 10847 7600
rect 10782 7474 10797 7557
rect 10782 7417 10797 7422
rect 10843 7417 10847 7557
rect 10782 7400 10847 7417
rect 10221 7250 10241 7315
rect 10221 7198 10222 7250
rect 10221 7175 10241 7198
rect 10221 7162 10287 7175
rect 10709 7315 10755 7334
rect 10709 7116 10755 7175
rect 10893 7315 10959 7648
rect 11361 7694 11407 7780
rect 12246 7734 12314 7780
rect 13170 7744 13216 7780
rect 11361 7608 11407 7648
rect 11565 7694 11631 7734
rect 11565 7648 11585 7694
rect 11454 7557 11519 7600
rect 11454 7474 11469 7557
rect 11454 7417 11469 7422
rect 11515 7417 11519 7557
rect 11454 7400 11519 7417
rect 10893 7250 10913 7315
rect 10893 7198 10894 7250
rect 10893 7175 10913 7198
rect 10893 7162 10959 7175
rect 11381 7315 11427 7334
rect 11381 7116 11427 7175
rect 11565 7315 11631 7648
rect 12020 7688 12033 7734
rect 12079 7688 12092 7734
rect 12246 7688 12257 7734
rect 12303 7688 12314 7734
rect 12464 7688 12481 7734
rect 12527 7688 13099 7734
rect 12020 7641 12092 7688
rect 12020 7595 12369 7641
rect 12415 7595 12586 7641
rect 12066 7487 12469 7500
rect 12066 7441 12121 7487
rect 12449 7441 12469 7487
rect 12066 7422 12350 7441
rect 12402 7422 12469 7441
rect 12066 7416 12469 7422
rect 12526 7359 12586 7595
rect 11565 7250 11585 7315
rect 11565 7198 11566 7250
rect 11565 7175 11585 7198
rect 11565 7162 11631 7175
rect 12033 7313 12529 7359
rect 12575 7313 12586 7359
rect 12632 7318 12678 7688
rect 12738 7596 12749 7642
rect 12795 7596 12806 7642
rect 12738 7410 12806 7596
rect 12890 7596 12901 7642
rect 12947 7596 12968 7642
rect 12738 7364 12840 7410
rect 12033 7241 12079 7313
rect 12632 7305 12748 7318
rect 12033 7162 12079 7195
rect 12237 7241 12283 7267
rect 12237 7116 12283 7195
rect 12441 7241 12487 7267
rect 12632 7259 12689 7305
rect 12735 7259 12748 7305
rect 12632 7258 12748 7259
rect 12794 7208 12840 7364
rect 12890 7362 12968 7596
rect 13053 7613 13099 7688
rect 13538 7734 13584 7780
rect 13170 7659 13216 7698
rect 13301 7688 13314 7734
rect 13360 7688 13371 7734
rect 13301 7613 13371 7688
rect 13538 7677 13584 7688
rect 13630 7688 13793 7734
rect 13839 7688 13852 7734
rect 13937 7694 13983 7780
rect 14640 7734 14686 7780
rect 15008 7744 15054 7780
rect 13630 7631 13676 7688
rect 13053 7575 13371 7613
rect 13099 7567 13371 7575
rect 13436 7611 13676 7631
rect 13937 7621 13983 7648
rect 14241 7694 14287 7734
rect 14372 7688 14385 7734
rect 14431 7688 14594 7734
rect 13053 7516 13099 7529
rect 12890 7319 12910 7362
rect 12890 7273 12903 7319
rect 12962 7310 12968 7362
rect 12949 7273 12968 7310
rect 12890 7254 12968 7273
rect 13014 7447 13060 7460
rect 13014 7333 13060 7401
rect 13014 7286 13380 7333
rect 13014 7208 13061 7286
rect 12487 7195 13061 7208
rect 12441 7162 13061 7195
rect 13107 7199 13153 7240
rect 13334 7224 13380 7286
rect 13482 7585 13676 7611
rect 13937 7529 14040 7575
rect 14180 7529 14192 7575
rect 13532 7517 13864 7528
rect 13532 7377 13672 7517
rect 13718 7474 13864 7517
rect 13718 7422 13806 7474
rect 13858 7422 13864 7474
rect 13718 7377 13864 7422
rect 13532 7365 13864 7377
rect 13937 7323 13983 7529
rect 14241 7448 14287 7648
rect 14548 7631 14594 7688
rect 14640 7677 14686 7688
rect 14853 7688 14864 7734
rect 14910 7688 14923 7734
rect 14548 7611 14788 7631
rect 14548 7585 14742 7611
rect 14034 7402 14048 7448
rect 14188 7402 14287 7448
rect 14360 7517 14692 7528
rect 14360 7377 14506 7517
rect 14552 7474 14692 7517
rect 14552 7422 14590 7474
rect 14642 7422 14692 7474
rect 14552 7377 14692 7422
rect 14360 7365 14692 7377
rect 13482 7283 13819 7310
rect 13436 7263 13819 7283
rect 13773 7224 13819 7263
rect 13334 7165 13380 7178
rect 13538 7206 13584 7217
rect 13107 7116 13153 7153
rect 13773 7165 13819 7178
rect 13937 7162 13983 7183
rect 14241 7323 14287 7342
rect 13538 7116 13584 7160
rect 14241 7116 14287 7183
rect 14405 7283 14742 7310
rect 14853 7613 14923 7688
rect 15910 7734 15978 7780
rect 15008 7659 15054 7698
rect 15125 7688 15697 7734
rect 15743 7688 15760 7734
rect 15910 7688 15921 7734
rect 15967 7688 15978 7734
rect 16132 7688 16145 7734
rect 16191 7688 16204 7734
rect 15125 7613 15171 7688
rect 14853 7575 15171 7613
rect 14853 7567 15125 7575
rect 15125 7516 15171 7529
rect 15256 7596 15277 7642
rect 15323 7596 15334 7642
rect 15164 7447 15210 7460
rect 15164 7333 15210 7401
rect 14405 7263 14788 7283
rect 14844 7286 15210 7333
rect 14405 7224 14451 7263
rect 14844 7224 14890 7286
rect 14405 7165 14451 7178
rect 14640 7206 14686 7217
rect 14844 7165 14890 7178
rect 15071 7199 15117 7240
rect 14640 7116 14686 7160
rect 15163 7208 15210 7286
rect 15256 7362 15334 7596
rect 15418 7596 15429 7642
rect 15475 7596 15486 7642
rect 15418 7410 15486 7596
rect 15256 7310 15262 7362
rect 15314 7319 15334 7362
rect 15256 7273 15275 7310
rect 15321 7273 15334 7319
rect 15256 7254 15334 7273
rect 15384 7364 15486 7410
rect 15384 7208 15430 7364
rect 15546 7318 15592 7688
rect 16132 7641 16204 7688
rect 15476 7305 15592 7318
rect 15638 7595 15809 7641
rect 15855 7595 16204 7641
rect 16513 7694 16559 7780
rect 17326 7761 17394 7780
rect 16513 7608 16559 7648
rect 16717 7698 16783 7734
rect 16717 7646 16718 7698
rect 16770 7694 16783 7698
rect 16770 7646 16783 7648
rect 15638 7359 15698 7595
rect 16606 7557 16671 7600
rect 15755 7487 16158 7500
rect 15755 7441 15775 7487
rect 16103 7441 16158 7487
rect 15755 7422 15822 7441
rect 15874 7422 16158 7441
rect 15755 7416 16158 7422
rect 16606 7474 16621 7557
rect 16606 7417 16621 7422
rect 16667 7417 16671 7557
rect 16606 7400 16671 7417
rect 15638 7313 15649 7359
rect 15695 7313 16191 7359
rect 15476 7259 15489 7305
rect 15535 7259 15592 7305
rect 15476 7258 15592 7259
rect 15737 7241 15783 7267
rect 15163 7195 15737 7208
rect 15163 7162 15783 7195
rect 15941 7241 15987 7267
rect 15071 7116 15117 7153
rect 15941 7116 15987 7195
rect 16145 7241 16191 7313
rect 16145 7162 16191 7195
rect 16533 7315 16579 7334
rect 16533 7116 16579 7175
rect 16717 7315 16783 7646
rect 17326 7614 17337 7761
rect 17383 7614 17394 7761
rect 17326 7603 17394 7614
rect 17633 7694 17679 7780
rect 18450 7761 18518 7780
rect 17633 7608 17679 7648
rect 17837 7698 17903 7734
rect 17837 7646 17838 7698
rect 17890 7694 17903 7698
rect 17890 7646 17903 7648
rect 17726 7557 17791 7600
rect 17726 7474 17741 7557
rect 16717 7175 16737 7315
rect 16717 7162 16783 7175
rect 17326 7443 17394 7454
rect 17326 7397 17337 7443
rect 17383 7397 17394 7443
rect 17726 7417 17741 7422
rect 17787 7417 17791 7557
rect 17726 7400 17791 7417
rect 17326 7315 17394 7397
rect 17326 7269 17337 7315
rect 17383 7269 17394 7315
rect 17326 7187 17394 7269
rect 17326 7141 17337 7187
rect 17383 7141 17394 7187
rect 17326 7116 17394 7141
rect 17653 7315 17699 7334
rect 17653 7116 17699 7175
rect 17837 7315 17903 7646
rect 18450 7614 18461 7761
rect 18507 7614 18518 7761
rect 18450 7602 18518 7614
rect 17837 7175 17857 7315
rect 17837 7162 17903 7175
rect 18450 7443 18518 7456
rect 18450 7397 18461 7443
rect 18507 7397 18518 7443
rect 18450 7315 18518 7397
rect 18450 7269 18461 7315
rect 18507 7269 18518 7315
rect 18450 7187 18518 7269
rect 18450 7141 18461 7187
rect 18507 7141 18518 7187
rect 18450 7116 18518 7141
rect 1344 7082 18592 7116
rect 1344 7030 3370 7082
rect 3630 7030 7682 7082
rect 7942 7030 11994 7082
rect 12254 7030 16306 7082
rect 16566 7030 18592 7082
rect 1344 6996 18592 7030
rect 1418 6971 1486 6996
rect 1418 6925 1429 6971
rect 1475 6925 1486 6971
rect 1418 6843 1486 6925
rect 1418 6797 1429 6843
rect 1475 6797 1486 6843
rect 1418 6715 1486 6797
rect 1418 6669 1429 6715
rect 1475 6669 1486 6715
rect 1418 6656 1486 6669
rect 1617 6929 1663 6950
rect 1617 6583 1663 6789
rect 1921 6929 1967 6996
rect 1921 6770 1967 6789
rect 2086 6937 2212 6941
rect 2086 6797 2106 6937
rect 2152 6914 2212 6937
rect 2152 6862 2158 6914
rect 2210 6862 2212 6914
rect 2152 6797 2212 6862
rect 2086 6730 2212 6797
rect 2310 6937 2356 6996
rect 3434 6959 3502 6996
rect 2310 6778 2356 6797
rect 2484 6914 2556 6941
rect 2484 6862 2494 6914
rect 2546 6862 2556 6914
rect 2484 6744 2556 6862
rect 1714 6664 1728 6710
rect 1868 6664 1967 6710
rect 1617 6537 1720 6583
rect 1860 6537 1872 6583
rect 1418 6498 1486 6510
rect 1418 6351 1429 6498
rect 1475 6351 1486 6498
rect 1418 6332 1486 6351
rect 1617 6464 1663 6491
rect 1617 6332 1663 6418
rect 1921 6464 1967 6664
rect 1921 6378 1967 6418
rect 2086 6480 2152 6730
rect 2484 6698 2494 6744
rect 2540 6698 2556 6744
rect 2484 6620 2556 6698
rect 2604 6898 2786 6944
rect 2832 6898 2845 6944
rect 3217 6937 3311 6948
rect 2205 6589 2376 6600
rect 2205 6543 2216 6589
rect 2262 6574 2376 6589
rect 2604 6574 2650 6898
rect 2262 6543 2650 6574
rect 2205 6528 2650 6543
rect 2086 6464 2239 6480
rect 2132 6418 2239 6464
rect 2086 6394 2239 6418
rect 2310 6423 2356 6442
rect 2571 6424 2650 6528
rect 2696 6736 2780 6848
rect 2696 6690 2698 6736
rect 2744 6690 2780 6736
rect 2696 6638 2718 6690
rect 2770 6638 2780 6690
rect 2696 6487 2780 6638
rect 3217 6797 3241 6937
rect 3287 6797 3311 6937
rect 3434 6913 3445 6959
rect 3491 6913 3502 6959
rect 3434 6898 3502 6913
rect 3682 6940 3759 6950
rect 3682 6894 3693 6940
rect 3739 6894 3759 6940
rect 3682 6835 3759 6894
rect 3217 6592 3311 6797
rect 3357 6788 3759 6835
rect 3357 6695 3414 6788
rect 3403 6649 3414 6695
rect 3357 6638 3414 6649
rect 3490 6669 3667 6710
rect 3490 6623 3587 6669
rect 3633 6623 3667 6669
rect 3490 6598 3667 6623
rect 3217 6578 3342 6592
rect 3217 6526 3278 6578
rect 3330 6526 3342 6578
rect 3217 6448 3342 6526
rect 2571 6378 2582 6424
rect 2628 6378 2650 6424
rect 2806 6424 2852 6437
rect 3217 6402 3221 6448
rect 3267 6402 3342 6448
rect 3564 6466 3667 6598
rect 3217 6387 3342 6402
rect 3445 6432 3491 6445
rect 2310 6332 2356 6377
rect 2806 6332 2852 6378
rect 3564 6414 3614 6466
rect 3666 6414 3667 6466
rect 3713 6491 3759 6788
rect 3857 6929 3903 6950
rect 3857 6583 3903 6789
rect 4161 6929 4207 6996
rect 4161 6770 4207 6789
rect 4305 6929 4351 6950
rect 3954 6664 3968 6710
rect 4108 6664 4207 6710
rect 3857 6537 3960 6583
rect 4100 6537 4112 6583
rect 3713 6432 3759 6445
rect 3857 6464 3903 6489
rect 3564 6402 3667 6414
rect 3445 6332 3491 6386
rect 3857 6332 3903 6418
rect 4161 6464 4207 6664
rect 4305 6583 4351 6789
rect 4609 6929 4655 6996
rect 4609 6770 4655 6789
rect 4753 6929 4799 6950
rect 4402 6664 4416 6710
rect 4556 6664 4655 6710
rect 4305 6537 4408 6583
rect 4548 6537 4560 6583
rect 4161 6378 4207 6418
rect 4305 6464 4351 6489
rect 4305 6332 4351 6418
rect 4609 6464 4655 6664
rect 4753 6583 4799 6789
rect 5057 6929 5103 6996
rect 5057 6770 5103 6789
rect 5342 6971 5410 6996
rect 5342 6925 5353 6971
rect 5399 6925 5410 6971
rect 5342 6843 5410 6925
rect 5342 6797 5353 6843
rect 5399 6797 5410 6843
rect 5342 6715 5410 6797
rect 4850 6664 4864 6710
rect 5004 6664 5103 6710
rect 4753 6537 4856 6583
rect 4996 6537 5008 6583
rect 4609 6378 4655 6418
rect 4753 6464 4799 6491
rect 4753 6332 4799 6418
rect 5057 6464 5103 6664
rect 5342 6669 5353 6715
rect 5399 6669 5410 6715
rect 5342 6658 5410 6669
rect 5537 6929 5583 6950
rect 5537 6583 5583 6789
rect 5841 6929 5887 6996
rect 5841 6770 5887 6789
rect 5985 6929 6031 6950
rect 5634 6664 5648 6710
rect 5788 6664 5887 6710
rect 5537 6537 5640 6583
rect 5780 6537 5792 6583
rect 5057 6378 5103 6418
rect 5342 6498 5410 6509
rect 5342 6351 5353 6498
rect 5399 6351 5410 6498
rect 5342 6332 5410 6351
rect 5537 6464 5583 6489
rect 5537 6332 5583 6418
rect 5841 6464 5887 6664
rect 5985 6583 6031 6789
rect 6289 6929 6335 6996
rect 6289 6770 6335 6789
rect 6852 6921 6924 6950
rect 6852 6802 6868 6921
rect 6852 6750 6862 6802
rect 6914 6750 6924 6921
rect 6852 6733 6924 6750
rect 7072 6921 7118 6996
rect 7072 6744 7118 6781
rect 7461 6937 7507 6996
rect 7461 6778 7507 6797
rect 7645 6937 7711 6950
rect 7645 6914 7665 6937
rect 7645 6862 7646 6914
rect 7645 6797 7665 6862
rect 6082 6664 6096 6710
rect 6236 6664 6335 6710
rect 5985 6537 6088 6583
rect 6228 6537 6240 6583
rect 5841 6378 5887 6418
rect 5985 6464 6031 6489
rect 5985 6332 6031 6418
rect 6289 6464 6335 6664
rect 7534 6695 7599 6712
rect 6289 6378 6335 6418
rect 6848 6540 6936 6586
rect 6982 6540 6993 6586
rect 6848 6539 6993 6540
rect 7534 6578 7549 6695
rect 7595 6555 7599 6695
rect 6848 6447 6894 6539
rect 7586 6526 7599 6555
rect 7534 6512 7599 6526
rect 6848 6378 6894 6401
rect 7072 6444 7118 6504
rect 7072 6332 7118 6398
rect 7441 6464 7487 6504
rect 7441 6332 7487 6418
rect 7645 6464 7711 6797
rect 8133 6937 8179 6996
rect 8133 6778 8179 6797
rect 8317 6937 8383 6950
rect 8317 6914 8337 6937
rect 8317 6862 8318 6914
rect 8317 6797 8337 6862
rect 8206 6695 8271 6712
rect 8206 6578 8221 6695
rect 8267 6555 8271 6695
rect 8258 6526 8271 6555
rect 8206 6512 8271 6526
rect 7645 6418 7665 6464
rect 7645 6378 7711 6418
rect 8113 6464 8159 6504
rect 8113 6332 8159 6418
rect 8317 6464 8383 6797
rect 8805 6937 8851 6996
rect 8805 6778 8851 6797
rect 8989 6937 9055 6950
rect 8989 6797 9009 6937
rect 8878 6695 8943 6712
rect 8878 6578 8893 6695
rect 8939 6555 8943 6695
rect 8930 6526 8943 6555
rect 8878 6512 8943 6526
rect 8317 6418 8337 6464
rect 8317 6378 8383 6418
rect 8785 6464 8831 6504
rect 8785 6332 8831 6418
rect 8989 6466 9055 6797
rect 9477 6937 9523 6996
rect 9477 6778 9523 6797
rect 9661 6937 9727 6950
rect 9661 6797 9681 6937
rect 9550 6695 9615 6712
rect 9550 6578 9565 6695
rect 9611 6555 9615 6695
rect 9602 6526 9615 6555
rect 9550 6512 9615 6526
rect 8989 6414 8990 6466
rect 9042 6464 9055 6466
rect 9042 6414 9055 6418
rect 8989 6378 9055 6414
rect 9457 6464 9503 6504
rect 9457 6332 9503 6418
rect 9661 6466 9727 6797
rect 10149 6937 10195 6996
rect 10149 6778 10195 6797
rect 10333 6937 10399 6950
rect 10333 6797 10353 6937
rect 10222 6695 10287 6712
rect 10222 6578 10237 6695
rect 10283 6555 10287 6695
rect 10274 6526 10287 6555
rect 10222 6512 10287 6526
rect 9661 6414 9662 6466
rect 9714 6464 9727 6466
rect 9714 6414 9727 6418
rect 9661 6378 9727 6414
rect 10129 6464 10175 6504
rect 10129 6332 10175 6418
rect 10333 6466 10399 6797
rect 10821 6937 10867 6996
rect 10821 6778 10867 6797
rect 11005 6937 11071 6950
rect 11005 6797 11025 6937
rect 10894 6695 10959 6712
rect 10894 6578 10909 6695
rect 10955 6555 10959 6695
rect 10946 6526 10959 6555
rect 10894 6512 10959 6526
rect 10333 6414 10334 6466
rect 10386 6464 10399 6466
rect 10386 6414 10399 6418
rect 10333 6378 10399 6414
rect 10801 6464 10847 6504
rect 10801 6332 10847 6418
rect 11005 6466 11071 6797
rect 11493 6937 11539 6996
rect 11493 6778 11539 6797
rect 11677 6937 11743 6950
rect 11677 6797 11697 6937
rect 11566 6695 11631 6712
rect 11566 6578 11581 6695
rect 11627 6555 11631 6695
rect 11618 6526 11631 6555
rect 11566 6512 11631 6526
rect 11005 6414 11006 6466
rect 11058 6464 11071 6466
rect 11058 6414 11071 6418
rect 11005 6378 11071 6414
rect 11473 6464 11519 6504
rect 11473 6332 11519 6418
rect 11677 6466 11743 6797
rect 12165 6937 12211 6996
rect 12165 6778 12211 6797
rect 12349 6937 12415 6950
rect 12349 6797 12369 6937
rect 12238 6695 12303 6712
rect 12238 6578 12253 6695
rect 12299 6555 12303 6695
rect 12290 6526 12303 6555
rect 12238 6512 12303 6526
rect 11677 6414 11678 6466
rect 11730 6464 11743 6466
rect 11730 6414 11743 6418
rect 11677 6378 11743 6414
rect 12145 6464 12191 6504
rect 12145 6332 12191 6418
rect 12349 6466 12415 6797
rect 12593 6929 12639 6950
rect 12593 6583 12639 6789
rect 12897 6929 12943 6996
rect 12897 6770 12943 6789
rect 13294 6971 13362 6996
rect 13294 6925 13305 6971
rect 13351 6925 13362 6971
rect 13294 6843 13362 6925
rect 13294 6797 13305 6843
rect 13351 6797 13362 6843
rect 13294 6715 13362 6797
rect 13621 6937 13667 6996
rect 13621 6778 13667 6797
rect 13805 6937 13871 6950
rect 13805 6797 13825 6937
rect 12690 6664 12704 6710
rect 12844 6664 12943 6710
rect 12593 6537 12696 6583
rect 12836 6537 12848 6583
rect 12349 6414 12350 6466
rect 12402 6464 12415 6466
rect 12402 6414 12415 6418
rect 12349 6378 12415 6414
rect 12593 6464 12639 6491
rect 12593 6332 12639 6418
rect 12897 6464 12943 6664
rect 13294 6669 13305 6715
rect 13351 6669 13362 6715
rect 13294 6658 13362 6669
rect 13694 6695 13759 6712
rect 13694 6690 13709 6695
rect 13694 6555 13709 6638
rect 13755 6555 13759 6695
rect 13694 6512 13759 6555
rect 12897 6378 12943 6418
rect 13294 6498 13362 6509
rect 13294 6351 13305 6498
rect 13351 6351 13362 6498
rect 13294 6332 13362 6351
rect 13601 6464 13647 6504
rect 13601 6332 13647 6418
rect 13805 6466 13871 6797
rect 14293 6937 14339 6996
rect 14293 6778 14339 6797
rect 14477 6937 14543 6950
rect 14477 6797 14497 6937
rect 14366 6695 14431 6712
rect 14366 6690 14381 6695
rect 14366 6555 14381 6638
rect 14427 6555 14431 6695
rect 14366 6512 14431 6555
rect 13805 6414 13806 6466
rect 13858 6464 13871 6466
rect 13858 6414 13871 6418
rect 13805 6378 13871 6414
rect 14273 6464 14319 6504
rect 14273 6332 14319 6418
rect 14477 6466 14543 6797
rect 14965 6937 15011 6996
rect 14965 6778 15011 6797
rect 15149 6937 15215 6950
rect 15149 6797 15169 6937
rect 15038 6695 15103 6712
rect 15038 6690 15053 6695
rect 15038 6555 15053 6638
rect 15099 6555 15103 6695
rect 15038 6512 15103 6555
rect 14477 6414 14478 6466
rect 14530 6464 14543 6466
rect 14530 6414 14543 6418
rect 14477 6378 14543 6414
rect 14945 6464 14991 6504
rect 14945 6332 14991 6418
rect 15149 6466 15215 6797
rect 15637 6937 15683 6996
rect 15637 6778 15683 6797
rect 15821 6937 15887 6950
rect 15821 6914 15841 6937
rect 15821 6862 15822 6914
rect 15821 6797 15841 6862
rect 15710 6695 15775 6712
rect 15710 6690 15725 6695
rect 15710 6555 15725 6638
rect 15771 6555 15775 6695
rect 15710 6512 15775 6555
rect 15149 6414 15150 6466
rect 15202 6464 15215 6466
rect 15202 6414 15215 6418
rect 15149 6378 15215 6414
rect 15617 6464 15663 6504
rect 15617 6332 15663 6418
rect 15821 6464 15887 6797
rect 16309 6937 16355 6996
rect 16309 6778 16355 6797
rect 16493 6937 16559 6950
rect 16493 6797 16513 6937
rect 16382 6695 16447 6712
rect 16382 6578 16397 6695
rect 16443 6555 16447 6695
rect 16434 6526 16447 6555
rect 16382 6512 16447 6526
rect 15821 6418 15841 6464
rect 15821 6378 15887 6418
rect 16289 6464 16335 6504
rect 16289 6332 16335 6418
rect 16493 6466 16559 6797
rect 16981 6937 17027 6996
rect 16981 6778 17027 6797
rect 17165 6937 17231 6950
rect 17165 6797 17185 6937
rect 17054 6695 17119 6712
rect 17054 6578 17069 6695
rect 17115 6555 17119 6695
rect 17106 6526 17119 6555
rect 17054 6512 17119 6526
rect 16493 6414 16494 6466
rect 16546 6464 16559 6466
rect 16546 6414 16559 6418
rect 16493 6378 16559 6414
rect 16961 6464 17007 6504
rect 16961 6332 17007 6418
rect 17165 6466 17231 6797
rect 17653 6937 17699 6996
rect 18450 6971 18518 6996
rect 17653 6778 17699 6797
rect 17837 6937 17903 6950
rect 17837 6797 17857 6937
rect 17726 6695 17791 6712
rect 17726 6578 17741 6695
rect 17787 6555 17791 6695
rect 17778 6526 17791 6555
rect 17726 6512 17791 6526
rect 17165 6414 17166 6466
rect 17218 6464 17231 6466
rect 17218 6414 17231 6418
rect 17165 6378 17231 6414
rect 17633 6464 17679 6504
rect 17633 6332 17679 6418
rect 17837 6466 17903 6797
rect 18450 6925 18461 6971
rect 18507 6925 18518 6971
rect 18450 6843 18518 6925
rect 18450 6797 18461 6843
rect 18507 6797 18518 6843
rect 18450 6715 18518 6797
rect 18450 6669 18461 6715
rect 18507 6669 18518 6715
rect 18450 6656 18518 6669
rect 17837 6414 17838 6466
rect 17890 6464 17903 6466
rect 17890 6414 17903 6418
rect 17837 6378 17903 6414
rect 18450 6498 18518 6510
rect 18450 6351 18461 6498
rect 18507 6351 18518 6498
rect 18450 6332 18518 6351
rect 1344 6298 18752 6332
rect 1344 6246 5526 6298
rect 5786 6246 9838 6298
rect 10098 6246 14150 6298
rect 14410 6246 18462 6298
rect 18722 6246 18752 6298
rect 1344 6212 18752 6246
rect 1418 6193 1486 6212
rect 1418 6046 1429 6193
rect 1475 6046 1486 6193
rect 2181 6176 2227 6212
rect 2181 6119 2227 6130
rect 2370 6130 2454 6161
rect 1418 6034 1486 6046
rect 1729 6100 1775 6111
rect 2370 6078 2382 6130
rect 2434 6100 2454 6130
rect 1775 6054 2315 6061
rect 1729 6014 2315 6054
rect 1812 5903 1884 5964
rect 1418 5875 1486 5888
rect 1418 5829 1429 5875
rect 1475 5829 1486 5875
rect 1418 5747 1486 5829
rect 1418 5701 1429 5747
rect 1475 5701 1486 5747
rect 1812 5857 1825 5903
rect 1871 5857 1884 5903
rect 1812 5794 1884 5857
rect 1812 5742 1822 5794
rect 1874 5742 1884 5794
rect 1812 5710 1884 5742
rect 1418 5619 1486 5701
rect 1933 5664 1979 6014
rect 1418 5573 1429 5619
rect 1475 5573 1486 5619
rect 1418 5548 1486 5573
rect 1729 5616 1775 5627
rect 1933 5607 1979 5618
rect 2036 5906 2108 5964
rect 2036 5854 2046 5906
rect 2098 5854 2108 5906
rect 2269 5956 2315 6014
rect 2269 5875 2315 5910
rect 2370 6054 2405 6078
rect 2451 6054 2454 6100
rect 2036 5598 2108 5854
rect 2201 5747 2247 5766
rect 1729 5548 1775 5570
rect 2201 5548 2247 5607
rect 2370 5747 2454 6054
rect 2849 6126 2895 6212
rect 2849 6040 2895 6080
rect 3053 6130 3119 6166
rect 3053 6078 3054 6130
rect 3106 6126 3119 6130
rect 3106 6078 3119 6080
rect 2942 5989 3007 6032
rect 2942 5906 2957 5989
rect 2942 5849 2957 5854
rect 3003 5849 3007 5989
rect 2942 5832 3007 5849
rect 2370 5607 2405 5747
rect 2451 5607 2454 5747
rect 2370 5596 2454 5607
rect 2869 5747 2915 5766
rect 2869 5548 2915 5607
rect 3053 5747 3119 6078
rect 3297 6126 3343 6212
rect 3297 6058 3343 6080
rect 3601 6126 3647 6166
rect 3053 5607 3073 5747
rect 3053 5594 3119 5607
rect 3297 5961 3400 6007
rect 3540 5961 3552 6007
rect 3297 5755 3343 5961
rect 3601 5880 3647 6080
rect 3745 6126 3791 6212
rect 3745 6058 3791 6080
rect 4049 6126 4095 6166
rect 3394 5834 3408 5880
rect 3548 5834 3647 5880
rect 3745 5961 3848 6007
rect 3988 5961 4000 6007
rect 3297 5594 3343 5615
rect 3601 5755 3647 5774
rect 3601 5548 3647 5615
rect 3745 5755 3791 5961
rect 4049 5880 4095 6080
rect 4193 6126 4239 6212
rect 4193 6058 4239 6080
rect 4497 6126 4543 6166
rect 3842 5834 3856 5880
rect 3996 5834 4095 5880
rect 4193 5961 4296 6007
rect 4436 5961 4448 6007
rect 3745 5594 3791 5615
rect 4049 5755 4095 5774
rect 4049 5548 4095 5615
rect 4193 5755 4239 5961
rect 4497 5880 4543 6080
rect 4641 6126 4687 6212
rect 4641 6058 4687 6080
rect 4945 6126 4991 6166
rect 4290 5834 4304 5880
rect 4444 5834 4543 5880
rect 4641 5961 4744 6007
rect 4884 5961 4896 6007
rect 4193 5594 4239 5615
rect 4497 5755 4543 5774
rect 4497 5548 4543 5615
rect 4641 5755 4687 5961
rect 4945 5880 4991 6080
rect 5426 6146 5472 6212
rect 5426 6040 5472 6100
rect 5650 6143 5696 6166
rect 5650 6005 5696 6097
rect 5551 6004 5696 6005
rect 5551 5958 5562 6004
rect 5608 5958 5696 6004
rect 6177 6126 6243 6166
rect 6223 6080 6243 6126
rect 4738 5834 4752 5880
rect 4892 5834 4991 5880
rect 6177 5906 6243 6080
rect 6401 6126 6447 6212
rect 6401 6040 6447 6080
rect 6849 6126 6915 6166
rect 6895 6080 6915 6126
rect 6177 5854 6190 5906
rect 6242 5854 6243 5906
rect 4641 5594 4687 5615
rect 4945 5755 4991 5774
rect 4945 5548 4991 5615
rect 5426 5763 5472 5800
rect 5426 5548 5472 5623
rect 5620 5794 5692 5811
rect 5620 5623 5630 5794
rect 5682 5742 5692 5794
rect 5676 5623 5692 5742
rect 5620 5594 5692 5623
rect 6177 5747 6243 5854
rect 6289 6018 6354 6032
rect 6289 5989 6302 6018
rect 6289 5849 6293 5989
rect 6339 5849 6354 5966
rect 6289 5832 6354 5849
rect 6849 5906 6915 6080
rect 7073 6126 7119 6212
rect 7073 6040 7119 6080
rect 7441 6126 7487 6212
rect 7441 6040 7487 6080
rect 7645 6126 7711 6166
rect 7645 6080 7665 6126
rect 6849 5854 6862 5906
rect 6914 5854 6915 5906
rect 6223 5607 6243 5747
rect 6177 5594 6243 5607
rect 6381 5747 6427 5766
rect 6381 5548 6427 5607
rect 6849 5747 6915 5854
rect 6961 5989 7026 6032
rect 6961 5849 6965 5989
rect 7011 5906 7026 5989
rect 7011 5849 7026 5854
rect 6961 5832 7026 5849
rect 7534 5989 7599 6032
rect 7534 5906 7549 5989
rect 7534 5849 7549 5854
rect 7595 5849 7599 5989
rect 7534 5832 7599 5849
rect 7645 5906 7711 6080
rect 8114 6146 8160 6212
rect 8114 6040 8160 6100
rect 8338 6143 8384 6166
rect 8338 6005 8384 6097
rect 8785 6126 8831 6212
rect 9374 6193 9442 6212
rect 8785 6040 8831 6080
rect 8989 6130 9055 6166
rect 8989 6078 8990 6130
rect 9042 6126 9055 6130
rect 9042 6078 9055 6080
rect 8239 6004 8384 6005
rect 8239 5958 8250 6004
rect 8296 5958 8384 6004
rect 8878 6018 8943 6032
rect 8930 5989 8943 6018
rect 7645 5854 7646 5906
rect 7698 5854 7711 5906
rect 6895 5607 6915 5747
rect 6849 5594 6915 5607
rect 7053 5747 7099 5766
rect 7053 5548 7099 5607
rect 7461 5747 7507 5766
rect 7461 5548 7507 5607
rect 7645 5747 7711 5854
rect 8878 5849 8893 5966
rect 8939 5849 8943 5989
rect 8878 5832 8943 5849
rect 7645 5607 7665 5747
rect 7645 5594 7711 5607
rect 8114 5763 8160 5800
rect 8114 5548 8160 5623
rect 8308 5763 8380 5811
rect 8308 5623 8318 5763
rect 8364 5682 8380 5763
rect 8370 5630 8380 5682
rect 8364 5623 8380 5630
rect 8308 5594 8380 5623
rect 8805 5747 8851 5766
rect 8805 5548 8851 5607
rect 8989 5747 9055 6078
rect 9374 6046 9385 6193
rect 9431 6046 9442 6193
rect 9569 6126 9615 6212
rect 9569 6053 9615 6080
rect 9873 6126 9919 6166
rect 9374 6035 9442 6046
rect 9569 5961 9672 6007
rect 9812 5961 9824 6007
rect 8989 5607 9009 5747
rect 8989 5594 9055 5607
rect 9374 5875 9442 5886
rect 9374 5829 9385 5875
rect 9431 5829 9442 5875
rect 9374 5747 9442 5829
rect 9374 5701 9385 5747
rect 9431 5701 9442 5747
rect 9374 5619 9442 5701
rect 9374 5573 9385 5619
rect 9431 5573 9442 5619
rect 9569 5755 9615 5961
rect 9873 5880 9919 6080
rect 10241 6126 10287 6212
rect 10241 6040 10287 6080
rect 10445 6126 10511 6166
rect 10445 6080 10465 6126
rect 9666 5834 9680 5880
rect 9820 5834 9919 5880
rect 10334 5989 10399 6032
rect 10334 5906 10349 5989
rect 10334 5849 10349 5854
rect 10395 5849 10399 5989
rect 10334 5832 10399 5849
rect 9569 5594 9615 5615
rect 9873 5755 9919 5774
rect 9374 5548 9442 5573
rect 9873 5548 9919 5615
rect 10261 5747 10307 5766
rect 10261 5548 10307 5607
rect 10445 5747 10511 6080
rect 10913 6126 10959 6212
rect 10913 6040 10959 6080
rect 11117 6130 11183 6166
rect 11117 6078 11118 6130
rect 11170 6126 11183 6130
rect 11170 6078 11183 6080
rect 11006 5989 11071 6032
rect 11006 5906 11021 5989
rect 11006 5849 11021 5854
rect 11067 5849 11071 5989
rect 11006 5832 11071 5849
rect 10445 5682 10465 5747
rect 10445 5630 10446 5682
rect 10445 5607 10465 5630
rect 10445 5594 10511 5607
rect 10933 5747 10979 5766
rect 10933 5548 10979 5607
rect 11117 5747 11183 6078
rect 11585 6126 11631 6212
rect 11585 6040 11631 6080
rect 11789 6126 11855 6166
rect 11789 6080 11809 6126
rect 11678 5989 11743 6032
rect 11678 5906 11693 5989
rect 11678 5849 11693 5854
rect 11739 5849 11743 5989
rect 11678 5832 11743 5849
rect 11117 5607 11137 5747
rect 11117 5594 11183 5607
rect 11605 5747 11651 5766
rect 11605 5548 11651 5607
rect 11789 5747 11855 6080
rect 12257 6126 12303 6212
rect 12257 6040 12303 6080
rect 12461 6126 12527 6166
rect 12461 6080 12481 6126
rect 12350 5989 12415 6032
rect 12350 5906 12365 5989
rect 12350 5849 12365 5854
rect 12411 5849 12415 5989
rect 12350 5832 12415 5849
rect 11789 5682 11809 5747
rect 11789 5630 11790 5682
rect 11789 5607 11809 5630
rect 11789 5594 11855 5607
rect 12277 5747 12323 5766
rect 12277 5548 12323 5607
rect 12461 5747 12527 6080
rect 12929 6126 12975 6212
rect 12929 6040 12975 6080
rect 13133 6126 13199 6166
rect 13133 6080 13153 6126
rect 13022 5989 13087 6032
rect 13022 5906 13037 5989
rect 13022 5849 13037 5854
rect 13083 5849 13087 5989
rect 13022 5832 13087 5849
rect 12461 5682 12481 5747
rect 12461 5630 12462 5682
rect 12461 5607 12481 5630
rect 12461 5594 12527 5607
rect 12949 5747 12995 5766
rect 12949 5548 12995 5607
rect 13133 5747 13199 6080
rect 13601 6126 13647 6212
rect 13601 6040 13647 6080
rect 13805 6126 13871 6166
rect 13805 6080 13825 6126
rect 13694 6018 13759 6032
rect 13746 5989 13759 6018
rect 13694 5849 13709 5966
rect 13755 5849 13759 5989
rect 13694 5832 13759 5849
rect 13133 5682 13153 5747
rect 13133 5630 13134 5682
rect 13133 5607 13153 5630
rect 13133 5594 13199 5607
rect 13621 5747 13667 5766
rect 13621 5548 13667 5607
rect 13805 5747 13871 6080
rect 14273 6126 14319 6212
rect 14273 6040 14319 6080
rect 14477 6130 14543 6166
rect 14477 6078 14478 6130
rect 14530 6126 14543 6130
rect 14530 6078 14543 6080
rect 14366 5989 14431 6032
rect 14366 5906 14381 5989
rect 14366 5849 14381 5854
rect 14427 5849 14431 5989
rect 14366 5832 14431 5849
rect 13805 5682 13825 5747
rect 13805 5630 13806 5682
rect 13805 5607 13825 5630
rect 13805 5594 13871 5607
rect 14293 5747 14339 5766
rect 14293 5548 14339 5607
rect 14477 5747 14543 6078
rect 14945 6126 14991 6212
rect 14945 6040 14991 6080
rect 15149 6126 15215 6166
rect 15149 6080 15169 6126
rect 15038 6018 15103 6032
rect 15090 5989 15103 6018
rect 15038 5849 15053 5966
rect 15099 5849 15103 5989
rect 15038 5832 15103 5849
rect 14477 5607 14497 5747
rect 14477 5594 14543 5607
rect 14965 5747 15011 5766
rect 14965 5548 15011 5607
rect 15149 5747 15215 6080
rect 15617 6126 15663 6212
rect 15617 6040 15663 6080
rect 15821 6130 15887 6166
rect 15821 6078 15822 6130
rect 15874 6126 15887 6130
rect 15874 6078 15887 6080
rect 15710 5989 15775 6032
rect 15710 5906 15725 5989
rect 15710 5849 15725 5854
rect 15771 5849 15775 5989
rect 15710 5832 15775 5849
rect 15149 5682 15169 5747
rect 15149 5630 15150 5682
rect 15149 5607 15169 5630
rect 15149 5594 15215 5607
rect 15637 5747 15683 5766
rect 15637 5548 15683 5607
rect 15821 5747 15887 6078
rect 16290 6146 16336 6212
rect 16290 6040 16336 6100
rect 16514 6143 16560 6166
rect 16514 6005 16560 6097
rect 16737 6126 16783 6212
rect 17326 6193 17394 6212
rect 16737 6053 16783 6080
rect 17041 6126 17087 6166
rect 16415 6004 16560 6005
rect 16415 5958 16426 6004
rect 16472 5958 16560 6004
rect 16737 5961 16840 6007
rect 16980 5961 16992 6007
rect 15821 5607 15841 5747
rect 15821 5594 15887 5607
rect 16290 5763 16336 5800
rect 16290 5548 16336 5623
rect 16484 5794 16556 5811
rect 16484 5623 16494 5794
rect 16546 5742 16556 5794
rect 16540 5623 16556 5742
rect 16484 5594 16556 5623
rect 16737 5755 16783 5961
rect 17041 5880 17087 6080
rect 17326 6046 17337 6193
rect 17383 6046 17394 6193
rect 17326 6035 17394 6046
rect 17712 6143 17758 6166
rect 17712 6005 17758 6097
rect 17936 6146 17982 6212
rect 17936 6040 17982 6100
rect 18450 6193 18518 6212
rect 18450 6046 18461 6193
rect 18507 6046 18518 6193
rect 18450 6034 18518 6046
rect 17712 6004 17857 6005
rect 17712 5958 17800 6004
rect 17846 5958 17857 6004
rect 16834 5834 16848 5880
rect 16988 5834 17087 5880
rect 17326 5875 17394 5886
rect 17326 5829 17337 5875
rect 17383 5829 17394 5875
rect 16737 5594 16783 5615
rect 17041 5755 17087 5774
rect 17041 5548 17087 5615
rect 17326 5747 17394 5829
rect 18450 5875 18518 5888
rect 18450 5829 18461 5875
rect 18507 5829 18518 5875
rect 17326 5701 17337 5747
rect 17383 5701 17394 5747
rect 17326 5619 17394 5701
rect 17326 5573 17337 5619
rect 17383 5573 17394 5619
rect 17716 5763 17788 5811
rect 17716 5682 17732 5763
rect 17716 5630 17726 5682
rect 17716 5623 17732 5630
rect 17778 5623 17788 5763
rect 17716 5594 17788 5623
rect 17936 5763 17982 5800
rect 17326 5548 17394 5573
rect 17936 5548 17982 5623
rect 18450 5747 18518 5829
rect 18450 5701 18461 5747
rect 18507 5701 18518 5747
rect 18450 5619 18518 5701
rect 18450 5573 18461 5619
rect 18507 5573 18518 5619
rect 18450 5548 18518 5573
rect 1344 5514 18592 5548
rect 1344 5462 3370 5514
rect 3630 5462 7682 5514
rect 7942 5462 11994 5514
rect 12254 5462 16306 5514
rect 16566 5462 18592 5514
rect 1344 5428 18592 5462
rect 1418 5403 1486 5428
rect 1418 5357 1429 5403
rect 1475 5357 1486 5403
rect 1418 5275 1486 5357
rect 1418 5229 1429 5275
rect 1475 5229 1486 5275
rect 1418 5147 1486 5229
rect 1418 5101 1429 5147
rect 1475 5101 1486 5147
rect 1418 5088 1486 5101
rect 1617 5361 1663 5382
rect 1617 5015 1663 5221
rect 1921 5361 1967 5428
rect 1921 5202 1967 5221
rect 2065 5361 2111 5382
rect 1714 5096 1728 5142
rect 1868 5096 1967 5142
rect 1617 4969 1720 5015
rect 1860 4969 1872 5015
rect 1418 4930 1486 4942
rect 1418 4783 1429 4930
rect 1475 4783 1486 4930
rect 1418 4764 1486 4783
rect 1617 4896 1663 4918
rect 1617 4764 1663 4850
rect 1921 4896 1967 5096
rect 2065 5015 2111 5221
rect 2369 5361 2415 5428
rect 2369 5202 2415 5221
rect 2513 5361 2559 5382
rect 2162 5096 2176 5142
rect 2316 5096 2415 5142
rect 2065 4969 2168 5015
rect 2308 4969 2320 5015
rect 1921 4810 1967 4850
rect 2065 4896 2111 4918
rect 2065 4764 2111 4850
rect 2369 4896 2415 5096
rect 2513 5015 2559 5221
rect 2817 5361 2863 5428
rect 2817 5202 2863 5221
rect 2961 5361 3007 5382
rect 2610 5096 2624 5142
rect 2764 5096 2863 5142
rect 2513 4969 2616 5015
rect 2756 4969 2768 5015
rect 2369 4810 2415 4850
rect 2513 4896 2559 4918
rect 2513 4764 2559 4850
rect 2817 4896 2863 5096
rect 2961 5015 3007 5221
rect 3265 5361 3311 5428
rect 3265 5202 3311 5221
rect 3409 5361 3455 5382
rect 3058 5096 3072 5142
rect 3212 5096 3311 5142
rect 2961 4969 3064 5015
rect 3204 4969 3216 5015
rect 2817 4810 2863 4850
rect 2961 4896 3007 4918
rect 2961 4764 3007 4850
rect 3265 4896 3311 5096
rect 3409 5015 3455 5221
rect 3713 5361 3759 5428
rect 3713 5202 3759 5221
rect 4082 5353 4128 5428
rect 4082 5176 4128 5213
rect 4276 5353 4348 5382
rect 4276 5182 4286 5353
rect 4332 5234 4348 5353
rect 4338 5182 4348 5234
rect 4276 5165 4348 5182
rect 4754 5353 4800 5428
rect 5342 5403 5410 5428
rect 4754 5176 4800 5213
rect 4948 5353 5020 5382
rect 4948 5213 4958 5353
rect 5004 5346 5020 5353
rect 5010 5294 5020 5346
rect 5004 5213 5020 5294
rect 4948 5165 5020 5213
rect 5342 5357 5353 5403
rect 5399 5357 5410 5403
rect 5342 5275 5410 5357
rect 5342 5229 5353 5275
rect 5399 5229 5410 5275
rect 5342 5147 5410 5229
rect 3506 5096 3520 5142
rect 3660 5096 3759 5142
rect 3409 4969 3512 5015
rect 3652 4969 3664 5015
rect 3265 4810 3311 4850
rect 3409 4896 3455 4923
rect 3409 4764 3455 4850
rect 3713 4896 3759 5096
rect 5342 5101 5353 5147
rect 5399 5101 5410 5147
rect 5342 5090 5410 5101
rect 5537 5361 5583 5382
rect 4207 4972 4218 5018
rect 4264 4972 4352 5018
rect 4207 4971 4352 4972
rect 4879 4972 4890 5018
rect 4936 4972 5024 5018
rect 4879 4971 5024 4972
rect 3713 4810 3759 4850
rect 4082 4876 4128 4936
rect 4082 4764 4128 4830
rect 4306 4879 4352 4971
rect 4306 4810 4352 4833
rect 4754 4876 4800 4936
rect 4754 4764 4800 4830
rect 4978 4879 5024 4971
rect 5537 5015 5583 5221
rect 5841 5361 5887 5428
rect 5841 5202 5887 5221
rect 6210 5353 6256 5428
rect 6210 5176 6256 5213
rect 6404 5353 6476 5382
rect 6404 5213 6414 5353
rect 6460 5346 6476 5353
rect 6466 5294 6476 5346
rect 6460 5213 6476 5294
rect 6404 5165 6476 5213
rect 6964 5353 7036 5382
rect 6964 5346 6980 5353
rect 6964 5294 6974 5346
rect 6964 5213 6980 5294
rect 7026 5213 7036 5353
rect 6964 5165 7036 5213
rect 7184 5353 7230 5428
rect 7184 5176 7230 5213
rect 7633 5369 7699 5382
rect 7679 5229 7699 5369
rect 5634 5096 5648 5142
rect 5788 5096 5887 5142
rect 5537 4969 5640 5015
rect 5780 4969 5792 5015
rect 4978 4810 5024 4833
rect 5342 4930 5410 4941
rect 5342 4783 5353 4930
rect 5399 4783 5410 4930
rect 5342 4764 5410 4783
rect 5537 4896 5583 4923
rect 5537 4764 5583 4850
rect 5841 4896 5887 5096
rect 7633 5122 7699 5229
rect 7837 5369 7883 5428
rect 7837 5210 7883 5229
rect 8226 5353 8272 5428
rect 8226 5176 8272 5213
rect 8420 5353 8492 5382
rect 8420 5182 8430 5353
rect 8476 5234 8492 5353
rect 8482 5182 8492 5234
rect 8917 5369 8963 5428
rect 8917 5210 8963 5229
rect 9101 5369 9167 5382
rect 9101 5234 9121 5369
rect 8420 5165 8492 5182
rect 9101 5182 9102 5234
rect 9154 5182 9167 5229
rect 9589 5369 9635 5428
rect 9589 5210 9635 5229
rect 9773 5369 9839 5382
rect 9773 5234 9793 5369
rect 7633 5070 7646 5122
rect 7698 5070 7699 5122
rect 6335 4972 6346 5018
rect 6392 4972 6480 5018
rect 6335 4971 6480 4972
rect 5841 4810 5887 4850
rect 6210 4876 6256 4936
rect 6210 4764 6256 4830
rect 6434 4879 6480 4971
rect 6434 4810 6480 4833
rect 6960 4972 7048 5018
rect 7094 4972 7105 5018
rect 6960 4971 7105 4972
rect 6960 4879 7006 4971
rect 6960 4810 7006 4833
rect 7184 4876 7230 4936
rect 7184 4764 7230 4830
rect 7633 4896 7699 5070
rect 7745 5127 7810 5144
rect 7745 4987 7749 5127
rect 7795 5010 7810 5127
rect 8990 5127 9055 5144
rect 8990 5122 9005 5127
rect 7745 4958 7758 4987
rect 8351 4972 8362 5018
rect 8408 4972 8496 5018
rect 8351 4971 8496 4972
rect 7745 4944 7810 4958
rect 7679 4850 7699 4896
rect 7633 4810 7699 4850
rect 7857 4896 7903 4936
rect 7857 4764 7903 4850
rect 8226 4876 8272 4936
rect 8226 4764 8272 4830
rect 8450 4879 8496 4971
rect 8990 4987 9005 5070
rect 9051 4987 9055 5127
rect 8990 4944 9055 4987
rect 8450 4810 8496 4833
rect 8897 4896 8943 4936
rect 8897 4764 8943 4850
rect 9101 4896 9167 5182
rect 9773 5182 9774 5234
rect 9826 5182 9839 5229
rect 10261 5369 10307 5428
rect 10261 5210 10307 5229
rect 10445 5369 10511 5382
rect 10445 5234 10465 5369
rect 9662 5127 9727 5144
rect 9662 5122 9677 5127
rect 9662 4987 9677 5070
rect 9723 4987 9727 5127
rect 9662 4944 9727 4987
rect 9101 4850 9121 4896
rect 9101 4810 9167 4850
rect 9569 4896 9615 4936
rect 9569 4764 9615 4850
rect 9773 4896 9839 5182
rect 10445 5182 10446 5234
rect 10498 5182 10511 5229
rect 10933 5369 10979 5428
rect 10933 5210 10979 5229
rect 11117 5369 11183 5382
rect 11117 5234 11137 5369
rect 10334 5127 10399 5144
rect 10334 5122 10349 5127
rect 10334 4987 10349 5070
rect 10395 4987 10399 5127
rect 10334 4944 10399 4987
rect 9773 4850 9793 4896
rect 9773 4810 9839 4850
rect 10241 4896 10287 4936
rect 10241 4764 10287 4850
rect 10445 4896 10511 5182
rect 11117 5182 11118 5234
rect 11170 5182 11183 5229
rect 11605 5369 11651 5428
rect 11605 5210 11651 5229
rect 11789 5369 11855 5382
rect 11789 5229 11809 5369
rect 11006 5127 11071 5144
rect 11006 5122 11021 5127
rect 11006 4987 11021 5070
rect 11067 4987 11071 5127
rect 11006 4944 11071 4987
rect 10445 4850 10465 4896
rect 10445 4810 10511 4850
rect 10913 4896 10959 4936
rect 10913 4764 10959 4850
rect 11117 4896 11183 5182
rect 11678 5127 11743 5144
rect 11678 5122 11693 5127
rect 11678 4987 11693 5070
rect 11739 4987 11743 5127
rect 11678 4944 11743 4987
rect 11117 4850 11137 4896
rect 11117 4810 11183 4850
rect 11585 4896 11631 4936
rect 11585 4764 11631 4850
rect 11789 4898 11855 5229
rect 12277 5369 12323 5428
rect 12277 5210 12323 5229
rect 12461 5369 12527 5382
rect 12461 5229 12481 5369
rect 12350 5127 12415 5144
rect 12350 5122 12365 5127
rect 12350 4987 12365 5070
rect 12411 4987 12415 5127
rect 12350 4944 12415 4987
rect 12461 5122 12527 5229
rect 12461 5070 12462 5122
rect 12514 5070 12527 5122
rect 11789 4846 11790 4898
rect 11842 4896 11855 4898
rect 11842 4846 11855 4850
rect 11789 4810 11855 4846
rect 12257 4896 12303 4936
rect 12257 4764 12303 4850
rect 12461 4896 12527 5070
rect 12705 5361 12751 5382
rect 12705 5015 12751 5221
rect 13009 5361 13055 5428
rect 13009 5202 13055 5221
rect 13294 5403 13362 5428
rect 13294 5357 13305 5403
rect 13351 5357 13362 5403
rect 13294 5275 13362 5357
rect 13294 5229 13305 5275
rect 13351 5229 13362 5275
rect 13294 5147 13362 5229
rect 13621 5369 13667 5428
rect 13621 5210 13667 5229
rect 13805 5369 13871 5382
rect 13805 5229 13825 5369
rect 12802 5096 12816 5142
rect 12956 5096 13055 5142
rect 12705 4969 12808 5015
rect 12948 4969 12960 5015
rect 12461 4850 12481 4896
rect 12461 4810 12527 4850
rect 12705 4896 12751 4923
rect 12705 4764 12751 4850
rect 13009 4896 13055 5096
rect 13294 5101 13305 5147
rect 13351 5101 13362 5147
rect 13294 5090 13362 5101
rect 13694 5127 13759 5144
rect 13694 5122 13709 5127
rect 13694 4987 13709 5070
rect 13755 4987 13759 5127
rect 13694 4944 13759 4987
rect 13805 5122 13871 5229
rect 14293 5369 14339 5428
rect 14293 5210 14339 5229
rect 14477 5369 14543 5382
rect 14477 5234 14497 5369
rect 14477 5182 14478 5234
rect 14530 5182 14543 5229
rect 13805 5070 13806 5122
rect 13858 5070 13871 5122
rect 13009 4810 13055 4850
rect 13294 4930 13362 4941
rect 13294 4783 13305 4930
rect 13351 4783 13362 4930
rect 13294 4764 13362 4783
rect 13601 4896 13647 4936
rect 13601 4764 13647 4850
rect 13805 4896 13871 5070
rect 14366 5127 14431 5144
rect 14366 5122 14381 5127
rect 14366 4987 14381 5070
rect 14427 4987 14431 5127
rect 14366 4944 14431 4987
rect 13805 4850 13825 4896
rect 13805 4810 13871 4850
rect 14273 4896 14319 4936
rect 14273 4764 14319 4850
rect 14477 4896 14543 5182
rect 14477 4850 14497 4896
rect 14477 4810 14543 4850
rect 15025 5369 15091 5382
rect 15071 5229 15091 5369
rect 15025 4898 15091 5229
rect 15229 5369 15275 5428
rect 15229 5210 15275 5229
rect 15700 5353 15772 5382
rect 15700 5234 15716 5353
rect 15700 5182 15710 5234
rect 15762 5182 15772 5353
rect 15700 5165 15772 5182
rect 15920 5353 15966 5428
rect 16656 5384 16702 5428
rect 16421 5366 16467 5379
rect 17087 5391 17133 5428
rect 16656 5327 16702 5338
rect 16860 5366 16906 5379
rect 16421 5281 16467 5320
rect 16421 5261 16804 5281
rect 16421 5234 16758 5261
rect 15920 5176 15966 5213
rect 16376 5167 16708 5179
rect 15137 5127 15202 5144
rect 15137 4987 15141 5127
rect 15187 5122 15202 5127
rect 15187 4987 15202 5070
rect 16376 5122 16522 5167
rect 16376 5070 16382 5122
rect 16434 5070 16522 5122
rect 16376 5027 16522 5070
rect 16568 5027 16708 5167
rect 15137 4944 15202 4987
rect 15696 4972 15784 5018
rect 15830 4972 15841 5018
rect 16376 5016 16708 5027
rect 15696 4971 15841 4972
rect 15025 4896 15038 4898
rect 15025 4846 15038 4850
rect 15090 4846 15091 4898
rect 15025 4810 15091 4846
rect 15249 4896 15295 4936
rect 15249 4764 15295 4850
rect 15696 4879 15742 4971
rect 15696 4810 15742 4833
rect 15920 4876 15966 4936
rect 16564 4933 16758 4959
rect 16860 5258 16906 5320
rect 17087 5304 17133 5345
rect 17179 5349 17799 5382
rect 17179 5336 17753 5349
rect 17179 5258 17226 5336
rect 16860 5211 17226 5258
rect 17180 5143 17226 5211
rect 17180 5084 17226 5097
rect 17272 5271 17350 5290
rect 17272 5225 17291 5271
rect 17337 5225 17350 5271
rect 17272 5122 17350 5225
rect 17400 5180 17446 5336
rect 17492 5285 17608 5286
rect 17492 5239 17505 5285
rect 17551 5239 17608 5285
rect 17753 5277 17799 5303
rect 17957 5349 18003 5428
rect 18450 5403 18518 5428
rect 17957 5277 18003 5303
rect 18161 5349 18207 5382
rect 17492 5226 17608 5239
rect 18161 5231 18207 5303
rect 17400 5134 17502 5180
rect 17272 5070 17278 5122
rect 17330 5070 17350 5122
rect 17141 5015 17187 5028
rect 16564 4913 16804 4933
rect 16869 4969 17141 4977
rect 16869 4931 17187 4969
rect 16564 4856 16610 4913
rect 15920 4764 15966 4830
rect 16388 4810 16401 4856
rect 16447 4810 16610 4856
rect 16656 4856 16702 4867
rect 16869 4856 16939 4931
rect 16869 4810 16880 4856
rect 16926 4810 16939 4856
rect 17024 4846 17070 4885
rect 16656 4764 16702 4810
rect 17141 4856 17187 4931
rect 17272 4948 17350 5070
rect 17272 4902 17293 4948
rect 17339 4902 17350 4948
rect 17434 4948 17502 5134
rect 17434 4902 17445 4948
rect 17491 4902 17502 4948
rect 17562 4856 17608 5226
rect 17654 5185 17665 5231
rect 17711 5185 18207 5231
rect 18450 5357 18461 5403
rect 18507 5357 18518 5403
rect 18450 5275 18518 5357
rect 18450 5229 18461 5275
rect 18507 5229 18518 5275
rect 17654 4949 17714 5185
rect 18450 5147 18518 5229
rect 17771 5122 18174 5128
rect 17771 5103 17838 5122
rect 17890 5103 18174 5122
rect 17771 5057 17791 5103
rect 18119 5057 18174 5103
rect 18450 5101 18461 5147
rect 18507 5101 18518 5147
rect 18450 5088 18518 5101
rect 17771 5044 18174 5057
rect 17654 4903 17825 4949
rect 17871 4903 18220 4949
rect 18148 4856 18220 4903
rect 17141 4810 17713 4856
rect 17759 4810 17776 4856
rect 17926 4810 17937 4856
rect 17983 4810 17994 4856
rect 18148 4810 18161 4856
rect 18207 4810 18220 4856
rect 18450 4930 18518 4942
rect 17024 4764 17070 4800
rect 17926 4764 17994 4810
rect 18450 4783 18461 4930
rect 18507 4783 18518 4930
rect 18450 4764 18518 4783
rect 1344 4730 18752 4764
rect 1344 4678 5526 4730
rect 5786 4678 9838 4730
rect 10098 4678 14150 4730
rect 14410 4678 18462 4730
rect 18722 4678 18752 4730
rect 1344 4644 18752 4678
rect 1418 4625 1486 4644
rect 1418 4478 1429 4625
rect 1475 4478 1486 4625
rect 1617 4558 1663 4644
rect 1617 4487 1663 4512
rect 1921 4558 1967 4598
rect 1418 4466 1486 4478
rect 1617 4393 1720 4439
rect 1860 4393 1872 4439
rect 1418 4307 1486 4320
rect 1418 4261 1429 4307
rect 1475 4261 1486 4307
rect 1418 4179 1486 4261
rect 1418 4133 1429 4179
rect 1475 4133 1486 4179
rect 1418 4051 1486 4133
rect 1418 4005 1429 4051
rect 1475 4005 1486 4051
rect 1617 4187 1663 4393
rect 1921 4312 1967 4512
rect 2065 4558 2111 4644
rect 2838 4598 2906 4644
rect 3762 4608 3808 4644
rect 2065 4487 2111 4512
rect 2369 4558 2415 4598
rect 1714 4266 1728 4312
rect 1868 4266 1967 4312
rect 2065 4393 2168 4439
rect 2308 4393 2320 4439
rect 1617 4026 1663 4047
rect 1921 4187 1967 4206
rect 1418 3980 1486 4005
rect 1921 3980 1967 4047
rect 2065 4187 2111 4393
rect 2369 4312 2415 4512
rect 2612 4552 2625 4598
rect 2671 4552 2684 4598
rect 2838 4552 2849 4598
rect 2895 4552 2906 4598
rect 3056 4552 3073 4598
rect 3119 4552 3691 4598
rect 2612 4505 2684 4552
rect 2612 4459 2961 4505
rect 3007 4459 3178 4505
rect 2162 4266 2176 4312
rect 2316 4266 2415 4312
rect 2658 4351 3061 4364
rect 2658 4305 2713 4351
rect 3041 4305 3061 4351
rect 2658 4286 2718 4305
rect 2770 4286 3061 4305
rect 2658 4280 3061 4286
rect 3118 4223 3178 4459
rect 2065 4026 2111 4047
rect 2369 4187 2415 4206
rect 2369 3980 2415 4047
rect 2625 4177 3121 4223
rect 3167 4177 3178 4223
rect 3224 4182 3270 4552
rect 3330 4460 3341 4506
rect 3387 4460 3398 4506
rect 3330 4274 3398 4460
rect 3482 4460 3493 4506
rect 3539 4460 3560 4506
rect 3482 4450 3560 4460
rect 3482 4398 3502 4450
rect 3554 4398 3560 4450
rect 3330 4228 3432 4274
rect 2625 4105 2671 4177
rect 3224 4169 3340 4182
rect 2625 4026 2671 4059
rect 2829 4105 2875 4131
rect 2829 3980 2875 4059
rect 3033 4105 3079 4131
rect 3224 4123 3281 4169
rect 3327 4123 3340 4169
rect 3224 4122 3340 4123
rect 3386 4072 3432 4228
rect 3482 4183 3560 4398
rect 3645 4477 3691 4552
rect 4130 4598 4176 4644
rect 3762 4523 3808 4562
rect 3893 4552 3906 4598
rect 3952 4552 3963 4598
rect 3893 4477 3963 4552
rect 4130 4541 4176 4552
rect 4222 4552 4385 4598
rect 4431 4552 4444 4598
rect 4529 4558 4575 4644
rect 4222 4495 4268 4552
rect 3645 4439 3963 4477
rect 3691 4431 3963 4439
rect 4028 4475 4268 4495
rect 4529 4485 4575 4512
rect 4833 4558 4879 4598
rect 3645 4380 3691 4393
rect 3482 4137 3495 4183
rect 3541 4137 3560 4183
rect 3482 4118 3560 4137
rect 3606 4311 3652 4324
rect 3606 4197 3652 4265
rect 3606 4150 3972 4197
rect 3606 4072 3653 4150
rect 3079 4059 3653 4072
rect 3033 4026 3653 4059
rect 3699 4063 3745 4104
rect 3926 4088 3972 4150
rect 4074 4449 4268 4475
rect 4529 4393 4632 4439
rect 4772 4393 4784 4439
rect 4124 4381 4456 4392
rect 4124 4241 4264 4381
rect 4310 4338 4456 4381
rect 4338 4286 4456 4338
rect 4310 4241 4456 4286
rect 4124 4229 4456 4241
rect 4529 4187 4575 4393
rect 4833 4312 4879 4512
rect 5090 4578 5136 4644
rect 5090 4472 5136 4532
rect 5314 4575 5360 4598
rect 5314 4437 5360 4529
rect 5762 4578 5808 4644
rect 5762 4472 5808 4532
rect 5986 4575 6032 4598
rect 5986 4437 6032 4529
rect 6434 4578 6480 4644
rect 7360 4598 7406 4644
rect 7728 4608 7774 4644
rect 6434 4472 6480 4532
rect 6658 4575 6704 4598
rect 7092 4552 7105 4598
rect 7151 4552 7314 4598
rect 6658 4437 6704 4529
rect 7268 4495 7314 4552
rect 7360 4541 7406 4552
rect 7573 4552 7584 4598
rect 7630 4552 7643 4598
rect 7268 4475 7508 4495
rect 7268 4449 7462 4475
rect 5215 4436 5360 4437
rect 5215 4390 5226 4436
rect 5272 4390 5360 4436
rect 5887 4436 6032 4437
rect 5887 4390 5898 4436
rect 5944 4390 6032 4436
rect 6559 4436 6704 4437
rect 6559 4390 6570 4436
rect 6616 4390 6704 4436
rect 4626 4266 4640 4312
rect 4780 4266 4879 4312
rect 7080 4381 7412 4392
rect 7080 4338 7226 4381
rect 7080 4286 7086 4338
rect 7138 4286 7226 4338
rect 4074 4147 4411 4174
rect 4028 4127 4411 4147
rect 4365 4088 4411 4127
rect 3926 4029 3972 4042
rect 4130 4070 4176 4081
rect 3699 3980 3745 4017
rect 4365 4029 4411 4042
rect 4529 4026 4575 4047
rect 4833 4187 4879 4206
rect 4130 3980 4176 4024
rect 4833 3980 4879 4047
rect 5090 4195 5136 4232
rect 5090 3980 5136 4055
rect 5284 4195 5356 4243
rect 5284 4055 5294 4195
rect 5340 4114 5356 4195
rect 5346 4062 5356 4114
rect 5340 4055 5356 4062
rect 5284 4026 5356 4055
rect 5762 4195 5808 4232
rect 5762 3980 5808 4055
rect 5956 4226 6028 4243
rect 5956 4055 5966 4226
rect 6018 4174 6028 4226
rect 6012 4055 6028 4174
rect 5956 4026 6028 4055
rect 6434 4195 6480 4232
rect 6434 3980 6480 4055
rect 6628 4226 6700 4243
rect 7080 4241 7226 4286
rect 7272 4241 7412 4381
rect 7080 4229 7412 4241
rect 6628 4055 6638 4226
rect 6690 4174 6700 4226
rect 6684 4055 6700 4174
rect 6628 4026 6700 4055
rect 7125 4147 7462 4174
rect 7573 4477 7643 4552
rect 8630 4598 8698 4644
rect 9374 4625 9442 4644
rect 7728 4523 7774 4562
rect 7845 4552 8417 4598
rect 8463 4552 8480 4598
rect 8630 4552 8641 4598
rect 8687 4552 8698 4598
rect 8852 4552 8865 4598
rect 8911 4552 8924 4598
rect 7845 4477 7891 4552
rect 7573 4439 7891 4477
rect 7573 4431 7845 4439
rect 7845 4380 7891 4393
rect 7976 4460 7997 4506
rect 8043 4460 8054 4506
rect 7976 4450 8054 4460
rect 7976 4398 7982 4450
rect 8034 4398 8054 4450
rect 7884 4311 7930 4324
rect 7884 4197 7930 4265
rect 7125 4127 7508 4147
rect 7564 4150 7930 4197
rect 7125 4088 7171 4127
rect 7564 4088 7610 4150
rect 7125 4029 7171 4042
rect 7360 4070 7406 4081
rect 7564 4029 7610 4042
rect 7791 4063 7837 4104
rect 7360 3980 7406 4024
rect 7883 4072 7930 4150
rect 7976 4183 8054 4398
rect 8138 4460 8149 4506
rect 8195 4460 8206 4506
rect 8138 4274 8206 4460
rect 7976 4137 7995 4183
rect 8041 4137 8054 4183
rect 7976 4118 8054 4137
rect 8104 4228 8206 4274
rect 8104 4072 8150 4228
rect 8266 4182 8312 4552
rect 8852 4505 8924 4552
rect 8196 4169 8312 4182
rect 8358 4459 8529 4505
rect 8575 4459 8924 4505
rect 9374 4478 9385 4625
rect 9431 4478 9442 4625
rect 9569 4558 9615 4644
rect 9569 4485 9615 4512
rect 9873 4558 9919 4598
rect 9374 4467 9442 4478
rect 8358 4223 8418 4459
rect 9569 4393 9672 4439
rect 9812 4393 9824 4439
rect 8475 4351 8878 4364
rect 8475 4305 8495 4351
rect 8823 4305 8878 4351
rect 8475 4286 8654 4305
rect 8706 4286 8878 4305
rect 8475 4280 8878 4286
rect 9374 4307 9442 4318
rect 9374 4261 9385 4307
rect 9431 4261 9442 4307
rect 8358 4177 8369 4223
rect 8415 4177 8911 4223
rect 8196 4123 8209 4169
rect 8255 4123 8312 4169
rect 8196 4122 8312 4123
rect 8457 4105 8503 4131
rect 7883 4059 8457 4072
rect 7883 4026 8503 4059
rect 8661 4105 8707 4131
rect 7791 3980 7837 4017
rect 8661 3980 8707 4059
rect 8865 4105 8911 4177
rect 8865 4026 8911 4059
rect 9374 4179 9442 4261
rect 9374 4133 9385 4179
rect 9431 4133 9442 4179
rect 9374 4051 9442 4133
rect 9374 4005 9385 4051
rect 9431 4005 9442 4051
rect 9569 4187 9615 4393
rect 9873 4312 9919 4512
rect 10018 4578 10064 4644
rect 10018 4472 10064 4532
rect 10242 4575 10288 4598
rect 10242 4437 10288 4529
rect 10143 4436 10288 4437
rect 10143 4390 10154 4436
rect 10200 4390 10288 4436
rect 10769 4562 10835 4598
rect 10769 4558 10782 4562
rect 10769 4510 10782 4512
rect 10834 4510 10835 4562
rect 9666 4266 9680 4312
rect 9820 4266 9919 4312
rect 9569 4026 9615 4047
rect 9873 4187 9919 4206
rect 9374 3980 9442 4005
rect 9873 3980 9919 4047
rect 10018 4195 10064 4232
rect 10018 3980 10064 4055
rect 10212 4195 10284 4243
rect 10212 4055 10222 4195
rect 10268 4114 10284 4195
rect 10274 4062 10284 4114
rect 10268 4055 10284 4062
rect 10212 4026 10284 4055
rect 10769 4179 10835 4510
rect 10993 4558 11039 4644
rect 10993 4472 11039 4512
rect 11441 4562 11507 4598
rect 11441 4558 11454 4562
rect 11441 4510 11454 4512
rect 11506 4510 11507 4562
rect 10881 4450 10946 4464
rect 10881 4421 10894 4450
rect 10881 4281 10885 4421
rect 10931 4281 10946 4398
rect 10881 4264 10946 4281
rect 10815 4039 10835 4179
rect 10769 4026 10835 4039
rect 10973 4179 11019 4198
rect 10973 3980 11019 4039
rect 11441 4179 11507 4510
rect 11665 4558 11711 4644
rect 12288 4598 12334 4644
rect 12656 4608 12702 4644
rect 12020 4552 12033 4598
rect 12079 4552 12242 4598
rect 11665 4472 11711 4512
rect 12196 4495 12242 4552
rect 12288 4541 12334 4552
rect 12501 4552 12512 4598
rect 12558 4552 12571 4598
rect 12196 4475 12436 4495
rect 11553 4450 11618 4464
rect 11553 4421 11566 4450
rect 12196 4449 12390 4475
rect 11553 4281 11557 4421
rect 11603 4281 11618 4398
rect 11553 4264 11618 4281
rect 12008 4381 12340 4392
rect 12008 4338 12154 4381
rect 12008 4286 12014 4338
rect 12066 4286 12154 4338
rect 12008 4241 12154 4286
rect 12200 4241 12340 4381
rect 12008 4229 12340 4241
rect 11487 4039 11507 4179
rect 11441 4026 11507 4039
rect 11645 4179 11691 4198
rect 11645 3980 11691 4039
rect 12053 4147 12390 4174
rect 12501 4477 12571 4552
rect 13558 4598 13626 4644
rect 12656 4523 12702 4562
rect 12773 4552 13345 4598
rect 13391 4552 13408 4598
rect 13558 4552 13569 4598
rect 13615 4552 13626 4598
rect 13780 4552 13793 4598
rect 13839 4552 13852 4598
rect 12773 4477 12819 4552
rect 12501 4439 12819 4477
rect 12501 4431 12773 4439
rect 12773 4380 12819 4393
rect 12904 4460 12925 4506
rect 12971 4460 12982 4506
rect 12904 4450 12982 4460
rect 12904 4398 12910 4450
rect 12962 4398 12982 4450
rect 12812 4311 12858 4324
rect 12812 4197 12858 4265
rect 12053 4127 12436 4147
rect 12492 4150 12858 4197
rect 12053 4088 12099 4127
rect 12492 4088 12538 4150
rect 12053 4029 12099 4042
rect 12288 4070 12334 4081
rect 12492 4029 12538 4042
rect 12719 4063 12765 4104
rect 12288 3980 12334 4024
rect 12811 4072 12858 4150
rect 12904 4183 12982 4398
rect 13066 4460 13077 4506
rect 13123 4460 13134 4506
rect 13066 4274 13134 4460
rect 12904 4137 12923 4183
rect 12969 4137 12982 4183
rect 12904 4118 12982 4137
rect 13032 4228 13134 4274
rect 13032 4072 13078 4228
rect 13194 4182 13240 4552
rect 13780 4505 13852 4552
rect 13124 4169 13240 4182
rect 13286 4459 13457 4505
rect 13503 4459 13852 4505
rect 14162 4578 14208 4644
rect 14162 4472 14208 4532
rect 14386 4575 14432 4598
rect 13286 4223 13346 4459
rect 14386 4437 14432 4529
rect 14833 4558 14879 4644
rect 14833 4472 14879 4512
rect 15037 4562 15103 4598
rect 15037 4510 15038 4562
rect 15090 4558 15103 4562
rect 15090 4510 15103 4512
rect 14287 4436 14432 4437
rect 14287 4390 14298 4436
rect 14344 4390 14432 4436
rect 14926 4450 14991 4464
rect 14978 4421 14991 4450
rect 13403 4351 13806 4364
rect 13403 4305 13423 4351
rect 13751 4305 13806 4351
rect 13403 4286 13470 4305
rect 13522 4286 13806 4305
rect 14466 4286 14478 4338
rect 14530 4335 14542 4338
rect 14802 4335 14814 4338
rect 14530 4289 14814 4335
rect 14530 4286 14542 4289
rect 14802 4286 14814 4289
rect 14866 4286 14878 4338
rect 13403 4280 13806 4286
rect 14926 4281 14941 4398
rect 14987 4281 14991 4421
rect 14926 4264 14991 4281
rect 13286 4177 13297 4223
rect 13343 4177 13839 4223
rect 13124 4123 13137 4169
rect 13183 4123 13240 4169
rect 13124 4122 13240 4123
rect 13385 4105 13431 4131
rect 12811 4059 13385 4072
rect 12811 4026 13431 4059
rect 13589 4105 13635 4131
rect 12719 3980 12765 4017
rect 13589 3980 13635 4059
rect 13793 4105 13839 4177
rect 13793 4026 13839 4059
rect 14162 4195 14208 4232
rect 14162 3980 14208 4055
rect 14356 4226 14428 4243
rect 14356 4055 14366 4226
rect 14418 4174 14428 4226
rect 14412 4055 14428 4174
rect 14356 4026 14428 4055
rect 14853 4179 14899 4198
rect 14853 3980 14899 4039
rect 15037 4179 15103 4510
rect 15505 4558 15551 4644
rect 15505 4472 15551 4512
rect 15709 4562 15775 4598
rect 15709 4510 15710 4562
rect 15762 4558 15775 4562
rect 15762 4510 15775 4512
rect 15598 4421 15663 4464
rect 15598 4338 15613 4421
rect 15598 4281 15613 4286
rect 15659 4281 15663 4421
rect 15598 4264 15663 4281
rect 15037 4039 15057 4179
rect 15037 4026 15103 4039
rect 15525 4179 15571 4198
rect 15525 3980 15571 4039
rect 15709 4179 15775 4510
rect 16177 4558 16223 4644
rect 16177 4472 16223 4512
rect 16381 4562 16447 4598
rect 16381 4510 16382 4562
rect 16434 4558 16447 4562
rect 16434 4510 16447 4512
rect 16270 4450 16335 4464
rect 16322 4421 16335 4450
rect 16270 4281 16285 4398
rect 16331 4281 16335 4421
rect 16270 4264 16335 4281
rect 15709 4039 15729 4179
rect 15709 4026 15775 4039
rect 16197 4179 16243 4198
rect 16197 3980 16243 4039
rect 16381 4179 16447 4510
rect 16625 4558 16671 4644
rect 17326 4625 17394 4644
rect 16625 4485 16671 4512
rect 16929 4558 16975 4598
rect 16381 4039 16401 4179
rect 16381 4026 16447 4039
rect 16625 4393 16728 4439
rect 16868 4393 16880 4439
rect 16625 4187 16671 4393
rect 16929 4312 16975 4512
rect 17326 4478 17337 4625
rect 17383 4478 17394 4625
rect 17326 4467 17394 4478
rect 17633 4558 17679 4644
rect 18450 4625 18518 4644
rect 17633 4472 17679 4512
rect 17837 4562 17903 4598
rect 17837 4510 17838 4562
rect 17890 4558 17903 4562
rect 17890 4510 17903 4512
rect 17726 4421 17791 4464
rect 17726 4338 17741 4421
rect 16722 4266 16736 4312
rect 16876 4266 16975 4312
rect 17326 4307 17394 4318
rect 17326 4261 17337 4307
rect 17383 4261 17394 4307
rect 17726 4281 17741 4286
rect 17787 4281 17791 4421
rect 17726 4264 17791 4281
rect 16625 4026 16671 4047
rect 16929 4187 16975 4206
rect 16929 3980 16975 4047
rect 17326 4179 17394 4261
rect 17326 4133 17337 4179
rect 17383 4133 17394 4179
rect 17326 4051 17394 4133
rect 17326 4005 17337 4051
rect 17383 4005 17394 4051
rect 17326 3980 17394 4005
rect 17653 4179 17699 4198
rect 17653 3980 17699 4039
rect 17837 4179 17903 4510
rect 18450 4478 18461 4625
rect 18507 4478 18518 4625
rect 18450 4466 18518 4478
rect 17837 4039 17857 4179
rect 17837 4026 17903 4039
rect 18450 4307 18518 4320
rect 18450 4261 18461 4307
rect 18507 4261 18518 4307
rect 18450 4179 18518 4261
rect 18450 4133 18461 4179
rect 18507 4133 18518 4179
rect 18450 4051 18518 4133
rect 18450 4005 18461 4051
rect 18507 4005 18518 4051
rect 18450 3980 18518 4005
rect 1344 3946 18592 3980
rect 1344 3894 3370 3946
rect 3630 3894 7682 3946
rect 7942 3894 11994 3946
rect 12254 3894 16306 3946
rect 16566 3894 18592 3946
rect 1344 3860 18592 3894
rect 1418 3835 1486 3860
rect 1418 3789 1429 3835
rect 1475 3789 1486 3835
rect 1418 3707 1486 3789
rect 1418 3661 1429 3707
rect 1475 3661 1486 3707
rect 1418 3579 1486 3661
rect 1954 3785 2000 3860
rect 2880 3816 2926 3860
rect 1954 3608 2000 3645
rect 2148 3785 2220 3814
rect 2148 3614 2158 3785
rect 2204 3666 2220 3785
rect 2645 3798 2691 3811
rect 3311 3823 3357 3860
rect 2880 3759 2926 3770
rect 3084 3798 3130 3811
rect 2645 3713 2691 3752
rect 2645 3693 3028 3713
rect 2645 3666 2982 3693
rect 2210 3614 2220 3666
rect 2148 3597 2220 3614
rect 2600 3599 2932 3611
rect 1418 3533 1429 3579
rect 1475 3533 1486 3579
rect 1418 3520 1486 3533
rect 2600 3554 2746 3599
rect 2600 3502 2606 3554
rect 2658 3502 2746 3554
rect 2600 3459 2746 3502
rect 2792 3459 2932 3599
rect 2079 3404 2090 3450
rect 2136 3404 2224 3450
rect 2600 3448 2932 3459
rect 2079 3403 2224 3404
rect 1418 3362 1486 3374
rect 1418 3215 1429 3362
rect 1475 3215 1486 3362
rect 1418 3196 1486 3215
rect 1954 3308 2000 3368
rect 1954 3196 2000 3262
rect 2178 3311 2224 3403
rect 2788 3365 2982 3391
rect 3084 3690 3130 3752
rect 3311 3736 3357 3777
rect 3403 3781 4023 3814
rect 3403 3768 3977 3781
rect 3403 3690 3450 3768
rect 3084 3643 3450 3690
rect 3404 3575 3450 3643
rect 3404 3516 3450 3529
rect 3496 3703 3574 3722
rect 3496 3666 3515 3703
rect 3496 3614 3502 3666
rect 3561 3657 3574 3703
rect 3554 3614 3574 3657
rect 3365 3447 3411 3460
rect 2788 3345 3028 3365
rect 3093 3401 3365 3409
rect 3093 3363 3411 3401
rect 2788 3288 2834 3345
rect 2178 3242 2224 3265
rect 2612 3242 2625 3288
rect 2671 3242 2834 3288
rect 2880 3288 2926 3299
rect 3093 3288 3163 3363
rect 3093 3242 3104 3288
rect 3150 3242 3163 3288
rect 3248 3278 3294 3317
rect 2880 3196 2926 3242
rect 3365 3288 3411 3363
rect 3496 3380 3574 3614
rect 3624 3612 3670 3768
rect 3716 3717 3832 3718
rect 3716 3671 3729 3717
rect 3775 3671 3832 3717
rect 3977 3709 4023 3735
rect 4181 3781 4227 3860
rect 4181 3709 4227 3735
rect 4385 3781 4431 3814
rect 3716 3658 3832 3671
rect 4385 3663 4431 3735
rect 3624 3566 3726 3612
rect 3496 3334 3517 3380
rect 3563 3334 3574 3380
rect 3658 3380 3726 3566
rect 3658 3334 3669 3380
rect 3715 3334 3726 3380
rect 3786 3288 3832 3658
rect 3878 3617 3889 3663
rect 3935 3617 4431 3663
rect 4754 3785 4800 3860
rect 5342 3835 5410 3860
rect 3878 3381 3938 3617
rect 4754 3608 4800 3645
rect 4948 3785 5020 3814
rect 4948 3614 4958 3785
rect 5004 3666 5020 3785
rect 5010 3614 5020 3666
rect 4948 3597 5020 3614
rect 5342 3789 5353 3835
rect 5399 3789 5410 3835
rect 5342 3707 5410 3789
rect 5342 3661 5353 3707
rect 5399 3661 5410 3707
rect 5342 3579 5410 3661
rect 5874 3785 5920 3860
rect 5874 3608 5920 3645
rect 6068 3785 6140 3814
rect 6068 3645 6078 3785
rect 6124 3778 6140 3785
rect 6130 3726 6140 3778
rect 6124 3645 6140 3726
rect 6068 3597 6140 3645
rect 6546 3785 6592 3860
rect 7472 3816 7518 3860
rect 6546 3608 6592 3645
rect 6740 3785 6812 3814
rect 6740 3614 6750 3785
rect 6796 3666 6812 3785
rect 7237 3798 7283 3811
rect 7903 3823 7949 3860
rect 7472 3759 7518 3770
rect 7676 3798 7722 3811
rect 7237 3713 7283 3752
rect 7237 3693 7620 3713
rect 7237 3666 7574 3693
rect 6802 3614 6812 3666
rect 6740 3597 6812 3614
rect 7192 3599 7524 3611
rect 3995 3554 4398 3560
rect 3995 3535 4062 3554
rect 4114 3535 4398 3554
rect 3995 3489 4015 3535
rect 4343 3489 4398 3535
rect 5342 3533 5353 3579
rect 5399 3533 5410 3579
rect 5342 3522 5410 3533
rect 7192 3554 7338 3599
rect 3995 3476 4398 3489
rect 7192 3502 7198 3554
rect 7250 3502 7338 3554
rect 7192 3459 7338 3502
rect 7384 3459 7524 3599
rect 4879 3404 4890 3450
rect 4936 3404 5024 3450
rect 4879 3403 5024 3404
rect 5999 3404 6010 3450
rect 6056 3404 6144 3450
rect 5999 3403 6144 3404
rect 6671 3404 6682 3450
rect 6728 3404 6816 3450
rect 7192 3448 7524 3459
rect 6671 3403 6816 3404
rect 3878 3335 4049 3381
rect 4095 3335 4444 3381
rect 4372 3288 4444 3335
rect 3365 3242 3937 3288
rect 3983 3242 4000 3288
rect 4150 3242 4161 3288
rect 4207 3242 4218 3288
rect 4372 3242 4385 3288
rect 4431 3242 4444 3288
rect 4754 3308 4800 3368
rect 3248 3196 3294 3232
rect 4150 3196 4218 3242
rect 4754 3196 4800 3262
rect 4978 3311 5024 3403
rect 4978 3242 5024 3265
rect 5342 3362 5410 3373
rect 5342 3215 5353 3362
rect 5399 3215 5410 3362
rect 5342 3196 5410 3215
rect 5874 3308 5920 3368
rect 5874 3196 5920 3262
rect 6098 3311 6144 3403
rect 6098 3242 6144 3265
rect 6546 3308 6592 3368
rect 6546 3196 6592 3262
rect 6770 3311 6816 3403
rect 7380 3365 7574 3391
rect 7676 3690 7722 3752
rect 7903 3736 7949 3777
rect 7995 3781 8615 3814
rect 7995 3768 8569 3781
rect 7995 3690 8042 3768
rect 7676 3643 8042 3690
rect 7996 3575 8042 3643
rect 7996 3516 8042 3529
rect 8088 3703 8166 3722
rect 8088 3666 8107 3703
rect 8088 3614 8094 3666
rect 8153 3657 8166 3703
rect 8146 3614 8166 3657
rect 7957 3447 8003 3460
rect 7380 3345 7620 3365
rect 7685 3401 7957 3409
rect 7685 3363 8003 3401
rect 7380 3288 7426 3345
rect 6770 3242 6816 3265
rect 7204 3242 7217 3288
rect 7263 3242 7426 3288
rect 7472 3288 7518 3299
rect 7685 3288 7755 3363
rect 7685 3242 7696 3288
rect 7742 3242 7755 3288
rect 7840 3278 7886 3317
rect 7472 3196 7518 3242
rect 7957 3288 8003 3363
rect 8088 3380 8166 3614
rect 8216 3612 8262 3768
rect 8308 3717 8424 3718
rect 8308 3671 8321 3717
rect 8367 3671 8424 3717
rect 8569 3709 8615 3735
rect 8773 3781 8819 3860
rect 9262 3835 9330 3860
rect 8773 3709 8819 3735
rect 8977 3781 9023 3814
rect 8308 3658 8424 3671
rect 8977 3663 9023 3735
rect 8216 3566 8318 3612
rect 8088 3334 8109 3380
rect 8155 3334 8166 3380
rect 8250 3380 8318 3566
rect 8250 3334 8261 3380
rect 8307 3334 8318 3380
rect 8378 3288 8424 3658
rect 8470 3617 8481 3663
rect 8527 3617 9023 3663
rect 9262 3789 9273 3835
rect 9319 3789 9330 3835
rect 9262 3707 9330 3789
rect 9262 3661 9273 3707
rect 9319 3661 9330 3707
rect 8470 3381 8530 3617
rect 9262 3579 9330 3661
rect 9794 3785 9840 3860
rect 9794 3608 9840 3645
rect 9988 3785 10060 3814
rect 9988 3645 9998 3785
rect 10044 3778 10060 3785
rect 10050 3726 10060 3778
rect 10044 3645 10060 3726
rect 9988 3597 10060 3645
rect 10466 3785 10512 3860
rect 11392 3816 11438 3860
rect 10466 3608 10512 3645
rect 10660 3785 10732 3814
rect 10660 3645 10670 3785
rect 10716 3778 10732 3785
rect 10722 3726 10732 3778
rect 10716 3645 10732 3726
rect 11157 3798 11203 3811
rect 11823 3823 11869 3860
rect 11392 3759 11438 3770
rect 11596 3798 11642 3811
rect 11157 3713 11203 3752
rect 11157 3693 11540 3713
rect 11157 3666 11494 3693
rect 10660 3597 10732 3645
rect 11112 3599 11444 3611
rect 8587 3554 8990 3560
rect 8587 3535 8654 3554
rect 8706 3535 8990 3554
rect 8587 3489 8607 3535
rect 8935 3489 8990 3535
rect 9262 3533 9273 3579
rect 9319 3533 9330 3579
rect 9262 3522 9330 3533
rect 11112 3554 11258 3599
rect 8587 3476 8990 3489
rect 11112 3502 11118 3554
rect 11170 3502 11258 3554
rect 11112 3459 11258 3502
rect 11304 3459 11444 3599
rect 9919 3404 9930 3450
rect 9976 3404 10064 3450
rect 9919 3403 10064 3404
rect 10591 3404 10602 3450
rect 10648 3404 10736 3450
rect 11112 3448 11444 3459
rect 10591 3403 10736 3404
rect 8470 3335 8641 3381
rect 8687 3335 9036 3381
rect 8964 3288 9036 3335
rect 7957 3242 8529 3288
rect 8575 3242 8592 3288
rect 8742 3242 8753 3288
rect 8799 3242 8810 3288
rect 8964 3242 8977 3288
rect 9023 3242 9036 3288
rect 9262 3362 9330 3373
rect 7840 3196 7886 3232
rect 8742 3196 8810 3242
rect 9262 3215 9273 3362
rect 9319 3215 9330 3362
rect 9262 3196 9330 3215
rect 9794 3308 9840 3368
rect 9794 3196 9840 3262
rect 10018 3311 10064 3403
rect 10018 3242 10064 3265
rect 10466 3308 10512 3368
rect 10466 3196 10512 3262
rect 10690 3311 10736 3403
rect 11300 3365 11494 3391
rect 11596 3690 11642 3752
rect 11823 3736 11869 3777
rect 11915 3781 12535 3814
rect 11915 3768 12489 3781
rect 11915 3690 11962 3768
rect 11596 3643 11962 3690
rect 11916 3575 11962 3643
rect 11916 3516 11962 3529
rect 12008 3703 12086 3722
rect 12008 3666 12027 3703
rect 12008 3614 12014 3666
rect 12073 3657 12086 3703
rect 12066 3614 12086 3657
rect 11877 3447 11923 3460
rect 11300 3345 11540 3365
rect 11605 3401 11877 3409
rect 11605 3363 11923 3401
rect 11300 3288 11346 3345
rect 10690 3242 10736 3265
rect 11124 3242 11137 3288
rect 11183 3242 11346 3288
rect 11392 3288 11438 3299
rect 11605 3288 11675 3363
rect 11605 3242 11616 3288
rect 11662 3242 11675 3288
rect 11760 3278 11806 3317
rect 11392 3196 11438 3242
rect 11877 3288 11923 3363
rect 12008 3380 12086 3614
rect 12136 3612 12182 3768
rect 12228 3717 12344 3718
rect 12228 3671 12241 3717
rect 12287 3671 12344 3717
rect 12489 3709 12535 3735
rect 12693 3781 12739 3860
rect 13182 3835 13250 3860
rect 12693 3709 12739 3735
rect 12897 3781 12943 3814
rect 12228 3658 12344 3671
rect 12897 3663 12943 3735
rect 12136 3566 12238 3612
rect 12008 3334 12029 3380
rect 12075 3334 12086 3380
rect 12170 3380 12238 3566
rect 12170 3334 12181 3380
rect 12227 3334 12238 3380
rect 12298 3288 12344 3658
rect 12390 3617 12401 3663
rect 12447 3617 12943 3663
rect 13182 3789 13193 3835
rect 13239 3789 13250 3835
rect 13182 3707 13250 3789
rect 13182 3661 13193 3707
rect 13239 3661 13250 3707
rect 12390 3381 12450 3617
rect 13182 3579 13250 3661
rect 12507 3554 12910 3560
rect 12507 3535 12574 3554
rect 12626 3535 12910 3554
rect 12507 3489 12527 3535
rect 12855 3489 12910 3535
rect 13182 3533 13193 3579
rect 13239 3533 13250 3579
rect 13182 3522 13250 3533
rect 13569 3801 13635 3814
rect 13615 3661 13635 3801
rect 12507 3476 12910 3489
rect 12390 3335 12561 3381
rect 12607 3335 12956 3381
rect 12884 3288 12956 3335
rect 11877 3242 12449 3288
rect 12495 3242 12512 3288
rect 12662 3242 12673 3288
rect 12719 3242 12730 3288
rect 12884 3242 12897 3288
rect 12943 3242 12956 3288
rect 13182 3362 13250 3373
rect 11760 3196 11806 3232
rect 12662 3196 12730 3242
rect 13182 3215 13193 3362
rect 13239 3215 13250 3362
rect 13569 3330 13635 3661
rect 13773 3801 13819 3860
rect 13773 3642 13819 3661
rect 14162 3785 14208 3860
rect 14162 3608 14208 3645
rect 14356 3785 14428 3814
rect 14356 3645 14366 3785
rect 14412 3778 14428 3785
rect 14418 3726 14428 3778
rect 14412 3645 14428 3726
rect 14356 3597 14428 3645
rect 14609 3793 14655 3814
rect 13681 3559 13746 3576
rect 13681 3419 13685 3559
rect 13731 3554 13746 3559
rect 13731 3419 13746 3502
rect 13681 3376 13746 3419
rect 14287 3404 14298 3450
rect 14344 3404 14432 3450
rect 14287 3403 14432 3404
rect 13569 3328 13582 3330
rect 13569 3278 13582 3282
rect 13634 3278 13635 3330
rect 13569 3242 13635 3278
rect 13793 3328 13839 3368
rect 13182 3196 13250 3215
rect 13793 3196 13839 3282
rect 14162 3308 14208 3368
rect 14162 3196 14208 3262
rect 14386 3311 14432 3403
rect 14609 3447 14655 3653
rect 14913 3793 14959 3860
rect 15312 3816 15358 3860
rect 15077 3798 15123 3811
rect 15743 3823 15789 3860
rect 15312 3759 15358 3770
rect 15516 3798 15562 3811
rect 15077 3713 15123 3752
rect 15077 3693 15460 3713
rect 15077 3666 15414 3693
rect 14913 3634 14959 3653
rect 15032 3599 15364 3611
rect 14706 3528 14720 3574
rect 14860 3528 14959 3574
rect 14609 3401 14712 3447
rect 14852 3401 14864 3447
rect 14386 3242 14432 3265
rect 14609 3328 14655 3355
rect 14609 3196 14655 3282
rect 14913 3328 14959 3528
rect 15032 3554 15178 3599
rect 15032 3502 15150 3554
rect 15032 3459 15178 3502
rect 15224 3459 15364 3599
rect 15032 3448 15364 3459
rect 15220 3365 15414 3391
rect 15516 3690 15562 3752
rect 15743 3736 15789 3777
rect 15835 3781 16455 3814
rect 15835 3768 16409 3781
rect 15835 3690 15882 3768
rect 15516 3643 15882 3690
rect 15836 3575 15882 3643
rect 15836 3516 15882 3529
rect 15928 3703 16006 3722
rect 15928 3666 15947 3703
rect 15928 3614 15934 3666
rect 15993 3657 16006 3703
rect 15986 3614 16006 3657
rect 15797 3447 15843 3460
rect 15220 3345 15460 3365
rect 15525 3401 15797 3409
rect 15525 3363 15843 3401
rect 15220 3288 15266 3345
rect 14913 3242 14959 3282
rect 15044 3242 15057 3288
rect 15103 3242 15266 3288
rect 15312 3288 15358 3299
rect 15525 3288 15595 3363
rect 15525 3242 15536 3288
rect 15582 3242 15595 3288
rect 15680 3278 15726 3317
rect 15312 3196 15358 3242
rect 15797 3288 15843 3363
rect 15928 3380 16006 3614
rect 16056 3612 16102 3768
rect 16148 3717 16264 3718
rect 16148 3671 16161 3717
rect 16207 3671 16264 3717
rect 16409 3709 16455 3735
rect 16613 3781 16659 3860
rect 17102 3835 17170 3860
rect 16613 3709 16659 3735
rect 16817 3781 16863 3814
rect 16148 3658 16264 3671
rect 16817 3663 16863 3735
rect 16056 3566 16158 3612
rect 15928 3334 15949 3380
rect 15995 3334 16006 3380
rect 16090 3380 16158 3566
rect 16090 3334 16101 3380
rect 16147 3334 16158 3380
rect 16218 3288 16264 3658
rect 16310 3617 16321 3663
rect 16367 3617 16863 3663
rect 17102 3789 17113 3835
rect 17159 3789 17170 3835
rect 17102 3707 17170 3789
rect 17102 3661 17113 3707
rect 17159 3661 17170 3707
rect 16310 3381 16370 3617
rect 17102 3579 17170 3661
rect 17492 3785 17564 3814
rect 17492 3778 17508 3785
rect 17492 3726 17502 3778
rect 17492 3645 17508 3726
rect 17554 3645 17564 3785
rect 17492 3597 17564 3645
rect 17712 3785 17758 3860
rect 17712 3608 17758 3645
rect 17857 3793 17903 3814
rect 16427 3554 16830 3560
rect 16427 3535 16718 3554
rect 16770 3535 16830 3554
rect 16427 3489 16447 3535
rect 16775 3489 16830 3535
rect 17102 3533 17113 3579
rect 17159 3533 17170 3579
rect 17102 3522 17170 3533
rect 16427 3476 16830 3489
rect 17488 3404 17576 3450
rect 17622 3404 17633 3450
rect 17488 3403 17633 3404
rect 17857 3447 17903 3653
rect 18161 3793 18207 3860
rect 18161 3634 18207 3653
rect 18450 3835 18518 3860
rect 18450 3789 18461 3835
rect 18507 3789 18518 3835
rect 18450 3707 18518 3789
rect 18450 3661 18461 3707
rect 18507 3661 18518 3707
rect 18450 3579 18518 3661
rect 17954 3528 17968 3574
rect 18108 3528 18207 3574
rect 16310 3335 16481 3381
rect 16527 3335 16876 3381
rect 16804 3288 16876 3335
rect 15797 3242 16369 3288
rect 16415 3242 16432 3288
rect 16582 3242 16593 3288
rect 16639 3242 16650 3288
rect 16804 3242 16817 3288
rect 16863 3242 16876 3288
rect 17102 3362 17170 3373
rect 15680 3196 15726 3232
rect 16582 3196 16650 3242
rect 17102 3215 17113 3362
rect 17159 3215 17170 3362
rect 17488 3311 17534 3403
rect 17857 3401 17960 3447
rect 18100 3401 18112 3447
rect 17488 3242 17534 3265
rect 17712 3308 17758 3368
rect 17102 3196 17170 3215
rect 17712 3196 17758 3262
rect 17857 3328 17903 3355
rect 17857 3196 17903 3282
rect 18161 3328 18207 3528
rect 18450 3533 18461 3579
rect 18507 3533 18518 3579
rect 18450 3520 18518 3533
rect 18161 3242 18207 3282
rect 18450 3362 18518 3374
rect 18450 3215 18461 3362
rect 18507 3215 18518 3362
rect 18450 3196 18518 3215
rect 1344 3162 18752 3196
rect 1344 3110 5526 3162
rect 5786 3110 9838 3162
rect 10098 3110 14150 3162
rect 14410 3110 18462 3162
rect 18722 3110 18752 3162
rect 1344 3076 18752 3110
<< via1 >>
rect 3370 8598 3630 8650
rect 7682 8598 7942 8650
rect 11994 8598 12254 8650
rect 16306 8598 16566 8650
rect 1822 8123 1837 8146
rect 1837 8123 1874 8146
rect 1822 8094 1874 8123
rect 2494 8239 2546 8258
rect 2494 8206 2546 8239
rect 1934 8032 1986 8034
rect 1934 7986 1953 8032
rect 1953 7986 1986 8032
rect 1934 7982 1986 7986
rect 3278 8094 3330 8146
rect 4174 8206 4226 8258
rect 4622 8094 4674 8146
rect 4958 7982 5010 8034
rect 7310 8239 7362 8258
rect 7310 8206 7362 8239
rect 6750 8123 6787 8146
rect 6787 8123 6802 8146
rect 6750 8094 6802 8123
rect 6638 8032 6690 8034
rect 6638 7986 6671 8032
rect 6671 7986 6690 8032
rect 6638 7982 6690 7986
rect 8094 8094 8146 8146
rect 8878 8206 8902 8258
rect 8902 8206 8930 8258
rect 9886 8206 9901 8258
rect 9901 8206 9938 8258
rect 9998 8032 10050 8034
rect 9998 7986 10017 8032
rect 10017 7986 10050 8032
rect 9998 7982 10050 7986
rect 10558 8365 10591 8370
rect 10591 8365 10610 8370
rect 10558 8318 10610 8365
rect 11342 8206 11394 8258
rect 10670 8123 10707 8146
rect 10707 8123 10722 8146
rect 10670 8094 10722 8123
rect 12014 8094 12066 8146
rect 12574 8239 12626 8258
rect 12574 8206 12626 8239
rect 14478 8206 14530 8258
rect 13694 8123 13731 8146
rect 13731 8123 13746 8146
rect 13694 8094 13746 8123
rect 13582 8032 13634 8034
rect 13582 7986 13615 8032
rect 13615 7986 13634 8032
rect 13582 7982 13634 7986
rect 15150 8094 15202 8146
rect 16606 8365 16625 8370
rect 16625 8365 16658 8370
rect 16606 8318 16658 8365
rect 15822 8239 15874 8258
rect 15822 8206 15874 8239
rect 16494 8123 16509 8146
rect 16509 8123 16546 8146
rect 16494 8094 16546 8123
rect 17502 8123 17517 8146
rect 17517 8123 17554 8146
rect 17502 8094 17554 8123
rect 17614 8032 17666 8034
rect 17614 7986 17633 8032
rect 17633 7986 17666 8032
rect 17614 7982 17666 7986
rect 5526 7814 5786 7866
rect 9838 7814 10098 7866
rect 14150 7814 14410 7866
rect 18462 7814 18722 7866
rect 1934 7694 1986 7698
rect 1934 7648 1953 7694
rect 1953 7648 1986 7694
rect 1934 7646 1986 7648
rect 1822 7422 1837 7474
rect 1837 7422 1874 7474
rect 2494 7441 2546 7474
rect 2494 7422 2546 7441
rect 3278 7422 3330 7474
rect 4174 7422 4226 7474
rect 4734 7422 4771 7474
rect 4771 7422 4786 7474
rect 4622 7198 4655 7250
rect 4655 7198 4674 7250
rect 7310 7441 7362 7474
rect 7310 7422 7362 7441
rect 8094 7319 8146 7362
rect 8094 7310 8133 7319
rect 8133 7310 8146 7319
rect 8878 7422 8902 7474
rect 8902 7422 8930 7474
rect 10110 7422 10125 7474
rect 10125 7422 10162 7474
rect 10782 7422 10797 7474
rect 10797 7422 10834 7474
rect 10222 7198 10241 7250
rect 10241 7198 10274 7250
rect 11454 7422 11469 7474
rect 11469 7422 11506 7474
rect 10894 7198 10913 7250
rect 10913 7198 10946 7250
rect 12350 7441 12402 7474
rect 12350 7422 12402 7441
rect 11566 7198 11585 7250
rect 11585 7198 11618 7250
rect 12910 7319 12962 7362
rect 12910 7310 12949 7319
rect 12949 7310 12962 7319
rect 13806 7422 13858 7474
rect 14590 7422 14642 7474
rect 15262 7319 15314 7362
rect 15262 7310 15275 7319
rect 15275 7310 15314 7319
rect 16718 7694 16770 7698
rect 16718 7648 16737 7694
rect 16737 7648 16770 7694
rect 16718 7646 16770 7648
rect 15822 7441 15874 7474
rect 15822 7422 15874 7441
rect 16606 7422 16621 7474
rect 16621 7422 16658 7474
rect 17838 7694 17890 7698
rect 17838 7648 17857 7694
rect 17857 7648 17890 7694
rect 17838 7646 17890 7648
rect 17726 7422 17741 7474
rect 17741 7422 17778 7474
rect 3370 7030 3630 7082
rect 7682 7030 7942 7082
rect 11994 7030 12254 7082
rect 16306 7030 16566 7082
rect 2158 6862 2210 6914
rect 2494 6862 2546 6914
rect 2718 6638 2770 6690
rect 3278 6526 3330 6578
rect 3614 6414 3666 6466
rect 6862 6781 6868 6802
rect 6868 6781 6914 6802
rect 6862 6750 6914 6781
rect 7646 6862 7665 6914
rect 7665 6862 7698 6914
rect 7534 6555 7549 6578
rect 7549 6555 7586 6578
rect 7534 6526 7586 6555
rect 8318 6862 8337 6914
rect 8337 6862 8370 6914
rect 8206 6555 8221 6578
rect 8221 6555 8258 6578
rect 8206 6526 8258 6555
rect 8878 6555 8893 6578
rect 8893 6555 8930 6578
rect 8878 6526 8930 6555
rect 9550 6555 9565 6578
rect 9565 6555 9602 6578
rect 9550 6526 9602 6555
rect 8990 6464 9042 6466
rect 8990 6418 9009 6464
rect 9009 6418 9042 6464
rect 8990 6414 9042 6418
rect 10222 6555 10237 6578
rect 10237 6555 10274 6578
rect 10222 6526 10274 6555
rect 9662 6464 9714 6466
rect 9662 6418 9681 6464
rect 9681 6418 9714 6464
rect 9662 6414 9714 6418
rect 10894 6555 10909 6578
rect 10909 6555 10946 6578
rect 10894 6526 10946 6555
rect 10334 6464 10386 6466
rect 10334 6418 10353 6464
rect 10353 6418 10386 6464
rect 10334 6414 10386 6418
rect 11566 6555 11581 6578
rect 11581 6555 11618 6578
rect 11566 6526 11618 6555
rect 11006 6464 11058 6466
rect 11006 6418 11025 6464
rect 11025 6418 11058 6464
rect 11006 6414 11058 6418
rect 12238 6555 12253 6578
rect 12253 6555 12290 6578
rect 12238 6526 12290 6555
rect 11678 6464 11730 6466
rect 11678 6418 11697 6464
rect 11697 6418 11730 6464
rect 11678 6414 11730 6418
rect 12350 6464 12402 6466
rect 12350 6418 12369 6464
rect 12369 6418 12402 6464
rect 12350 6414 12402 6418
rect 13694 6638 13709 6690
rect 13709 6638 13746 6690
rect 14366 6638 14381 6690
rect 14381 6638 14418 6690
rect 13806 6464 13858 6466
rect 13806 6418 13825 6464
rect 13825 6418 13858 6464
rect 13806 6414 13858 6418
rect 15038 6638 15053 6690
rect 15053 6638 15090 6690
rect 14478 6464 14530 6466
rect 14478 6418 14497 6464
rect 14497 6418 14530 6464
rect 14478 6414 14530 6418
rect 15822 6862 15841 6914
rect 15841 6862 15874 6914
rect 15710 6638 15725 6690
rect 15725 6638 15762 6690
rect 15150 6464 15202 6466
rect 15150 6418 15169 6464
rect 15169 6418 15202 6464
rect 15150 6414 15202 6418
rect 16382 6555 16397 6578
rect 16397 6555 16434 6578
rect 16382 6526 16434 6555
rect 17054 6555 17069 6578
rect 17069 6555 17106 6578
rect 17054 6526 17106 6555
rect 16494 6464 16546 6466
rect 16494 6418 16513 6464
rect 16513 6418 16546 6464
rect 16494 6414 16546 6418
rect 17726 6555 17741 6578
rect 17741 6555 17778 6578
rect 17726 6526 17778 6555
rect 17166 6464 17218 6466
rect 17166 6418 17185 6464
rect 17185 6418 17218 6464
rect 17166 6414 17218 6418
rect 17838 6464 17890 6466
rect 17838 6418 17857 6464
rect 17857 6418 17890 6464
rect 17838 6414 17890 6418
rect 5526 6246 5786 6298
rect 9838 6246 10098 6298
rect 14150 6246 14410 6298
rect 18462 6246 18722 6298
rect 2382 6100 2434 6130
rect 2382 6078 2405 6100
rect 2405 6078 2434 6100
rect 1822 5742 1874 5794
rect 2046 5903 2098 5906
rect 2046 5857 2049 5903
rect 2049 5857 2095 5903
rect 2095 5857 2098 5903
rect 2046 5854 2098 5857
rect 3054 6126 3106 6130
rect 3054 6080 3073 6126
rect 3073 6080 3106 6126
rect 3054 6078 3106 6080
rect 2942 5854 2957 5906
rect 2957 5854 2994 5906
rect 6190 5854 6242 5906
rect 5630 5763 5682 5794
rect 5630 5742 5676 5763
rect 5676 5742 5682 5763
rect 6302 5989 6354 6018
rect 6302 5966 6339 5989
rect 6339 5966 6354 5989
rect 6862 5854 6914 5906
rect 6974 5854 7011 5906
rect 7011 5854 7026 5906
rect 7534 5854 7549 5906
rect 7549 5854 7586 5906
rect 8990 6126 9042 6130
rect 8990 6080 9009 6126
rect 9009 6080 9042 6126
rect 8990 6078 9042 6080
rect 8878 5989 8930 6018
rect 8878 5966 8893 5989
rect 8893 5966 8930 5989
rect 7646 5854 7698 5906
rect 8318 5630 8364 5682
rect 8364 5630 8370 5682
rect 10334 5854 10349 5906
rect 10349 5854 10386 5906
rect 11118 6126 11170 6130
rect 11118 6080 11137 6126
rect 11137 6080 11170 6126
rect 11118 6078 11170 6080
rect 11006 5854 11021 5906
rect 11021 5854 11058 5906
rect 10446 5630 10465 5682
rect 10465 5630 10498 5682
rect 11678 5854 11693 5906
rect 11693 5854 11730 5906
rect 12350 5854 12365 5906
rect 12365 5854 12402 5906
rect 11790 5630 11809 5682
rect 11809 5630 11842 5682
rect 13022 5854 13037 5906
rect 13037 5854 13074 5906
rect 12462 5630 12481 5682
rect 12481 5630 12514 5682
rect 13694 5989 13746 6018
rect 13694 5966 13709 5989
rect 13709 5966 13746 5989
rect 13134 5630 13153 5682
rect 13153 5630 13186 5682
rect 14478 6126 14530 6130
rect 14478 6080 14497 6126
rect 14497 6080 14530 6126
rect 14478 6078 14530 6080
rect 14366 5854 14381 5906
rect 14381 5854 14418 5906
rect 13806 5630 13825 5682
rect 13825 5630 13858 5682
rect 15038 5989 15090 6018
rect 15038 5966 15053 5989
rect 15053 5966 15090 5989
rect 15822 6126 15874 6130
rect 15822 6080 15841 6126
rect 15841 6080 15874 6126
rect 15822 6078 15874 6080
rect 15710 5854 15725 5906
rect 15725 5854 15762 5906
rect 15150 5630 15169 5682
rect 15169 5630 15202 5682
rect 16494 5763 16546 5794
rect 16494 5742 16540 5763
rect 16540 5742 16546 5763
rect 17726 5630 17732 5682
rect 17732 5630 17778 5682
rect 3370 5462 3630 5514
rect 7682 5462 7942 5514
rect 11994 5462 12254 5514
rect 16306 5462 16566 5514
rect 4286 5213 4332 5234
rect 4332 5213 4338 5234
rect 4286 5182 4338 5213
rect 4958 5294 5004 5346
rect 5004 5294 5010 5346
rect 6414 5294 6460 5346
rect 6460 5294 6466 5346
rect 6974 5294 6980 5346
rect 6980 5294 7026 5346
rect 8430 5213 8476 5234
rect 8476 5213 8482 5234
rect 8430 5182 8482 5213
rect 9102 5229 9121 5234
rect 9121 5229 9154 5234
rect 9102 5182 9154 5229
rect 7646 5070 7698 5122
rect 8990 5070 9005 5122
rect 9005 5070 9042 5122
rect 7758 4987 7795 5010
rect 7795 4987 7810 5010
rect 7758 4958 7810 4987
rect 9774 5229 9793 5234
rect 9793 5229 9826 5234
rect 9774 5182 9826 5229
rect 9662 5070 9677 5122
rect 9677 5070 9714 5122
rect 10446 5229 10465 5234
rect 10465 5229 10498 5234
rect 10446 5182 10498 5229
rect 10334 5070 10349 5122
rect 10349 5070 10386 5122
rect 11118 5229 11137 5234
rect 11137 5229 11170 5234
rect 11118 5182 11170 5229
rect 11006 5070 11021 5122
rect 11021 5070 11058 5122
rect 11678 5070 11693 5122
rect 11693 5070 11730 5122
rect 12350 5070 12365 5122
rect 12365 5070 12402 5122
rect 12462 5070 12514 5122
rect 11790 4896 11842 4898
rect 11790 4850 11809 4896
rect 11809 4850 11842 4896
rect 11790 4846 11842 4850
rect 13694 5070 13709 5122
rect 13709 5070 13746 5122
rect 14478 5229 14497 5234
rect 14497 5229 14530 5234
rect 14478 5182 14530 5229
rect 13806 5070 13858 5122
rect 14366 5070 14381 5122
rect 14381 5070 14418 5122
rect 15710 5213 15716 5234
rect 15716 5213 15762 5234
rect 15710 5182 15762 5213
rect 15150 5070 15187 5122
rect 15187 5070 15202 5122
rect 16382 5070 16434 5122
rect 15038 4896 15090 4898
rect 15038 4850 15071 4896
rect 15071 4850 15090 4896
rect 15038 4846 15090 4850
rect 17278 5070 17330 5122
rect 17838 5103 17890 5122
rect 17838 5070 17890 5103
rect 5526 4678 5786 4730
rect 9838 4678 10098 4730
rect 14150 4678 14410 4730
rect 18462 4678 18722 4730
rect 2718 4305 2770 4338
rect 2718 4286 2770 4305
rect 3502 4398 3554 4450
rect 4286 4286 4310 4338
rect 4310 4286 4338 4338
rect 7086 4286 7138 4338
rect 5294 4062 5340 4114
rect 5340 4062 5346 4114
rect 5966 4195 6018 4226
rect 5966 4174 6012 4195
rect 6012 4174 6018 4195
rect 6638 4195 6690 4226
rect 6638 4174 6684 4195
rect 6684 4174 6690 4195
rect 7982 4398 8034 4450
rect 8654 4305 8706 4338
rect 8654 4286 8706 4305
rect 10782 4558 10834 4562
rect 10782 4512 10815 4558
rect 10815 4512 10834 4558
rect 10782 4510 10834 4512
rect 10222 4062 10268 4114
rect 10268 4062 10274 4114
rect 11454 4558 11506 4562
rect 11454 4512 11487 4558
rect 11487 4512 11506 4558
rect 11454 4510 11506 4512
rect 10894 4421 10946 4450
rect 10894 4398 10931 4421
rect 10931 4398 10946 4421
rect 11566 4421 11618 4450
rect 11566 4398 11603 4421
rect 11603 4398 11618 4421
rect 12014 4286 12066 4338
rect 12910 4398 12962 4450
rect 15038 4558 15090 4562
rect 15038 4512 15057 4558
rect 15057 4512 15090 4558
rect 15038 4510 15090 4512
rect 14926 4421 14978 4450
rect 14926 4398 14941 4421
rect 14941 4398 14978 4421
rect 13470 4305 13522 4338
rect 13470 4286 13522 4305
rect 14478 4286 14530 4338
rect 14814 4286 14866 4338
rect 14366 4195 14418 4226
rect 14366 4174 14412 4195
rect 14412 4174 14418 4195
rect 15710 4558 15762 4562
rect 15710 4512 15729 4558
rect 15729 4512 15762 4558
rect 15710 4510 15762 4512
rect 15598 4286 15613 4338
rect 15613 4286 15650 4338
rect 16382 4558 16434 4562
rect 16382 4512 16401 4558
rect 16401 4512 16434 4558
rect 16382 4510 16434 4512
rect 16270 4421 16322 4450
rect 16270 4398 16285 4421
rect 16285 4398 16322 4421
rect 17838 4558 17890 4562
rect 17838 4512 17857 4558
rect 17857 4512 17890 4558
rect 17838 4510 17890 4512
rect 17726 4286 17741 4338
rect 17741 4286 17778 4338
rect 3370 3894 3630 3946
rect 7682 3894 7942 3946
rect 11994 3894 12254 3946
rect 16306 3894 16566 3946
rect 2158 3645 2204 3666
rect 2204 3645 2210 3666
rect 2158 3614 2210 3645
rect 2606 3502 2658 3554
rect 3502 3657 3515 3666
rect 3515 3657 3554 3666
rect 3502 3614 3554 3657
rect 4958 3645 5004 3666
rect 5004 3645 5010 3666
rect 4958 3614 5010 3645
rect 6078 3726 6124 3778
rect 6124 3726 6130 3778
rect 6750 3645 6796 3666
rect 6796 3645 6802 3666
rect 6750 3614 6802 3645
rect 4062 3535 4114 3554
rect 4062 3502 4114 3535
rect 7198 3502 7250 3554
rect 8094 3657 8107 3666
rect 8107 3657 8146 3666
rect 8094 3614 8146 3657
rect 9998 3726 10044 3778
rect 10044 3726 10050 3778
rect 10670 3726 10716 3778
rect 10716 3726 10722 3778
rect 8654 3535 8706 3554
rect 8654 3502 8706 3535
rect 11118 3502 11170 3554
rect 12014 3657 12027 3666
rect 12027 3657 12066 3666
rect 12014 3614 12066 3657
rect 12574 3535 12626 3554
rect 12574 3502 12626 3535
rect 14366 3726 14412 3778
rect 14412 3726 14418 3778
rect 13694 3502 13731 3554
rect 13731 3502 13746 3554
rect 13582 3328 13634 3330
rect 13582 3282 13615 3328
rect 13615 3282 13634 3328
rect 13582 3278 13634 3282
rect 15150 3502 15178 3554
rect 15178 3502 15202 3554
rect 15934 3657 15947 3666
rect 15947 3657 15986 3666
rect 15934 3614 15986 3657
rect 17502 3726 17508 3778
rect 17508 3726 17554 3778
rect 16718 3535 16770 3554
rect 16718 3502 16770 3535
rect 5526 3110 5786 3162
rect 9838 3110 10098 3162
rect 14150 3110 14410 3162
rect 18462 3110 18722 3162
<< metal2 >>
rect 2464 11200 2576 12000
rect 7392 11200 7504 12000
rect 12320 11200 12432 12000
rect 17248 11200 17360 12000
rect 2044 8372 2100 8382
rect 1820 8148 1876 8158
rect 1820 8054 1876 8092
rect 1932 8034 1988 8046
rect 1932 7982 1934 8034
rect 1986 7982 1988 8034
rect 1932 7924 1988 7982
rect 1932 7858 1988 7868
rect 1932 7700 1988 7710
rect 1932 7606 1988 7644
rect 1820 7474 1876 7486
rect 1820 7422 1822 7474
rect 1874 7422 1876 7474
rect 1820 6580 1876 7422
rect 1820 6514 1876 6524
rect 2044 7476 2100 8316
rect 2492 8258 2548 11200
rect 3368 8652 3632 8662
rect 3368 8586 3632 8596
rect 7420 8428 7476 11200
rect 7680 8652 7944 8662
rect 7680 8586 7944 8596
rect 11992 8652 12256 8662
rect 11992 8586 12256 8596
rect 7308 8372 7476 8428
rect 10556 8372 10612 8382
rect 2492 8206 2494 8258
rect 2546 8206 2548 8258
rect 2044 5906 2100 7420
rect 2156 8036 2212 8046
rect 2156 6914 2212 7980
rect 2492 7474 2548 8206
rect 4172 8258 4228 8270
rect 4172 8206 4174 8258
rect 4226 8206 4228 8258
rect 3276 8146 3332 8158
rect 3276 8094 3278 8146
rect 3330 8094 3332 8146
rect 3276 7700 3332 8094
rect 2492 7422 2494 7474
rect 2546 7422 2548 7474
rect 2492 7410 2548 7422
rect 3164 7644 3276 7700
rect 3052 7364 3108 7374
rect 2716 7252 2772 7262
rect 2156 6862 2158 6914
rect 2210 6862 2212 6914
rect 2156 6850 2212 6862
rect 2492 6916 2548 6926
rect 2492 6822 2548 6860
rect 2716 6690 2772 7196
rect 2716 6638 2718 6690
rect 2770 6638 2772 6690
rect 2716 6626 2772 6638
rect 3052 6916 3108 7308
rect 2380 6132 2436 6142
rect 2380 6038 2436 6076
rect 3052 6130 3108 6860
rect 3052 6078 3054 6130
rect 3106 6078 3108 6130
rect 3052 6066 3108 6078
rect 2044 5854 2046 5906
rect 2098 5854 2100 5906
rect 2044 5842 2100 5854
rect 2940 5906 2996 5918
rect 2940 5854 2942 5906
rect 2994 5854 2996 5906
rect 1820 5794 1876 5806
rect 1820 5742 1822 5794
rect 1874 5742 1876 5794
rect 1820 5012 1876 5742
rect 1820 2996 1876 4956
rect 2940 5012 2996 5854
rect 3164 5908 3220 7644
rect 3276 7634 3332 7644
rect 3388 7924 3444 7934
rect 3276 7476 3332 7486
rect 3388 7476 3444 7868
rect 3276 7474 3444 7476
rect 3276 7422 3278 7474
rect 3330 7422 3444 7474
rect 3276 7420 3444 7422
rect 3724 7924 3780 7934
rect 3276 7410 3332 7420
rect 3368 7084 3632 7094
rect 3368 7018 3632 7028
rect 3276 6580 3332 6590
rect 3276 6486 3332 6524
rect 3612 6466 3668 6478
rect 3612 6414 3614 6466
rect 3666 6414 3668 6466
rect 3612 6132 3668 6414
rect 3612 6066 3668 6076
rect 3164 5348 3220 5852
rect 3368 5516 3632 5526
rect 3368 5450 3632 5460
rect 3164 5292 3556 5348
rect 2940 4946 2996 4956
rect 3500 4450 3556 5292
rect 3500 4398 3502 4450
rect 3554 4398 3556 4450
rect 3500 4386 3556 4398
rect 2716 4338 2772 4350
rect 2716 4286 2718 4338
rect 2770 4286 2772 4338
rect 2156 3666 2212 3678
rect 2156 3614 2158 3666
rect 2210 3614 2212 3666
rect 2156 3556 2212 3614
rect 2604 3556 2660 3566
rect 2156 3554 2660 3556
rect 2156 3502 2606 3554
rect 2658 3502 2660 3554
rect 2156 3500 2660 3502
rect 2604 3490 2660 3500
rect 2716 3556 2772 4286
rect 3368 3948 3632 3958
rect 3368 3882 3632 3892
rect 3500 3668 3556 3678
rect 3724 3668 3780 7868
rect 4172 7474 4228 8206
rect 7308 8258 7364 8372
rect 10556 8370 10948 8372
rect 10556 8318 10558 8370
rect 10610 8318 10948 8370
rect 10556 8316 10948 8318
rect 10556 8306 10612 8316
rect 7308 8206 7310 8258
rect 7362 8206 7364 8258
rect 4620 8148 4676 8158
rect 4620 8054 4676 8092
rect 6748 8146 6804 8158
rect 6748 8094 6750 8146
rect 6802 8094 6804 8146
rect 4956 8036 5012 8046
rect 4956 7942 5012 7980
rect 6636 8036 6692 8046
rect 6636 7942 6692 7980
rect 5524 7868 5788 7878
rect 5524 7802 5788 7812
rect 4172 7422 4174 7474
rect 4226 7422 4228 7474
rect 4172 7364 4228 7422
rect 4732 7476 4788 7486
rect 4732 7382 4788 7420
rect 4172 7298 4228 7308
rect 6748 7364 6804 8094
rect 7308 7474 7364 8206
rect 8876 8258 8932 8270
rect 8876 8206 8878 8258
rect 8930 8206 8932 8258
rect 8092 8146 8148 8158
rect 8092 8094 8094 8146
rect 8146 8094 8148 8146
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 7308 7410 7364 7422
rect 7532 8036 7588 8046
rect 4620 7252 4676 7262
rect 4620 7158 4676 7196
rect 6300 6804 6356 6814
rect 4956 6692 5012 6702
rect 4956 5346 5012 6636
rect 5524 6300 5788 6310
rect 5524 6234 5788 6244
rect 6300 6018 6356 6748
rect 6748 6580 6804 7308
rect 7532 6916 7588 7980
rect 8092 8036 8148 8094
rect 8092 7970 8148 7980
rect 8876 7474 8932 8206
rect 9884 8260 9940 8270
rect 9884 8258 10388 8260
rect 9884 8206 9886 8258
rect 9938 8206 10388 8258
rect 9884 8204 10388 8206
rect 9884 8194 9940 8204
rect 10332 8148 10388 8204
rect 10668 8148 10724 8158
rect 10332 8146 10836 8148
rect 10332 8094 10670 8146
rect 10722 8094 10836 8146
rect 10332 8092 10836 8094
rect 10668 8082 10724 8092
rect 9996 8036 10052 8046
rect 9996 8034 10388 8036
rect 9996 7982 9998 8034
rect 10050 7982 10388 8034
rect 9996 7980 10388 7982
rect 9996 7970 10052 7980
rect 9836 7868 10100 7878
rect 9836 7802 10100 7812
rect 8876 7422 8878 7474
rect 8930 7422 8932 7474
rect 8092 7362 8148 7374
rect 8092 7310 8094 7362
rect 8146 7310 8148 7362
rect 7680 7084 7944 7094
rect 7680 7018 7944 7028
rect 7644 6916 7700 6926
rect 7532 6860 7644 6916
rect 6860 6804 6916 6814
rect 7644 6784 7700 6860
rect 6860 6710 6916 6748
rect 6748 6514 6804 6524
rect 7532 6580 7588 6590
rect 7532 6486 7588 6524
rect 6300 5966 6302 6018
rect 6354 5966 6356 6018
rect 6300 5954 6356 5966
rect 6188 5908 6244 5918
rect 6188 5814 6244 5852
rect 6860 5908 6916 5918
rect 6860 5814 6916 5852
rect 6972 5906 7028 5918
rect 6972 5854 6974 5906
rect 7026 5854 7028 5906
rect 5628 5796 5684 5806
rect 5628 5702 5684 5740
rect 4956 5294 4958 5346
rect 5010 5294 5012 5346
rect 4956 5282 5012 5294
rect 6412 5348 6468 5358
rect 6412 5254 6468 5292
rect 6972 5346 7028 5854
rect 6972 5294 6974 5346
rect 7026 5294 7028 5346
rect 6972 5282 7028 5294
rect 7420 5908 7476 5918
rect 4284 5234 4340 5246
rect 4284 5182 4286 5234
rect 4338 5182 4340 5234
rect 4284 4338 4340 5182
rect 7420 5124 7476 5852
rect 7532 5906 7588 5918
rect 7532 5854 7534 5906
rect 7586 5854 7588 5906
rect 7532 5348 7588 5854
rect 7644 5908 7700 5918
rect 7644 5814 7700 5852
rect 8092 5908 8148 7310
rect 8316 6916 8372 6926
rect 8204 6580 8260 6590
rect 8204 6486 8260 6524
rect 8316 6468 8372 6860
rect 8316 5908 8372 6412
rect 8876 6580 8932 7422
rect 10108 7474 10164 7486
rect 10108 7422 10110 7474
rect 10162 7422 10164 7474
rect 8876 6018 8932 6524
rect 9548 6580 9604 6590
rect 9548 6486 9604 6524
rect 10108 6580 10164 7422
rect 10220 7252 10276 7262
rect 10332 7252 10388 7980
rect 10220 7250 10388 7252
rect 10220 7198 10222 7250
rect 10274 7198 10388 7250
rect 10220 7196 10388 7198
rect 10220 7186 10276 7196
rect 10220 6580 10276 6590
rect 10164 6578 10276 6580
rect 10164 6526 10222 6578
rect 10274 6526 10276 6578
rect 10164 6524 10276 6526
rect 8988 6468 9044 6478
rect 8988 6132 9044 6412
rect 8988 6038 9044 6076
rect 9660 6466 9716 6478
rect 9660 6414 9662 6466
rect 9714 6414 9716 6466
rect 10108 6448 10164 6524
rect 9660 6132 9716 6414
rect 9836 6300 10100 6310
rect 9836 6234 10100 6244
rect 9660 6066 9716 6076
rect 8876 5966 8878 6018
rect 8930 5966 8932 6018
rect 8876 5954 8932 5966
rect 8092 5684 8148 5852
rect 8092 5618 8148 5628
rect 8204 5852 8372 5908
rect 10220 5908 10276 6524
rect 10332 6468 10388 7196
rect 10780 7474 10836 8092
rect 10780 7422 10782 7474
rect 10834 7422 10836 7474
rect 10780 6580 10836 7422
rect 10892 7252 10948 8316
rect 11340 8260 11396 8270
rect 12348 8260 12404 11200
rect 16304 8652 16568 8662
rect 16304 8586 16568 8596
rect 15260 8372 15316 8382
rect 12572 8260 12628 8270
rect 11340 8258 11508 8260
rect 11340 8206 11342 8258
rect 11394 8206 11508 8258
rect 11340 8204 11508 8206
rect 11340 8194 11396 8204
rect 11452 7474 11508 8204
rect 12348 8258 12628 8260
rect 12348 8206 12574 8258
rect 12626 8206 12628 8258
rect 12348 8204 12628 8206
rect 11452 7422 11454 7474
rect 11506 7422 11508 7474
rect 10892 7250 11172 7252
rect 10892 7198 10894 7250
rect 10946 7198 11172 7250
rect 10892 7196 11172 7198
rect 10892 7186 10948 7196
rect 10892 6580 10948 6590
rect 10780 6578 10948 6580
rect 10780 6526 10894 6578
rect 10946 6526 10948 6578
rect 10780 6524 10948 6526
rect 10332 6374 10388 6412
rect 10668 6020 10724 6030
rect 10332 5908 10388 5918
rect 10220 5852 10332 5908
rect 7680 5516 7944 5526
rect 7680 5450 7944 5460
rect 7532 5282 7588 5292
rect 7644 5124 7700 5134
rect 7420 5122 7700 5124
rect 7420 5070 7646 5122
rect 7698 5070 7700 5122
rect 7420 5068 7700 5070
rect 7644 4788 7700 5068
rect 7756 5012 7812 5022
rect 7756 5010 8148 5012
rect 7756 4958 7758 5010
rect 7810 4958 8148 5010
rect 7756 4956 8148 4958
rect 7756 4946 7812 4956
rect 5524 4732 5788 4742
rect 7644 4732 8036 4788
rect 5524 4666 5788 4676
rect 7980 4450 8036 4732
rect 7980 4398 7982 4450
rect 8034 4398 8036 4450
rect 7980 4386 8036 4398
rect 4284 4286 4286 4338
rect 4338 4286 4340 4338
rect 4284 4274 4340 4286
rect 5964 4340 6020 4350
rect 5964 4226 6020 4284
rect 7084 4340 7140 4350
rect 7084 4246 7140 4284
rect 5964 4174 5966 4226
rect 6018 4174 6020 4226
rect 5964 4162 6020 4174
rect 6636 4228 6692 4238
rect 6636 4134 6692 4172
rect 5292 4116 5348 4126
rect 5292 4022 5348 4060
rect 7680 3948 7944 3958
rect 7680 3882 7944 3892
rect 8092 3892 8148 4956
rect 8092 3826 8148 3836
rect 6076 3780 6132 3790
rect 6076 3686 6132 3724
rect 3500 3666 3780 3668
rect 3500 3614 3502 3666
rect 3554 3614 3780 3666
rect 3500 3612 3780 3614
rect 4956 3668 5012 3678
rect 3500 3602 3556 3612
rect 4956 3574 5012 3612
rect 6748 3666 6804 3678
rect 6748 3614 6750 3666
rect 6802 3614 6804 3666
rect 1820 2930 1876 2940
rect 2716 2660 2772 3500
rect 4060 3556 4116 3566
rect 4060 3462 4116 3500
rect 6748 3444 6804 3614
rect 7196 3668 7252 3678
rect 7196 3554 7252 3612
rect 8092 3668 8148 3678
rect 8204 3668 8260 5852
rect 8316 5682 8372 5694
rect 8316 5630 8318 5682
rect 8370 5630 8372 5682
rect 8316 5348 8372 5630
rect 8316 5282 8372 5292
rect 9100 5684 9156 5694
rect 8428 5236 8484 5246
rect 9100 5236 9156 5628
rect 8428 5234 9044 5236
rect 8428 5182 8430 5234
rect 8482 5182 9044 5234
rect 8428 5180 9044 5182
rect 8428 5170 8484 5180
rect 8988 5122 9044 5180
rect 9100 5142 9156 5180
rect 9772 5236 9828 5246
rect 9772 5142 9828 5180
rect 8988 5070 8990 5122
rect 9042 5070 9044 5122
rect 8988 5058 9044 5070
rect 9660 5124 9716 5134
rect 9660 5030 9716 5068
rect 10332 5124 10388 5852
rect 10444 5682 10500 5694
rect 10444 5630 10446 5682
rect 10498 5630 10500 5682
rect 10444 5236 10500 5630
rect 10444 5142 10500 5180
rect 10332 4992 10388 5068
rect 9836 4732 10100 4742
rect 9836 4666 10100 4676
rect 9996 4452 10052 4462
rect 8092 3666 8260 3668
rect 8092 3614 8094 3666
rect 8146 3614 8260 3666
rect 8092 3612 8260 3614
rect 8652 4338 8708 4350
rect 8652 4286 8654 4338
rect 8706 4286 8708 4338
rect 8092 3602 8148 3612
rect 7196 3502 7198 3554
rect 7250 3502 7252 3554
rect 7196 3490 7252 3502
rect 7420 3556 7476 3566
rect 6748 3378 6804 3388
rect 5524 3164 5788 3174
rect 5524 3098 5788 3108
rect 2492 2604 2772 2660
rect 2492 800 2548 2604
rect 7420 800 7476 3500
rect 8652 3556 8708 4286
rect 9884 4116 9940 4126
rect 9884 3668 9940 4060
rect 9996 3778 10052 4396
rect 10220 4116 10276 4126
rect 10220 4022 10276 4060
rect 9996 3726 9998 3778
rect 10050 3726 10052 3778
rect 9996 3714 10052 3726
rect 10668 3778 10724 5964
rect 10892 5908 10948 6524
rect 11004 6468 11060 6478
rect 11004 6374 11060 6412
rect 11116 6132 11172 7196
rect 11452 6580 11508 7422
rect 12012 8146 12068 8158
rect 12012 8094 12014 8146
rect 12066 8094 12068 8146
rect 11564 7252 11620 7262
rect 12012 7252 12068 8094
rect 12348 7474 12404 8204
rect 12572 8194 12628 8204
rect 14476 8258 14532 8270
rect 14476 8206 14478 8258
rect 14530 8206 14532 8258
rect 13692 8146 13748 8158
rect 13692 8094 13694 8146
rect 13746 8094 13748 8146
rect 12348 7422 12350 7474
rect 12402 7422 12404 7474
rect 12348 7410 12404 7422
rect 13580 8034 13636 8046
rect 13580 7982 13582 8034
rect 13634 7982 13636 8034
rect 12908 7364 12964 7374
rect 13580 7364 13636 7982
rect 13692 7476 13748 8094
rect 14148 7868 14412 7878
rect 14148 7802 14412 7812
rect 13804 7476 13860 7486
rect 13692 7420 13804 7476
rect 12908 7362 13636 7364
rect 12908 7310 12910 7362
rect 12962 7310 13636 7362
rect 12908 7308 13636 7310
rect 11564 7250 11732 7252
rect 11564 7198 11566 7250
rect 11618 7198 11732 7250
rect 11564 7196 11732 7198
rect 12012 7196 12404 7252
rect 11564 7186 11620 7196
rect 11564 6580 11620 6590
rect 11452 6578 11620 6580
rect 11452 6526 11566 6578
rect 11618 6526 11620 6578
rect 11452 6524 11620 6526
rect 11116 6038 11172 6076
rect 11004 5908 11060 5918
rect 10892 5852 11004 5908
rect 11564 5908 11620 6524
rect 11676 6468 11732 7196
rect 11992 7084 12256 7094
rect 11992 7018 12256 7028
rect 12236 6578 12292 6590
rect 12236 6526 12238 6578
rect 12290 6526 12292 6578
rect 11676 6466 11844 6468
rect 11676 6414 11678 6466
rect 11730 6414 11844 6466
rect 11676 6412 11844 6414
rect 11676 6402 11732 6412
rect 11788 6132 11844 6412
rect 11676 5908 11732 5918
rect 11564 5852 11676 5908
rect 10780 5236 10836 5246
rect 10780 4562 10836 5180
rect 10780 4510 10782 4562
rect 10834 4510 10836 4562
rect 10780 4498 10836 4510
rect 11004 5122 11060 5852
rect 11116 5236 11172 5246
rect 11116 5142 11172 5180
rect 11452 5236 11508 5246
rect 11004 5070 11006 5122
rect 11058 5070 11060 5122
rect 10892 4452 10948 4462
rect 11004 4452 11060 5070
rect 11452 4562 11508 5180
rect 11452 4510 11454 4562
rect 11506 4510 11508 4562
rect 11452 4498 11508 4510
rect 11676 5122 11732 5852
rect 11676 5070 11678 5122
rect 11730 5070 11732 5122
rect 10892 4450 11060 4452
rect 10892 4398 10894 4450
rect 10946 4398 11060 4450
rect 10892 4396 11060 4398
rect 11564 4452 11620 4462
rect 11676 4452 11732 5070
rect 11788 5682 11844 6076
rect 12236 5908 12292 6526
rect 12348 6468 12404 7196
rect 12404 6412 12516 6468
rect 12348 6336 12404 6412
rect 12348 5908 12404 5918
rect 12236 5852 12348 5908
rect 11788 5630 11790 5682
rect 11842 5630 11844 5682
rect 11788 5124 11844 5630
rect 11992 5516 12256 5526
rect 11992 5450 12256 5460
rect 11788 5058 11844 5068
rect 11900 5236 11956 5246
rect 11788 4900 11844 4910
rect 11900 4900 11956 5180
rect 12348 5122 12404 5852
rect 12460 5684 12516 6412
rect 12908 5684 12964 7308
rect 13692 6692 13748 6702
rect 13804 6692 13860 7420
rect 14476 7476 14532 8206
rect 15148 8146 15204 8158
rect 15148 8094 15150 8146
rect 15202 8094 15204 8146
rect 14588 7476 14644 7486
rect 14476 7420 14588 7476
rect 13692 6690 13860 6692
rect 13692 6638 13694 6690
rect 13746 6638 13860 6690
rect 13692 6636 13860 6638
rect 14364 6692 14420 6702
rect 14476 6692 14532 7420
rect 14588 7382 14644 7420
rect 14364 6690 14532 6692
rect 14364 6638 14366 6690
rect 14418 6638 14532 6690
rect 14364 6636 14532 6638
rect 15036 6804 15092 6814
rect 15036 6690 15092 6748
rect 15036 6638 15038 6690
rect 15090 6638 15092 6690
rect 13692 6018 13748 6636
rect 14364 6626 14420 6636
rect 14812 6580 14868 6590
rect 13692 5966 13694 6018
rect 13746 5966 13748 6018
rect 13020 5908 13076 5918
rect 13020 5814 13076 5852
rect 13692 5908 13748 5966
rect 13132 5684 13188 5694
rect 12460 5682 12628 5684
rect 12460 5630 12462 5682
rect 12514 5630 12628 5682
rect 12460 5628 12628 5630
rect 12908 5682 13188 5684
rect 12908 5630 13134 5682
rect 13186 5630 13188 5682
rect 12908 5628 13188 5630
rect 12460 5618 12516 5628
rect 12572 5236 12628 5628
rect 12572 5170 12628 5180
rect 12908 5236 12964 5246
rect 12348 5070 12350 5122
rect 12402 5070 12404 5122
rect 12348 5058 12404 5070
rect 12460 5124 12516 5134
rect 11788 4898 11956 4900
rect 11788 4846 11790 4898
rect 11842 4846 11956 4898
rect 11788 4844 11956 4846
rect 11788 4834 11844 4844
rect 11564 4450 11732 4452
rect 11564 4398 11566 4450
rect 11618 4398 11732 4450
rect 11564 4396 11732 4398
rect 10892 4386 10948 4396
rect 11564 4386 11620 4396
rect 12012 4340 12068 4350
rect 11788 4338 12068 4340
rect 11788 4286 12014 4338
rect 12066 4286 12068 4338
rect 11788 4284 12068 4286
rect 10668 3726 10670 3778
rect 10722 3726 10724 3778
rect 10668 3714 10724 3726
rect 11116 3780 11172 3790
rect 9884 3602 9940 3612
rect 8652 3424 8708 3500
rect 11116 3554 11172 3724
rect 11116 3502 11118 3554
rect 11170 3502 11172 3554
rect 11116 3490 11172 3502
rect 11788 3444 11844 4284
rect 12012 4274 12068 4284
rect 11992 3948 12256 3958
rect 11992 3882 12256 3892
rect 12460 3780 12516 5068
rect 12908 4450 12964 5180
rect 13132 5124 13188 5628
rect 13132 5058 13188 5068
rect 13580 5684 13636 5694
rect 12908 4398 12910 4450
rect 12962 4398 12964 4450
rect 12908 4386 12964 4398
rect 12012 3724 12516 3780
rect 12572 4340 12628 4350
rect 12012 3666 12068 3724
rect 12012 3614 12014 3666
rect 12066 3614 12068 3666
rect 12012 3602 12068 3614
rect 12572 3556 12628 4284
rect 13468 4340 13524 4350
rect 13468 4246 13524 4284
rect 11788 3378 11844 3388
rect 12348 3554 12628 3556
rect 12348 3502 12574 3554
rect 12626 3502 12628 3554
rect 12348 3500 12628 3502
rect 13580 3556 13636 5628
rect 13692 5122 13748 5852
rect 13804 6466 13860 6478
rect 13804 6414 13806 6466
rect 13858 6414 13860 6466
rect 13804 5684 13860 6414
rect 14476 6468 14532 6478
rect 14148 6300 14412 6310
rect 14148 6234 14412 6244
rect 14476 6130 14532 6412
rect 14476 6078 14478 6130
rect 14530 6078 14532 6130
rect 14476 6066 14532 6078
rect 14364 5908 14420 5918
rect 13804 5682 13972 5684
rect 13804 5630 13806 5682
rect 13858 5630 13972 5682
rect 13804 5628 13972 5630
rect 13804 5618 13860 5628
rect 13916 5236 13972 5628
rect 13916 5170 13972 5180
rect 13692 5070 13694 5122
rect 13746 5070 13748 5122
rect 13692 5058 13748 5070
rect 13804 5124 13860 5134
rect 13692 3556 13748 3566
rect 13580 3554 13748 3556
rect 13580 3502 13694 3554
rect 13746 3502 13748 3554
rect 13580 3500 13748 3502
rect 9836 3164 10100 3174
rect 9836 3098 10100 3108
rect 12348 800 12404 3500
rect 12572 3490 12628 3500
rect 13692 3490 13748 3500
rect 13580 3332 13636 3342
rect 13804 3332 13860 5068
rect 14364 5122 14420 5852
rect 14588 5908 14644 5918
rect 14476 5236 14532 5246
rect 14476 5142 14532 5180
rect 14364 5070 14366 5122
rect 14418 5070 14420 5122
rect 14364 5058 14420 5070
rect 14148 4732 14412 4742
rect 14148 4666 14412 4676
rect 14476 4338 14532 4350
rect 14476 4286 14478 4338
rect 14530 4286 14532 4338
rect 14364 4228 14420 4238
rect 14476 4228 14532 4286
rect 14364 4226 14532 4228
rect 14364 4174 14366 4226
rect 14418 4174 14532 4226
rect 14364 4172 14532 4174
rect 14364 4162 14420 4172
rect 14588 3892 14644 5852
rect 14812 4338 14868 6524
rect 15036 6018 15092 6638
rect 15148 6468 15204 8094
rect 15148 6374 15204 6412
rect 15260 7362 15316 8316
rect 15932 8372 15988 8382
rect 15820 8260 15876 8270
rect 15260 7310 15262 7362
rect 15314 7310 15316 7362
rect 15036 5966 15038 6018
rect 15090 5966 15092 6018
rect 15036 5954 15092 5966
rect 15148 5684 15204 5694
rect 15260 5684 15316 7310
rect 15708 7476 15764 7486
rect 15708 6804 15764 7420
rect 15820 7474 15876 8204
rect 15820 7422 15822 7474
rect 15874 7422 15876 7474
rect 15820 7410 15876 7422
rect 15820 6916 15876 6926
rect 15932 6916 15988 8316
rect 16604 8372 16660 8382
rect 16492 8148 16548 8158
rect 16492 7476 16548 8092
rect 16604 7700 16660 8316
rect 17276 8260 17332 11200
rect 17276 8194 17332 8204
rect 17836 8932 17892 8942
rect 17836 8484 17892 8876
rect 17500 8148 17556 8158
rect 17500 8054 17556 8092
rect 17612 8034 17668 8046
rect 17612 7982 17614 8034
rect 17666 7982 17668 8034
rect 16716 7700 16772 7710
rect 16604 7698 16772 7700
rect 16604 7646 16718 7698
rect 16770 7646 16772 7698
rect 16604 7644 16772 7646
rect 16716 7634 16772 7644
rect 17612 7588 17668 7982
rect 17836 7698 17892 8428
rect 18460 7868 18724 7878
rect 18460 7802 18724 7812
rect 17836 7646 17838 7698
rect 17890 7646 17892 7698
rect 17836 7634 17892 7646
rect 17500 7532 17668 7588
rect 16604 7476 16660 7486
rect 16548 7474 16660 7476
rect 16548 7422 16606 7474
rect 16658 7422 16660 7474
rect 16548 7420 16660 7422
rect 16492 7344 16548 7420
rect 16604 7410 16660 7420
rect 16304 7084 16568 7094
rect 16304 7018 16568 7028
rect 15820 6914 15988 6916
rect 15820 6862 15822 6914
rect 15874 6862 15988 6914
rect 15820 6860 15988 6862
rect 15820 6850 15876 6860
rect 15708 6690 15764 6748
rect 15708 6638 15710 6690
rect 15762 6638 15764 6690
rect 15708 6626 15764 6638
rect 16380 6580 16436 6590
rect 16380 6486 16436 6524
rect 17052 6578 17108 6590
rect 17052 6526 17054 6578
rect 17106 6526 17108 6578
rect 15820 6468 15876 6478
rect 15820 6130 15876 6412
rect 16492 6468 16548 6478
rect 16492 6374 16548 6412
rect 15820 6078 15822 6130
rect 15874 6078 15876 6130
rect 15708 5908 15764 5918
rect 15708 5814 15764 5852
rect 15148 5682 15316 5684
rect 15148 5630 15150 5682
rect 15202 5630 15316 5682
rect 15148 5628 15316 5630
rect 15148 5460 15204 5628
rect 15148 5394 15204 5404
rect 14924 5348 14980 5358
rect 14924 4450 14980 5292
rect 15708 5236 15764 5246
rect 15148 5234 15764 5236
rect 15148 5182 15710 5234
rect 15762 5182 15764 5234
rect 15148 5180 15764 5182
rect 15036 5124 15092 5134
rect 15036 4898 15092 5068
rect 15148 5122 15204 5180
rect 15708 5170 15764 5180
rect 15148 5070 15150 5122
rect 15202 5070 15204 5122
rect 15148 5058 15204 5070
rect 15036 4846 15038 4898
rect 15090 4846 15092 4898
rect 15036 4564 15092 4846
rect 15708 4564 15764 4574
rect 15820 4564 15876 6078
rect 16156 5796 16212 5806
rect 16156 5124 16212 5740
rect 16492 5796 16548 5806
rect 16492 5702 16548 5740
rect 17052 5796 17108 6526
rect 17164 6468 17220 6478
rect 17276 6468 17332 6478
rect 17164 6466 17276 6468
rect 17164 6414 17166 6466
rect 17218 6414 17276 6466
rect 17164 6412 17276 6414
rect 17164 6402 17220 6412
rect 17052 5730 17108 5740
rect 16304 5516 16568 5526
rect 16304 5450 16568 5460
rect 16380 5124 16436 5134
rect 16156 5122 16436 5124
rect 16156 5070 16382 5122
rect 16434 5070 16436 5122
rect 16156 5068 16436 5070
rect 16380 5058 16436 5068
rect 16492 5124 16548 5134
rect 15036 4562 15876 4564
rect 15036 4510 15038 4562
rect 15090 4510 15710 4562
rect 15762 4510 15876 4562
rect 15036 4508 15876 4510
rect 16380 4564 16436 4574
rect 16492 4564 16548 5068
rect 17276 5122 17332 6412
rect 17500 6468 17556 7532
rect 17724 7476 17780 7486
rect 17612 7474 17780 7476
rect 17612 7422 17726 7474
rect 17778 7422 17780 7474
rect 17612 7420 17780 7422
rect 17612 6692 17668 7420
rect 17724 7410 17780 7420
rect 17612 6626 17668 6636
rect 17500 6402 17556 6412
rect 17724 6578 17780 6590
rect 17724 6526 17726 6578
rect 17778 6526 17780 6578
rect 17724 6020 17780 6526
rect 17836 6468 17892 6478
rect 17836 6374 17892 6412
rect 18460 6300 18724 6310
rect 18460 6234 18724 6244
rect 17724 5954 17780 5964
rect 17724 5684 17780 5694
rect 17724 5590 17780 5628
rect 17276 5070 17278 5122
rect 17330 5070 17332 5122
rect 16380 4562 16548 4564
rect 16380 4510 16382 4562
rect 16434 4510 16548 4562
rect 16380 4508 16548 4510
rect 16828 5012 16884 5022
rect 15036 4498 15092 4508
rect 15708 4498 15764 4508
rect 14924 4398 14926 4450
rect 14978 4398 14980 4450
rect 14924 4386 14980 4398
rect 16268 4452 16324 4462
rect 16268 4358 16324 4396
rect 14812 4286 14814 4338
rect 14866 4286 14868 4338
rect 14812 4274 14868 4286
rect 15596 4338 15652 4350
rect 15596 4286 15598 4338
rect 15650 4286 15652 4338
rect 15596 4116 15652 4286
rect 16380 4116 16436 4508
rect 15596 4050 15652 4060
rect 15932 4060 16436 4116
rect 14364 3836 14644 3892
rect 14364 3778 14420 3836
rect 14364 3726 14366 3778
rect 14418 3726 14420 3778
rect 14364 3714 14420 3726
rect 15148 3668 15204 3678
rect 15148 3554 15204 3612
rect 15932 3666 15988 4060
rect 16304 3948 16568 3958
rect 16304 3882 16568 3892
rect 15932 3614 15934 3666
rect 15986 3614 15988 3666
rect 15932 3602 15988 3614
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3490 15204 3502
rect 16716 3556 16772 3566
rect 16828 3556 16884 4956
rect 16716 3554 16884 3556
rect 16716 3502 16718 3554
rect 16770 3502 16884 3554
rect 16716 3500 16884 3502
rect 16716 3490 16772 3500
rect 13580 3330 13860 3332
rect 13580 3278 13582 3330
rect 13634 3278 13860 3330
rect 13580 3276 13860 3278
rect 13580 3266 13636 3276
rect 14148 3164 14412 3174
rect 14148 3098 14412 3108
rect 16828 2772 16884 3500
rect 17276 2996 17332 5070
rect 17724 5124 17780 5134
rect 17724 4788 17780 5068
rect 17836 5122 17892 5134
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5012 17892 5070
rect 17836 4946 17892 4956
rect 17724 4732 17892 4788
rect 17836 4562 17892 4732
rect 18460 4732 18724 4742
rect 18460 4666 18724 4676
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 17724 4338 17780 4350
rect 17724 4286 17726 4338
rect 17778 4286 17780 4338
rect 17724 4228 17780 4286
rect 17724 4162 17780 4172
rect 17500 3780 17556 3790
rect 17500 3686 17556 3724
rect 18460 3164 18724 3174
rect 18460 3098 18724 3108
rect 17276 2930 17332 2940
rect 16828 2716 17332 2772
rect 17276 800 17332 2716
rect 2464 0 2576 800
rect 7392 0 7504 800
rect 12320 0 12432 800
rect 17248 0 17360 800
<< via2 >>
rect 2044 8316 2100 8372
rect 1820 8146 1876 8148
rect 1820 8094 1822 8146
rect 1822 8094 1874 8146
rect 1874 8094 1876 8146
rect 1820 8092 1876 8094
rect 1932 7868 1988 7924
rect 1932 7698 1988 7700
rect 1932 7646 1934 7698
rect 1934 7646 1986 7698
rect 1986 7646 1988 7698
rect 1932 7644 1988 7646
rect 1820 6524 1876 6580
rect 3368 8650 3632 8652
rect 3368 8598 3370 8650
rect 3370 8598 3630 8650
rect 3630 8598 3632 8650
rect 3368 8596 3632 8598
rect 7680 8650 7944 8652
rect 7680 8598 7682 8650
rect 7682 8598 7942 8650
rect 7942 8598 7944 8650
rect 7680 8596 7944 8598
rect 11992 8650 12256 8652
rect 11992 8598 11994 8650
rect 11994 8598 12254 8650
rect 12254 8598 12256 8650
rect 11992 8596 12256 8598
rect 2044 7420 2100 7476
rect 2156 7980 2212 8036
rect 3276 7644 3332 7700
rect 3052 7308 3108 7364
rect 2716 7196 2772 7252
rect 2492 6914 2548 6916
rect 2492 6862 2494 6914
rect 2494 6862 2546 6914
rect 2546 6862 2548 6914
rect 2492 6860 2548 6862
rect 3052 6860 3108 6916
rect 2380 6130 2436 6132
rect 2380 6078 2382 6130
rect 2382 6078 2434 6130
rect 2434 6078 2436 6130
rect 2380 6076 2436 6078
rect 1820 4956 1876 5012
rect 3388 7868 3444 7924
rect 3724 7868 3780 7924
rect 3368 7082 3632 7084
rect 3368 7030 3370 7082
rect 3370 7030 3630 7082
rect 3630 7030 3632 7082
rect 3368 7028 3632 7030
rect 3276 6578 3332 6580
rect 3276 6526 3278 6578
rect 3278 6526 3330 6578
rect 3330 6526 3332 6578
rect 3276 6524 3332 6526
rect 3612 6076 3668 6132
rect 3164 5852 3220 5908
rect 3368 5514 3632 5516
rect 3368 5462 3370 5514
rect 3370 5462 3630 5514
rect 3630 5462 3632 5514
rect 3368 5460 3632 5462
rect 2940 4956 2996 5012
rect 3368 3946 3632 3948
rect 3368 3894 3370 3946
rect 3370 3894 3630 3946
rect 3630 3894 3632 3946
rect 3368 3892 3632 3894
rect 4620 8146 4676 8148
rect 4620 8094 4622 8146
rect 4622 8094 4674 8146
rect 4674 8094 4676 8146
rect 4620 8092 4676 8094
rect 4956 8034 5012 8036
rect 4956 7982 4958 8034
rect 4958 7982 5010 8034
rect 5010 7982 5012 8034
rect 4956 7980 5012 7982
rect 6636 8034 6692 8036
rect 6636 7982 6638 8034
rect 6638 7982 6690 8034
rect 6690 7982 6692 8034
rect 6636 7980 6692 7982
rect 5524 7866 5788 7868
rect 5524 7814 5526 7866
rect 5526 7814 5786 7866
rect 5786 7814 5788 7866
rect 5524 7812 5788 7814
rect 4732 7474 4788 7476
rect 4732 7422 4734 7474
rect 4734 7422 4786 7474
rect 4786 7422 4788 7474
rect 4732 7420 4788 7422
rect 4172 7308 4228 7364
rect 7532 7980 7588 8036
rect 6748 7308 6804 7364
rect 4620 7250 4676 7252
rect 4620 7198 4622 7250
rect 4622 7198 4674 7250
rect 4674 7198 4676 7250
rect 4620 7196 4676 7198
rect 6300 6748 6356 6804
rect 4956 6636 5012 6692
rect 5524 6298 5788 6300
rect 5524 6246 5526 6298
rect 5526 6246 5786 6298
rect 5786 6246 5788 6298
rect 5524 6244 5788 6246
rect 8092 7980 8148 8036
rect 9836 7866 10100 7868
rect 9836 7814 9838 7866
rect 9838 7814 10098 7866
rect 10098 7814 10100 7866
rect 9836 7812 10100 7814
rect 7680 7082 7944 7084
rect 7680 7030 7682 7082
rect 7682 7030 7942 7082
rect 7942 7030 7944 7082
rect 7680 7028 7944 7030
rect 7644 6914 7700 6916
rect 7644 6862 7646 6914
rect 7646 6862 7698 6914
rect 7698 6862 7700 6914
rect 7644 6860 7700 6862
rect 6860 6802 6916 6804
rect 6860 6750 6862 6802
rect 6862 6750 6914 6802
rect 6914 6750 6916 6802
rect 6860 6748 6916 6750
rect 6748 6524 6804 6580
rect 7532 6578 7588 6580
rect 7532 6526 7534 6578
rect 7534 6526 7586 6578
rect 7586 6526 7588 6578
rect 7532 6524 7588 6526
rect 6188 5906 6244 5908
rect 6188 5854 6190 5906
rect 6190 5854 6242 5906
rect 6242 5854 6244 5906
rect 6188 5852 6244 5854
rect 6860 5906 6916 5908
rect 6860 5854 6862 5906
rect 6862 5854 6914 5906
rect 6914 5854 6916 5906
rect 6860 5852 6916 5854
rect 5628 5794 5684 5796
rect 5628 5742 5630 5794
rect 5630 5742 5682 5794
rect 5682 5742 5684 5794
rect 5628 5740 5684 5742
rect 6412 5346 6468 5348
rect 6412 5294 6414 5346
rect 6414 5294 6466 5346
rect 6466 5294 6468 5346
rect 6412 5292 6468 5294
rect 7420 5852 7476 5908
rect 7644 5906 7700 5908
rect 7644 5854 7646 5906
rect 7646 5854 7698 5906
rect 7698 5854 7700 5906
rect 7644 5852 7700 5854
rect 8316 6914 8372 6916
rect 8316 6862 8318 6914
rect 8318 6862 8370 6914
rect 8370 6862 8372 6914
rect 8316 6860 8372 6862
rect 8204 6578 8260 6580
rect 8204 6526 8206 6578
rect 8206 6526 8258 6578
rect 8258 6526 8260 6578
rect 8204 6524 8260 6526
rect 8316 6412 8372 6468
rect 8876 6578 8932 6580
rect 8876 6526 8878 6578
rect 8878 6526 8930 6578
rect 8930 6526 8932 6578
rect 8876 6524 8932 6526
rect 9548 6578 9604 6580
rect 9548 6526 9550 6578
rect 9550 6526 9602 6578
rect 9602 6526 9604 6578
rect 9548 6524 9604 6526
rect 10108 6524 10164 6580
rect 8988 6466 9044 6468
rect 8988 6414 8990 6466
rect 8990 6414 9042 6466
rect 9042 6414 9044 6466
rect 8988 6412 9044 6414
rect 8988 6130 9044 6132
rect 8988 6078 8990 6130
rect 8990 6078 9042 6130
rect 9042 6078 9044 6130
rect 8988 6076 9044 6078
rect 9836 6298 10100 6300
rect 9836 6246 9838 6298
rect 9838 6246 10098 6298
rect 10098 6246 10100 6298
rect 9836 6244 10100 6246
rect 9660 6076 9716 6132
rect 8092 5852 8148 5908
rect 8092 5628 8148 5684
rect 16304 8650 16568 8652
rect 16304 8598 16306 8650
rect 16306 8598 16566 8650
rect 16566 8598 16568 8650
rect 16304 8596 16568 8598
rect 15260 8316 15316 8372
rect 10332 6466 10388 6468
rect 10332 6414 10334 6466
rect 10334 6414 10386 6466
rect 10386 6414 10388 6466
rect 10332 6412 10388 6414
rect 10668 5964 10724 6020
rect 10332 5906 10388 5908
rect 10332 5854 10334 5906
rect 10334 5854 10386 5906
rect 10386 5854 10388 5906
rect 10332 5852 10388 5854
rect 7680 5514 7944 5516
rect 7680 5462 7682 5514
rect 7682 5462 7942 5514
rect 7942 5462 7944 5514
rect 7680 5460 7944 5462
rect 7532 5292 7588 5348
rect 5524 4730 5788 4732
rect 5524 4678 5526 4730
rect 5526 4678 5786 4730
rect 5786 4678 5788 4730
rect 5524 4676 5788 4678
rect 5964 4284 6020 4340
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 6636 4226 6692 4228
rect 6636 4174 6638 4226
rect 6638 4174 6690 4226
rect 6690 4174 6692 4226
rect 6636 4172 6692 4174
rect 5292 4114 5348 4116
rect 5292 4062 5294 4114
rect 5294 4062 5346 4114
rect 5346 4062 5348 4114
rect 5292 4060 5348 4062
rect 7680 3946 7944 3948
rect 7680 3894 7682 3946
rect 7682 3894 7942 3946
rect 7942 3894 7944 3946
rect 7680 3892 7944 3894
rect 8092 3836 8148 3892
rect 6076 3778 6132 3780
rect 6076 3726 6078 3778
rect 6078 3726 6130 3778
rect 6130 3726 6132 3778
rect 6076 3724 6132 3726
rect 4956 3666 5012 3668
rect 4956 3614 4958 3666
rect 4958 3614 5010 3666
rect 5010 3614 5012 3666
rect 4956 3612 5012 3614
rect 2716 3500 2772 3556
rect 1820 2940 1876 2996
rect 4060 3554 4116 3556
rect 4060 3502 4062 3554
rect 4062 3502 4114 3554
rect 4114 3502 4116 3554
rect 4060 3500 4116 3502
rect 7196 3612 7252 3668
rect 8316 5292 8372 5348
rect 9100 5628 9156 5684
rect 9100 5234 9156 5236
rect 9100 5182 9102 5234
rect 9102 5182 9154 5234
rect 9154 5182 9156 5234
rect 9100 5180 9156 5182
rect 9772 5234 9828 5236
rect 9772 5182 9774 5234
rect 9774 5182 9826 5234
rect 9826 5182 9828 5234
rect 9772 5180 9828 5182
rect 9660 5122 9716 5124
rect 9660 5070 9662 5122
rect 9662 5070 9714 5122
rect 9714 5070 9716 5122
rect 9660 5068 9716 5070
rect 10444 5234 10500 5236
rect 10444 5182 10446 5234
rect 10446 5182 10498 5234
rect 10498 5182 10500 5234
rect 10444 5180 10500 5182
rect 10332 5122 10388 5124
rect 10332 5070 10334 5122
rect 10334 5070 10386 5122
rect 10386 5070 10388 5122
rect 10332 5068 10388 5070
rect 9836 4730 10100 4732
rect 9836 4678 9838 4730
rect 9838 4678 10098 4730
rect 10098 4678 10100 4730
rect 9836 4676 10100 4678
rect 9996 4396 10052 4452
rect 7420 3500 7476 3556
rect 6748 3388 6804 3444
rect 5524 3162 5788 3164
rect 5524 3110 5526 3162
rect 5526 3110 5786 3162
rect 5786 3110 5788 3162
rect 5524 3108 5788 3110
rect 9884 4060 9940 4116
rect 10220 4114 10276 4116
rect 10220 4062 10222 4114
rect 10222 4062 10274 4114
rect 10274 4062 10276 4114
rect 10220 4060 10276 4062
rect 11004 6466 11060 6468
rect 11004 6414 11006 6466
rect 11006 6414 11058 6466
rect 11058 6414 11060 6466
rect 11004 6412 11060 6414
rect 14148 7866 14412 7868
rect 14148 7814 14150 7866
rect 14150 7814 14410 7866
rect 14410 7814 14412 7866
rect 14148 7812 14412 7814
rect 13804 7474 13860 7476
rect 13804 7422 13806 7474
rect 13806 7422 13858 7474
rect 13858 7422 13860 7474
rect 13804 7420 13860 7422
rect 11116 6130 11172 6132
rect 11116 6078 11118 6130
rect 11118 6078 11170 6130
rect 11170 6078 11172 6130
rect 11116 6076 11172 6078
rect 11004 5906 11060 5908
rect 11004 5854 11006 5906
rect 11006 5854 11058 5906
rect 11058 5854 11060 5906
rect 11004 5852 11060 5854
rect 11992 7082 12256 7084
rect 11992 7030 11994 7082
rect 11994 7030 12254 7082
rect 12254 7030 12256 7082
rect 11992 7028 12256 7030
rect 11788 6076 11844 6132
rect 11676 5906 11732 5908
rect 11676 5854 11678 5906
rect 11678 5854 11730 5906
rect 11730 5854 11732 5906
rect 11676 5852 11732 5854
rect 10780 5180 10836 5236
rect 11116 5234 11172 5236
rect 11116 5182 11118 5234
rect 11118 5182 11170 5234
rect 11170 5182 11172 5234
rect 11116 5180 11172 5182
rect 11452 5180 11508 5236
rect 12348 6466 12404 6468
rect 12348 6414 12350 6466
rect 12350 6414 12402 6466
rect 12402 6414 12404 6466
rect 12348 6412 12404 6414
rect 12348 5906 12404 5908
rect 12348 5854 12350 5906
rect 12350 5854 12402 5906
rect 12402 5854 12404 5906
rect 12348 5852 12404 5854
rect 11992 5514 12256 5516
rect 11992 5462 11994 5514
rect 11994 5462 12254 5514
rect 12254 5462 12256 5514
rect 11992 5460 12256 5462
rect 11788 5068 11844 5124
rect 11900 5180 11956 5236
rect 14588 7474 14644 7476
rect 14588 7422 14590 7474
rect 14590 7422 14642 7474
rect 14642 7422 14644 7474
rect 14588 7420 14644 7422
rect 15036 6748 15092 6804
rect 14812 6524 14868 6580
rect 13020 5906 13076 5908
rect 13020 5854 13022 5906
rect 13022 5854 13074 5906
rect 13074 5854 13076 5906
rect 13020 5852 13076 5854
rect 13692 5852 13748 5908
rect 12572 5180 12628 5236
rect 12908 5180 12964 5236
rect 12460 5122 12516 5124
rect 12460 5070 12462 5122
rect 12462 5070 12514 5122
rect 12514 5070 12516 5122
rect 12460 5068 12516 5070
rect 11116 3724 11172 3780
rect 9884 3612 9940 3668
rect 8652 3554 8708 3556
rect 8652 3502 8654 3554
rect 8654 3502 8706 3554
rect 8706 3502 8708 3554
rect 8652 3500 8708 3502
rect 11992 3946 12256 3948
rect 11992 3894 11994 3946
rect 11994 3894 12254 3946
rect 12254 3894 12256 3946
rect 11992 3892 12256 3894
rect 13132 5068 13188 5124
rect 13580 5628 13636 5684
rect 12572 4284 12628 4340
rect 13468 4338 13524 4340
rect 13468 4286 13470 4338
rect 13470 4286 13522 4338
rect 13522 4286 13524 4338
rect 13468 4284 13524 4286
rect 11788 3388 11844 3444
rect 14476 6466 14532 6468
rect 14476 6414 14478 6466
rect 14478 6414 14530 6466
rect 14530 6414 14532 6466
rect 14476 6412 14532 6414
rect 14148 6298 14412 6300
rect 14148 6246 14150 6298
rect 14150 6246 14410 6298
rect 14410 6246 14412 6298
rect 14148 6244 14412 6246
rect 14364 5906 14420 5908
rect 14364 5854 14366 5906
rect 14366 5854 14418 5906
rect 14418 5854 14420 5906
rect 14364 5852 14420 5854
rect 13916 5180 13972 5236
rect 13804 5122 13860 5124
rect 13804 5070 13806 5122
rect 13806 5070 13858 5122
rect 13858 5070 13860 5122
rect 13804 5068 13860 5070
rect 9836 3162 10100 3164
rect 9836 3110 9838 3162
rect 9838 3110 10098 3162
rect 10098 3110 10100 3162
rect 9836 3108 10100 3110
rect 14588 5852 14644 5908
rect 14476 5234 14532 5236
rect 14476 5182 14478 5234
rect 14478 5182 14530 5234
rect 14530 5182 14532 5234
rect 14476 5180 14532 5182
rect 14148 4730 14412 4732
rect 14148 4678 14150 4730
rect 14150 4678 14410 4730
rect 14410 4678 14412 4730
rect 14148 4676 14412 4678
rect 15148 6466 15204 6468
rect 15148 6414 15150 6466
rect 15150 6414 15202 6466
rect 15202 6414 15204 6466
rect 15148 6412 15204 6414
rect 15932 8316 15988 8372
rect 15820 8258 15876 8260
rect 15820 8206 15822 8258
rect 15822 8206 15874 8258
rect 15874 8206 15876 8258
rect 15820 8204 15876 8206
rect 15708 7420 15764 7476
rect 16604 8370 16660 8372
rect 16604 8318 16606 8370
rect 16606 8318 16658 8370
rect 16658 8318 16660 8370
rect 16604 8316 16660 8318
rect 16492 8146 16548 8148
rect 16492 8094 16494 8146
rect 16494 8094 16546 8146
rect 16546 8094 16548 8146
rect 16492 8092 16548 8094
rect 17276 8204 17332 8260
rect 17836 8876 17892 8932
rect 17836 8428 17892 8484
rect 17500 8146 17556 8148
rect 17500 8094 17502 8146
rect 17502 8094 17554 8146
rect 17554 8094 17556 8146
rect 17500 8092 17556 8094
rect 18460 7866 18724 7868
rect 18460 7814 18462 7866
rect 18462 7814 18722 7866
rect 18722 7814 18724 7866
rect 18460 7812 18724 7814
rect 16492 7420 16548 7476
rect 16304 7082 16568 7084
rect 16304 7030 16306 7082
rect 16306 7030 16566 7082
rect 16566 7030 16568 7082
rect 16304 7028 16568 7030
rect 15708 6748 15764 6804
rect 16380 6578 16436 6580
rect 16380 6526 16382 6578
rect 16382 6526 16434 6578
rect 16434 6526 16436 6578
rect 16380 6524 16436 6526
rect 15820 6412 15876 6468
rect 16492 6466 16548 6468
rect 16492 6414 16494 6466
rect 16494 6414 16546 6466
rect 16546 6414 16548 6466
rect 16492 6412 16548 6414
rect 15708 5906 15764 5908
rect 15708 5854 15710 5906
rect 15710 5854 15762 5906
rect 15762 5854 15764 5906
rect 15708 5852 15764 5854
rect 15148 5404 15204 5460
rect 14924 5292 14980 5348
rect 15036 5068 15092 5124
rect 16156 5740 16212 5796
rect 16492 5794 16548 5796
rect 16492 5742 16494 5794
rect 16494 5742 16546 5794
rect 16546 5742 16548 5794
rect 16492 5740 16548 5742
rect 17276 6412 17332 6468
rect 17052 5740 17108 5796
rect 16304 5514 16568 5516
rect 16304 5462 16306 5514
rect 16306 5462 16566 5514
rect 16566 5462 16568 5514
rect 16304 5460 16568 5462
rect 16492 5068 16548 5124
rect 17612 6636 17668 6692
rect 17500 6412 17556 6468
rect 17836 6466 17892 6468
rect 17836 6414 17838 6466
rect 17838 6414 17890 6466
rect 17890 6414 17892 6466
rect 17836 6412 17892 6414
rect 18460 6298 18724 6300
rect 18460 6246 18462 6298
rect 18462 6246 18722 6298
rect 18722 6246 18724 6298
rect 18460 6244 18724 6246
rect 17724 5964 17780 6020
rect 17724 5682 17780 5684
rect 17724 5630 17726 5682
rect 17726 5630 17778 5682
rect 17778 5630 17780 5682
rect 17724 5628 17780 5630
rect 16828 4956 16884 5012
rect 16268 4450 16324 4452
rect 16268 4398 16270 4450
rect 16270 4398 16322 4450
rect 16322 4398 16324 4450
rect 16268 4396 16324 4398
rect 15596 4060 15652 4116
rect 15148 3612 15204 3668
rect 16304 3946 16568 3948
rect 16304 3894 16306 3946
rect 16306 3894 16566 3946
rect 16566 3894 16568 3946
rect 16304 3892 16568 3894
rect 14148 3162 14412 3164
rect 14148 3110 14150 3162
rect 14150 3110 14410 3162
rect 14410 3110 14412 3162
rect 14148 3108 14412 3110
rect 17724 5068 17780 5124
rect 17836 4956 17892 5012
rect 18460 4730 18724 4732
rect 18460 4678 18462 4730
rect 18462 4678 18722 4730
rect 18722 4678 18724 4730
rect 18460 4676 18724 4678
rect 17724 4172 17780 4228
rect 17500 3778 17556 3780
rect 17500 3726 17502 3778
rect 17502 3726 17554 3778
rect 17554 3726 17556 3778
rect 17500 3724 17556 3726
rect 18460 3162 18724 3164
rect 18460 3110 18462 3162
rect 18462 3110 18722 3162
rect 18722 3110 18724 3162
rect 18460 3108 18724 3110
rect 17276 2940 17332 2996
<< metal3 >>
rect 0 8932 800 8960
rect 19200 8932 20000 8960
rect 0 8876 2100 8932
rect 17826 8876 17836 8932
rect 17892 8876 20000 8932
rect 0 8848 800 8876
rect 2044 8372 2100 8876
rect 19200 8848 20000 8876
rect 3358 8596 3368 8652
rect 3632 8596 3642 8652
rect 7670 8596 7680 8652
rect 7944 8596 7954 8652
rect 11982 8596 11992 8652
rect 12256 8596 12266 8652
rect 16294 8596 16304 8652
rect 16568 8596 16578 8652
rect 15260 8428 17836 8484
rect 17892 8428 17902 8484
rect 15260 8372 15316 8428
rect 15820 8372 15876 8428
rect 16716 8372 16772 8428
rect 2034 8316 2044 8372
rect 2100 8316 2110 8372
rect 15250 8316 15260 8372
rect 15316 8316 15326 8372
rect 15820 8316 15932 8372
rect 15988 8316 15998 8372
rect 16594 8316 16604 8372
rect 16660 8316 16772 8372
rect 15810 8204 15820 8260
rect 15876 8204 17276 8260
rect 17332 8204 17342 8260
rect 1810 8092 1820 8148
rect 1876 8092 4620 8148
rect 4676 8092 4686 8148
rect 16482 8092 16492 8148
rect 16548 8092 17500 8148
rect 17556 8092 17566 8148
rect 2146 7980 2156 8036
rect 2212 7980 4956 8036
rect 5012 7980 5022 8036
rect 5292 7980 6636 8036
rect 6692 7980 7532 8036
rect 7588 7980 8092 8036
rect 8148 7980 8158 8036
rect 5292 7924 5348 7980
rect 1922 7868 1932 7924
rect 1988 7868 3388 7924
rect 3444 7868 3724 7924
rect 3780 7868 5348 7924
rect 5514 7812 5524 7868
rect 5788 7812 5798 7868
rect 9826 7812 9836 7868
rect 10100 7812 10110 7868
rect 14138 7812 14148 7868
rect 14412 7812 14422 7868
rect 18450 7812 18460 7868
rect 18724 7812 18734 7868
rect 1922 7644 1932 7700
rect 1988 7644 3276 7700
rect 3332 7644 3342 7700
rect 2034 7420 2044 7476
rect 2100 7420 4732 7476
rect 4788 7420 4798 7476
rect 13794 7420 13804 7476
rect 13860 7420 14588 7476
rect 14644 7420 15708 7476
rect 15764 7420 16492 7476
rect 16548 7420 16558 7476
rect 3042 7308 3052 7364
rect 3108 7308 4172 7364
rect 4228 7308 6748 7364
rect 6804 7308 6814 7364
rect 2706 7196 2716 7252
rect 2772 7196 4620 7252
rect 4676 7196 4686 7252
rect 3358 7028 3368 7084
rect 3632 7028 3642 7084
rect 7670 7028 7680 7084
rect 7944 7028 7954 7084
rect 11982 7028 11992 7084
rect 12256 7028 12266 7084
rect 16294 7028 16304 7084
rect 16568 7028 16578 7084
rect 2482 6860 2492 6916
rect 2548 6860 3052 6916
rect 3108 6860 3118 6916
rect 7634 6860 7644 6916
rect 7700 6860 8316 6916
rect 8372 6860 8382 6916
rect 6290 6748 6300 6804
rect 6356 6748 6860 6804
rect 6916 6748 6926 6804
rect 15026 6748 15036 6804
rect 15092 6748 15708 6804
rect 15764 6748 15774 6804
rect 4946 6636 4956 6692
rect 5012 6636 17612 6692
rect 17668 6636 17678 6692
rect 1810 6524 1820 6580
rect 1876 6524 3276 6580
rect 3332 6524 3342 6580
rect 6738 6524 6748 6580
rect 6804 6524 7532 6580
rect 7588 6524 8204 6580
rect 8260 6524 8876 6580
rect 8932 6524 9548 6580
rect 9604 6524 10108 6580
rect 10164 6524 10174 6580
rect 14802 6524 14812 6580
rect 14868 6524 16380 6580
rect 16436 6524 16446 6580
rect 8306 6412 8316 6468
rect 8372 6412 8988 6468
rect 9044 6412 9054 6468
rect 10322 6412 10332 6468
rect 10388 6412 11004 6468
rect 11060 6412 12348 6468
rect 12404 6412 12414 6468
rect 14466 6412 14476 6468
rect 14532 6412 15148 6468
rect 15204 6412 15820 6468
rect 15876 6412 16492 6468
rect 16548 6412 17276 6468
rect 17332 6412 17500 6468
rect 17556 6412 17836 6468
rect 17892 6412 17902 6468
rect 5514 6244 5524 6300
rect 5788 6244 5798 6300
rect 9826 6244 9836 6300
rect 10100 6244 10110 6300
rect 14138 6244 14148 6300
rect 14412 6244 14422 6300
rect 18450 6244 18460 6300
rect 18724 6244 18734 6300
rect 2370 6076 2380 6132
rect 2436 6076 3612 6132
rect 3668 6076 3678 6132
rect 8978 6076 8988 6132
rect 9044 6076 9660 6132
rect 9716 6076 11116 6132
rect 11172 6076 11788 6132
rect 11844 6076 11854 6132
rect 10658 5964 10668 6020
rect 10724 5964 17724 6020
rect 17780 5964 17790 6020
rect 3154 5852 3164 5908
rect 3220 5852 6188 5908
rect 6244 5852 6860 5908
rect 6916 5852 7420 5908
rect 7476 5852 7644 5908
rect 7700 5852 8092 5908
rect 8148 5852 8158 5908
rect 10322 5852 10332 5908
rect 10388 5852 11004 5908
rect 11060 5852 11676 5908
rect 11732 5852 12348 5908
rect 12404 5852 13020 5908
rect 13076 5852 13692 5908
rect 13748 5852 14364 5908
rect 14420 5852 14430 5908
rect 14578 5852 14588 5908
rect 14644 5852 15708 5908
rect 15764 5852 15774 5908
rect 5618 5740 5628 5796
rect 5684 5740 16156 5796
rect 16212 5740 16222 5796
rect 16482 5740 16492 5796
rect 16548 5740 17052 5796
rect 17108 5740 17118 5796
rect 8082 5628 8092 5684
rect 8148 5628 9100 5684
rect 9156 5628 9166 5684
rect 13570 5628 13580 5684
rect 13636 5628 17724 5684
rect 17780 5628 17790 5684
rect 3358 5460 3368 5516
rect 3632 5460 3642 5516
rect 7670 5460 7680 5516
rect 7944 5460 7954 5516
rect 11982 5460 11992 5516
rect 12256 5460 12266 5516
rect 16294 5460 16304 5516
rect 16568 5460 16578 5516
rect 15138 5404 15148 5460
rect 15204 5404 15214 5460
rect 6402 5292 6412 5348
rect 6468 5292 7532 5348
rect 7588 5292 7598 5348
rect 8306 5292 8316 5348
rect 8372 5292 14924 5348
rect 14980 5292 14990 5348
rect 15148 5236 15204 5404
rect 9090 5180 9100 5236
rect 9156 5180 9772 5236
rect 9828 5180 10444 5236
rect 10500 5180 10780 5236
rect 10836 5180 11116 5236
rect 11172 5180 11452 5236
rect 11508 5180 11900 5236
rect 11956 5180 12572 5236
rect 12628 5180 12908 5236
rect 12964 5180 13916 5236
rect 13972 5180 14476 5236
rect 14532 5180 16548 5236
rect 16492 5124 16548 5180
rect 9650 5068 9660 5124
rect 9716 5068 10332 5124
rect 10388 5068 10398 5124
rect 11778 5068 11788 5124
rect 11844 5068 12460 5124
rect 12516 5068 13132 5124
rect 13188 5068 13804 5124
rect 13860 5068 15036 5124
rect 15092 5068 15102 5124
rect 16482 5068 16492 5124
rect 16548 5068 17724 5124
rect 17780 5068 17790 5124
rect 1810 4956 1820 5012
rect 1876 4956 2940 5012
rect 2996 4956 3006 5012
rect 16818 4956 16828 5012
rect 16884 4956 17836 5012
rect 17892 4956 17902 5012
rect 5514 4676 5524 4732
rect 5788 4676 5798 4732
rect 9826 4676 9836 4732
rect 10100 4676 10110 4732
rect 14138 4676 14148 4732
rect 14412 4676 14422 4732
rect 18450 4676 18460 4732
rect 18724 4676 18734 4732
rect 9986 4396 9996 4452
rect 10052 4396 16268 4452
rect 16324 4396 16334 4452
rect 5954 4284 5964 4340
rect 6020 4284 7084 4340
rect 7140 4284 7150 4340
rect 12562 4284 12572 4340
rect 12628 4284 13468 4340
rect 13524 4284 13534 4340
rect 6626 4172 6636 4228
rect 6692 4172 17724 4228
rect 17780 4172 17790 4228
rect 5282 4060 5292 4116
rect 5348 4060 9884 4116
rect 9940 4060 9950 4116
rect 10210 4060 10220 4116
rect 10276 4060 15596 4116
rect 15652 4060 15662 4116
rect 8372 3948 11844 4004
rect 3358 3892 3368 3948
rect 3632 3892 3642 3948
rect 7670 3892 7680 3948
rect 7944 3892 7954 3948
rect 8372 3892 8428 3948
rect 8082 3836 8092 3892
rect 8148 3836 8428 3892
rect 11788 3780 11844 3948
rect 11982 3892 11992 3948
rect 12256 3892 12266 3948
rect 16294 3892 16304 3948
rect 16568 3892 16578 3948
rect 6066 3724 6076 3780
rect 6132 3724 11116 3780
rect 11172 3724 11182 3780
rect 11788 3724 17500 3780
rect 17556 3724 17566 3780
rect 4946 3612 4956 3668
rect 5012 3612 7196 3668
rect 7252 3612 7262 3668
rect 9874 3612 9884 3668
rect 9940 3612 15148 3668
rect 15204 3612 15214 3668
rect 2706 3500 2716 3556
rect 2772 3500 4060 3556
rect 4116 3500 4126 3556
rect 7410 3500 7420 3556
rect 7476 3500 8652 3556
rect 8708 3500 8718 3556
rect 6738 3388 6748 3444
rect 6804 3388 11788 3444
rect 11844 3388 11854 3444
rect 5514 3108 5524 3164
rect 5788 3108 5798 3164
rect 9826 3108 9836 3164
rect 10100 3108 10110 3164
rect 14138 3108 14148 3164
rect 14412 3108 14422 3164
rect 18450 3108 18460 3164
rect 18724 3108 18734 3164
rect 0 2996 800 3024
rect 19200 2996 20000 3024
rect 0 2940 1820 2996
rect 1876 2940 1886 2996
rect 17266 2940 17276 2996
rect 17332 2940 20000 2996
rect 0 2912 800 2940
rect 19200 2912 20000 2940
<< via3 >>
rect 3368 8596 3632 8652
rect 7680 8596 7944 8652
rect 11992 8596 12256 8652
rect 16304 8596 16568 8652
rect 5524 7812 5788 7868
rect 9836 7812 10100 7868
rect 14148 7812 14412 7868
rect 18460 7812 18724 7868
rect 3368 7028 3632 7084
rect 7680 7028 7944 7084
rect 11992 7028 12256 7084
rect 16304 7028 16568 7084
rect 5524 6244 5788 6300
rect 9836 6244 10100 6300
rect 14148 6244 14412 6300
rect 18460 6244 18724 6300
rect 3368 5460 3632 5516
rect 7680 5460 7944 5516
rect 11992 5460 12256 5516
rect 16304 5460 16568 5516
rect 5524 4676 5788 4732
rect 9836 4676 10100 4732
rect 14148 4676 14412 4732
rect 18460 4676 18724 4732
rect 3368 3892 3632 3948
rect 7680 3892 7944 3948
rect 11992 3892 12256 3948
rect 16304 3892 16568 3948
rect 5524 3108 5788 3164
rect 9836 3108 10100 3164
rect 14148 3108 14412 3164
rect 18460 3108 18724 3164
<< metal4 >>
rect 3340 8652 3660 8684
rect 3340 8596 3368 8652
rect 3632 8596 3660 8652
rect 3340 7084 3660 8596
rect 3340 7028 3368 7084
rect 3632 7028 3660 7084
rect 3340 5516 3660 7028
rect 3340 5460 3368 5516
rect 3632 5460 3660 5516
rect 3340 3948 3660 5460
rect 3340 3892 3368 3948
rect 3632 3892 3660 3948
rect 3340 3076 3660 3892
rect 5496 7868 5816 8684
rect 5496 7812 5524 7868
rect 5788 7812 5816 7868
rect 5496 6300 5816 7812
rect 5496 6244 5524 6300
rect 5788 6244 5816 6300
rect 5496 4732 5816 6244
rect 5496 4676 5524 4732
rect 5788 4676 5816 4732
rect 5496 3164 5816 4676
rect 5496 3108 5524 3164
rect 5788 3108 5816 3164
rect 5496 3076 5816 3108
rect 7652 8652 7972 8684
rect 7652 8596 7680 8652
rect 7944 8596 7972 8652
rect 7652 7084 7972 8596
rect 7652 7028 7680 7084
rect 7944 7028 7972 7084
rect 7652 5516 7972 7028
rect 7652 5460 7680 5516
rect 7944 5460 7972 5516
rect 7652 3948 7972 5460
rect 7652 3892 7680 3948
rect 7944 3892 7972 3948
rect 7652 3076 7972 3892
rect 9808 7868 10128 8684
rect 9808 7812 9836 7868
rect 10100 7812 10128 7868
rect 9808 6300 10128 7812
rect 9808 6244 9836 6300
rect 10100 6244 10128 6300
rect 9808 4732 10128 6244
rect 9808 4676 9836 4732
rect 10100 4676 10128 4732
rect 9808 3164 10128 4676
rect 9808 3108 9836 3164
rect 10100 3108 10128 3164
rect 9808 3076 10128 3108
rect 11964 8652 12284 8684
rect 11964 8596 11992 8652
rect 12256 8596 12284 8652
rect 11964 7084 12284 8596
rect 11964 7028 11992 7084
rect 12256 7028 12284 7084
rect 11964 5516 12284 7028
rect 11964 5460 11992 5516
rect 12256 5460 12284 5516
rect 11964 3948 12284 5460
rect 11964 3892 11992 3948
rect 12256 3892 12284 3948
rect 11964 3076 12284 3892
rect 14120 7868 14440 8684
rect 14120 7812 14148 7868
rect 14412 7812 14440 7868
rect 14120 6300 14440 7812
rect 14120 6244 14148 6300
rect 14412 6244 14440 6300
rect 14120 4732 14440 6244
rect 14120 4676 14148 4732
rect 14412 4676 14440 4732
rect 14120 3164 14440 4676
rect 14120 3108 14148 3164
rect 14412 3108 14440 3164
rect 14120 3076 14440 3108
rect 16276 8652 16596 8684
rect 16276 8596 16304 8652
rect 16568 8596 16596 8652
rect 16276 7084 16596 8596
rect 16276 7028 16304 7084
rect 16568 7028 16596 7084
rect 16276 5516 16596 7028
rect 16276 5460 16304 5516
rect 16568 5460 16596 5516
rect 16276 3948 16596 5460
rect 16276 3892 16304 3948
rect 16568 3892 16596 3948
rect 16276 3076 16596 3892
rect 18432 7868 18752 8684
rect 18432 7812 18460 7868
rect 18724 7812 18752 7868
rect 18432 6300 18752 7812
rect 18432 6244 18460 6300
rect 18724 6244 18752 6300
rect 18432 4732 18752 6244
rect 18432 4676 18460 4732
rect 18724 4676 18752 4732
rect 18432 3164 18752 4676
rect 18432 3108 18460 3164
rect 18724 3108 18752 3164
rect 18432 3076 18752 3108
<< labels >>
rlabel metal1 s 9968 8624 9968 8624 4 vdd
rlabel metal2 s 10048 7840 10048 7840 4 vss
rlabel metal3 s 7896 6552 7896 6552 4 _00_
rlabel metal3 s 3248 8120 3248 8120 4 _01_
rlabel metal3 s 2576 6552 2576 6552 4 _02_
rlabel metal3 s 3024 6104 3024 6104 4 _03_
rlabel metal2 s 2184 7448 2184 7448 4 _04_
rlabel metal2 s 10024 4088 10024 4088 4 _05_
rlabel metal2 s 14448 4200 14448 4200 4 _06_
rlabel metal2 s 8120 4424 8120 4424 4 _07_
rlabel metal2 s 8344 5488 8344 5488 4 _08_
rlabel metal3 s 7000 5320 7000 5320 4 _09_
rlabel metal3 s 12936 4088 12936 4088 4 _10_
rlabel metal2 s 7000 5600 7000 5600 4 _11_
rlabel metal3 s 16800 5768 16800 5768 4 _12_
rlabel metal2 s 9016 5152 9016 5152 4 _13_
rlabel metal2 s 15176 5152 15176 5152 4 _14_
rlabel metal2 s 6328 6384 6328 6384 4 _15_
rlabel metal2 s 10696 4872 10696 4872 4 _16_
rlabel metal2 s 4984 5992 4984 5992 4 _17_
rlabel metal2 s 14392 3808 14392 3808 4 _18_
rlabel metal2 s 17752 4256 17752 4256 4 _19_
rlabel metal2 s 13664 3528 13664 3528 4 _20_
rlabel metal2 s 4312 4760 4312 4760 4 _21_
rlabel metal2 s 2184 3584 2184 3584 4 _22_
rlabel metal2 s 5992 4256 5992 4256 4 _23_
rlabel metal3 s 6104 3640 6104 3640 4 _24_
rlabel metal2 s 6776 3528 6776 3528 4 _25_
rlabel metal2 s 11144 3640 11144 3640 4 _26_
rlabel metal2 s 9912 3864 9912 3864 4 _27_
rlabel metal2 s 16184 5432 16184 5432 4 _28_
rlabel metal2 s 1848 4368 1848 4368 4 enable
rlabel metal2 s 3304 7896 3304 7896 4 outn
rlabel metal2 s 3360 7448 3360 7448 4 outp
rlabel metal2 s 2072 7112 2072 7112 4 signal
rlabel metal2 s 2744 6944 2744 6944 4 signal_n
rlabel metal2 s 2744 3472 2744 3472 4 trim_n[0]
rlabel metal2 s 7448 2142 7448 2142 4 trim_n[1]
rlabel metal2 s 12488 3528 12488 3528 4 trim_n[2]
rlabel metal2 s 16800 3528 16800 3528 4 trim_n[3]
rlabel metal2 s 2520 7840 2520 7840 4 trim_p[0]
rlabel metal2 s 7336 7840 7336 7840 4 trim_p[1]
rlabel metal2 s 12488 8232 12488 8232 4 trim_p[2]
rlabel metal3 s 16576 8232 16576 8232 4 trim_p[3]
flabel metal3 s 0 2912 800 3024 0 FreeSans 560 0 0 0 enable
port 1 nsew
flabel metal3 s 19200 8848 20000 8960 0 FreeSans 560 0 0 0 outn
port 2 nsew
flabel metal3 s 19200 2912 20000 3024 0 FreeSans 560 0 0 0 outp
port 3 nsew
flabel metal3 s 0 8848 800 8960 0 FreeSans 560 0 0 0 signal
port 4 nsew
flabel metal2 s 2464 0 2576 800 0 FreeSans 560 90 0 0 trim_n[0]
port 5 nsew
flabel metal2 s 7392 0 7504 800 0 FreeSans 560 90 0 0 trim_n[1]
port 6 nsew
flabel metal2 s 12320 0 12432 800 0 FreeSans 560 90 0 0 trim_n[2]
port 7 nsew
flabel metal2 s 17248 0 17360 800 0 FreeSans 560 90 0 0 trim_n[3]
port 8 nsew
flabel metal2 s 2464 11200 2576 12000 0 FreeSans 560 90 0 0 trim_p[0]
port 9 nsew
flabel metal2 s 7392 11200 7504 12000 0 FreeSans 560 90 0 0 trim_p[1]
port 10 nsew
flabel metal2 s 12320 11200 12432 12000 0 FreeSans 560 90 0 0 trim_p[2]
port 11 nsew
flabel metal2 s 17248 11200 17360 12000 0 FreeSans 560 90 0 0 trim_p[3]
port 12 nsew
flabel metal4 s 3340 3076 3660 8684 0 FreeSans 1600 90 0 0 vdd
port 13 nsew
flabel metal4 s 7652 3076 7972 8684 0 FreeSans 1600 90 0 0 vdd
port 13 nsew
flabel metal4 s 11964 3076 12284 8684 0 FreeSans 1600 90 0 0 vdd
port 13 nsew
flabel metal4 s 16276 3076 16596 8684 0 FreeSans 1600 90 0 0 vdd
port 13 nsew
flabel metal4 s 5496 3076 5816 8684 0 FreeSans 1600 90 0 0 vss
port 14 nsew
flabel metal4 s 9808 3076 10128 8684 0 FreeSans 1600 90 0 0 vss
port 14 nsew
flabel metal4 s 14120 3076 14440 8684 0 FreeSans 1600 90 0 0 vss
port 14 nsew
flabel metal4 s 18432 3076 18752 8684 0 FreeSans 1600 90 0 0 vss
port 14 nsew
<< end >>