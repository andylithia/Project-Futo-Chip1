magic
tech gf180mcuC
magscale 1 5
timestamp 1669701303
<< metal1 >>
rect 672 4325 9296 4342
rect 672 4299 1685 4325
rect 1711 4299 1737 4325
rect 1763 4299 1789 4325
rect 1815 4299 3841 4325
rect 3867 4299 3893 4325
rect 3919 4299 3945 4325
rect 3971 4299 5997 4325
rect 6023 4299 6049 4325
rect 6075 4299 6101 4325
rect 6127 4299 8153 4325
rect 8179 4299 8205 4325
rect 8231 4299 8257 4325
rect 8283 4299 9296 4325
rect 672 4282 9296 4299
rect 8079 4129 8105 4135
rect 8079 4097 8105 4103
rect 8695 4129 8721 4135
rect 8695 4097 8721 4103
rect 8863 4129 8889 4135
rect 8863 4097 8889 4103
rect 8975 4129 9001 4135
rect 8975 4097 9001 4103
rect 1191 4073 1217 4079
rect 1191 4041 1217 4047
rect 1303 4073 1329 4079
rect 1303 4041 1329 4047
rect 1471 4073 1497 4079
rect 1471 4041 1497 4047
rect 1751 4073 1777 4079
rect 1751 4041 1777 4047
rect 1919 4073 1945 4079
rect 1919 4041 1945 4047
rect 2031 4073 2057 4079
rect 2031 4041 2057 4047
rect 7911 4073 7937 4079
rect 7911 4041 7937 4047
rect 8191 4073 8217 4079
rect 8191 4041 8217 4047
rect 672 3933 9376 3950
rect 672 3907 2763 3933
rect 2789 3907 2815 3933
rect 2841 3907 2867 3933
rect 2893 3907 4919 3933
rect 4945 3907 4971 3933
rect 4997 3907 5023 3933
rect 5049 3907 7075 3933
rect 7101 3907 7127 3933
rect 7153 3907 7179 3933
rect 7205 3907 9231 3933
rect 9257 3907 9283 3933
rect 9309 3907 9335 3933
rect 9361 3907 9376 3933
rect 672 3890 9376 3907
rect 1191 3793 1217 3799
rect 1191 3761 1217 3767
rect 1359 3737 1385 3743
rect 1359 3705 1385 3711
rect 1471 3737 1497 3743
rect 1471 3705 1497 3711
rect 1751 3737 1777 3743
rect 1751 3705 1777 3711
rect 1863 3737 1889 3743
rect 1863 3705 1889 3711
rect 1975 3737 2001 3743
rect 1975 3705 2001 3711
rect 2311 3737 2337 3743
rect 2311 3705 2337 3711
rect 2423 3737 2449 3743
rect 2423 3705 2449 3711
rect 2535 3737 2561 3743
rect 2535 3705 2561 3711
rect 7239 3737 7265 3743
rect 7239 3705 7265 3711
rect 7351 3737 7377 3743
rect 7351 3705 7377 3711
rect 7519 3737 7545 3743
rect 7519 3705 7545 3711
rect 7799 3737 7825 3743
rect 7799 3705 7825 3711
rect 7911 3737 7937 3743
rect 7911 3705 7937 3711
rect 8023 3737 8049 3743
rect 8023 3705 8049 3711
rect 672 3541 9296 3558
rect 672 3515 1685 3541
rect 1711 3515 1737 3541
rect 1763 3515 1789 3541
rect 1815 3515 3841 3541
rect 3867 3515 3893 3541
rect 3919 3515 3945 3541
rect 3971 3515 5997 3541
rect 6023 3515 6049 3541
rect 6075 3515 6101 3541
rect 6127 3515 8153 3541
rect 8179 3515 8205 3541
rect 8231 3515 8257 3541
rect 8283 3515 9296 3541
rect 672 3498 9296 3515
rect 1079 3345 1105 3351
rect 1079 3313 1105 3319
rect 1639 3345 1665 3351
rect 1639 3313 1665 3319
rect 1975 3345 2001 3351
rect 1975 3313 2001 3319
rect 2199 3345 2225 3351
rect 2199 3313 2225 3319
rect 2367 3345 2393 3351
rect 2367 3313 2393 3319
rect 3487 3345 3513 3351
rect 3487 3313 3513 3319
rect 3599 3345 3625 3351
rect 3599 3313 3625 3319
rect 7071 3345 7097 3351
rect 7071 3313 7097 3319
rect 7183 3345 7209 3351
rect 7183 3313 7209 3319
rect 7351 3345 7377 3351
rect 7351 3313 7377 3319
rect 7855 3345 7881 3351
rect 7855 3313 7881 3319
rect 8247 3345 8273 3351
rect 8247 3313 8273 3319
rect 8415 3345 8441 3351
rect 8415 3313 8441 3319
rect 8975 3345 9001 3351
rect 8975 3313 9001 3319
rect 1191 3289 1217 3295
rect 1191 3257 1217 3263
rect 1359 3289 1385 3295
rect 1359 3257 1385 3263
rect 1751 3289 1777 3295
rect 1751 3257 1777 3263
rect 2479 3289 2505 3295
rect 2479 3257 2505 3263
rect 3375 3289 3401 3295
rect 3375 3257 3401 3263
rect 7575 3289 7601 3295
rect 7575 3257 7601 3263
rect 7743 3289 7769 3295
rect 7743 3257 7769 3263
rect 8135 3289 8161 3295
rect 8135 3257 8161 3263
rect 8695 3289 8721 3295
rect 8695 3257 8721 3263
rect 8863 3289 8889 3295
rect 8863 3257 8889 3263
rect 672 3149 9376 3166
rect 672 3123 2763 3149
rect 2789 3123 2815 3149
rect 2841 3123 2867 3149
rect 2893 3123 4919 3149
rect 4945 3123 4971 3149
rect 4997 3123 5023 3149
rect 5049 3123 7075 3149
rect 7101 3123 7127 3149
rect 7153 3123 7179 3149
rect 7205 3123 9231 3149
rect 9257 3123 9283 3149
rect 9309 3123 9335 3149
rect 9361 3123 9376 3149
rect 672 3106 9376 3123
rect 1415 3009 1441 3015
rect 1415 2977 1441 2983
rect 1975 3009 2001 3015
rect 1975 2977 2001 2983
rect 2535 3009 2561 3015
rect 2535 2977 2561 2983
rect 4495 3009 4521 3015
rect 4495 2977 4521 2983
rect 7015 3009 7041 3015
rect 7015 2977 7041 2983
rect 7575 3009 7601 3015
rect 7575 2977 7601 2983
rect 8135 3009 8161 3015
rect 8135 2977 8161 2983
rect 1583 2953 1609 2959
rect 1583 2921 1609 2927
rect 1751 2953 1777 2959
rect 1751 2921 1777 2927
rect 2143 2953 2169 2959
rect 2143 2921 2169 2927
rect 2255 2953 2281 2959
rect 2255 2921 2281 2927
rect 2703 2953 2729 2959
rect 2703 2921 2729 2927
rect 2871 2953 2897 2959
rect 2871 2921 2897 2927
rect 3095 2953 3121 2959
rect 3095 2921 3121 2927
rect 3263 2953 3289 2959
rect 3263 2921 3289 2927
rect 3375 2953 3401 2959
rect 3375 2921 3401 2927
rect 3655 2953 3681 2959
rect 3655 2921 3681 2927
rect 3823 2953 3849 2959
rect 3823 2921 3849 2927
rect 3991 2953 4017 2959
rect 3991 2921 4017 2927
rect 4215 2953 4241 2959
rect 4215 2921 4241 2927
rect 4383 2953 4409 2959
rect 4383 2921 4409 2927
rect 4831 2953 4857 2959
rect 4831 2921 4857 2927
rect 4999 2953 5025 2959
rect 4999 2921 5025 2927
rect 5167 2953 5193 2959
rect 5167 2921 5193 2927
rect 6735 2953 6761 2959
rect 6735 2921 6761 2927
rect 6847 2953 6873 2959
rect 6847 2921 6873 2927
rect 7239 2953 7265 2959
rect 7239 2921 7265 2927
rect 7407 2953 7433 2959
rect 7407 2921 7433 2927
rect 7799 2953 7825 2959
rect 7799 2921 7825 2927
rect 7967 2953 7993 2959
rect 7967 2921 7993 2927
rect 672 2757 9296 2774
rect 672 2731 1685 2757
rect 1711 2731 1737 2757
rect 1763 2731 1789 2757
rect 1815 2731 3841 2757
rect 3867 2731 3893 2757
rect 3919 2731 3945 2757
rect 3971 2731 5997 2757
rect 6023 2731 6049 2757
rect 6075 2731 6101 2757
rect 6127 2731 8153 2757
rect 8179 2731 8205 2757
rect 8231 2731 8257 2757
rect 8283 2731 9296 2757
rect 672 2714 9296 2731
rect 1079 2561 1105 2567
rect 1079 2529 1105 2535
rect 1639 2561 1665 2567
rect 1639 2529 1665 2535
rect 2199 2561 2225 2567
rect 2199 2529 2225 2535
rect 3039 2561 3065 2567
rect 3039 2529 3065 2535
rect 3599 2561 3625 2567
rect 3599 2529 3625 2535
rect 4215 2561 4241 2567
rect 4215 2529 4241 2535
rect 7071 2561 7097 2567
rect 7071 2529 7097 2535
rect 7687 2561 7713 2567
rect 7687 2529 7713 2535
rect 8247 2561 8273 2567
rect 8247 2529 8273 2535
rect 8751 2561 8777 2567
rect 8751 2529 8777 2535
rect 1191 2505 1217 2511
rect 1191 2473 1217 2479
rect 1359 2505 1385 2511
rect 1359 2473 1385 2479
rect 1751 2505 1777 2511
rect 1751 2473 1777 2479
rect 1919 2505 1945 2511
rect 1919 2473 1945 2479
rect 2311 2505 2337 2511
rect 2311 2473 2337 2479
rect 2479 2505 2505 2511
rect 2479 2473 2505 2479
rect 3151 2505 3177 2511
rect 3151 2473 3177 2479
rect 3319 2505 3345 2511
rect 3319 2473 3345 2479
rect 3711 2505 3737 2511
rect 3711 2473 3737 2479
rect 3879 2505 3905 2511
rect 3879 2473 3905 2479
rect 4271 2505 4297 2511
rect 4271 2473 4297 2479
rect 4439 2505 4465 2511
rect 4439 2473 4465 2479
rect 4719 2505 4745 2511
rect 4719 2473 4745 2479
rect 4831 2505 4857 2511
rect 4831 2473 4857 2479
rect 4999 2505 5025 2511
rect 4999 2473 5025 2479
rect 5279 2505 5305 2511
rect 5279 2473 5305 2479
rect 5447 2505 5473 2511
rect 5447 2473 5473 2479
rect 5559 2505 5585 2511
rect 5559 2473 5585 2479
rect 6063 2505 6089 2511
rect 6063 2473 6089 2479
rect 6231 2505 6257 2511
rect 6231 2473 6257 2479
rect 6343 2505 6369 2511
rect 6343 2473 6369 2479
rect 6847 2505 6873 2511
rect 6847 2473 6873 2479
rect 7015 2505 7041 2511
rect 7015 2473 7041 2479
rect 7407 2505 7433 2511
rect 7407 2473 7433 2479
rect 7575 2505 7601 2511
rect 7575 2473 7601 2479
rect 7967 2505 7993 2511
rect 7967 2473 7993 2479
rect 8135 2505 8161 2511
rect 8135 2473 8161 2479
rect 8527 2505 8553 2511
rect 8527 2473 8553 2479
rect 8695 2505 8721 2511
rect 8695 2473 8721 2479
rect 672 2365 9376 2382
rect 672 2339 2763 2365
rect 2789 2339 2815 2365
rect 2841 2339 2867 2365
rect 2893 2339 4919 2365
rect 4945 2339 4971 2365
rect 4997 2339 5023 2365
rect 5049 2339 7075 2365
rect 7101 2339 7127 2365
rect 7153 2339 7179 2365
rect 7205 2339 9231 2365
rect 9257 2339 9283 2365
rect 9309 2339 9335 2365
rect 9361 2339 9376 2365
rect 672 2322 9376 2339
rect 1415 2225 1441 2231
rect 1415 2193 1441 2199
rect 1975 2225 2001 2231
rect 1975 2193 2001 2199
rect 2535 2225 2561 2231
rect 2535 2193 2561 2199
rect 3095 2225 3121 2231
rect 3095 2193 3121 2199
rect 3655 2225 3681 2231
rect 3655 2193 3681 2199
rect 4215 2225 4241 2231
rect 4215 2193 4241 2199
rect 5055 2225 5081 2231
rect 5055 2193 5081 2199
rect 5895 2225 5921 2231
rect 5895 2193 5921 2199
rect 6455 2225 6481 2231
rect 6455 2193 6481 2199
rect 7575 2225 7601 2231
rect 7575 2193 7601 2199
rect 8135 2225 8161 2231
rect 8135 2193 8161 2199
rect 1583 2169 1609 2175
rect 1583 2137 1609 2143
rect 1751 2169 1777 2175
rect 1751 2137 1777 2143
rect 2087 2169 2113 2175
rect 2087 2137 2113 2143
rect 2311 2169 2337 2175
rect 2311 2137 2337 2143
rect 2703 2169 2729 2175
rect 2703 2137 2729 2143
rect 2871 2169 2897 2175
rect 2871 2137 2897 2143
rect 3263 2169 3289 2175
rect 3263 2137 3289 2143
rect 3375 2169 3401 2175
rect 3375 2137 3401 2143
rect 3823 2169 3849 2175
rect 3823 2137 3849 2143
rect 3991 2169 4017 2175
rect 3991 2137 4017 2143
rect 4327 2169 4353 2175
rect 4327 2137 4353 2143
rect 4551 2169 4577 2175
rect 4551 2137 4577 2143
rect 5223 2169 5249 2175
rect 5223 2137 5249 2143
rect 5391 2169 5417 2175
rect 5391 2137 5417 2143
rect 5615 2169 5641 2175
rect 5615 2137 5641 2143
rect 5727 2169 5753 2175
rect 5727 2137 5753 2143
rect 6119 2169 6145 2175
rect 6119 2137 6145 2143
rect 6287 2169 6313 2175
rect 6287 2137 6313 2143
rect 6735 2169 6761 2175
rect 6735 2137 6761 2143
rect 6903 2169 6929 2175
rect 6903 2137 6929 2143
rect 6959 2169 6985 2175
rect 6959 2137 6985 2143
rect 7295 2169 7321 2175
rect 7295 2137 7321 2143
rect 7463 2169 7489 2175
rect 7463 2137 7489 2143
rect 7799 2169 7825 2175
rect 7799 2137 7825 2143
rect 7967 2169 7993 2175
rect 7967 2137 7993 2143
rect 672 1973 9296 1990
rect 672 1947 1685 1973
rect 1711 1947 1737 1973
rect 1763 1947 1789 1973
rect 1815 1947 3841 1973
rect 3867 1947 3893 1973
rect 3919 1947 3945 1973
rect 3971 1947 5997 1973
rect 6023 1947 6049 1973
rect 6075 1947 6101 1973
rect 6127 1947 8153 1973
rect 8179 1947 8205 1973
rect 8231 1947 8257 1973
rect 8283 1947 9296 1973
rect 672 1930 9296 1947
rect 1079 1777 1105 1783
rect 1079 1745 1105 1751
rect 1639 1777 1665 1783
rect 1639 1745 1665 1751
rect 1807 1777 1833 1783
rect 1807 1745 1833 1751
rect 1919 1777 1945 1783
rect 1919 1745 1945 1751
rect 2199 1777 2225 1783
rect 2199 1745 2225 1751
rect 2311 1777 2337 1783
rect 2311 1745 2337 1751
rect 2479 1777 2505 1783
rect 2479 1745 2505 1751
rect 3039 1777 3065 1783
rect 3039 1745 3065 1751
rect 3207 1777 3233 1783
rect 3207 1745 3233 1751
rect 3319 1777 3345 1783
rect 3319 1745 3345 1751
rect 3599 1777 3625 1783
rect 3599 1745 3625 1751
rect 3767 1777 3793 1783
rect 3767 1745 3793 1751
rect 3935 1777 3961 1783
rect 3935 1745 3961 1751
rect 4159 1777 4185 1783
rect 4159 1745 4185 1751
rect 5167 1777 5193 1783
rect 5167 1745 5193 1751
rect 5335 1777 5361 1783
rect 5335 1745 5361 1751
rect 5503 1777 5529 1783
rect 5503 1745 5529 1751
rect 5839 1777 5865 1783
rect 5839 1745 5865 1751
rect 6007 1777 6033 1783
rect 6007 1745 6033 1751
rect 7071 1777 7097 1783
rect 7071 1745 7097 1751
rect 7295 1777 7321 1783
rect 7295 1745 7321 1751
rect 7463 1777 7489 1783
rect 7463 1745 7489 1751
rect 7631 1777 7657 1783
rect 7631 1745 7657 1751
rect 7855 1777 7881 1783
rect 7855 1745 7881 1751
rect 8023 1777 8049 1783
rect 8023 1745 8049 1751
rect 8135 1777 8161 1783
rect 8135 1745 8161 1751
rect 8975 1777 9001 1783
rect 8975 1745 9001 1751
rect 1191 1721 1217 1727
rect 1191 1689 1217 1695
rect 1359 1721 1385 1727
rect 1359 1689 1385 1695
rect 4271 1721 4297 1727
rect 4271 1689 4297 1695
rect 4439 1721 4465 1727
rect 4439 1689 4465 1695
rect 5727 1721 5753 1727
rect 5727 1689 5753 1695
rect 6791 1721 6817 1727
rect 6791 1689 6817 1695
rect 6959 1721 6985 1727
rect 6959 1689 6985 1695
rect 8751 1721 8777 1727
rect 8751 1689 8777 1695
rect 8919 1721 8945 1727
rect 8919 1689 8945 1695
rect 672 1581 9376 1598
rect 672 1555 2763 1581
rect 2789 1555 2815 1581
rect 2841 1555 2867 1581
rect 2893 1555 4919 1581
rect 4945 1555 4971 1581
rect 4997 1555 5023 1581
rect 5049 1555 7075 1581
rect 7101 1555 7127 1581
rect 7153 1555 7179 1581
rect 7205 1555 9231 1581
rect 9257 1555 9283 1581
rect 9309 1555 9335 1581
rect 9361 1555 9376 1581
rect 672 1538 9376 1555
<< via1 >>
rect 1685 4299 1711 4325
rect 1737 4299 1763 4325
rect 1789 4299 1815 4325
rect 3841 4299 3867 4325
rect 3893 4299 3919 4325
rect 3945 4299 3971 4325
rect 5997 4299 6023 4325
rect 6049 4299 6075 4325
rect 6101 4299 6127 4325
rect 8153 4299 8179 4325
rect 8205 4299 8231 4325
rect 8257 4299 8283 4325
rect 8079 4103 8105 4129
rect 8695 4103 8721 4129
rect 8863 4103 8889 4129
rect 8975 4103 9001 4129
rect 1191 4047 1217 4073
rect 1303 4047 1329 4073
rect 1471 4047 1497 4073
rect 1751 4047 1777 4073
rect 1919 4047 1945 4073
rect 2031 4047 2057 4073
rect 7911 4047 7937 4073
rect 8191 4047 8217 4073
rect 2763 3907 2789 3933
rect 2815 3907 2841 3933
rect 2867 3907 2893 3933
rect 4919 3907 4945 3933
rect 4971 3907 4997 3933
rect 5023 3907 5049 3933
rect 7075 3907 7101 3933
rect 7127 3907 7153 3933
rect 7179 3907 7205 3933
rect 9231 3907 9257 3933
rect 9283 3907 9309 3933
rect 9335 3907 9361 3933
rect 1191 3767 1217 3793
rect 1359 3711 1385 3737
rect 1471 3711 1497 3737
rect 1751 3711 1777 3737
rect 1863 3711 1889 3737
rect 1975 3711 2001 3737
rect 2311 3711 2337 3737
rect 2423 3711 2449 3737
rect 2535 3711 2561 3737
rect 7239 3711 7265 3737
rect 7351 3711 7377 3737
rect 7519 3711 7545 3737
rect 7799 3711 7825 3737
rect 7911 3711 7937 3737
rect 8023 3711 8049 3737
rect 1685 3515 1711 3541
rect 1737 3515 1763 3541
rect 1789 3515 1815 3541
rect 3841 3515 3867 3541
rect 3893 3515 3919 3541
rect 3945 3515 3971 3541
rect 5997 3515 6023 3541
rect 6049 3515 6075 3541
rect 6101 3515 6127 3541
rect 8153 3515 8179 3541
rect 8205 3515 8231 3541
rect 8257 3515 8283 3541
rect 1079 3319 1105 3345
rect 1639 3319 1665 3345
rect 1975 3319 2001 3345
rect 2199 3319 2225 3345
rect 2367 3319 2393 3345
rect 3487 3319 3513 3345
rect 3599 3319 3625 3345
rect 7071 3319 7097 3345
rect 7183 3319 7209 3345
rect 7351 3319 7377 3345
rect 7855 3319 7881 3345
rect 8247 3319 8273 3345
rect 8415 3319 8441 3345
rect 8975 3319 9001 3345
rect 1191 3263 1217 3289
rect 1359 3263 1385 3289
rect 1751 3263 1777 3289
rect 2479 3263 2505 3289
rect 3375 3263 3401 3289
rect 7575 3263 7601 3289
rect 7743 3263 7769 3289
rect 8135 3263 8161 3289
rect 8695 3263 8721 3289
rect 8863 3263 8889 3289
rect 2763 3123 2789 3149
rect 2815 3123 2841 3149
rect 2867 3123 2893 3149
rect 4919 3123 4945 3149
rect 4971 3123 4997 3149
rect 5023 3123 5049 3149
rect 7075 3123 7101 3149
rect 7127 3123 7153 3149
rect 7179 3123 7205 3149
rect 9231 3123 9257 3149
rect 9283 3123 9309 3149
rect 9335 3123 9361 3149
rect 1415 2983 1441 3009
rect 1975 2983 2001 3009
rect 2535 2983 2561 3009
rect 4495 2983 4521 3009
rect 7015 2983 7041 3009
rect 7575 2983 7601 3009
rect 8135 2983 8161 3009
rect 1583 2927 1609 2953
rect 1751 2927 1777 2953
rect 2143 2927 2169 2953
rect 2255 2927 2281 2953
rect 2703 2927 2729 2953
rect 2871 2927 2897 2953
rect 3095 2927 3121 2953
rect 3263 2927 3289 2953
rect 3375 2927 3401 2953
rect 3655 2927 3681 2953
rect 3823 2927 3849 2953
rect 3991 2927 4017 2953
rect 4215 2927 4241 2953
rect 4383 2927 4409 2953
rect 4831 2927 4857 2953
rect 4999 2927 5025 2953
rect 5167 2927 5193 2953
rect 6735 2927 6761 2953
rect 6847 2927 6873 2953
rect 7239 2927 7265 2953
rect 7407 2927 7433 2953
rect 7799 2927 7825 2953
rect 7967 2927 7993 2953
rect 1685 2731 1711 2757
rect 1737 2731 1763 2757
rect 1789 2731 1815 2757
rect 3841 2731 3867 2757
rect 3893 2731 3919 2757
rect 3945 2731 3971 2757
rect 5997 2731 6023 2757
rect 6049 2731 6075 2757
rect 6101 2731 6127 2757
rect 8153 2731 8179 2757
rect 8205 2731 8231 2757
rect 8257 2731 8283 2757
rect 1079 2535 1105 2561
rect 1639 2535 1665 2561
rect 2199 2535 2225 2561
rect 3039 2535 3065 2561
rect 3599 2535 3625 2561
rect 4215 2535 4241 2561
rect 7071 2535 7097 2561
rect 7687 2535 7713 2561
rect 8247 2535 8273 2561
rect 8751 2535 8777 2561
rect 1191 2479 1217 2505
rect 1359 2479 1385 2505
rect 1751 2479 1777 2505
rect 1919 2479 1945 2505
rect 2311 2479 2337 2505
rect 2479 2479 2505 2505
rect 3151 2479 3177 2505
rect 3319 2479 3345 2505
rect 3711 2479 3737 2505
rect 3879 2479 3905 2505
rect 4271 2479 4297 2505
rect 4439 2479 4465 2505
rect 4719 2479 4745 2505
rect 4831 2479 4857 2505
rect 4999 2479 5025 2505
rect 5279 2479 5305 2505
rect 5447 2479 5473 2505
rect 5559 2479 5585 2505
rect 6063 2479 6089 2505
rect 6231 2479 6257 2505
rect 6343 2479 6369 2505
rect 6847 2479 6873 2505
rect 7015 2479 7041 2505
rect 7407 2479 7433 2505
rect 7575 2479 7601 2505
rect 7967 2479 7993 2505
rect 8135 2479 8161 2505
rect 8527 2479 8553 2505
rect 8695 2479 8721 2505
rect 2763 2339 2789 2365
rect 2815 2339 2841 2365
rect 2867 2339 2893 2365
rect 4919 2339 4945 2365
rect 4971 2339 4997 2365
rect 5023 2339 5049 2365
rect 7075 2339 7101 2365
rect 7127 2339 7153 2365
rect 7179 2339 7205 2365
rect 9231 2339 9257 2365
rect 9283 2339 9309 2365
rect 9335 2339 9361 2365
rect 1415 2199 1441 2225
rect 1975 2199 2001 2225
rect 2535 2199 2561 2225
rect 3095 2199 3121 2225
rect 3655 2199 3681 2225
rect 4215 2199 4241 2225
rect 5055 2199 5081 2225
rect 5895 2199 5921 2225
rect 6455 2199 6481 2225
rect 7575 2199 7601 2225
rect 8135 2199 8161 2225
rect 1583 2143 1609 2169
rect 1751 2143 1777 2169
rect 2087 2143 2113 2169
rect 2311 2143 2337 2169
rect 2703 2143 2729 2169
rect 2871 2143 2897 2169
rect 3263 2143 3289 2169
rect 3375 2143 3401 2169
rect 3823 2143 3849 2169
rect 3991 2143 4017 2169
rect 4327 2143 4353 2169
rect 4551 2143 4577 2169
rect 5223 2143 5249 2169
rect 5391 2143 5417 2169
rect 5615 2143 5641 2169
rect 5727 2143 5753 2169
rect 6119 2143 6145 2169
rect 6287 2143 6313 2169
rect 6735 2143 6761 2169
rect 6903 2143 6929 2169
rect 6959 2143 6985 2169
rect 7295 2143 7321 2169
rect 7463 2143 7489 2169
rect 7799 2143 7825 2169
rect 7967 2143 7993 2169
rect 1685 1947 1711 1973
rect 1737 1947 1763 1973
rect 1789 1947 1815 1973
rect 3841 1947 3867 1973
rect 3893 1947 3919 1973
rect 3945 1947 3971 1973
rect 5997 1947 6023 1973
rect 6049 1947 6075 1973
rect 6101 1947 6127 1973
rect 8153 1947 8179 1973
rect 8205 1947 8231 1973
rect 8257 1947 8283 1973
rect 1079 1751 1105 1777
rect 1639 1751 1665 1777
rect 1807 1751 1833 1777
rect 1919 1751 1945 1777
rect 2199 1751 2225 1777
rect 2311 1751 2337 1777
rect 2479 1751 2505 1777
rect 3039 1751 3065 1777
rect 3207 1751 3233 1777
rect 3319 1751 3345 1777
rect 3599 1751 3625 1777
rect 3767 1751 3793 1777
rect 3935 1751 3961 1777
rect 4159 1751 4185 1777
rect 5167 1751 5193 1777
rect 5335 1751 5361 1777
rect 5503 1751 5529 1777
rect 5839 1751 5865 1777
rect 6007 1751 6033 1777
rect 7071 1751 7097 1777
rect 7295 1751 7321 1777
rect 7463 1751 7489 1777
rect 7631 1751 7657 1777
rect 7855 1751 7881 1777
rect 8023 1751 8049 1777
rect 8135 1751 8161 1777
rect 8975 1751 9001 1777
rect 1191 1695 1217 1721
rect 1359 1695 1385 1721
rect 4271 1695 4297 1721
rect 4439 1695 4465 1721
rect 5727 1695 5753 1721
rect 6791 1695 6817 1721
rect 6959 1695 6985 1721
rect 8751 1695 8777 1721
rect 8919 1695 8945 1721
rect 2763 1555 2789 1581
rect 2815 1555 2841 1581
rect 2867 1555 2893 1581
rect 4919 1555 4945 1581
rect 4971 1555 4997 1581
rect 5023 1555 5049 1581
rect 7075 1555 7101 1581
rect 7127 1555 7153 1581
rect 7179 1555 7205 1581
rect 9231 1555 9257 1581
rect 9283 1555 9309 1581
rect 9335 1555 9361 1581
<< metal2 >>
rect 4928 5600 4984 6000
rect 1684 4326 1816 4331
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1684 4293 1816 4298
rect 3840 4326 3972 4331
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3840 4293 3972 4298
rect 4942 4214 4970 5600
rect 5996 4326 6128 4331
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 5996 4293 6128 4298
rect 8152 4326 8284 4331
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8152 4293 8284 4298
rect 4830 4186 4970 4214
rect 1190 4073 1218 4079
rect 1190 4047 1191 4073
rect 1217 4047 1218 4073
rect 1190 3794 1218 4047
rect 1078 3793 1218 3794
rect 1078 3767 1191 3793
rect 1217 3767 1218 3793
rect 1078 3766 1218 3767
rect 1078 3346 1106 3766
rect 1190 3761 1218 3766
rect 1302 4074 1330 4079
rect 1470 4074 1498 4079
rect 1302 4073 1498 4074
rect 1302 4047 1303 4073
rect 1329 4047 1471 4073
rect 1497 4047 1498 4073
rect 1302 4046 1498 4047
rect 1302 3458 1330 4046
rect 1470 4041 1498 4046
rect 1750 4074 1778 4079
rect 1918 4074 1946 4079
rect 1750 4073 1946 4074
rect 1750 4047 1751 4073
rect 1777 4047 1919 4073
rect 1945 4047 1946 4073
rect 1750 4046 1946 4047
rect 1750 4041 1778 4046
rect 1918 3850 1946 4046
rect 1918 3817 1946 3822
rect 2030 4073 2058 4079
rect 2030 4047 2031 4073
rect 2057 4047 2058 4073
rect 1358 3738 1386 3743
rect 1470 3738 1498 3743
rect 1750 3738 1778 3743
rect 1862 3738 1890 3743
rect 1974 3738 2002 3743
rect 2030 3738 2058 4047
rect 2762 3934 2894 3939
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2762 3901 2894 3906
rect 1358 3737 1610 3738
rect 1358 3711 1359 3737
rect 1385 3711 1471 3737
rect 1497 3711 1610 3737
rect 1358 3710 1610 3711
rect 1358 3705 1386 3710
rect 1470 3705 1498 3710
rect 1582 3458 1610 3710
rect 1750 3737 1890 3738
rect 1750 3711 1751 3737
rect 1777 3711 1863 3737
rect 1889 3711 1890 3737
rect 1750 3710 1890 3711
rect 1750 3705 1778 3710
rect 1684 3542 1816 3547
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1684 3509 1816 3514
rect 1862 3458 1890 3710
rect 1302 3430 1498 3458
rect 1078 2562 1106 3318
rect 1414 3346 1442 3351
rect 1190 3290 1218 3295
rect 1358 3290 1386 3295
rect 1078 1777 1106 2534
rect 1134 3289 1386 3290
rect 1134 3263 1191 3289
rect 1217 3263 1359 3289
rect 1385 3263 1386 3289
rect 1134 3262 1386 3263
rect 1134 1834 1162 3262
rect 1190 3257 1218 3262
rect 1358 3257 1386 3262
rect 1414 3010 1442 3318
rect 1414 2944 1442 2982
rect 1414 2562 1442 2567
rect 1190 2506 1218 2511
rect 1358 2506 1386 2511
rect 1190 2505 1386 2506
rect 1190 2479 1191 2505
rect 1217 2479 1359 2505
rect 1385 2479 1386 2505
rect 1190 2478 1386 2479
rect 1190 2473 1218 2478
rect 1358 2282 1386 2478
rect 1358 2249 1386 2254
rect 1134 1801 1162 1806
rect 1414 2225 1442 2534
rect 1414 2199 1415 2225
rect 1441 2199 1442 2225
rect 1078 1751 1079 1777
rect 1105 1751 1106 1777
rect 1078 1745 1106 1751
rect 1414 1778 1442 2199
rect 1414 1745 1442 1750
rect 1190 1722 1218 1741
rect 1190 1689 1218 1694
rect 1358 1722 1386 1741
rect 1470 1694 1498 3430
rect 1358 1689 1386 1694
rect 1414 1666 1498 1694
rect 1526 3430 1610 3458
rect 1806 3430 1890 3458
rect 1918 3737 2058 3738
rect 1918 3711 1975 3737
rect 2001 3711 2058 3737
rect 1918 3710 2058 3711
rect 2086 3850 2114 3855
rect 1414 400 1442 1666
rect 1526 400 1554 3430
rect 1638 3346 1666 3351
rect 1638 3299 1666 3318
rect 1750 3290 1778 3295
rect 1750 3243 1778 3262
rect 1806 3234 1834 3430
rect 1918 3346 1946 3710
rect 1974 3705 2002 3710
rect 1918 3313 1946 3318
rect 1974 3346 2002 3351
rect 1974 3345 2058 3346
rect 1974 3319 1975 3345
rect 2001 3319 2058 3345
rect 1974 3318 2058 3319
rect 1974 3290 2002 3318
rect 1974 3257 2002 3262
rect 1806 3206 1890 3234
rect 1582 2953 1610 2959
rect 1582 2927 1583 2953
rect 1609 2927 1610 2953
rect 1582 2842 1610 2927
rect 1582 2809 1610 2814
rect 1750 2953 1778 2959
rect 1750 2927 1751 2953
rect 1777 2927 1778 2953
rect 1750 2842 1778 2927
rect 1750 2809 1778 2814
rect 1684 2758 1816 2763
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1684 2725 1816 2730
rect 1638 2562 1666 2567
rect 1638 2515 1666 2534
rect 1750 2506 1778 2511
rect 1750 2459 1778 2478
rect 1582 2170 1610 2175
rect 1582 2123 1610 2142
rect 1750 2170 1778 2175
rect 1750 2058 1778 2142
rect 1750 2025 1778 2030
rect 1684 1974 1816 1979
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1684 1941 1816 1946
rect 1582 1890 1610 1895
rect 1582 1666 1610 1862
rect 1694 1834 1722 1839
rect 1638 1778 1666 1783
rect 1638 1731 1666 1750
rect 1582 1638 1666 1666
rect 1638 400 1666 1638
rect 1694 1610 1722 1806
rect 1806 1778 1834 1783
rect 1806 1731 1834 1750
rect 1694 1582 1778 1610
rect 1750 400 1778 1582
rect 1862 400 1890 3206
rect 1974 3010 2002 3015
rect 1974 2963 2002 2982
rect 1974 2562 2002 2567
rect 1918 2506 1946 2511
rect 1918 2459 1946 2478
rect 1974 2225 2002 2534
rect 1974 2199 1975 2225
rect 2001 2199 2002 2225
rect 1974 2193 2002 2199
rect 2030 2114 2058 3318
rect 2086 2842 2114 3822
rect 2310 3738 2338 3743
rect 2422 3738 2450 3743
rect 2310 3737 2450 3738
rect 2310 3711 2311 3737
rect 2337 3711 2423 3737
rect 2449 3711 2450 3737
rect 2310 3710 2450 3711
rect 2198 3346 2226 3351
rect 2198 3299 2226 3318
rect 2142 2954 2170 2959
rect 2254 2954 2282 2959
rect 2142 2953 2282 2954
rect 2142 2927 2143 2953
rect 2169 2927 2255 2953
rect 2281 2927 2282 2953
rect 2142 2926 2282 2927
rect 2142 2921 2170 2926
rect 2086 2814 2170 2842
rect 2086 2170 2114 2175
rect 2086 2123 2114 2142
rect 1918 2086 2058 2114
rect 1918 1890 1946 2086
rect 2142 1890 2170 2814
rect 1918 1862 2002 1890
rect 1918 1778 1946 1783
rect 1918 1731 1946 1750
rect 1974 400 2002 1862
rect 2142 1857 2170 1862
rect 2198 2562 2226 2567
rect 2086 1834 2114 1839
rect 2086 400 2114 1806
rect 2198 1777 2226 2534
rect 2254 2394 2282 2926
rect 2310 2618 2338 3710
rect 2422 3705 2450 3710
rect 2534 3737 2562 3743
rect 2534 3711 2535 3737
rect 2561 3711 2562 3737
rect 2366 3346 2394 3351
rect 2366 3345 2450 3346
rect 2366 3319 2367 3345
rect 2393 3319 2450 3345
rect 2366 3318 2450 3319
rect 2366 3313 2394 3318
rect 2422 3290 2450 3318
rect 2478 3290 2506 3295
rect 2422 3289 2506 3290
rect 2422 3263 2479 3289
rect 2505 3263 2506 3289
rect 2422 3262 2506 3263
rect 2310 2590 2394 2618
rect 2310 2506 2338 2511
rect 2310 2459 2338 2478
rect 2254 2361 2282 2366
rect 2198 1751 2199 1777
rect 2225 1751 2226 1777
rect 2198 1745 2226 1751
rect 2254 2282 2282 2287
rect 2254 1610 2282 2254
rect 2310 2170 2338 2175
rect 2310 2123 2338 2142
rect 2310 1890 2338 1895
rect 2310 1777 2338 1862
rect 2310 1751 2311 1777
rect 2337 1751 2338 1777
rect 2310 1745 2338 1751
rect 2366 1610 2394 2590
rect 2198 1582 2282 1610
rect 2310 1582 2394 1610
rect 2198 400 2226 1582
rect 2310 400 2338 1582
rect 2422 400 2450 3262
rect 2478 3257 2506 3262
rect 2534 3010 2562 3711
rect 3840 3542 3972 3547
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3840 3509 3972 3514
rect 3486 3346 3514 3351
rect 3430 3345 3514 3346
rect 3430 3319 3487 3345
rect 3513 3319 3514 3345
rect 3430 3318 3514 3319
rect 3374 3290 3402 3295
rect 3430 3290 3458 3318
rect 3486 3313 3514 3318
rect 3598 3345 3626 3351
rect 3598 3319 3599 3345
rect 3625 3319 3626 3345
rect 3374 3289 3458 3290
rect 3374 3263 3375 3289
rect 3401 3263 3458 3289
rect 3374 3262 3458 3263
rect 3374 3257 3402 3262
rect 2762 3150 2894 3155
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2762 3117 2894 3122
rect 2534 2562 2562 2982
rect 2702 2954 2730 2959
rect 2870 2954 2898 2959
rect 2702 2953 2898 2954
rect 2702 2927 2703 2953
rect 2729 2927 2871 2953
rect 2897 2927 2898 2953
rect 2702 2926 2898 2927
rect 2702 2921 2730 2926
rect 2870 2842 2898 2926
rect 3094 2953 3122 2959
rect 3094 2927 3095 2953
rect 3121 2927 3122 2953
rect 2870 2814 3010 2842
rect 2478 2506 2506 2525
rect 2478 2473 2506 2478
rect 2478 2394 2506 2399
rect 2478 2058 2506 2366
rect 2534 2225 2562 2534
rect 2926 2506 2954 2511
rect 2534 2199 2535 2225
rect 2561 2199 2562 2225
rect 2534 2193 2562 2199
rect 2646 2450 2674 2455
rect 2478 2030 2562 2058
rect 2478 1890 2506 1895
rect 2478 1777 2506 1862
rect 2478 1751 2479 1777
rect 2505 1751 2506 1777
rect 2478 1745 2506 1751
rect 2534 400 2562 2030
rect 2646 400 2674 2422
rect 2762 2366 2894 2371
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2762 2333 2894 2338
rect 2702 2170 2730 2175
rect 2870 2170 2898 2175
rect 2702 2169 2898 2170
rect 2702 2143 2703 2169
rect 2729 2143 2871 2169
rect 2897 2143 2898 2169
rect 2702 2142 2898 2143
rect 2702 2137 2730 2142
rect 2702 2058 2730 2063
rect 2702 1498 2730 2030
rect 2870 2058 2898 2142
rect 2870 2025 2898 2030
rect 2926 1834 2954 2478
rect 2926 1801 2954 1806
rect 2926 1722 2954 1727
rect 2762 1582 2894 1587
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2762 1549 2894 1554
rect 2702 1470 2786 1498
rect 2758 400 2786 1470
rect 2926 1218 2954 1694
rect 2870 1190 2954 1218
rect 2870 400 2898 1190
rect 2982 400 3010 2814
rect 3038 2562 3066 2567
rect 3094 2562 3122 2927
rect 3262 2954 3290 2959
rect 3262 2907 3290 2926
rect 3374 2954 3402 2959
rect 3374 2907 3402 2926
rect 3066 2534 3122 2562
rect 3038 2515 3066 2534
rect 3094 2226 3122 2534
rect 3150 2506 3178 2511
rect 3318 2506 3346 2511
rect 3150 2505 3346 2506
rect 3150 2479 3151 2505
rect 3177 2479 3319 2505
rect 3345 2479 3346 2505
rect 3150 2478 3346 2479
rect 3150 2473 3178 2478
rect 3318 2394 3346 2478
rect 3318 2361 3346 2366
rect 3038 2225 3122 2226
rect 3038 2199 3095 2225
rect 3121 2199 3122 2225
rect 3038 2198 3122 2199
rect 3038 1777 3066 2198
rect 3094 2193 3122 2198
rect 3150 2170 3178 2175
rect 3038 1751 3039 1777
rect 3065 1751 3066 1777
rect 3038 1745 3066 1751
rect 3094 1834 3122 1839
rect 3094 400 3122 1806
rect 3150 1554 3178 2142
rect 3262 2170 3290 2175
rect 3262 2123 3290 2142
rect 3374 2170 3402 2175
rect 3374 2123 3402 2142
rect 3318 1834 3346 1839
rect 3206 1778 3234 1783
rect 3318 1778 3346 1806
rect 3206 1777 3346 1778
rect 3206 1751 3207 1777
rect 3233 1751 3319 1777
rect 3345 1751 3346 1777
rect 3206 1750 3346 1751
rect 3206 1745 3234 1750
rect 3318 1745 3346 1750
rect 3206 1666 3234 1671
rect 3234 1638 3290 1666
rect 3206 1633 3234 1638
rect 3150 1526 3234 1554
rect 3206 400 3234 1526
rect 3262 1274 3290 1638
rect 3262 1246 3346 1274
rect 3318 400 3346 1246
rect 3430 400 3458 3262
rect 3542 2954 3570 2959
rect 3542 400 3570 2926
rect 3598 2954 3626 3319
rect 4494 3234 4522 3239
rect 4494 3009 4522 3206
rect 4830 3234 4858 4186
rect 8078 4129 8106 4135
rect 8694 4130 8722 4135
rect 8862 4130 8890 4135
rect 8078 4103 8079 4129
rect 8105 4103 8106 4129
rect 7910 4074 7938 4079
rect 7854 4073 7938 4074
rect 7854 4047 7911 4073
rect 7937 4047 7938 4073
rect 7854 4046 7938 4047
rect 4918 3934 5050 3939
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 4918 3901 5050 3906
rect 7074 3934 7206 3939
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7074 3901 7206 3906
rect 7238 3738 7266 3743
rect 7070 3710 7238 3738
rect 5996 3542 6128 3547
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 5996 3509 6128 3514
rect 7070 3346 7098 3710
rect 7238 3691 7266 3710
rect 7350 3738 7378 3743
rect 7518 3738 7546 3743
rect 7350 3737 7546 3738
rect 7350 3711 7351 3737
rect 7377 3711 7519 3737
rect 7545 3711 7546 3737
rect 7350 3710 7546 3711
rect 7350 3705 7378 3710
rect 7014 3345 7098 3346
rect 7014 3319 7071 3345
rect 7097 3319 7098 3345
rect 7014 3318 7098 3319
rect 4858 3206 5138 3234
rect 4830 3168 4858 3206
rect 4918 3150 5050 3155
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 4918 3117 5050 3122
rect 4494 2983 4495 3009
rect 4521 2983 4522 3009
rect 4494 2977 4522 2983
rect 3654 2954 3682 2959
rect 3598 2953 3682 2954
rect 3598 2927 3655 2953
rect 3681 2927 3682 2953
rect 3598 2926 3682 2927
rect 3598 2562 3626 2926
rect 3654 2921 3682 2926
rect 3822 2954 3850 2959
rect 3990 2954 4018 2959
rect 4214 2954 4242 2959
rect 4382 2954 4410 2959
rect 3822 2953 4074 2954
rect 3822 2927 3823 2953
rect 3849 2927 3991 2953
rect 4017 2927 4074 2953
rect 3822 2926 4074 2927
rect 3822 2921 3850 2926
rect 3990 2921 4018 2926
rect 3840 2758 3972 2763
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3840 2725 3972 2730
rect 3598 2226 3626 2534
rect 3710 2506 3738 2511
rect 3878 2506 3906 2511
rect 3710 2505 3906 2506
rect 3710 2479 3711 2505
rect 3737 2479 3879 2505
rect 3905 2479 3906 2505
rect 3710 2478 3906 2479
rect 3710 2473 3738 2478
rect 3710 2394 3738 2399
rect 3654 2226 3682 2231
rect 3598 2225 3682 2226
rect 3598 2199 3655 2225
rect 3681 2199 3682 2225
rect 3598 2198 3682 2199
rect 3598 1777 3626 2198
rect 3654 2193 3682 2198
rect 3598 1751 3599 1777
rect 3625 1751 3626 1777
rect 3598 1745 3626 1751
rect 3654 2058 3682 2063
rect 3654 400 3682 2030
rect 3710 1666 3738 2366
rect 3822 2169 3850 2175
rect 3822 2143 3823 2169
rect 3849 2143 3850 2169
rect 3822 2114 3850 2143
rect 3822 2081 3850 2086
rect 3878 2058 3906 2478
rect 3990 2169 4018 2175
rect 3990 2143 3991 2169
rect 4017 2143 4018 2169
rect 3990 2114 4018 2143
rect 3990 2081 4018 2086
rect 3878 2025 3906 2030
rect 3840 1974 3972 1979
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3840 1941 3972 1946
rect 3878 1890 3906 1895
rect 4046 1890 4074 2926
rect 4214 2953 4410 2954
rect 4214 2927 4215 2953
rect 4241 2927 4383 2953
rect 4409 2927 4410 2953
rect 4214 2926 4410 2927
rect 4214 2921 4242 2926
rect 4214 2562 4242 2567
rect 4214 2226 4242 2534
rect 4270 2506 4298 2511
rect 4270 2459 4298 2478
rect 4158 2198 4214 2226
rect 3766 1778 3794 1783
rect 3766 1731 3794 1750
rect 3710 1638 3794 1666
rect 3766 400 3794 1638
rect 3878 400 3906 1862
rect 3990 1862 4074 1890
rect 4102 2170 4130 2175
rect 3934 1778 3962 1783
rect 3934 1731 3962 1750
rect 3990 400 4018 1862
rect 4102 400 4130 2142
rect 4158 1777 4186 2198
rect 4214 2179 4242 2198
rect 4326 2170 4354 2175
rect 4326 2123 4354 2142
rect 4158 1751 4159 1777
rect 4185 1751 4186 1777
rect 4158 1745 4186 1751
rect 4214 2058 4242 2063
rect 4214 400 4242 2030
rect 4382 2002 4410 2926
rect 4830 2954 4858 2959
rect 4998 2954 5026 2959
rect 4830 2953 5026 2954
rect 4830 2927 4831 2953
rect 4857 2927 4999 2953
rect 5025 2927 5026 2953
rect 4830 2926 5026 2927
rect 5110 2954 5138 3206
rect 7014 3010 7042 3318
rect 7070 3313 7098 3318
rect 7182 3346 7210 3351
rect 7182 3299 7210 3318
rect 7350 3346 7378 3351
rect 7350 3299 7378 3318
rect 7518 3178 7546 3710
rect 7798 3738 7826 3743
rect 7854 3738 7882 4046
rect 7910 4041 7938 4046
rect 8078 4074 8106 4103
rect 8470 4129 8890 4130
rect 8470 4103 8695 4129
rect 8721 4103 8863 4129
rect 8889 4103 8890 4129
rect 8470 4102 8890 4103
rect 8190 4074 8218 4079
rect 8078 4073 8218 4074
rect 8078 4047 8191 4073
rect 8217 4047 8218 4073
rect 8078 4046 8218 4047
rect 7826 3710 7882 3738
rect 7798 3672 7826 3710
rect 7854 3346 7882 3710
rect 7910 3738 7938 3743
rect 8022 3738 8050 3743
rect 7910 3737 8050 3738
rect 7910 3711 7911 3737
rect 7937 3711 8023 3737
rect 8049 3711 8050 3737
rect 7910 3710 8050 3711
rect 7910 3705 7938 3710
rect 7574 3290 7602 3295
rect 7742 3290 7770 3295
rect 7574 3289 7770 3290
rect 7574 3263 7575 3289
rect 7601 3263 7743 3289
rect 7769 3263 7770 3289
rect 7574 3262 7770 3263
rect 7574 3257 7602 3262
rect 7074 3150 7206 3155
rect 7518 3150 7658 3178
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7074 3117 7206 3122
rect 7574 3066 7602 3071
rect 7014 3009 7098 3010
rect 7014 2983 7015 3009
rect 7041 2983 7098 3009
rect 7014 2982 7098 2983
rect 7014 2977 7042 2982
rect 5166 2954 5194 2959
rect 5110 2953 5194 2954
rect 5110 2927 5167 2953
rect 5193 2927 5194 2953
rect 5110 2926 5194 2927
rect 4494 2842 4522 2847
rect 4438 2506 4466 2511
rect 4438 2459 4466 2478
rect 4326 1974 4410 2002
rect 4270 1722 4298 1727
rect 4270 1675 4298 1694
rect 4326 400 4354 1974
rect 4438 1722 4466 1727
rect 4438 1675 4466 1694
rect 4494 1610 4522 2814
rect 4830 2842 4858 2926
rect 4998 2921 5026 2926
rect 4830 2809 4858 2814
rect 4718 2505 4746 2511
rect 4718 2479 4719 2505
rect 4745 2479 4746 2505
rect 4718 2226 4746 2479
rect 4718 2193 4746 2198
rect 4774 2506 4802 2511
rect 4550 2170 4578 2175
rect 4578 2142 4634 2170
rect 4550 2104 4578 2142
rect 4438 1582 4522 1610
rect 4550 1834 4578 1839
rect 4438 400 4466 1582
rect 4550 400 4578 1806
rect 4606 1442 4634 2142
rect 4606 1409 4634 1414
rect 4662 2114 4690 2119
rect 4662 400 4690 2086
rect 4774 400 4802 2478
rect 4830 2506 4858 2511
rect 4998 2506 5026 2511
rect 4830 2505 5138 2506
rect 4830 2479 4831 2505
rect 4857 2479 4999 2505
rect 5025 2479 5138 2505
rect 4830 2478 5138 2479
rect 4830 2473 4858 2478
rect 4998 2473 5026 2478
rect 4918 2366 5050 2371
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 4918 2333 5050 2338
rect 5054 2226 5082 2231
rect 5054 2179 5082 2198
rect 4830 1778 4858 1783
rect 4830 882 4858 1750
rect 4918 1582 5050 1587
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 4918 1549 5050 1554
rect 4998 1442 5026 1447
rect 4830 854 4914 882
rect 4886 400 4914 854
rect 4998 400 5026 1414
rect 5110 400 5138 2478
rect 5166 2226 5194 2926
rect 6734 2954 6762 2959
rect 6846 2954 6874 2959
rect 6734 2953 6874 2954
rect 6734 2927 6735 2953
rect 6761 2927 6847 2953
rect 6873 2927 6874 2953
rect 6734 2926 6874 2927
rect 5996 2758 6128 2763
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 5996 2725 6128 2730
rect 5166 1777 5194 2198
rect 5278 2506 5306 2511
rect 5446 2506 5474 2511
rect 5278 2505 5474 2506
rect 5278 2479 5279 2505
rect 5305 2479 5447 2505
rect 5473 2479 5474 2505
rect 5278 2478 5474 2479
rect 5222 2170 5250 2175
rect 5222 2123 5250 2142
rect 5166 1751 5167 1777
rect 5193 1751 5194 1777
rect 5166 1745 5194 1751
rect 5222 1722 5250 1727
rect 5222 400 5250 1694
rect 5278 1666 5306 2478
rect 5446 2473 5474 2478
rect 5558 2505 5586 2511
rect 5558 2479 5559 2505
rect 5585 2479 5586 2505
rect 5558 2226 5586 2479
rect 6062 2506 6090 2511
rect 6230 2506 6258 2511
rect 6062 2505 6258 2506
rect 6062 2479 6063 2505
rect 6089 2479 6231 2505
rect 6257 2479 6258 2505
rect 6062 2478 6258 2479
rect 6062 2473 6090 2478
rect 5558 2193 5586 2198
rect 5894 2226 5922 2231
rect 5894 2179 5922 2198
rect 6174 2226 6202 2231
rect 5390 2170 5418 2175
rect 5614 2170 5642 2175
rect 5726 2170 5754 2175
rect 5418 2142 5474 2170
rect 5390 2104 5418 2142
rect 5334 1778 5362 1783
rect 5334 1731 5362 1750
rect 5278 1638 5362 1666
rect 5334 400 5362 1638
rect 5446 400 5474 2142
rect 5614 2169 5754 2170
rect 5614 2143 5615 2169
rect 5641 2143 5727 2169
rect 5753 2143 5754 2169
rect 5614 2142 5754 2143
rect 5614 2137 5642 2142
rect 5502 1778 5530 1783
rect 5530 1750 5586 1778
rect 5502 1712 5530 1750
rect 5558 400 5586 1750
rect 5670 400 5698 2142
rect 5726 2137 5754 2142
rect 6118 2170 6146 2175
rect 6118 2058 6146 2142
rect 5894 2030 6146 2058
rect 5838 1778 5866 1783
rect 5782 1777 5866 1778
rect 5782 1751 5839 1777
rect 5865 1751 5866 1777
rect 5782 1750 5866 1751
rect 5726 1722 5754 1727
rect 5782 1722 5810 1750
rect 5838 1745 5866 1750
rect 5726 1721 5810 1722
rect 5726 1695 5727 1721
rect 5753 1695 5810 1721
rect 5726 1694 5810 1695
rect 5726 1689 5754 1694
rect 5782 400 5810 1694
rect 5894 400 5922 2030
rect 5996 1974 6128 1979
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 5996 1941 6128 1946
rect 6174 1890 6202 2198
rect 6006 1862 6202 1890
rect 6006 1777 6034 1862
rect 6006 1751 6007 1777
rect 6033 1751 6034 1777
rect 6006 1745 6034 1751
rect 6062 1722 6090 1727
rect 6062 1274 6090 1694
rect 6230 1666 6258 2478
rect 6342 2506 6370 2511
rect 6510 2506 6538 2511
rect 6342 2505 6482 2506
rect 6342 2479 6343 2505
rect 6369 2479 6482 2505
rect 6342 2478 6482 2479
rect 6342 2473 6370 2478
rect 6454 2226 6482 2478
rect 6454 2179 6482 2198
rect 6286 2170 6314 2175
rect 6286 2123 6314 2142
rect 6006 1246 6090 1274
rect 6118 1638 6258 1666
rect 6286 2058 6314 2063
rect 6510 2058 6538 2478
rect 6734 2282 6762 2926
rect 6846 2921 6874 2926
rect 7070 2618 7098 2982
rect 7574 3009 7602 3038
rect 7574 2983 7575 3009
rect 7601 2983 7602 3009
rect 7574 2977 7602 2983
rect 6958 2590 7098 2618
rect 6846 2506 6874 2511
rect 6846 2459 6874 2478
rect 6734 2254 6874 2282
rect 6006 400 6034 1246
rect 6118 400 6146 1638
rect 6286 1610 6314 2030
rect 6454 2030 6538 2058
rect 6566 2170 6594 2175
rect 6230 1582 6314 1610
rect 6342 1778 6370 1783
rect 6230 400 6258 1582
rect 6342 400 6370 1750
rect 6454 400 6482 2030
rect 6566 400 6594 2142
rect 6734 2169 6762 2175
rect 6734 2143 6735 2169
rect 6761 2143 6762 2169
rect 6734 2058 6762 2143
rect 6734 2025 6762 2030
rect 6678 1834 6706 1839
rect 6678 400 6706 1806
rect 6790 1722 6818 1727
rect 6790 1675 6818 1694
rect 6846 1610 6874 2254
rect 6958 2226 6986 2590
rect 7070 2561 7098 2590
rect 7070 2535 7071 2561
rect 7097 2535 7098 2561
rect 7070 2529 7098 2535
rect 7238 2954 7266 2959
rect 7406 2954 7434 2959
rect 7238 2953 7434 2954
rect 7238 2927 7239 2953
rect 7265 2927 7407 2953
rect 7433 2927 7434 2953
rect 7238 2926 7434 2927
rect 7014 2506 7042 2511
rect 7014 2459 7042 2478
rect 7074 2366 7206 2371
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7074 2333 7206 2338
rect 6902 2169 6930 2175
rect 6902 2143 6903 2169
rect 6929 2143 6930 2169
rect 6902 2058 6930 2143
rect 6958 2170 6986 2198
rect 6958 2169 7098 2170
rect 6958 2143 6959 2169
rect 6985 2143 7098 2169
rect 6958 2142 7098 2143
rect 6958 2137 6986 2142
rect 6902 2025 6930 2030
rect 7014 2058 7042 2063
rect 6790 1582 6874 1610
rect 6902 1946 6930 1951
rect 6790 400 6818 1582
rect 6902 400 6930 1918
rect 6958 1722 6986 1727
rect 6958 1675 6986 1694
rect 7014 400 7042 2030
rect 7070 1777 7098 2142
rect 7070 1751 7071 1777
rect 7097 1751 7098 1777
rect 7070 1745 7098 1751
rect 7074 1582 7206 1587
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7074 1549 7206 1554
rect 7238 1498 7266 2926
rect 7406 2921 7434 2926
rect 7350 2842 7378 2847
rect 7294 2170 7322 2175
rect 7294 2123 7322 2142
rect 7350 1946 7378 2814
rect 7406 2506 7434 2511
rect 7574 2506 7602 2511
rect 7406 2505 7602 2506
rect 7406 2479 7407 2505
rect 7433 2479 7575 2505
rect 7601 2479 7602 2505
rect 7406 2478 7602 2479
rect 7406 2058 7434 2478
rect 7574 2473 7602 2478
rect 7518 2394 7546 2399
rect 7462 2170 7490 2175
rect 7462 2123 7490 2142
rect 7406 2025 7434 2030
rect 7350 1918 7434 1946
rect 7294 1778 7322 1783
rect 7294 1731 7322 1750
rect 7126 1470 7266 1498
rect 7350 1722 7378 1727
rect 7126 400 7154 1470
rect 7350 1386 7378 1694
rect 7406 1666 7434 1918
rect 7462 1778 7490 1783
rect 7462 1731 7490 1750
rect 7406 1638 7490 1666
rect 7238 1358 7378 1386
rect 7238 400 7266 1358
rect 7462 1330 7490 1638
rect 7462 1297 7490 1302
rect 7518 1218 7546 2366
rect 7574 2226 7602 2231
rect 7574 2179 7602 2198
rect 7350 1190 7546 1218
rect 7574 2058 7602 2063
rect 7350 400 7378 1190
rect 7462 1050 7490 1055
rect 7462 400 7490 1022
rect 7574 400 7602 2030
rect 7630 1890 7658 3150
rect 7630 1857 7658 1862
rect 7686 3066 7714 3071
rect 7686 2561 7714 3038
rect 7686 2535 7687 2561
rect 7713 2535 7714 2561
rect 7686 2450 7714 2535
rect 7686 2226 7714 2422
rect 7630 1778 7658 1783
rect 7686 1778 7714 2198
rect 7630 1777 7686 1778
rect 7630 1751 7631 1777
rect 7657 1751 7686 1777
rect 7630 1750 7686 1751
rect 7630 1745 7658 1750
rect 7686 1745 7714 1750
rect 7742 1694 7770 3262
rect 7854 3066 7882 3318
rect 7854 3033 7882 3038
rect 7798 2954 7826 2959
rect 7966 2954 7994 2959
rect 7798 2953 7994 2954
rect 7798 2927 7799 2953
rect 7825 2927 7967 2953
rect 7993 2927 7994 2953
rect 7798 2926 7994 2927
rect 7798 2842 7826 2926
rect 7966 2921 7994 2926
rect 7798 2809 7826 2814
rect 7910 2842 7938 2847
rect 7798 2170 7826 2175
rect 7798 1946 7826 2142
rect 7798 1913 7826 1918
rect 7854 1834 7882 1839
rect 7854 1777 7882 1806
rect 7854 1751 7855 1777
rect 7881 1751 7882 1777
rect 7854 1745 7882 1751
rect 7910 1694 7938 2814
rect 7966 2506 7994 2511
rect 7966 2459 7994 2478
rect 7966 2170 7994 2175
rect 7966 2123 7994 2142
rect 8022 2058 8050 3710
rect 7686 1666 7770 1694
rect 7798 1666 7938 1694
rect 7966 2030 8050 2058
rect 7686 400 7714 1666
rect 7798 400 7826 1666
rect 7966 1610 7994 2030
rect 8022 1834 8050 1839
rect 8022 1777 8050 1806
rect 8022 1751 8023 1777
rect 8049 1751 8050 1777
rect 8022 1745 8050 1751
rect 8078 1694 8106 4046
rect 8190 4041 8218 4046
rect 8152 3542 8284 3547
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8152 3509 8284 3514
rect 8246 3346 8274 3351
rect 8190 3345 8274 3346
rect 8190 3319 8247 3345
rect 8273 3319 8274 3345
rect 8190 3318 8274 3319
rect 8134 3290 8162 3295
rect 8190 3290 8218 3318
rect 8246 3313 8274 3318
rect 8414 3346 8442 3351
rect 8414 3299 8442 3318
rect 8134 3289 8218 3290
rect 8134 3263 8135 3289
rect 8161 3263 8218 3289
rect 8134 3262 8218 3263
rect 8134 3257 8162 3262
rect 8134 3066 8162 3071
rect 8134 3009 8162 3038
rect 8134 2983 8135 3009
rect 8161 2983 8162 3009
rect 8134 2977 8162 2983
rect 8190 2842 8218 3262
rect 8190 2809 8218 2814
rect 8358 3290 8386 3295
rect 8152 2758 8284 2763
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8152 2725 8284 2730
rect 8246 2562 8274 2567
rect 8246 2561 8330 2562
rect 8246 2535 8247 2561
rect 8273 2535 8330 2561
rect 8246 2534 8330 2535
rect 8246 2529 8274 2534
rect 8134 2506 8162 2511
rect 8134 2459 8162 2478
rect 8302 2450 8330 2534
rect 8302 2417 8330 2422
rect 8134 2394 8162 2399
rect 8134 2225 8162 2366
rect 8134 2199 8135 2225
rect 8161 2199 8162 2225
rect 8134 2193 8162 2199
rect 8152 1974 8284 1979
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8152 1941 8284 1946
rect 8302 1890 8330 1895
rect 8134 1778 8162 1797
rect 8134 1745 8162 1750
rect 7910 1582 7994 1610
rect 8022 1666 8050 1671
rect 8078 1666 8162 1694
rect 7910 400 7938 1582
rect 8022 400 8050 1638
rect 8134 400 8162 1666
rect 8246 1610 8274 1615
rect 8246 400 8274 1582
rect 8302 1554 8330 1862
rect 8358 1666 8386 3262
rect 8358 1633 8386 1638
rect 8302 1526 8386 1554
rect 8358 400 8386 1526
rect 8470 400 8498 4102
rect 8694 4097 8722 4102
rect 8862 4097 8890 4102
rect 8974 4129 9002 4135
rect 8974 4103 8975 4129
rect 9001 4103 9002 4129
rect 8974 3346 9002 4103
rect 9230 3934 9362 3939
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9230 3901 9362 3906
rect 8694 3290 8722 3295
rect 8694 3243 8722 3262
rect 8862 3290 8890 3295
rect 8974 3280 9002 3318
rect 8862 3243 8890 3262
rect 9230 3150 9362 3155
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9230 3117 9362 3122
rect 8750 2561 8778 2567
rect 8750 2535 8751 2561
rect 8777 2535 8778 2561
rect 8526 2506 8554 2511
rect 8694 2506 8722 2511
rect 8526 2505 8722 2506
rect 8526 2479 8527 2505
rect 8553 2479 8695 2505
rect 8721 2479 8722 2505
rect 8526 2478 8722 2479
rect 8526 2058 8554 2478
rect 8694 2473 8722 2478
rect 8750 2450 8778 2535
rect 8750 2417 8778 2422
rect 9230 2366 9362 2371
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9230 2333 9362 2338
rect 8526 2025 8554 2030
rect 8974 1778 9002 1783
rect 8750 1722 8778 1741
rect 8750 1689 8778 1694
rect 8918 1722 8946 1741
rect 8974 1731 9002 1750
rect 8918 1689 8946 1694
rect 9230 1582 9362 1587
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9230 1549 9362 1554
rect 1400 0 1456 400
rect 1512 0 1568 400
rect 1624 0 1680 400
rect 1736 0 1792 400
rect 1848 0 1904 400
rect 1960 0 2016 400
rect 2072 0 2128 400
rect 2184 0 2240 400
rect 2296 0 2352 400
rect 2408 0 2464 400
rect 2520 0 2576 400
rect 2632 0 2688 400
rect 2744 0 2800 400
rect 2856 0 2912 400
rect 2968 0 3024 400
rect 3080 0 3136 400
rect 3192 0 3248 400
rect 3304 0 3360 400
rect 3416 0 3472 400
rect 3528 0 3584 400
rect 3640 0 3696 400
rect 3752 0 3808 400
rect 3864 0 3920 400
rect 3976 0 4032 400
rect 4088 0 4144 400
rect 4200 0 4256 400
rect 4312 0 4368 400
rect 4424 0 4480 400
rect 4536 0 4592 400
rect 4648 0 4704 400
rect 4760 0 4816 400
rect 4872 0 4928 400
rect 4984 0 5040 400
rect 5096 0 5152 400
rect 5208 0 5264 400
rect 5320 0 5376 400
rect 5432 0 5488 400
rect 5544 0 5600 400
rect 5656 0 5712 400
rect 5768 0 5824 400
rect 5880 0 5936 400
rect 5992 0 6048 400
rect 6104 0 6160 400
rect 6216 0 6272 400
rect 6328 0 6384 400
rect 6440 0 6496 400
rect 6552 0 6608 400
rect 6664 0 6720 400
rect 6776 0 6832 400
rect 6888 0 6944 400
rect 7000 0 7056 400
rect 7112 0 7168 400
rect 7224 0 7280 400
rect 7336 0 7392 400
rect 7448 0 7504 400
rect 7560 0 7616 400
rect 7672 0 7728 400
rect 7784 0 7840 400
rect 7896 0 7952 400
rect 8008 0 8064 400
rect 8120 0 8176 400
rect 8232 0 8288 400
rect 8344 0 8400 400
rect 8456 0 8512 400
<< via2 >>
rect 1684 4325 1712 4326
rect 1684 4299 1685 4325
rect 1685 4299 1711 4325
rect 1711 4299 1712 4325
rect 1684 4298 1712 4299
rect 1736 4325 1764 4326
rect 1736 4299 1737 4325
rect 1737 4299 1763 4325
rect 1763 4299 1764 4325
rect 1736 4298 1764 4299
rect 1788 4325 1816 4326
rect 1788 4299 1789 4325
rect 1789 4299 1815 4325
rect 1815 4299 1816 4325
rect 1788 4298 1816 4299
rect 3840 4325 3868 4326
rect 3840 4299 3841 4325
rect 3841 4299 3867 4325
rect 3867 4299 3868 4325
rect 3840 4298 3868 4299
rect 3892 4325 3920 4326
rect 3892 4299 3893 4325
rect 3893 4299 3919 4325
rect 3919 4299 3920 4325
rect 3892 4298 3920 4299
rect 3944 4325 3972 4326
rect 3944 4299 3945 4325
rect 3945 4299 3971 4325
rect 3971 4299 3972 4325
rect 3944 4298 3972 4299
rect 5996 4325 6024 4326
rect 5996 4299 5997 4325
rect 5997 4299 6023 4325
rect 6023 4299 6024 4325
rect 5996 4298 6024 4299
rect 6048 4325 6076 4326
rect 6048 4299 6049 4325
rect 6049 4299 6075 4325
rect 6075 4299 6076 4325
rect 6048 4298 6076 4299
rect 6100 4325 6128 4326
rect 6100 4299 6101 4325
rect 6101 4299 6127 4325
rect 6127 4299 6128 4325
rect 6100 4298 6128 4299
rect 8152 4325 8180 4326
rect 8152 4299 8153 4325
rect 8153 4299 8179 4325
rect 8179 4299 8180 4325
rect 8152 4298 8180 4299
rect 8204 4325 8232 4326
rect 8204 4299 8205 4325
rect 8205 4299 8231 4325
rect 8231 4299 8232 4325
rect 8204 4298 8232 4299
rect 8256 4325 8284 4326
rect 8256 4299 8257 4325
rect 8257 4299 8283 4325
rect 8283 4299 8284 4325
rect 8256 4298 8284 4299
rect 1918 3822 1946 3850
rect 2762 3933 2790 3934
rect 2762 3907 2763 3933
rect 2763 3907 2789 3933
rect 2789 3907 2790 3933
rect 2762 3906 2790 3907
rect 2814 3933 2842 3934
rect 2814 3907 2815 3933
rect 2815 3907 2841 3933
rect 2841 3907 2842 3933
rect 2814 3906 2842 3907
rect 2866 3933 2894 3934
rect 2866 3907 2867 3933
rect 2867 3907 2893 3933
rect 2893 3907 2894 3933
rect 2866 3906 2894 3907
rect 1684 3541 1712 3542
rect 1684 3515 1685 3541
rect 1685 3515 1711 3541
rect 1711 3515 1712 3541
rect 1684 3514 1712 3515
rect 1736 3541 1764 3542
rect 1736 3515 1737 3541
rect 1737 3515 1763 3541
rect 1763 3515 1764 3541
rect 1736 3514 1764 3515
rect 1788 3541 1816 3542
rect 1788 3515 1789 3541
rect 1789 3515 1815 3541
rect 1815 3515 1816 3541
rect 1788 3514 1816 3515
rect 1078 3345 1106 3346
rect 1078 3319 1079 3345
rect 1079 3319 1105 3345
rect 1105 3319 1106 3345
rect 1078 3318 1106 3319
rect 1414 3318 1442 3346
rect 1078 2561 1106 2562
rect 1078 2535 1079 2561
rect 1079 2535 1105 2561
rect 1105 2535 1106 2561
rect 1078 2534 1106 2535
rect 1414 3009 1442 3010
rect 1414 2983 1415 3009
rect 1415 2983 1441 3009
rect 1441 2983 1442 3009
rect 1414 2982 1442 2983
rect 1414 2534 1442 2562
rect 1358 2254 1386 2282
rect 1134 1806 1162 1834
rect 1414 1750 1442 1778
rect 1190 1721 1218 1722
rect 1190 1695 1191 1721
rect 1191 1695 1217 1721
rect 1217 1695 1218 1721
rect 1190 1694 1218 1695
rect 1358 1721 1386 1722
rect 1358 1695 1359 1721
rect 1359 1695 1385 1721
rect 1385 1695 1386 1721
rect 1358 1694 1386 1695
rect 2086 3822 2114 3850
rect 1638 3345 1666 3346
rect 1638 3319 1639 3345
rect 1639 3319 1665 3345
rect 1665 3319 1666 3345
rect 1638 3318 1666 3319
rect 1750 3289 1778 3290
rect 1750 3263 1751 3289
rect 1751 3263 1777 3289
rect 1777 3263 1778 3289
rect 1750 3262 1778 3263
rect 1918 3318 1946 3346
rect 1974 3262 2002 3290
rect 1582 2814 1610 2842
rect 1750 2814 1778 2842
rect 1684 2757 1712 2758
rect 1684 2731 1685 2757
rect 1685 2731 1711 2757
rect 1711 2731 1712 2757
rect 1684 2730 1712 2731
rect 1736 2757 1764 2758
rect 1736 2731 1737 2757
rect 1737 2731 1763 2757
rect 1763 2731 1764 2757
rect 1736 2730 1764 2731
rect 1788 2757 1816 2758
rect 1788 2731 1789 2757
rect 1789 2731 1815 2757
rect 1815 2731 1816 2757
rect 1788 2730 1816 2731
rect 1638 2561 1666 2562
rect 1638 2535 1639 2561
rect 1639 2535 1665 2561
rect 1665 2535 1666 2561
rect 1638 2534 1666 2535
rect 1750 2505 1778 2506
rect 1750 2479 1751 2505
rect 1751 2479 1777 2505
rect 1777 2479 1778 2505
rect 1750 2478 1778 2479
rect 1582 2169 1610 2170
rect 1582 2143 1583 2169
rect 1583 2143 1609 2169
rect 1609 2143 1610 2169
rect 1582 2142 1610 2143
rect 1750 2169 1778 2170
rect 1750 2143 1751 2169
rect 1751 2143 1777 2169
rect 1777 2143 1778 2169
rect 1750 2142 1778 2143
rect 1750 2030 1778 2058
rect 1684 1973 1712 1974
rect 1684 1947 1685 1973
rect 1685 1947 1711 1973
rect 1711 1947 1712 1973
rect 1684 1946 1712 1947
rect 1736 1973 1764 1974
rect 1736 1947 1737 1973
rect 1737 1947 1763 1973
rect 1763 1947 1764 1973
rect 1736 1946 1764 1947
rect 1788 1973 1816 1974
rect 1788 1947 1789 1973
rect 1789 1947 1815 1973
rect 1815 1947 1816 1973
rect 1788 1946 1816 1947
rect 1582 1862 1610 1890
rect 1694 1806 1722 1834
rect 1638 1777 1666 1778
rect 1638 1751 1639 1777
rect 1639 1751 1665 1777
rect 1665 1751 1666 1777
rect 1638 1750 1666 1751
rect 1806 1777 1834 1778
rect 1806 1751 1807 1777
rect 1807 1751 1833 1777
rect 1833 1751 1834 1777
rect 1806 1750 1834 1751
rect 1974 3009 2002 3010
rect 1974 2983 1975 3009
rect 1975 2983 2001 3009
rect 2001 2983 2002 3009
rect 1974 2982 2002 2983
rect 1974 2534 2002 2562
rect 1918 2505 1946 2506
rect 1918 2479 1919 2505
rect 1919 2479 1945 2505
rect 1945 2479 1946 2505
rect 1918 2478 1946 2479
rect 2198 3345 2226 3346
rect 2198 3319 2199 3345
rect 2199 3319 2225 3345
rect 2225 3319 2226 3345
rect 2198 3318 2226 3319
rect 2086 2169 2114 2170
rect 2086 2143 2087 2169
rect 2087 2143 2113 2169
rect 2113 2143 2114 2169
rect 2086 2142 2114 2143
rect 1918 1777 1946 1778
rect 1918 1751 1919 1777
rect 1919 1751 1945 1777
rect 1945 1751 1946 1777
rect 1918 1750 1946 1751
rect 2142 1862 2170 1890
rect 2198 2561 2226 2562
rect 2198 2535 2199 2561
rect 2199 2535 2225 2561
rect 2225 2535 2226 2561
rect 2198 2534 2226 2535
rect 2086 1806 2114 1834
rect 2310 2505 2338 2506
rect 2310 2479 2311 2505
rect 2311 2479 2337 2505
rect 2337 2479 2338 2505
rect 2310 2478 2338 2479
rect 2254 2366 2282 2394
rect 2254 2254 2282 2282
rect 2310 2169 2338 2170
rect 2310 2143 2311 2169
rect 2311 2143 2337 2169
rect 2337 2143 2338 2169
rect 2310 2142 2338 2143
rect 2310 1862 2338 1890
rect 3840 3541 3868 3542
rect 3840 3515 3841 3541
rect 3841 3515 3867 3541
rect 3867 3515 3868 3541
rect 3840 3514 3868 3515
rect 3892 3541 3920 3542
rect 3892 3515 3893 3541
rect 3893 3515 3919 3541
rect 3919 3515 3920 3541
rect 3892 3514 3920 3515
rect 3944 3541 3972 3542
rect 3944 3515 3945 3541
rect 3945 3515 3971 3541
rect 3971 3515 3972 3541
rect 3944 3514 3972 3515
rect 2762 3149 2790 3150
rect 2762 3123 2763 3149
rect 2763 3123 2789 3149
rect 2789 3123 2790 3149
rect 2762 3122 2790 3123
rect 2814 3149 2842 3150
rect 2814 3123 2815 3149
rect 2815 3123 2841 3149
rect 2841 3123 2842 3149
rect 2814 3122 2842 3123
rect 2866 3149 2894 3150
rect 2866 3123 2867 3149
rect 2867 3123 2893 3149
rect 2893 3123 2894 3149
rect 2866 3122 2894 3123
rect 2534 3009 2562 3010
rect 2534 2983 2535 3009
rect 2535 2983 2561 3009
rect 2561 2983 2562 3009
rect 2534 2982 2562 2983
rect 2534 2534 2562 2562
rect 2478 2505 2506 2506
rect 2478 2479 2479 2505
rect 2479 2479 2505 2505
rect 2505 2479 2506 2505
rect 2478 2478 2506 2479
rect 2478 2366 2506 2394
rect 2926 2478 2954 2506
rect 2646 2422 2674 2450
rect 2478 1862 2506 1890
rect 2762 2365 2790 2366
rect 2762 2339 2763 2365
rect 2763 2339 2789 2365
rect 2789 2339 2790 2365
rect 2762 2338 2790 2339
rect 2814 2365 2842 2366
rect 2814 2339 2815 2365
rect 2815 2339 2841 2365
rect 2841 2339 2842 2365
rect 2814 2338 2842 2339
rect 2866 2365 2894 2366
rect 2866 2339 2867 2365
rect 2867 2339 2893 2365
rect 2893 2339 2894 2365
rect 2866 2338 2894 2339
rect 2702 2030 2730 2058
rect 2870 2030 2898 2058
rect 2926 1806 2954 1834
rect 2926 1694 2954 1722
rect 2762 1581 2790 1582
rect 2762 1555 2763 1581
rect 2763 1555 2789 1581
rect 2789 1555 2790 1581
rect 2762 1554 2790 1555
rect 2814 1581 2842 1582
rect 2814 1555 2815 1581
rect 2815 1555 2841 1581
rect 2841 1555 2842 1581
rect 2814 1554 2842 1555
rect 2866 1581 2894 1582
rect 2866 1555 2867 1581
rect 2867 1555 2893 1581
rect 2893 1555 2894 1581
rect 2866 1554 2894 1555
rect 3262 2953 3290 2954
rect 3262 2927 3263 2953
rect 3263 2927 3289 2953
rect 3289 2927 3290 2953
rect 3262 2926 3290 2927
rect 3374 2953 3402 2954
rect 3374 2927 3375 2953
rect 3375 2927 3401 2953
rect 3401 2927 3402 2953
rect 3374 2926 3402 2927
rect 3038 2561 3066 2562
rect 3038 2535 3039 2561
rect 3039 2535 3065 2561
rect 3065 2535 3066 2561
rect 3038 2534 3066 2535
rect 3318 2366 3346 2394
rect 3150 2142 3178 2170
rect 3094 1806 3122 1834
rect 3262 2169 3290 2170
rect 3262 2143 3263 2169
rect 3263 2143 3289 2169
rect 3289 2143 3290 2169
rect 3262 2142 3290 2143
rect 3374 2169 3402 2170
rect 3374 2143 3375 2169
rect 3375 2143 3401 2169
rect 3401 2143 3402 2169
rect 3374 2142 3402 2143
rect 3318 1806 3346 1834
rect 3206 1638 3234 1666
rect 3542 2926 3570 2954
rect 4494 3206 4522 3234
rect 4918 3933 4946 3934
rect 4918 3907 4919 3933
rect 4919 3907 4945 3933
rect 4945 3907 4946 3933
rect 4918 3906 4946 3907
rect 4970 3933 4998 3934
rect 4970 3907 4971 3933
rect 4971 3907 4997 3933
rect 4997 3907 4998 3933
rect 4970 3906 4998 3907
rect 5022 3933 5050 3934
rect 5022 3907 5023 3933
rect 5023 3907 5049 3933
rect 5049 3907 5050 3933
rect 5022 3906 5050 3907
rect 7074 3933 7102 3934
rect 7074 3907 7075 3933
rect 7075 3907 7101 3933
rect 7101 3907 7102 3933
rect 7074 3906 7102 3907
rect 7126 3933 7154 3934
rect 7126 3907 7127 3933
rect 7127 3907 7153 3933
rect 7153 3907 7154 3933
rect 7126 3906 7154 3907
rect 7178 3933 7206 3934
rect 7178 3907 7179 3933
rect 7179 3907 7205 3933
rect 7205 3907 7206 3933
rect 7178 3906 7206 3907
rect 7238 3737 7266 3738
rect 7238 3711 7239 3737
rect 7239 3711 7265 3737
rect 7265 3711 7266 3737
rect 7238 3710 7266 3711
rect 5996 3541 6024 3542
rect 5996 3515 5997 3541
rect 5997 3515 6023 3541
rect 6023 3515 6024 3541
rect 5996 3514 6024 3515
rect 6048 3541 6076 3542
rect 6048 3515 6049 3541
rect 6049 3515 6075 3541
rect 6075 3515 6076 3541
rect 6048 3514 6076 3515
rect 6100 3541 6128 3542
rect 6100 3515 6101 3541
rect 6101 3515 6127 3541
rect 6127 3515 6128 3541
rect 6100 3514 6128 3515
rect 4830 3206 4858 3234
rect 4918 3149 4946 3150
rect 4918 3123 4919 3149
rect 4919 3123 4945 3149
rect 4945 3123 4946 3149
rect 4918 3122 4946 3123
rect 4970 3149 4998 3150
rect 4970 3123 4971 3149
rect 4971 3123 4997 3149
rect 4997 3123 4998 3149
rect 4970 3122 4998 3123
rect 5022 3149 5050 3150
rect 5022 3123 5023 3149
rect 5023 3123 5049 3149
rect 5049 3123 5050 3149
rect 5022 3122 5050 3123
rect 3840 2757 3868 2758
rect 3840 2731 3841 2757
rect 3841 2731 3867 2757
rect 3867 2731 3868 2757
rect 3840 2730 3868 2731
rect 3892 2757 3920 2758
rect 3892 2731 3893 2757
rect 3893 2731 3919 2757
rect 3919 2731 3920 2757
rect 3892 2730 3920 2731
rect 3944 2757 3972 2758
rect 3944 2731 3945 2757
rect 3945 2731 3971 2757
rect 3971 2731 3972 2757
rect 3944 2730 3972 2731
rect 3598 2561 3626 2562
rect 3598 2535 3599 2561
rect 3599 2535 3625 2561
rect 3625 2535 3626 2561
rect 3598 2534 3626 2535
rect 3710 2366 3738 2394
rect 3654 2030 3682 2058
rect 3822 2086 3850 2114
rect 3990 2086 4018 2114
rect 3878 2030 3906 2058
rect 3840 1973 3868 1974
rect 3840 1947 3841 1973
rect 3841 1947 3867 1973
rect 3867 1947 3868 1973
rect 3840 1946 3868 1947
rect 3892 1973 3920 1974
rect 3892 1947 3893 1973
rect 3893 1947 3919 1973
rect 3919 1947 3920 1973
rect 3892 1946 3920 1947
rect 3944 1973 3972 1974
rect 3944 1947 3945 1973
rect 3945 1947 3971 1973
rect 3971 1947 3972 1973
rect 3944 1946 3972 1947
rect 4214 2561 4242 2562
rect 4214 2535 4215 2561
rect 4215 2535 4241 2561
rect 4241 2535 4242 2561
rect 4214 2534 4242 2535
rect 4270 2505 4298 2506
rect 4270 2479 4271 2505
rect 4271 2479 4297 2505
rect 4297 2479 4298 2505
rect 4270 2478 4298 2479
rect 4214 2225 4242 2226
rect 4214 2199 4215 2225
rect 4215 2199 4241 2225
rect 4241 2199 4242 2225
rect 4214 2198 4242 2199
rect 3878 1862 3906 1890
rect 3766 1777 3794 1778
rect 3766 1751 3767 1777
rect 3767 1751 3793 1777
rect 3793 1751 3794 1777
rect 3766 1750 3794 1751
rect 4102 2142 4130 2170
rect 3934 1777 3962 1778
rect 3934 1751 3935 1777
rect 3935 1751 3961 1777
rect 3961 1751 3962 1777
rect 3934 1750 3962 1751
rect 4326 2169 4354 2170
rect 4326 2143 4327 2169
rect 4327 2143 4353 2169
rect 4353 2143 4354 2169
rect 4326 2142 4354 2143
rect 4214 2030 4242 2058
rect 7182 3345 7210 3346
rect 7182 3319 7183 3345
rect 7183 3319 7209 3345
rect 7209 3319 7210 3345
rect 7182 3318 7210 3319
rect 7350 3345 7378 3346
rect 7350 3319 7351 3345
rect 7351 3319 7377 3345
rect 7377 3319 7378 3345
rect 7350 3318 7378 3319
rect 7798 3737 7826 3738
rect 7798 3711 7799 3737
rect 7799 3711 7825 3737
rect 7825 3711 7826 3737
rect 7798 3710 7826 3711
rect 7854 3345 7882 3346
rect 7854 3319 7855 3345
rect 7855 3319 7881 3345
rect 7881 3319 7882 3345
rect 7854 3318 7882 3319
rect 7074 3149 7102 3150
rect 7074 3123 7075 3149
rect 7075 3123 7101 3149
rect 7101 3123 7102 3149
rect 7074 3122 7102 3123
rect 7126 3149 7154 3150
rect 7126 3123 7127 3149
rect 7127 3123 7153 3149
rect 7153 3123 7154 3149
rect 7126 3122 7154 3123
rect 7178 3149 7206 3150
rect 7178 3123 7179 3149
rect 7179 3123 7205 3149
rect 7205 3123 7206 3149
rect 7178 3122 7206 3123
rect 7574 3038 7602 3066
rect 4494 2814 4522 2842
rect 4438 2505 4466 2506
rect 4438 2479 4439 2505
rect 4439 2479 4465 2505
rect 4465 2479 4466 2505
rect 4438 2478 4466 2479
rect 4270 1721 4298 1722
rect 4270 1695 4271 1721
rect 4271 1695 4297 1721
rect 4297 1695 4298 1721
rect 4270 1694 4298 1695
rect 4438 1721 4466 1722
rect 4438 1695 4439 1721
rect 4439 1695 4465 1721
rect 4465 1695 4466 1721
rect 4438 1694 4466 1695
rect 4830 2814 4858 2842
rect 4718 2198 4746 2226
rect 4774 2478 4802 2506
rect 4550 2169 4578 2170
rect 4550 2143 4551 2169
rect 4551 2143 4577 2169
rect 4577 2143 4578 2169
rect 4550 2142 4578 2143
rect 4550 1806 4578 1834
rect 4606 1414 4634 1442
rect 4662 2086 4690 2114
rect 4918 2365 4946 2366
rect 4918 2339 4919 2365
rect 4919 2339 4945 2365
rect 4945 2339 4946 2365
rect 4918 2338 4946 2339
rect 4970 2365 4998 2366
rect 4970 2339 4971 2365
rect 4971 2339 4997 2365
rect 4997 2339 4998 2365
rect 4970 2338 4998 2339
rect 5022 2365 5050 2366
rect 5022 2339 5023 2365
rect 5023 2339 5049 2365
rect 5049 2339 5050 2365
rect 5022 2338 5050 2339
rect 5054 2225 5082 2226
rect 5054 2199 5055 2225
rect 5055 2199 5081 2225
rect 5081 2199 5082 2225
rect 5054 2198 5082 2199
rect 4830 1750 4858 1778
rect 4918 1581 4946 1582
rect 4918 1555 4919 1581
rect 4919 1555 4945 1581
rect 4945 1555 4946 1581
rect 4918 1554 4946 1555
rect 4970 1581 4998 1582
rect 4970 1555 4971 1581
rect 4971 1555 4997 1581
rect 4997 1555 4998 1581
rect 4970 1554 4998 1555
rect 5022 1581 5050 1582
rect 5022 1555 5023 1581
rect 5023 1555 5049 1581
rect 5049 1555 5050 1581
rect 5022 1554 5050 1555
rect 4998 1414 5026 1442
rect 5996 2757 6024 2758
rect 5996 2731 5997 2757
rect 5997 2731 6023 2757
rect 6023 2731 6024 2757
rect 5996 2730 6024 2731
rect 6048 2757 6076 2758
rect 6048 2731 6049 2757
rect 6049 2731 6075 2757
rect 6075 2731 6076 2757
rect 6048 2730 6076 2731
rect 6100 2757 6128 2758
rect 6100 2731 6101 2757
rect 6101 2731 6127 2757
rect 6127 2731 6128 2757
rect 6100 2730 6128 2731
rect 5166 2198 5194 2226
rect 5222 2169 5250 2170
rect 5222 2143 5223 2169
rect 5223 2143 5249 2169
rect 5249 2143 5250 2169
rect 5222 2142 5250 2143
rect 5222 1694 5250 1722
rect 5558 2198 5586 2226
rect 5894 2225 5922 2226
rect 5894 2199 5895 2225
rect 5895 2199 5921 2225
rect 5921 2199 5922 2225
rect 5894 2198 5922 2199
rect 6174 2198 6202 2226
rect 5390 2169 5418 2170
rect 5390 2143 5391 2169
rect 5391 2143 5417 2169
rect 5417 2143 5418 2169
rect 5390 2142 5418 2143
rect 5334 1777 5362 1778
rect 5334 1751 5335 1777
rect 5335 1751 5361 1777
rect 5361 1751 5362 1777
rect 5334 1750 5362 1751
rect 5502 1777 5530 1778
rect 5502 1751 5503 1777
rect 5503 1751 5529 1777
rect 5529 1751 5530 1777
rect 5502 1750 5530 1751
rect 6118 2169 6146 2170
rect 6118 2143 6119 2169
rect 6119 2143 6145 2169
rect 6145 2143 6146 2169
rect 6118 2142 6146 2143
rect 5996 1973 6024 1974
rect 5996 1947 5997 1973
rect 5997 1947 6023 1973
rect 6023 1947 6024 1973
rect 5996 1946 6024 1947
rect 6048 1973 6076 1974
rect 6048 1947 6049 1973
rect 6049 1947 6075 1973
rect 6075 1947 6076 1973
rect 6048 1946 6076 1947
rect 6100 1973 6128 1974
rect 6100 1947 6101 1973
rect 6101 1947 6127 1973
rect 6127 1947 6128 1973
rect 6100 1946 6128 1947
rect 6062 1694 6090 1722
rect 6454 2225 6482 2226
rect 6454 2199 6455 2225
rect 6455 2199 6481 2225
rect 6481 2199 6482 2225
rect 6454 2198 6482 2199
rect 6510 2478 6538 2506
rect 6286 2169 6314 2170
rect 6286 2143 6287 2169
rect 6287 2143 6313 2169
rect 6313 2143 6314 2169
rect 6286 2142 6314 2143
rect 6846 2505 6874 2506
rect 6846 2479 6847 2505
rect 6847 2479 6873 2505
rect 6873 2479 6874 2505
rect 6846 2478 6874 2479
rect 6286 2030 6314 2058
rect 6566 2142 6594 2170
rect 6342 1750 6370 1778
rect 6734 2030 6762 2058
rect 6678 1806 6706 1834
rect 6790 1721 6818 1722
rect 6790 1695 6791 1721
rect 6791 1695 6817 1721
rect 6817 1695 6818 1721
rect 6790 1694 6818 1695
rect 7014 2505 7042 2506
rect 7014 2479 7015 2505
rect 7015 2479 7041 2505
rect 7041 2479 7042 2505
rect 7014 2478 7042 2479
rect 7074 2365 7102 2366
rect 7074 2339 7075 2365
rect 7075 2339 7101 2365
rect 7101 2339 7102 2365
rect 7074 2338 7102 2339
rect 7126 2365 7154 2366
rect 7126 2339 7127 2365
rect 7127 2339 7153 2365
rect 7153 2339 7154 2365
rect 7126 2338 7154 2339
rect 7178 2365 7206 2366
rect 7178 2339 7179 2365
rect 7179 2339 7205 2365
rect 7205 2339 7206 2365
rect 7178 2338 7206 2339
rect 6958 2198 6986 2226
rect 6902 2030 6930 2058
rect 7014 2030 7042 2058
rect 6902 1918 6930 1946
rect 6958 1721 6986 1722
rect 6958 1695 6959 1721
rect 6959 1695 6985 1721
rect 6985 1695 6986 1721
rect 6958 1694 6986 1695
rect 7074 1581 7102 1582
rect 7074 1555 7075 1581
rect 7075 1555 7101 1581
rect 7101 1555 7102 1581
rect 7074 1554 7102 1555
rect 7126 1581 7154 1582
rect 7126 1555 7127 1581
rect 7127 1555 7153 1581
rect 7153 1555 7154 1581
rect 7126 1554 7154 1555
rect 7178 1581 7206 1582
rect 7178 1555 7179 1581
rect 7179 1555 7205 1581
rect 7205 1555 7206 1581
rect 7178 1554 7206 1555
rect 7350 2814 7378 2842
rect 7294 2169 7322 2170
rect 7294 2143 7295 2169
rect 7295 2143 7321 2169
rect 7321 2143 7322 2169
rect 7294 2142 7322 2143
rect 7518 2366 7546 2394
rect 7462 2169 7490 2170
rect 7462 2143 7463 2169
rect 7463 2143 7489 2169
rect 7489 2143 7490 2169
rect 7462 2142 7490 2143
rect 7406 2030 7434 2058
rect 7294 1777 7322 1778
rect 7294 1751 7295 1777
rect 7295 1751 7321 1777
rect 7321 1751 7322 1777
rect 7294 1750 7322 1751
rect 7350 1694 7378 1722
rect 7462 1777 7490 1778
rect 7462 1751 7463 1777
rect 7463 1751 7489 1777
rect 7489 1751 7490 1777
rect 7462 1750 7490 1751
rect 7462 1302 7490 1330
rect 7574 2225 7602 2226
rect 7574 2199 7575 2225
rect 7575 2199 7601 2225
rect 7601 2199 7602 2225
rect 7574 2198 7602 2199
rect 7574 2030 7602 2058
rect 7462 1022 7490 1050
rect 7630 1862 7658 1890
rect 7686 3038 7714 3066
rect 7686 2422 7714 2450
rect 7686 2198 7714 2226
rect 7686 1750 7714 1778
rect 7854 3038 7882 3066
rect 7798 2814 7826 2842
rect 7910 2814 7938 2842
rect 7798 2169 7826 2170
rect 7798 2143 7799 2169
rect 7799 2143 7825 2169
rect 7825 2143 7826 2169
rect 7798 2142 7826 2143
rect 7798 1918 7826 1946
rect 7854 1806 7882 1834
rect 7966 2505 7994 2506
rect 7966 2479 7967 2505
rect 7967 2479 7993 2505
rect 7993 2479 7994 2505
rect 7966 2478 7994 2479
rect 7966 2169 7994 2170
rect 7966 2143 7967 2169
rect 7967 2143 7993 2169
rect 7993 2143 7994 2169
rect 7966 2142 7994 2143
rect 8022 1806 8050 1834
rect 8152 3541 8180 3542
rect 8152 3515 8153 3541
rect 8153 3515 8179 3541
rect 8179 3515 8180 3541
rect 8152 3514 8180 3515
rect 8204 3541 8232 3542
rect 8204 3515 8205 3541
rect 8205 3515 8231 3541
rect 8231 3515 8232 3541
rect 8204 3514 8232 3515
rect 8256 3541 8284 3542
rect 8256 3515 8257 3541
rect 8257 3515 8283 3541
rect 8283 3515 8284 3541
rect 8256 3514 8284 3515
rect 8414 3345 8442 3346
rect 8414 3319 8415 3345
rect 8415 3319 8441 3345
rect 8441 3319 8442 3345
rect 8414 3318 8442 3319
rect 8134 3038 8162 3066
rect 8190 2814 8218 2842
rect 8358 3262 8386 3290
rect 8152 2757 8180 2758
rect 8152 2731 8153 2757
rect 8153 2731 8179 2757
rect 8179 2731 8180 2757
rect 8152 2730 8180 2731
rect 8204 2757 8232 2758
rect 8204 2731 8205 2757
rect 8205 2731 8231 2757
rect 8231 2731 8232 2757
rect 8204 2730 8232 2731
rect 8256 2757 8284 2758
rect 8256 2731 8257 2757
rect 8257 2731 8283 2757
rect 8283 2731 8284 2757
rect 8256 2730 8284 2731
rect 8134 2505 8162 2506
rect 8134 2479 8135 2505
rect 8135 2479 8161 2505
rect 8161 2479 8162 2505
rect 8134 2478 8162 2479
rect 8302 2422 8330 2450
rect 8134 2366 8162 2394
rect 8152 1973 8180 1974
rect 8152 1947 8153 1973
rect 8153 1947 8179 1973
rect 8179 1947 8180 1973
rect 8152 1946 8180 1947
rect 8204 1973 8232 1974
rect 8204 1947 8205 1973
rect 8205 1947 8231 1973
rect 8231 1947 8232 1973
rect 8204 1946 8232 1947
rect 8256 1973 8284 1974
rect 8256 1947 8257 1973
rect 8257 1947 8283 1973
rect 8283 1947 8284 1973
rect 8256 1946 8284 1947
rect 8302 1862 8330 1890
rect 8134 1777 8162 1778
rect 8134 1751 8135 1777
rect 8135 1751 8161 1777
rect 8161 1751 8162 1777
rect 8134 1750 8162 1751
rect 8022 1638 8050 1666
rect 8246 1582 8274 1610
rect 8358 1638 8386 1666
rect 9230 3933 9258 3934
rect 9230 3907 9231 3933
rect 9231 3907 9257 3933
rect 9257 3907 9258 3933
rect 9230 3906 9258 3907
rect 9282 3933 9310 3934
rect 9282 3907 9283 3933
rect 9283 3907 9309 3933
rect 9309 3907 9310 3933
rect 9282 3906 9310 3907
rect 9334 3933 9362 3934
rect 9334 3907 9335 3933
rect 9335 3907 9361 3933
rect 9361 3907 9362 3933
rect 9334 3906 9362 3907
rect 8974 3345 9002 3346
rect 8974 3319 8975 3345
rect 8975 3319 9001 3345
rect 9001 3319 9002 3345
rect 8974 3318 9002 3319
rect 8694 3289 8722 3290
rect 8694 3263 8695 3289
rect 8695 3263 8721 3289
rect 8721 3263 8722 3289
rect 8694 3262 8722 3263
rect 8862 3289 8890 3290
rect 8862 3263 8863 3289
rect 8863 3263 8889 3289
rect 8889 3263 8890 3289
rect 8862 3262 8890 3263
rect 9230 3149 9258 3150
rect 9230 3123 9231 3149
rect 9231 3123 9257 3149
rect 9257 3123 9258 3149
rect 9230 3122 9258 3123
rect 9282 3149 9310 3150
rect 9282 3123 9283 3149
rect 9283 3123 9309 3149
rect 9309 3123 9310 3149
rect 9282 3122 9310 3123
rect 9334 3149 9362 3150
rect 9334 3123 9335 3149
rect 9335 3123 9361 3149
rect 9361 3123 9362 3149
rect 9334 3122 9362 3123
rect 8750 2422 8778 2450
rect 9230 2365 9258 2366
rect 9230 2339 9231 2365
rect 9231 2339 9257 2365
rect 9257 2339 9258 2365
rect 9230 2338 9258 2339
rect 9282 2365 9310 2366
rect 9282 2339 9283 2365
rect 9283 2339 9309 2365
rect 9309 2339 9310 2365
rect 9282 2338 9310 2339
rect 9334 2365 9362 2366
rect 9334 2339 9335 2365
rect 9335 2339 9361 2365
rect 9361 2339 9362 2365
rect 9334 2338 9362 2339
rect 8526 2030 8554 2058
rect 8974 1777 9002 1778
rect 8974 1751 8975 1777
rect 8975 1751 9001 1777
rect 9001 1751 9002 1777
rect 8974 1750 9002 1751
rect 8750 1721 8778 1722
rect 8750 1695 8751 1721
rect 8751 1695 8777 1721
rect 8777 1695 8778 1721
rect 8750 1694 8778 1695
rect 8918 1721 8946 1722
rect 8918 1695 8919 1721
rect 8919 1695 8945 1721
rect 8945 1695 8946 1721
rect 8918 1694 8946 1695
rect 9230 1581 9258 1582
rect 9230 1555 9231 1581
rect 9231 1555 9257 1581
rect 9257 1555 9258 1581
rect 9230 1554 9258 1555
rect 9282 1581 9310 1582
rect 9282 1555 9283 1581
rect 9283 1555 9309 1581
rect 9309 1555 9310 1581
rect 9282 1554 9310 1555
rect 9334 1581 9362 1582
rect 9334 1555 9335 1581
rect 9335 1555 9361 1581
rect 9361 1555 9362 1581
rect 9334 1554 9362 1555
<< metal3 >>
rect 1679 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1821 4326
rect 3835 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3977 4326
rect 5991 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6133 4326
rect 8147 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8289 4326
rect 2757 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2899 3934
rect 4913 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5055 3934
rect 7069 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7211 3934
rect 9225 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9367 3934
rect 1913 3822 1918 3850
rect 1946 3822 2086 3850
rect 2114 3822 2119 3850
rect 7233 3710 7238 3738
rect 7266 3710 7798 3738
rect 7826 3710 7831 3738
rect 1679 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1821 3542
rect 3835 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3977 3542
rect 5991 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6133 3542
rect 8147 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8289 3542
rect 1073 3318 1078 3346
rect 1106 3318 1414 3346
rect 1442 3318 1638 3346
rect 1666 3318 1918 3346
rect 1946 3318 2198 3346
rect 2226 3318 2231 3346
rect 7177 3318 7182 3346
rect 7210 3318 7350 3346
rect 7378 3318 7383 3346
rect 7849 3318 7854 3346
rect 7882 3318 8414 3346
rect 8442 3318 8974 3346
rect 9002 3318 9007 3346
rect 1745 3262 1750 3290
rect 1778 3262 1974 3290
rect 2002 3262 2007 3290
rect 8353 3262 8358 3290
rect 8386 3262 8694 3290
rect 8722 3262 8862 3290
rect 8890 3262 8895 3290
rect 4489 3206 4494 3234
rect 4522 3206 4830 3234
rect 4858 3206 4863 3234
rect 2757 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2899 3150
rect 4913 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5055 3150
rect 7069 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7211 3150
rect 9225 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9367 3150
rect 7569 3038 7574 3066
rect 7602 3038 7686 3066
rect 7714 3038 7854 3066
rect 7882 3038 8134 3066
rect 8162 3038 8167 3066
rect 1409 2982 1414 3010
rect 1442 2982 1974 3010
rect 2002 2982 2534 3010
rect 2562 2982 2567 3010
rect 3257 2926 3262 2954
rect 3290 2926 3374 2954
rect 3402 2926 3542 2954
rect 3570 2926 3575 2954
rect 1577 2814 1582 2842
rect 1610 2814 1750 2842
rect 1778 2814 2086 2842
rect 2114 2814 2119 2842
rect 4489 2814 4494 2842
rect 4522 2814 4830 2842
rect 4858 2814 4863 2842
rect 7345 2814 7350 2842
rect 7378 2814 7798 2842
rect 7826 2814 7831 2842
rect 7905 2814 7910 2842
rect 7938 2814 8190 2842
rect 8218 2814 8223 2842
rect 1679 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1821 2758
rect 3835 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3977 2758
rect 5991 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6133 2758
rect 8147 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8289 2758
rect 1073 2534 1078 2562
rect 1106 2534 1414 2562
rect 1442 2534 1638 2562
rect 1666 2534 1974 2562
rect 2002 2534 2198 2562
rect 2226 2534 2231 2562
rect 2529 2534 2534 2562
rect 2562 2534 3038 2562
rect 3066 2534 3598 2562
rect 3626 2534 4214 2562
rect 4242 2534 4247 2562
rect 1745 2478 1750 2506
rect 1778 2478 1918 2506
rect 1946 2478 1951 2506
rect 2305 2478 2310 2506
rect 2338 2478 2478 2506
rect 2506 2478 2926 2506
rect 2954 2478 2959 2506
rect 4265 2478 4270 2506
rect 4298 2478 4438 2506
rect 4466 2478 4774 2506
rect 4802 2478 4807 2506
rect 6505 2478 6510 2506
rect 6538 2478 6846 2506
rect 6874 2478 7014 2506
rect 7042 2478 7047 2506
rect 7518 2478 7966 2506
rect 7994 2478 8134 2506
rect 8162 2478 8167 2506
rect 1918 2450 1946 2478
rect 1918 2422 2646 2450
rect 2674 2422 2679 2450
rect 7518 2394 7546 2478
rect 7681 2422 7686 2450
rect 7714 2422 8302 2450
rect 8330 2422 8750 2450
rect 8778 2422 8783 2450
rect 8134 2394 8162 2422
rect 2249 2366 2254 2394
rect 2282 2366 2478 2394
rect 2506 2366 2511 2394
rect 3313 2366 3318 2394
rect 3346 2366 3710 2394
rect 3738 2366 3743 2394
rect 7513 2366 7518 2394
rect 7546 2366 7551 2394
rect 8129 2366 8134 2394
rect 8162 2366 8167 2394
rect 2757 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2899 2366
rect 4913 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5055 2366
rect 7069 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7211 2366
rect 9225 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9367 2366
rect 1353 2254 1358 2282
rect 1386 2254 2254 2282
rect 2282 2254 2287 2282
rect 4209 2198 4214 2226
rect 4242 2198 4718 2226
rect 4746 2198 5054 2226
rect 5082 2198 5166 2226
rect 5194 2198 5558 2226
rect 5586 2198 5894 2226
rect 5922 2198 6174 2226
rect 6202 2198 6454 2226
rect 6482 2198 6958 2226
rect 6986 2198 6991 2226
rect 7569 2198 7574 2226
rect 7602 2198 7686 2226
rect 7714 2198 7719 2226
rect 1577 2142 1582 2170
rect 1610 2142 1750 2170
rect 1778 2142 1783 2170
rect 2081 2142 2086 2170
rect 2114 2142 2310 2170
rect 2338 2142 3150 2170
rect 3178 2142 3183 2170
rect 3257 2142 3262 2170
rect 3290 2142 3374 2170
rect 3402 2142 4102 2170
rect 4130 2142 4135 2170
rect 4321 2142 4326 2170
rect 4354 2142 4550 2170
rect 4578 2142 4583 2170
rect 5217 2142 5222 2170
rect 5250 2142 5390 2170
rect 5418 2142 5423 2170
rect 6113 2142 6118 2170
rect 6146 2142 6286 2170
rect 6314 2142 6319 2170
rect 6561 2142 6566 2170
rect 6594 2142 7294 2170
rect 7322 2142 7462 2170
rect 7490 2142 7495 2170
rect 7793 2142 7798 2170
rect 7826 2142 7966 2170
rect 7994 2142 7999 2170
rect 3817 2086 3822 2114
rect 3850 2086 3990 2114
rect 4018 2086 4662 2114
rect 4690 2086 4695 2114
rect 1745 2030 1750 2058
rect 1778 2030 2702 2058
rect 2730 2030 2735 2058
rect 2865 2030 2870 2058
rect 2898 2030 3654 2058
rect 3682 2030 3687 2058
rect 3873 2030 3878 2058
rect 3906 2030 4214 2058
rect 4242 2030 4247 2058
rect 6281 2030 6286 2058
rect 6314 2030 6734 2058
rect 6762 2030 6902 2058
rect 6930 2030 6935 2058
rect 7009 2030 7014 2058
rect 7042 2030 7406 2058
rect 7434 2030 7439 2058
rect 7569 2030 7574 2058
rect 7602 2030 8526 2058
rect 8554 2030 8559 2058
rect 1679 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1821 1974
rect 3835 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3977 1974
rect 5991 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6133 1974
rect 8147 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8289 1974
rect 6897 1918 6902 1946
rect 6930 1918 7798 1946
rect 7826 1918 7831 1946
rect 1577 1862 1582 1890
rect 1610 1862 2142 1890
rect 2170 1862 2175 1890
rect 2305 1862 2310 1890
rect 2338 1862 2478 1890
rect 2506 1862 3878 1890
rect 3906 1862 3911 1890
rect 7625 1862 7630 1890
rect 7658 1862 8302 1890
rect 8330 1862 8335 1890
rect 1129 1806 1134 1834
rect 1162 1806 1694 1834
rect 1722 1806 1727 1834
rect 2067 1806 2086 1834
rect 2114 1806 2119 1834
rect 2921 1806 2926 1834
rect 2954 1806 3094 1834
rect 3122 1806 3127 1834
rect 3313 1806 3318 1834
rect 3346 1806 4550 1834
rect 4578 1806 4583 1834
rect 6673 1806 6678 1834
rect 6706 1806 7854 1834
rect 7882 1806 8022 1834
rect 8050 1806 8055 1834
rect 1409 1750 1414 1778
rect 1442 1750 1638 1778
rect 1666 1750 1671 1778
rect 1801 1750 1806 1778
rect 1834 1750 1918 1778
rect 1946 1750 3122 1778
rect 3761 1750 3766 1778
rect 3794 1750 3934 1778
rect 3962 1750 4830 1778
rect 4858 1750 4863 1778
rect 5329 1750 5334 1778
rect 5362 1750 5502 1778
rect 5530 1750 5535 1778
rect 6337 1750 6342 1778
rect 6370 1750 7294 1778
rect 7322 1750 7462 1778
rect 7490 1750 7495 1778
rect 7681 1750 7686 1778
rect 7714 1750 8134 1778
rect 8162 1750 8974 1778
rect 9002 1750 9007 1778
rect 1185 1694 1190 1722
rect 1218 1694 1358 1722
rect 1386 1694 2926 1722
rect 2954 1694 2959 1722
rect 3094 1666 3122 1750
rect 4265 1694 4270 1722
rect 4298 1694 4438 1722
rect 4466 1694 5222 1722
rect 5250 1694 5255 1722
rect 6057 1694 6062 1722
rect 6090 1694 6790 1722
rect 6818 1694 6958 1722
rect 6986 1694 6991 1722
rect 7345 1694 7350 1722
rect 7378 1694 8750 1722
rect 8778 1694 8918 1722
rect 8946 1694 8951 1722
rect 3094 1638 3206 1666
rect 3234 1638 3239 1666
rect 8017 1638 8022 1666
rect 8050 1638 8358 1666
rect 8386 1638 8391 1666
rect 7345 1582 7350 1610
rect 7378 1582 8246 1610
rect 8274 1582 8279 1610
rect 2757 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2899 1582
rect 4913 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5055 1582
rect 7069 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7211 1582
rect 9225 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9367 1582
rect 4601 1414 4606 1442
rect 4634 1414 4998 1442
rect 5026 1414 5031 1442
rect 7457 1302 7462 1330
rect 7490 1302 7495 1330
rect 7462 1050 7490 1302
rect 7457 1022 7462 1050
rect 7490 1022 7495 1050
<< via3 >>
rect 1684 4298 1712 4326
rect 1736 4298 1764 4326
rect 1788 4298 1816 4326
rect 3840 4298 3868 4326
rect 3892 4298 3920 4326
rect 3944 4298 3972 4326
rect 5996 4298 6024 4326
rect 6048 4298 6076 4326
rect 6100 4298 6128 4326
rect 8152 4298 8180 4326
rect 8204 4298 8232 4326
rect 8256 4298 8284 4326
rect 2762 3906 2790 3934
rect 2814 3906 2842 3934
rect 2866 3906 2894 3934
rect 4918 3906 4946 3934
rect 4970 3906 4998 3934
rect 5022 3906 5050 3934
rect 7074 3906 7102 3934
rect 7126 3906 7154 3934
rect 7178 3906 7206 3934
rect 9230 3906 9258 3934
rect 9282 3906 9310 3934
rect 9334 3906 9362 3934
rect 1684 3514 1712 3542
rect 1736 3514 1764 3542
rect 1788 3514 1816 3542
rect 3840 3514 3868 3542
rect 3892 3514 3920 3542
rect 3944 3514 3972 3542
rect 5996 3514 6024 3542
rect 6048 3514 6076 3542
rect 6100 3514 6128 3542
rect 8152 3514 8180 3542
rect 8204 3514 8232 3542
rect 8256 3514 8284 3542
rect 7350 3318 7378 3346
rect 2762 3122 2790 3150
rect 2814 3122 2842 3150
rect 2866 3122 2894 3150
rect 4918 3122 4946 3150
rect 4970 3122 4998 3150
rect 5022 3122 5050 3150
rect 7074 3122 7102 3150
rect 7126 3122 7154 3150
rect 7178 3122 7206 3150
rect 9230 3122 9258 3150
rect 9282 3122 9310 3150
rect 9334 3122 9362 3150
rect 2086 2814 2114 2842
rect 1684 2730 1712 2758
rect 1736 2730 1764 2758
rect 1788 2730 1816 2758
rect 3840 2730 3868 2758
rect 3892 2730 3920 2758
rect 3944 2730 3972 2758
rect 5996 2730 6024 2758
rect 6048 2730 6076 2758
rect 6100 2730 6128 2758
rect 8152 2730 8180 2758
rect 8204 2730 8232 2758
rect 8256 2730 8284 2758
rect 2762 2338 2790 2366
rect 2814 2338 2842 2366
rect 2866 2338 2894 2366
rect 4918 2338 4946 2366
rect 4970 2338 4998 2366
rect 5022 2338 5050 2366
rect 7074 2338 7102 2366
rect 7126 2338 7154 2366
rect 7178 2338 7206 2366
rect 9230 2338 9258 2366
rect 9282 2338 9310 2366
rect 9334 2338 9362 2366
rect 1684 1946 1712 1974
rect 1736 1946 1764 1974
rect 1788 1946 1816 1974
rect 3840 1946 3868 1974
rect 3892 1946 3920 1974
rect 3944 1946 3972 1974
rect 5996 1946 6024 1974
rect 6048 1946 6076 1974
rect 6100 1946 6128 1974
rect 8152 1946 8180 1974
rect 8204 1946 8232 1974
rect 8256 1946 8284 1974
rect 2086 1806 2114 1834
rect 7350 1582 7378 1610
rect 2762 1554 2790 1582
rect 2814 1554 2842 1582
rect 2866 1554 2894 1582
rect 4918 1554 4946 1582
rect 4970 1554 4998 1582
rect 5022 1554 5050 1582
rect 7074 1554 7102 1582
rect 7126 1554 7154 1582
rect 7178 1554 7206 1582
rect 9230 1554 9258 1582
rect 9282 1554 9310 1582
rect 9334 1554 9362 1582
<< metal4 >>
rect 1670 4326 1830 4342
rect 1670 4298 1684 4326
rect 1712 4298 1736 4326
rect 1764 4298 1788 4326
rect 1816 4298 1830 4326
rect 1670 3542 1830 4298
rect 1670 3514 1684 3542
rect 1712 3514 1736 3542
rect 1764 3514 1788 3542
rect 1816 3514 1830 3542
rect 1670 2758 1830 3514
rect 2748 3934 2908 4342
rect 2748 3906 2762 3934
rect 2790 3906 2814 3934
rect 2842 3906 2866 3934
rect 2894 3906 2908 3934
rect 2748 3150 2908 3906
rect 2748 3122 2762 3150
rect 2790 3122 2814 3150
rect 2842 3122 2866 3150
rect 2894 3122 2908 3150
rect 1670 2730 1684 2758
rect 1712 2730 1736 2758
rect 1764 2730 1788 2758
rect 1816 2730 1830 2758
rect 1670 1974 1830 2730
rect 1670 1946 1684 1974
rect 1712 1946 1736 1974
rect 1764 1946 1788 1974
rect 1816 1946 1830 1974
rect 1670 1538 1830 1946
rect 2086 2842 2114 2847
rect 2086 1834 2114 2814
rect 2086 1801 2114 1806
rect 2748 2366 2908 3122
rect 2748 2338 2762 2366
rect 2790 2338 2814 2366
rect 2842 2338 2866 2366
rect 2894 2338 2908 2366
rect 2748 1582 2908 2338
rect 2748 1554 2762 1582
rect 2790 1554 2814 1582
rect 2842 1554 2866 1582
rect 2894 1554 2908 1582
rect 2748 1538 2908 1554
rect 3826 4326 3986 4342
rect 3826 4298 3840 4326
rect 3868 4298 3892 4326
rect 3920 4298 3944 4326
rect 3972 4298 3986 4326
rect 3826 3542 3986 4298
rect 3826 3514 3840 3542
rect 3868 3514 3892 3542
rect 3920 3514 3944 3542
rect 3972 3514 3986 3542
rect 3826 2758 3986 3514
rect 3826 2730 3840 2758
rect 3868 2730 3892 2758
rect 3920 2730 3944 2758
rect 3972 2730 3986 2758
rect 3826 1974 3986 2730
rect 3826 1946 3840 1974
rect 3868 1946 3892 1974
rect 3920 1946 3944 1974
rect 3972 1946 3986 1974
rect 3826 1538 3986 1946
rect 4904 3934 5064 4342
rect 4904 3906 4918 3934
rect 4946 3906 4970 3934
rect 4998 3906 5022 3934
rect 5050 3906 5064 3934
rect 4904 3150 5064 3906
rect 4904 3122 4918 3150
rect 4946 3122 4970 3150
rect 4998 3122 5022 3150
rect 5050 3122 5064 3150
rect 4904 2366 5064 3122
rect 4904 2338 4918 2366
rect 4946 2338 4970 2366
rect 4998 2338 5022 2366
rect 5050 2338 5064 2366
rect 4904 1582 5064 2338
rect 4904 1554 4918 1582
rect 4946 1554 4970 1582
rect 4998 1554 5022 1582
rect 5050 1554 5064 1582
rect 4904 1538 5064 1554
rect 5982 4326 6142 4342
rect 5982 4298 5996 4326
rect 6024 4298 6048 4326
rect 6076 4298 6100 4326
rect 6128 4298 6142 4326
rect 5982 3542 6142 4298
rect 5982 3514 5996 3542
rect 6024 3514 6048 3542
rect 6076 3514 6100 3542
rect 6128 3514 6142 3542
rect 5982 2758 6142 3514
rect 5982 2730 5996 2758
rect 6024 2730 6048 2758
rect 6076 2730 6100 2758
rect 6128 2730 6142 2758
rect 5982 1974 6142 2730
rect 5982 1946 5996 1974
rect 6024 1946 6048 1974
rect 6076 1946 6100 1974
rect 6128 1946 6142 1974
rect 5982 1538 6142 1946
rect 7060 3934 7220 4342
rect 7060 3906 7074 3934
rect 7102 3906 7126 3934
rect 7154 3906 7178 3934
rect 7206 3906 7220 3934
rect 7060 3150 7220 3906
rect 8138 4326 8298 4342
rect 8138 4298 8152 4326
rect 8180 4298 8204 4326
rect 8232 4298 8256 4326
rect 8284 4298 8298 4326
rect 8138 3542 8298 4298
rect 8138 3514 8152 3542
rect 8180 3514 8204 3542
rect 8232 3514 8256 3542
rect 8284 3514 8298 3542
rect 7060 3122 7074 3150
rect 7102 3122 7126 3150
rect 7154 3122 7178 3150
rect 7206 3122 7220 3150
rect 7060 2366 7220 3122
rect 7060 2338 7074 2366
rect 7102 2338 7126 2366
rect 7154 2338 7178 2366
rect 7206 2338 7220 2366
rect 7060 1582 7220 2338
rect 7060 1554 7074 1582
rect 7102 1554 7126 1582
rect 7154 1554 7178 1582
rect 7206 1554 7220 1582
rect 7350 3346 7378 3351
rect 7350 1610 7378 3318
rect 7350 1577 7378 1582
rect 8138 2758 8298 3514
rect 8138 2730 8152 2758
rect 8180 2730 8204 2758
rect 8232 2730 8256 2758
rect 8284 2730 8298 2758
rect 8138 1974 8298 2730
rect 8138 1946 8152 1974
rect 8180 1946 8204 1974
rect 8232 1946 8256 1974
rect 8284 1946 8298 1974
rect 7060 1538 7220 1554
rect 8138 1538 8298 1946
rect 9216 3934 9376 4342
rect 9216 3906 9230 3934
rect 9258 3906 9282 3934
rect 9310 3906 9334 3934
rect 9362 3906 9376 3934
rect 9216 3150 9376 3906
rect 9216 3122 9230 3150
rect 9258 3122 9282 3150
rect 9310 3122 9334 3150
rect 9362 3122 9376 3150
rect 9216 2366 9376 3122
rect 9216 2338 9230 2366
rect 9258 2338 9282 2366
rect 9310 2338 9334 2366
rect 9362 2338 9376 2366
rect 9216 1582 9376 2338
rect 9216 1554 9230 1582
rect 9258 1554 9282 1582
rect 9310 1554 9334 1582
rect 9362 1554 9376 1582
rect 9216 1538 9376 1554
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 1456 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24
timestamp 1667941163
transform 1 0 2016 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49
timestamp 1667941163
transform 1 0 3416 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59
timestamp 1667941163
transform 1 0 3976 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 4536 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76
timestamp 1667941163
transform 1 0 4928 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78
timestamp 1667941163
transform 1 0 5040 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87
timestamp 1667941163
transform 1 0 5544 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 6104 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1667941163
transform 1 0 6664 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116
timestamp 1667941163
transform 1 0 7168 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_126
timestamp 1667941163
transform 1 0 7728 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_136
timestamp 1667941163
transform 1 0 8288 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1667941163
transform 1 0 8624 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_151
timestamp 1667941163
transform 1 0 9128 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2
timestamp 1667941163
transform 1 0 784 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_10
timestamp 1667941163
transform 1 0 1232 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_20
timestamp 1667941163
transform 1 0 1792 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_30
timestamp 1667941163
transform 1 0 2352 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_40
timestamp 1667941163
transform 1 0 2912 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_50
timestamp 1667941163
transform 1 0 3472 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_60
timestamp 1667941163
transform 1 0 4032 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_85
timestamp 1667941163
transform 1 0 5432 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_95
timestamp 1667941163
transform 1 0 5992 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_105
timestamp 1667941163
transform 1 0 6552 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_115
timestamp 1667941163
transform 1 0 7112 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_125
timestamp 1667941163
transform 1 0 7672 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_135
timestamp 1667941163
transform 1 0 8232 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_139
timestamp 1667941163
transform 1 0 8456 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 8568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_144
timestamp 1667941163
transform 1 0 8736 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_14
timestamp 1667941163
transform 1 0 1456 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_24
timestamp 1667941163
transform 1 0 2016 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_49
timestamp 1667941163
transform 1 0 3416 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_59
timestamp 1667941163
transform 1 0 3976 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_69
timestamp 1667941163
transform 1 0 4536 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_79
timestamp 1667941163
transform 1 0 5096 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_89
timestamp 1667941163
transform 1 0 5656 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_93
timestamp 1667941163
transform 1 0 5880 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_103
timestamp 1667941163
transform 1 0 6440 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1667941163
transform 1 0 6720 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_117
timestamp 1667941163
transform 1 0 7224 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_127
timestamp 1667941163
transform 1 0 7784 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_137
timestamp 1667941163
transform 1 0 8344 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_147
timestamp 1667941163
transform 1 0 8904 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_151
timestamp 1667941163
transform 1 0 9128 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_10
timestamp 1667941163
transform 1 0 1232 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_20
timestamp 1667941163
transform 1 0 1792 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_30
timestamp 1667941163
transform 1 0 2352 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_40
timestamp 1667941163
transform 1 0 2912 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_50
timestamp 1667941163
transform 1 0 3472 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_60
timestamp 1667941163
transform 1 0 4032 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_82 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5264 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_98
timestamp 1667941163
transform 1 0 6160 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_106
timestamp 1667941163
transform 1 0 6608 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_115
timestamp 1667941163
transform 1 0 7112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_125
timestamp 1667941163
transform 1 0 7672 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_135
timestamp 1667941163
transform 1 0 8232 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_139
timestamp 1667941163
transform 1 0 8456 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 8568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_144
timestamp 1667941163
transform 1 0 8736 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1667941163
transform 1 0 1456 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_24
timestamp 1667941163
transform 1 0 2016 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_45
timestamp 1667941163
transform 1 0 3192 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_55 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 3752 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_87
timestamp 1667941163
transform 1 0 5544 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_103
timestamp 1667941163
transform 1 0 6440 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_108
timestamp 1667941163
transform 1 0 6720 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_120
timestamp 1667941163
transform 1 0 7392 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_130
timestamp 1667941163
transform 1 0 7952 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_140
timestamp 1667941163
transform 1 0 8512 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_150
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_6
timestamp 1667941163
transform 1 0 1008 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_16
timestamp 1667941163
transform 1 0 1568 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_26
timestamp 1667941163
transform 1 0 2128 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_36
timestamp 1667941163
transform 1 0 2688 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_68
timestamp 1667941163
transform 1 0 4480 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_105
timestamp 1667941163
transform 1 0 6552 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 7000 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_123
timestamp 1667941163
transform 1 0 7560 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_133
timestamp 1667941163
transform 1 0 8120 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 8568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_144
timestamp 1667941163
transform 1 0 8736 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_6
timestamp 1667941163
transform 1 0 1008 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_16
timestamp 1667941163
transform 1 0 1568 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_26
timestamp 1667941163
transform 1 0 2128 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_69
timestamp 1667941163
transform 1 0 4536 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_72
timestamp 1667941163
transform 1 0 4704 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1667941163
transform 1 0 6496 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_107
timestamp 1667941163
transform 1 0 6664 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_123
timestamp 1667941163
transform 1 0 7560 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_127
timestamp 1667941163
transform 1 0 7784 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_136
timestamp 1667941163
transform 1 0 8288 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_142
timestamp 1667941163
transform 1 0 8624 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_151
timestamp 1667941163
transform 1 0 9128 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 9296 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 9296 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 9296 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 9296 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 9296 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 9296 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 9296 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_14 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_15
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_16
timestamp 1667941163
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_17
timestamp 1667941163
transform 1 0 8512 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_18
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_19
timestamp 1667941163
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_20
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_21
timestamp 1667941163
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_22
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_23
timestamp 1667941163
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1667941163
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1667941163
transform 1 0 8624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1667941163
transform 1 0 4592 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1667941163
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1667941163
transform 1 0 8512 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[0\].u_cap pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 1568 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[1\].u_cap
timestamp 1667941163
transform -1 0 1568 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[2\].u_cap
timestamp 1667941163
transform 1 0 1680 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[3\].u_cap
timestamp 1667941163
transform -1 0 1456 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[4\].u_cap
timestamp 1667941163
transform 1 0 1680 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[5\].u_cap
timestamp 1667941163
transform -1 0 2016 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[6\].u_cap
timestamp 1667941163
transform -1 0 1792 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[7\].u_cap
timestamp 1667941163
transform -1 0 1456 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[8\].u_cap
timestamp 1667941163
transform 1 0 2240 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[9\].u_cap
timestamp 1667941163
transform -1 0 2576 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[10\].u_cap
timestamp 1667941163
transform -1 0 2352 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[11\].u_cap
timestamp 1667941163
transform -1 0 2016 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[12\].u_cap
timestamp 1667941163
transform -1 0 1792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[13\].u_cap
timestamp 1667941163
transform -1 0 1456 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[14\].u_cap
timestamp 1667941163
transform -1 0 2912 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[15\].u_cap
timestamp 1667941163
transform -1 0 2576 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[16\].u_cap
timestamp 1667941163
transform -1 0 2352 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[17\].u_cap
timestamp 1667941163
transform -1 0 2016 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[18\].u_cap
timestamp 1667941163
transform 1 0 3304 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[19\].u_cap
timestamp 1667941163
transform -1 0 3472 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[20\].u_cap
timestamp 1667941163
transform -1 0 2912 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[21\].u_cap
timestamp 1667941163
transform -1 0 3416 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[22\].u_cap
timestamp 1667941163
transform -1 0 2576 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[23\].u_cap
timestamp 1667941163
transform -1 0 4032 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[24\].u_cap
timestamp 1667941163
transform -1 0 3472 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[25\].u_cap
timestamp 1667941163
transform -1 0 3976 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[26\].u_cap
timestamp 1667941163
transform 1 0 4144 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[27\].u_cap
timestamp 1667941163
transform 1 0 4816 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[28\].u_cap
timestamp 1667941163
transform -1 0 3416 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[29\].u_cap
timestamp 1667941163
transform -1 0 4032 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[30\].u_cap
timestamp 1667941163
transform -1 0 4536 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[31\].u_cap
timestamp 1667941163
transform -1 0 3976 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[32\].u_cap
timestamp 1667941163
transform -1 0 4592 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[33\].u_cap
timestamp 1667941163
transform -1 0 5096 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[34\].u_cap
timestamp 1667941163
transform -1 0 4536 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[35\].u_cap
timestamp 1667941163
transform 1 0 5208 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[36\].u_cap
timestamp 1667941163
transform -1 0 5432 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[37\].u_cap
timestamp 1667941163
transform -1 0 5544 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[38\].u_cap
timestamp 1667941163
transform 1 0 5544 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[39\].u_cap
timestamp 1667941163
transform 1 0 5656 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[40\].u_cap
timestamp 1667941163
transform 1 0 6104 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[41\].u_cap
timestamp 1667941163
transform 1 0 6720 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[42\].u_cap
timestamp 1667941163
transform 1 0 5992 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[43\].u_cap
timestamp 1667941163
transform 1 0 6664 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[44\].u_cap
timestamp 1667941163
transform 1 0 7280 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[45\].u_cap
timestamp 1667941163
transform 1 0 6776 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[46\].u_cap
timestamp 1667941163
transform 1 0 7224 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[47\].u_cap
timestamp 1667941163
transform 1 0 7840 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[48\].u_cap
timestamp 1667941163
transform 1 0 6664 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[49\].u_cap
timestamp 1667941163
transform 1 0 7784 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[50\].u_cap
timestamp 1667941163
transform 1 0 7336 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[51\].u_cap
timestamp 1667941163
transform 1 0 7224 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[52\].u_cap
timestamp 1667941163
transform 1 0 8680 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[53\].u_cap
timestamp 1667941163
transform 1 0 7896 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[54\].u_cap
timestamp 1667941163
transform 1 0 7784 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[55\].u_cap
timestamp 1667941163
transform 1 0 8456 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[56\].u_cap
timestamp 1667941163
transform 1 0 7504 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[57\].u_cap
timestamp 1667941163
transform 1 0 8064 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[58\].u_cap
timestamp 1667941163
transform -1 0 8120 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[59\].u_cap
timestamp 1667941163
transform 1 0 8624 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[60\].u_cap
timestamp 1667941163
transform -1 0 8288 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[61\].u_cap
timestamp 1667941163
transform -1 0 7392 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[62\].u_cap
timestamp 1667941163
transform -1 0 7560 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_cap\[63\].u_cap
timestamp 1667941163
transform 1 0 8680 0 1 3920
box -43 -43 491 435
<< labels >>
flabel metal2 s 4928 5600 4984 6000 0 FreeSans 224 90 0 0 cap
port 0 nsew signal bidirectional
flabel metal2 s 1400 0 1456 400 0 FreeSans 224 90 0 0 tune[0]
port 1 nsew signal input
flabel metal2 s 2520 0 2576 400 0 FreeSans 224 90 0 0 tune[10]
port 2 nsew signal input
flabel metal2 s 2632 0 2688 400 0 FreeSans 224 90 0 0 tune[11]
port 3 nsew signal input
flabel metal2 s 2744 0 2800 400 0 FreeSans 224 90 0 0 tune[12]
port 4 nsew signal input
flabel metal2 s 2856 0 2912 400 0 FreeSans 224 90 0 0 tune[13]
port 5 nsew signal input
flabel metal2 s 2968 0 3024 400 0 FreeSans 224 90 0 0 tune[14]
port 6 nsew signal input
flabel metal2 s 3080 0 3136 400 0 FreeSans 224 90 0 0 tune[15]
port 7 nsew signal input
flabel metal2 s 3192 0 3248 400 0 FreeSans 224 90 0 0 tune[16]
port 8 nsew signal input
flabel metal2 s 3304 0 3360 400 0 FreeSans 224 90 0 0 tune[17]
port 9 nsew signal input
flabel metal2 s 3416 0 3472 400 0 FreeSans 224 90 0 0 tune[18]
port 10 nsew signal input
flabel metal2 s 3528 0 3584 400 0 FreeSans 224 90 0 0 tune[19]
port 11 nsew signal input
flabel metal2 s 1512 0 1568 400 0 FreeSans 224 90 0 0 tune[1]
port 12 nsew signal input
flabel metal2 s 3640 0 3696 400 0 FreeSans 224 90 0 0 tune[20]
port 13 nsew signal input
flabel metal2 s 3752 0 3808 400 0 FreeSans 224 90 0 0 tune[21]
port 14 nsew signal input
flabel metal2 s 3864 0 3920 400 0 FreeSans 224 90 0 0 tune[22]
port 15 nsew signal input
flabel metal2 s 3976 0 4032 400 0 FreeSans 224 90 0 0 tune[23]
port 16 nsew signal input
flabel metal2 s 4088 0 4144 400 0 FreeSans 224 90 0 0 tune[24]
port 17 nsew signal input
flabel metal2 s 4200 0 4256 400 0 FreeSans 224 90 0 0 tune[25]
port 18 nsew signal input
flabel metal2 s 4312 0 4368 400 0 FreeSans 224 90 0 0 tune[26]
port 19 nsew signal input
flabel metal2 s 4424 0 4480 400 0 FreeSans 224 90 0 0 tune[27]
port 20 nsew signal input
flabel metal2 s 4536 0 4592 400 0 FreeSans 224 90 0 0 tune[28]
port 21 nsew signal input
flabel metal2 s 4648 0 4704 400 0 FreeSans 224 90 0 0 tune[29]
port 22 nsew signal input
flabel metal2 s 1624 0 1680 400 0 FreeSans 224 90 0 0 tune[2]
port 23 nsew signal input
flabel metal2 s 4760 0 4816 400 0 FreeSans 224 90 0 0 tune[30]
port 24 nsew signal input
flabel metal2 s 4872 0 4928 400 0 FreeSans 224 90 0 0 tune[31]
port 25 nsew signal input
flabel metal2 s 4984 0 5040 400 0 FreeSans 224 90 0 0 tune[32]
port 26 nsew signal input
flabel metal2 s 5096 0 5152 400 0 FreeSans 224 90 0 0 tune[33]
port 27 nsew signal input
flabel metal2 s 5208 0 5264 400 0 FreeSans 224 90 0 0 tune[34]
port 28 nsew signal input
flabel metal2 s 5320 0 5376 400 0 FreeSans 224 90 0 0 tune[35]
port 29 nsew signal input
flabel metal2 s 5432 0 5488 400 0 FreeSans 224 90 0 0 tune[36]
port 30 nsew signal input
flabel metal2 s 5544 0 5600 400 0 FreeSans 224 90 0 0 tune[37]
port 31 nsew signal input
flabel metal2 s 5656 0 5712 400 0 FreeSans 224 90 0 0 tune[38]
port 32 nsew signal input
flabel metal2 s 5768 0 5824 400 0 FreeSans 224 90 0 0 tune[39]
port 33 nsew signal input
flabel metal2 s 1736 0 1792 400 0 FreeSans 224 90 0 0 tune[3]
port 34 nsew signal input
flabel metal2 s 5880 0 5936 400 0 FreeSans 224 90 0 0 tune[40]
port 35 nsew signal input
flabel metal2 s 5992 0 6048 400 0 FreeSans 224 90 0 0 tune[41]
port 36 nsew signal input
flabel metal2 s 6104 0 6160 400 0 FreeSans 224 90 0 0 tune[42]
port 37 nsew signal input
flabel metal2 s 6216 0 6272 400 0 FreeSans 224 90 0 0 tune[43]
port 38 nsew signal input
flabel metal2 s 6328 0 6384 400 0 FreeSans 224 90 0 0 tune[44]
port 39 nsew signal input
flabel metal2 s 6440 0 6496 400 0 FreeSans 224 90 0 0 tune[45]
port 40 nsew signal input
flabel metal2 s 6552 0 6608 400 0 FreeSans 224 90 0 0 tune[46]
port 41 nsew signal input
flabel metal2 s 6664 0 6720 400 0 FreeSans 224 90 0 0 tune[47]
port 42 nsew signal input
flabel metal2 s 6776 0 6832 400 0 FreeSans 224 90 0 0 tune[48]
port 43 nsew signal input
flabel metal2 s 6888 0 6944 400 0 FreeSans 224 90 0 0 tune[49]
port 44 nsew signal input
flabel metal2 s 1848 0 1904 400 0 FreeSans 224 90 0 0 tune[4]
port 45 nsew signal input
flabel metal2 s 7000 0 7056 400 0 FreeSans 224 90 0 0 tune[50]
port 46 nsew signal input
flabel metal2 s 7112 0 7168 400 0 FreeSans 224 90 0 0 tune[51]
port 47 nsew signal input
flabel metal2 s 7224 0 7280 400 0 FreeSans 224 90 0 0 tune[52]
port 48 nsew signal input
flabel metal2 s 7336 0 7392 400 0 FreeSans 224 90 0 0 tune[53]
port 49 nsew signal input
flabel metal2 s 7448 0 7504 400 0 FreeSans 224 90 0 0 tune[54]
port 50 nsew signal input
flabel metal2 s 7560 0 7616 400 0 FreeSans 224 90 0 0 tune[55]
port 51 nsew signal input
flabel metal2 s 7672 0 7728 400 0 FreeSans 224 90 0 0 tune[56]
port 52 nsew signal input
flabel metal2 s 7784 0 7840 400 0 FreeSans 224 90 0 0 tune[57]
port 53 nsew signal input
flabel metal2 s 7896 0 7952 400 0 FreeSans 224 90 0 0 tune[58]
port 54 nsew signal input
flabel metal2 s 8008 0 8064 400 0 FreeSans 224 90 0 0 tune[59]
port 55 nsew signal input
flabel metal2 s 1960 0 2016 400 0 FreeSans 224 90 0 0 tune[5]
port 56 nsew signal input
flabel metal2 s 8120 0 8176 400 0 FreeSans 224 90 0 0 tune[60]
port 57 nsew signal input
flabel metal2 s 8232 0 8288 400 0 FreeSans 224 90 0 0 tune[61]
port 58 nsew signal input
flabel metal2 s 8344 0 8400 400 0 FreeSans 224 90 0 0 tune[62]
port 59 nsew signal input
flabel metal2 s 8456 0 8512 400 0 FreeSans 224 90 0 0 tune[63]
port 60 nsew signal input
flabel metal2 s 2072 0 2128 400 0 FreeSans 224 90 0 0 tune[6]
port 61 nsew signal input
flabel metal2 s 2184 0 2240 400 0 FreeSans 224 90 0 0 tune[7]
port 62 nsew signal input
flabel metal2 s 2296 0 2352 400 0 FreeSans 224 90 0 0 tune[8]
port 63 nsew signal input
flabel metal2 s 2408 0 2464 400 0 FreeSans 224 90 0 0 tune[9]
port 64 nsew signal input
flabel metal4 s 1670 1538 1830 4342 0 FreeSans 640 90 0 0 vdd
port 65 nsew power bidirectional
flabel metal4 s 3826 1538 3986 4342 0 FreeSans 640 90 0 0 vdd
port 65 nsew power bidirectional
flabel metal4 s 5982 1538 6142 4342 0 FreeSans 640 90 0 0 vdd
port 65 nsew power bidirectional
flabel metal4 s 8138 1538 8298 4342 0 FreeSans 640 90 0 0 vdd
port 65 nsew power bidirectional
flabel metal4 s 2748 1538 2908 4342 0 FreeSans 640 90 0 0 vss
port 66 nsew ground bidirectional
flabel metal4 s 4904 1538 5064 4342 0 FreeSans 640 90 0 0 vss
port 66 nsew ground bidirectional
flabel metal4 s 7060 1538 7220 4342 0 FreeSans 640 90 0 0 vss
port 66 nsew ground bidirectional
flabel metal4 s 9216 1538 9376 4342 0 FreeSans 640 90 0 0 vss
port 66 nsew ground bidirectional
rlabel metal1 4984 4312 4984 4312 0 vdd
rlabel via1 5024 3920 5024 3920 0 vss
rlabel metal2 1960 3724 1960 3724 0 cap
rlabel metal2 1428 1029 1428 1029 0 tune[0]
rlabel metal2 2268 2660 2268 2660 0 tune[10]
rlabel metal3 1932 2464 1932 2464 0 tune[11]
rlabel metal2 1764 2100 1764 2100 0 tune[12]
rlabel metal2 2940 1456 2940 1456 0 tune[13]
rlabel metal2 2884 2884 2884 2884 0 tune[14]
rlabel metal3 2716 2492 2716 2492 0 tune[15]
rlabel metal3 2744 2156 2744 2156 0 tune[16]
rlabel metal3 2520 1764 2520 1764 0 tune[17]
rlabel metal2 3416 3276 3416 3276 0 tune[18]
rlabel metal3 3472 2940 3472 2940 0 tune[19]
rlabel metal2 1540 3724 1540 3724 0 tune[1]
rlabel metal2 2884 2100 2884 2100 0 tune[20]
rlabel metal2 3332 2436 3332 2436 0 tune[21]
rlabel metal2 2492 1820 2492 1820 0 tune[22]
rlabel metal2 4032 2940 4032 2940 0 tune[23]
rlabel metal3 3752 2156 3752 2156 0 tune[24]
rlabel metal2 3892 2268 3892 2268 0 tune[25]
rlabel metal2 4396 2464 4396 2464 0 tune[26]
rlabel metal2 4844 2884 4844 2884 0 tune[27]
rlabel metal2 3332 1792 3332 1792 0 tune[28]
rlabel metal2 4004 2128 4004 2128 0 tune[29]
rlabel metal2 1932 3948 1932 3948 0 tune[2]
rlabel metal3 4620 2492 4620 2492 0 tune[30]
rlabel metal3 3864 1764 3864 1764 0 tune[31]
rlabel metal2 4592 2156 4592 2156 0 tune[32]
rlabel metal2 5068 2492 5068 2492 0 tune[33]
rlabel metal3 4844 1708 4844 1708 0 tune[34]
rlabel metal2 5292 2072 5292 2072 0 tune[35]
rlabel metal2 5432 2156 5432 2156 0 tune[36]
rlabel metal2 5544 1764 5544 1764 0 tune[37]
rlabel metal2 5656 2156 5656 2156 0 tune[38]
rlabel metal2 5768 1708 5768 1708 0 tune[39]
rlabel metal2 1708 1708 1708 1708 0 tune[3]
rlabel metal2 6132 2100 6132 2100 0 tune[40]
rlabel metal3 6440 1708 6440 1708 0 tune[41]
rlabel metal2 6244 2072 6244 2072 0 tune[42]
rlabel metal2 6748 2100 6748 2100 0 tune[43]
rlabel metal3 6832 1764 6832 1764 0 tune[44]
rlabel metal3 6692 2492 6692 2492 0 tune[45]
rlabel metal3 6944 2156 6944 2156 0 tune[46]
rlabel metal2 6692 1099 6692 1099 0 tune[47]
rlabel metal2 6748 2604 6748 2604 0 tune[48]
rlabel metal2 6916 1155 6916 1155 0 tune[49]
rlabel metal2 1876 3584 1876 3584 0 tune[4]
rlabel metal2 7420 2268 7420 2268 0 tune[50]
rlabel metal2 7252 2212 7252 2212 0 tune[51]
rlabel metal2 7364 1540 7364 1540 0 tune[52]
rlabel metal3 7532 2436 7532 2436 0 tune[53]
rlabel metal2 7364 2380 7364 2380 0 tune[54]
rlabel metal2 8540 2268 8540 2268 0 tune[55]
rlabel metal2 7700 1029 7700 1029 0 tune[56]
rlabel metal2 7812 1029 7812 1029 0 tune[57]
rlabel metal2 7952 1596 7952 1596 0 tune[58]
rlabel metal3 8204 1652 8204 1652 0 tune[59]
rlabel metal2 2016 3332 2016 3332 0 tune[5]
rlabel metal2 8148 1029 8148 1029 0 tune[60]
rlabel metal4 7364 2464 7364 2464 0 tune[61]
rlabel metal2 7532 3444 7532 3444 0 tune[62]
rlabel metal2 8596 4116 8596 4116 0 tune[63]
rlabel metal2 1764 2884 1764 2884 0 tune[6]
rlabel metal2 2268 1932 2268 1932 0 tune[7]
rlabel metal2 2324 3164 2324 3164 0 tune[8]
rlabel metal2 2464 3276 2464 3276 0 tune[9]
<< properties >>
string FIXED_BBOX 0 0 10000 6000
<< end >>
