magic
tech gf180mcuC
magscale 1 10
timestamp 1669565339
<< nwell >>
rect 132 1758 668 3714
rect 132 710 668 1268
<< pwell >>
rect 132 3714 668 4260
rect 132 1268 668 1758
rect 132 164 668 710
<< mvnmos >>
rect 270 3922 510 4062
rect 330 1393 470 1633
rect 270 362 510 502
<< mvpmos >>
rect 340 1936 460 3536
rect 340 888 460 1088
<< mvndiff >>
rect 270 4137 510 4150
rect 270 4091 283 4137
rect 497 4091 510 4137
rect 270 4062 510 4091
rect 270 3893 510 3922
rect 270 3847 283 3893
rect 497 3847 510 3893
rect 270 3834 510 3847
rect 242 1620 330 1633
rect 242 1406 255 1620
rect 301 1406 330 1620
rect 242 1393 330 1406
rect 470 1620 558 1633
rect 470 1406 499 1620
rect 545 1406 558 1620
rect 470 1393 558 1406
rect 270 577 510 590
rect 270 531 283 577
rect 497 531 510 577
rect 270 502 510 531
rect 270 333 510 362
rect 270 287 283 333
rect 497 287 510 333
rect 270 274 510 287
<< mvpdiff >>
rect 252 3523 340 3536
rect 252 1949 265 3523
rect 311 1949 340 3523
rect 252 1936 340 1949
rect 460 3523 548 3536
rect 460 1949 489 3523
rect 535 1949 548 3523
rect 460 1936 548 1949
rect 252 1075 340 1088
rect 252 901 265 1075
rect 311 901 340 1075
rect 252 888 340 901
rect 460 1075 548 1088
rect 460 901 489 1075
rect 535 901 548 1075
rect 460 888 548 901
<< mvndiffc >>
rect 283 4091 497 4137
rect 283 3847 497 3893
rect 255 1406 301 1620
rect 499 1406 545 1620
rect 283 531 497 577
rect 283 287 497 333
<< mvpdiffc >>
rect 265 1949 311 3523
rect 489 1949 535 3523
rect 265 901 311 1075
rect 489 901 535 1075
<< polysilicon >>
rect 178 4049 270 4062
rect 178 3935 191 4049
rect 237 3935 270 4049
rect 178 3922 270 3935
rect 510 4049 602 4062
rect 510 3935 543 4049
rect 589 3935 602 4049
rect 510 3922 602 3935
rect 340 3615 460 3628
rect 340 3569 353 3615
rect 447 3569 460 3615
rect 340 3536 460 3569
rect 340 1903 460 1936
rect 340 1857 353 1903
rect 447 1857 460 1903
rect 340 1844 460 1857
rect 330 1712 470 1725
rect 330 1666 343 1712
rect 457 1666 470 1712
rect 330 1633 470 1666
rect 330 1360 470 1393
rect 330 1314 343 1360
rect 457 1314 470 1360
rect 330 1301 470 1314
rect 340 1167 460 1180
rect 340 1121 353 1167
rect 447 1121 460 1167
rect 340 1088 460 1121
rect 340 855 460 888
rect 340 809 353 855
rect 447 809 460 855
rect 340 796 460 809
rect 178 489 270 502
rect 178 375 191 489
rect 237 375 270 489
rect 178 362 270 375
rect 510 489 602 502
rect 510 375 543 489
rect 589 375 602 489
rect 510 362 602 375
<< polycontact >>
rect 191 3935 237 4049
rect 543 3935 589 4049
rect 353 3569 447 3615
rect 353 1857 447 1903
rect 343 1666 457 1712
rect 343 1314 457 1360
rect 353 1121 447 1167
rect 353 809 447 855
rect 191 375 237 489
rect 543 375 589 489
<< metal1 >>
rect 296 4174 484 4176
rect 296 4137 308 4174
rect 364 4137 416 4174
rect 472 4137 484 4174
rect 154 4084 214 4096
rect 272 4091 283 4137
rect 497 4091 508 4137
rect 154 4028 156 4084
rect 212 4060 214 4084
rect 566 4084 626 4096
rect 566 4060 568 4084
rect 212 4049 237 4060
rect 154 3956 191 4028
rect 154 3900 156 3956
rect 212 3924 237 3935
rect 543 4049 568 4060
rect 624 4028 626 4084
rect 589 3956 626 4028
rect 543 3924 568 3935
rect 212 3900 214 3924
rect 154 3888 214 3900
rect 566 3900 568 3924
rect 624 3900 626 3956
rect 272 3847 283 3893
rect 497 3847 508 3893
rect 566 3888 626 3900
rect 296 3808 508 3847
rect 296 3748 682 3808
rect 296 3650 504 3652
rect 296 3594 308 3650
rect 364 3615 436 3650
rect 492 3594 504 3650
rect 296 3592 353 3594
rect 342 3569 353 3592
rect 447 3592 504 3594
rect 447 3569 458 3592
rect 265 3523 311 3534
rect 226 3466 265 3478
rect 226 3410 228 3466
rect 226 3358 265 3410
rect 226 3302 228 3358
rect 226 3250 265 3302
rect 226 3194 228 3250
rect 226 3142 265 3194
rect 226 3086 228 3142
rect 226 3034 265 3086
rect 226 2978 228 3034
rect 226 2926 265 2978
rect 226 2870 228 2926
rect 226 2818 265 2870
rect 226 2762 228 2818
rect 226 2710 265 2762
rect 226 2654 228 2710
rect 226 2602 265 2654
rect 226 2546 228 2602
rect 226 2494 265 2546
rect 226 2438 228 2494
rect 226 2386 265 2438
rect 226 2330 228 2386
rect 226 2278 265 2330
rect 226 2222 228 2278
rect 226 2170 265 2222
rect 226 2114 228 2170
rect 226 2062 265 2114
rect 226 2006 228 2062
rect 226 1994 265 2006
rect 265 1938 311 1949
rect 489 3523 535 3534
rect 535 3466 574 3478
rect 572 3410 574 3466
rect 535 3358 574 3410
rect 572 3302 574 3358
rect 535 3250 574 3302
rect 572 3194 574 3250
rect 535 3142 574 3194
rect 572 3086 574 3142
rect 535 3034 574 3086
rect 572 2978 574 3034
rect 535 2926 574 2978
rect 572 2870 574 2926
rect 535 2818 574 2870
rect 572 2762 574 2818
rect 535 2710 574 2762
rect 572 2654 574 2710
rect 535 2602 574 2654
rect 572 2546 574 2602
rect 535 2494 574 2546
rect 572 2438 574 2494
rect 535 2386 574 2438
rect 572 2330 574 2386
rect 535 2278 574 2330
rect 572 2222 574 2278
rect 535 2170 574 2222
rect 572 2114 574 2170
rect 535 2062 574 2114
rect 572 2006 574 2062
rect 535 1994 574 2006
rect 489 1938 535 1949
rect 342 1880 353 1903
rect 296 1878 353 1880
rect 447 1880 458 1903
rect 447 1878 504 1880
rect 296 1822 308 1878
rect 364 1822 436 1857
rect 492 1822 504 1878
rect 296 1820 504 1822
rect 296 1747 504 1749
rect 296 1691 308 1747
rect 364 1712 436 1747
rect 492 1691 504 1747
rect 296 1689 343 1691
rect 332 1666 343 1689
rect 457 1689 504 1691
rect 457 1666 468 1689
rect 621 1631 682 3748
rect 255 1620 301 1631
rect 107 1406 255 1478
rect 107 1395 301 1406
rect 499 1620 682 1631
rect 545 1548 682 1620
rect 499 1395 545 1406
rect 107 676 167 1395
rect 332 1337 343 1360
rect 296 1335 343 1337
rect 457 1337 468 1360
rect 457 1335 504 1337
rect 296 1279 308 1335
rect 364 1279 436 1314
rect 492 1279 504 1335
rect 296 1277 504 1279
rect 296 1202 504 1204
rect 296 1146 308 1202
rect 364 1167 436 1202
rect 492 1146 504 1202
rect 296 1144 353 1146
rect 342 1121 353 1144
rect 447 1144 504 1146
rect 447 1121 458 1144
rect 265 1082 311 1086
rect 226 1075 311 1082
rect 226 1070 265 1075
rect 226 1014 228 1070
rect 226 962 265 1014
rect 226 906 228 962
rect 226 901 265 906
rect 226 894 311 901
rect 265 890 311 894
rect 489 1082 535 1086
rect 489 1075 574 1082
rect 535 1070 574 1075
rect 572 1014 574 1070
rect 535 962 574 1014
rect 572 906 574 962
rect 535 901 574 906
rect 489 894 574 901
rect 489 890 535 894
rect 342 832 353 855
rect 296 830 353 832
rect 447 832 458 855
rect 447 830 504 832
rect 296 774 308 830
rect 364 774 436 809
rect 492 774 504 830
rect 296 772 504 774
rect 107 616 484 676
rect 272 577 484 616
rect 154 524 214 536
rect 272 531 283 577
rect 497 531 508 577
rect 154 468 156 524
rect 212 500 214 524
rect 566 524 626 536
rect 566 500 568 524
rect 212 489 237 500
rect 154 396 191 468
rect 154 340 156 396
rect 212 364 237 375
rect 543 489 568 500
rect 624 468 626 524
rect 589 396 626 468
rect 543 364 568 375
rect 212 340 214 364
rect 154 328 214 340
rect 566 340 568 364
rect 624 340 626 396
rect 272 287 283 333
rect 497 287 508 333
rect 566 328 626 340
rect 296 250 308 287
rect 364 250 416 287
rect 472 250 484 287
rect 296 248 484 250
<< via1 >>
rect 308 4137 364 4174
rect 416 4137 472 4174
rect 308 4118 364 4137
rect 416 4118 472 4137
rect 156 4049 212 4084
rect 156 4028 191 4049
rect 191 4028 212 4049
rect 156 3935 191 3956
rect 191 3935 212 3956
rect 156 3900 212 3935
rect 568 4049 624 4084
rect 568 4028 589 4049
rect 589 4028 624 4049
rect 568 3935 589 3956
rect 589 3935 624 3956
rect 568 3900 624 3935
rect 308 3615 364 3650
rect 436 3615 492 3650
rect 308 3594 353 3615
rect 353 3594 364 3615
rect 436 3594 447 3615
rect 447 3594 492 3615
rect 228 3410 265 3466
rect 265 3410 284 3466
rect 228 3302 265 3358
rect 265 3302 284 3358
rect 228 3194 265 3250
rect 265 3194 284 3250
rect 228 3086 265 3142
rect 265 3086 284 3142
rect 228 2978 265 3034
rect 265 2978 284 3034
rect 228 2870 265 2926
rect 265 2870 284 2926
rect 228 2762 265 2818
rect 265 2762 284 2818
rect 228 2654 265 2710
rect 265 2654 284 2710
rect 228 2546 265 2602
rect 265 2546 284 2602
rect 228 2438 265 2494
rect 265 2438 284 2494
rect 228 2330 265 2386
rect 265 2330 284 2386
rect 228 2222 265 2278
rect 265 2222 284 2278
rect 228 2114 265 2170
rect 265 2114 284 2170
rect 228 2006 265 2062
rect 265 2006 284 2062
rect 516 3410 535 3466
rect 535 3410 572 3466
rect 516 3302 535 3358
rect 535 3302 572 3358
rect 516 3194 535 3250
rect 535 3194 572 3250
rect 516 3086 535 3142
rect 535 3086 572 3142
rect 516 2978 535 3034
rect 535 2978 572 3034
rect 516 2870 535 2926
rect 535 2870 572 2926
rect 516 2762 535 2818
rect 535 2762 572 2818
rect 516 2654 535 2710
rect 535 2654 572 2710
rect 516 2546 535 2602
rect 535 2546 572 2602
rect 516 2438 535 2494
rect 535 2438 572 2494
rect 516 2330 535 2386
rect 535 2330 572 2386
rect 516 2222 535 2278
rect 535 2222 572 2278
rect 516 2114 535 2170
rect 535 2114 572 2170
rect 516 2006 535 2062
rect 535 2006 572 2062
rect 308 1857 353 1878
rect 353 1857 364 1878
rect 436 1857 447 1878
rect 447 1857 492 1878
rect 308 1822 364 1857
rect 436 1822 492 1857
rect 308 1712 364 1747
rect 436 1712 492 1747
rect 308 1691 343 1712
rect 343 1691 364 1712
rect 436 1691 457 1712
rect 457 1691 492 1712
rect 308 1314 343 1335
rect 343 1314 364 1335
rect 436 1314 457 1335
rect 457 1314 492 1335
rect 308 1279 364 1314
rect 436 1279 492 1314
rect 308 1167 364 1202
rect 436 1167 492 1202
rect 308 1146 353 1167
rect 353 1146 364 1167
rect 436 1146 447 1167
rect 447 1146 492 1167
rect 228 1014 265 1070
rect 265 1014 284 1070
rect 228 906 265 962
rect 265 906 284 962
rect 516 1014 535 1070
rect 535 1014 572 1070
rect 516 906 535 962
rect 535 906 572 962
rect 308 809 353 830
rect 353 809 364 830
rect 436 809 447 830
rect 447 809 492 830
rect 308 774 364 809
rect 436 774 492 809
rect 156 489 212 524
rect 156 468 191 489
rect 191 468 212 489
rect 156 375 191 396
rect 191 375 212 396
rect 156 340 212 375
rect 568 489 624 524
rect 568 468 589 489
rect 589 468 624 489
rect 568 375 589 396
rect 589 375 624 396
rect 568 340 624 375
rect 308 287 364 306
rect 416 287 472 306
rect 308 250 364 287
rect 416 250 472 287
<< metal2 >>
rect 296 4174 484 4176
rect 296 4118 308 4174
rect 364 4118 416 4174
rect 472 4118 484 4174
rect 296 4116 484 4118
rect 132 4084 214 4096
rect 132 4028 156 4084
rect 212 4060 214 4084
rect 566 4084 673 4096
rect 566 4060 568 4084
rect 212 4028 568 4060
rect 624 4028 673 4084
rect 132 3956 673 4028
rect 132 3900 156 3956
rect 212 3924 568 3956
rect 212 3900 214 3924
rect 132 3888 214 3900
rect 566 3900 568 3924
rect 624 3900 673 3956
rect 566 3888 673 3900
rect 296 3650 504 3652
rect 296 3594 308 3650
rect 364 3594 436 3650
rect 492 3594 504 3650
rect 296 3592 504 3594
rect 226 3466 286 3478
rect 226 3408 228 3466
rect 284 3408 286 3466
rect 226 3360 286 3408
rect 226 3302 228 3360
rect 284 3302 286 3360
rect 226 3250 286 3302
rect 226 3192 228 3250
rect 284 3192 286 3250
rect 226 3144 286 3192
rect 226 3086 228 3144
rect 284 3086 286 3144
rect 226 3034 286 3086
rect 226 2976 228 3034
rect 284 2976 286 3034
rect 226 2928 286 2976
rect 226 2870 228 2928
rect 284 2870 286 2928
rect 226 2818 286 2870
rect 226 2760 228 2818
rect 284 2760 286 2818
rect 226 2712 286 2760
rect 226 2654 228 2712
rect 284 2654 286 2712
rect 226 2602 286 2654
rect 226 2544 228 2602
rect 284 2544 286 2602
rect 226 2496 286 2544
rect 226 2438 228 2496
rect 284 2438 286 2496
rect 226 2386 286 2438
rect 226 2328 228 2386
rect 284 2328 286 2386
rect 226 2280 286 2328
rect 226 2222 228 2280
rect 284 2222 286 2280
rect 226 2170 286 2222
rect 226 2112 228 2170
rect 284 2112 286 2170
rect 226 2064 286 2112
rect 226 2006 228 2064
rect 284 2006 286 2064
rect 226 1994 286 2006
rect 342 1880 458 3592
rect 514 3466 574 3478
rect 514 3408 516 3466
rect 572 3408 574 3466
rect 514 3360 574 3408
rect 514 3302 516 3360
rect 572 3302 574 3360
rect 514 3250 574 3302
rect 514 3192 516 3250
rect 572 3192 574 3250
rect 514 3144 574 3192
rect 514 3086 516 3144
rect 572 3086 574 3144
rect 514 3034 574 3086
rect 514 2976 516 3034
rect 572 2976 574 3034
rect 514 2928 574 2976
rect 514 2870 516 2928
rect 572 2870 574 2928
rect 514 2818 574 2870
rect 514 2760 516 2818
rect 572 2760 574 2818
rect 514 2712 574 2760
rect 514 2654 516 2712
rect 572 2654 574 2712
rect 514 2602 574 2654
rect 514 2544 516 2602
rect 572 2544 574 2602
rect 514 2496 574 2544
rect 514 2438 516 2496
rect 572 2438 574 2496
rect 514 2386 574 2438
rect 514 2328 516 2386
rect 572 2328 574 2386
rect 514 2280 574 2328
rect 514 2222 516 2280
rect 572 2222 574 2280
rect 514 2170 574 2222
rect 514 2112 516 2170
rect 572 2112 574 2170
rect 514 2064 574 2112
rect 514 2006 516 2064
rect 572 2006 574 2064
rect 514 1994 574 2006
rect 296 1878 504 1880
rect 296 1822 308 1878
rect 364 1822 436 1878
rect 492 1822 504 1878
rect 296 1747 504 1822
rect 296 1691 308 1747
rect 364 1691 436 1747
rect 492 1691 504 1747
rect 296 1689 504 1691
rect 332 1337 468 1689
rect 296 1335 504 1337
rect 296 1279 308 1335
rect 364 1279 436 1335
rect 492 1279 504 1335
rect 296 1202 504 1279
rect 296 1146 308 1202
rect 364 1146 436 1202
rect 492 1146 504 1202
rect 296 1144 504 1146
rect 226 1070 286 1082
rect 226 1012 228 1070
rect 284 1012 286 1070
rect 226 964 286 1012
rect 226 906 228 964
rect 284 906 286 964
rect 226 894 286 906
rect 342 832 458 1144
rect 514 1070 574 1082
rect 514 1012 516 1070
rect 572 1012 574 1070
rect 514 964 574 1012
rect 514 906 516 964
rect 572 906 574 964
rect 514 894 574 906
rect 296 830 504 832
rect 296 774 308 830
rect 364 774 436 830
rect 492 774 504 830
rect 296 772 504 774
rect 333 764 469 772
rect 107 524 214 536
rect 107 468 156 524
rect 212 500 214 524
rect 566 524 648 536
rect 566 500 568 524
rect 212 468 568 500
rect 624 468 648 524
rect 107 396 648 468
rect 107 340 156 396
rect 212 364 568 396
rect 212 340 214 364
rect 107 328 214 340
rect 566 340 568 364
rect 624 340 648 396
rect 566 328 648 340
rect 296 306 484 308
rect 296 250 308 306
rect 364 250 416 306
rect 472 250 484 306
rect 296 248 484 250
<< via2 >>
rect 228 3410 284 3464
rect 228 3408 284 3410
rect 228 3358 284 3360
rect 228 3304 284 3358
rect 228 3194 284 3248
rect 228 3192 284 3194
rect 228 3142 284 3144
rect 228 3088 284 3142
rect 228 2978 284 3032
rect 228 2976 284 2978
rect 228 2926 284 2928
rect 228 2872 284 2926
rect 228 2762 284 2816
rect 228 2760 284 2762
rect 228 2710 284 2712
rect 228 2656 284 2710
rect 228 2546 284 2600
rect 228 2544 284 2546
rect 228 2494 284 2496
rect 228 2440 284 2494
rect 228 2330 284 2384
rect 228 2328 284 2330
rect 228 2278 284 2280
rect 228 2224 284 2278
rect 228 2114 284 2168
rect 228 2112 284 2114
rect 228 2062 284 2064
rect 228 2008 284 2062
rect 516 3410 572 3464
rect 516 3408 572 3410
rect 516 3358 572 3360
rect 516 3304 572 3358
rect 516 3194 572 3248
rect 516 3192 572 3194
rect 516 3142 572 3144
rect 516 3088 572 3142
rect 516 2978 572 3032
rect 516 2976 572 2978
rect 516 2926 572 2928
rect 516 2872 572 2926
rect 516 2762 572 2816
rect 516 2760 572 2762
rect 516 2710 572 2712
rect 516 2656 572 2710
rect 516 2546 572 2600
rect 516 2544 572 2546
rect 516 2494 572 2496
rect 516 2440 572 2494
rect 516 2330 572 2384
rect 516 2328 572 2330
rect 516 2278 572 2280
rect 516 2224 572 2278
rect 516 2114 572 2168
rect 516 2112 572 2114
rect 516 2062 572 2064
rect 516 2008 572 2062
rect 228 1014 284 1068
rect 228 1012 284 1014
rect 228 962 284 964
rect 228 908 284 962
rect 516 1014 572 1068
rect 516 1012 572 1014
rect 516 962 572 964
rect 516 908 572 962
<< metal3 >>
rect 226 3464 286 3478
rect 226 3408 228 3464
rect 284 3408 286 3464
rect 226 3360 286 3408
rect 226 3304 228 3360
rect 284 3304 286 3360
rect 226 3248 286 3304
rect 226 3192 228 3248
rect 284 3192 286 3248
rect 226 3144 286 3192
rect 226 3088 228 3144
rect 284 3088 286 3144
rect 226 3032 286 3088
rect 226 2976 228 3032
rect 284 2976 286 3032
rect 226 2928 286 2976
rect 226 2872 228 2928
rect 284 2872 286 2928
rect 226 2819 286 2872
rect 514 3464 574 3478
rect 514 3408 516 3464
rect 572 3408 574 3464
rect 514 3360 574 3408
rect 514 3304 516 3360
rect 572 3304 574 3360
rect 514 3248 574 3304
rect 514 3192 516 3248
rect 572 3192 574 3248
rect 514 3144 574 3192
rect 514 3088 516 3144
rect 572 3088 574 3144
rect 514 3032 574 3088
rect 514 2976 516 3032
rect 572 2976 574 3032
rect 514 2928 574 2976
rect 514 2872 516 2928
rect 572 2872 574 2928
rect 514 2819 574 2872
rect 132 2816 673 2819
rect 132 2760 228 2816
rect 284 2760 516 2816
rect 572 2760 673 2816
rect 132 2712 673 2760
rect 132 2656 228 2712
rect 284 2656 516 2712
rect 572 2656 673 2712
rect 132 2654 673 2656
rect 226 2600 286 2654
rect 226 2544 228 2600
rect 284 2544 286 2600
rect 226 2496 286 2544
rect 226 2440 228 2496
rect 284 2440 286 2496
rect 226 2384 286 2440
rect 226 2328 228 2384
rect 284 2328 286 2384
rect 226 2280 286 2328
rect 226 2224 228 2280
rect 284 2224 286 2280
rect 226 2168 286 2224
rect 226 2112 228 2168
rect 284 2112 286 2168
rect 226 2064 286 2112
rect 226 2008 228 2064
rect 284 2008 286 2064
rect 226 1994 286 2008
rect 514 2600 574 2654
rect 514 2544 516 2600
rect 572 2544 574 2600
rect 514 2496 574 2544
rect 514 2440 516 2496
rect 572 2440 574 2496
rect 514 2384 574 2440
rect 514 2328 516 2384
rect 572 2328 574 2384
rect 514 2280 574 2328
rect 514 2224 516 2280
rect 572 2224 574 2280
rect 514 2168 574 2224
rect 514 2112 516 2168
rect 572 2112 574 2168
rect 514 2064 574 2112
rect 514 2008 516 2064
rect 572 2008 574 2064
rect 514 1994 574 2008
rect 112 1068 648 1082
rect 112 1012 228 1068
rect 284 1012 516 1068
rect 572 1012 648 1068
rect 112 964 648 1012
rect 112 908 228 964
rect 284 908 516 964
rect 572 908 648 964
rect 112 894 648 908
<< end >>
