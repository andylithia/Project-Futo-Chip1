// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire net215;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net144;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net145;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net146;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net106;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net107;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net108;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net103;
 wire net104;
 wire net105;
 wire net41;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net42;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net43;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net44;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net45;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net46;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire \u_inj.outn ;
 wire \u_inj.outp ;
 wire \u_inj.signal_n ;
 wire \u_inj.trim_n_r[0] ;
 wire \u_inj.trim_n_r[1] ;
 wire \u_inj.trim_n_r[2] ;
 wire \u_inj.trim_n_r[3] ;
 wire \u_inj.trim_p_r[0] ;
 wire \u_inj.trim_p_r[1] ;
 wire \u_inj.trim_p_r[2] ;
 wire \u_inj.trim_p_r[3] ;
 wire net182;
 wire net183;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net184;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net185;
 wire net213;
 wire net214;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _030_ (.I(net1),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _031_ (.A1(net14),
    .A2(\u_inj.signal_n ),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _032_ (.I(_002_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _033_ (.D(net2),
    .CLK(net10),
    .Q(\u_inj.trim_p_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _034_ (.D(net3),
    .CLK(net10),
    .Q(\u_inj.trim_p_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _035_ (.D(net4),
    .CLK(net10),
    .Q(\u_inj.trim_p_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _036_ (.D(net5),
    .CLK(net10),
    .Q(\u_inj.trim_p_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _037_ (.D(net6),
    .CLK(net10),
    .Q(\u_inj.trim_n_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _038_ (.D(net7),
    .CLK(net10),
    .Q(\u_inj.trim_n_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _039_ (.D(net8),
    .CLK(net10),
    .Q(\u_inj.trim_n_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _040_ (.D(net9),
    .CLK(net10),
    .Q(\u_inj.trim_n_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh \u_inj.psijn_215  (.Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[0].pdp_16  (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[1].pdn_17  (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[1].pdp_18  (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[2].pdn_19  (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[2].pdp_20  (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[3].pdn_21  (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[3].pdp_22  (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[4].pdn_23  (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[4].pdp_24  (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[5].pdn_25  (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[5].pdp_26  (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[6].pdn_27  (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[6].pdp_28  (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[7].pdn_29  (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[7].pdp_30  (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[0].ntrimn_31  (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[0].ntrimp_32  (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[1].ntrimn_33  (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[1].ntrimp_34  (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[2].ntrimn_35  (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[2].ntrimp_36  (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[3].ntrimn_37  (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_TRIM[3].ntrimp_38  (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.siginv_39  (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tieh \u_inj.nsijp_214  (.Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _242_ (.I(\u_inj.outp ),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _243_ (.I(\u_inj.outn ),
    .Z(la_data_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[0].pdn  (.I(net15),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[0].pdp  (.I(net16),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[1].pdn  (.I(net17),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[1].pdp  (.I(net18),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[2].pdn  (.I(net19),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[2].pdp  (.I(net20),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[3].pdn  (.I(net21),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[3].pdp  (.I(net22),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[4].pdn  (.I(net23),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[4].pdp  (.I(net24),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[5].pdn  (.I(net25),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[5].pdp  (.I(net26),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[6].pdn  (.I(net27),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[6].pdp  (.I(net28),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[7].pdn  (.I(net29),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.gen_PD[7].pdp  (.I(net30),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[0].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[0].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[10].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[10].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[11].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[11].pup  (.I(net13),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[12].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[12].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[13].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[13].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[14].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[14].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[15].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[15].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[16].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[16].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[17].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[17].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[18].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[18].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[1].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[1].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[2].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[2].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[3].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[3].pup  (.I(net13),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[4].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[4].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[5].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[5].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[6].pun  (.I(net12),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[6].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[7].pun  (.I(net13),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[7].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[8].pun  (.I(net13),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[8].pup  (.I(net11),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[9].pun  (.I(net13),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \u_inj.gen_PU[9].pup  (.I(net13),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[0].ntrimn  (.EN(\u_inj.trim_n_r[0] ),
    .I(net31),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[0].ntrimp  (.EN(\u_inj.trim_n_r[0] ),
    .I(net32),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[0].ptrimn  (.EN(\u_inj.trim_p_r[0] ),
    .I(net14),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[0].ptrimp  (.EN(\u_inj.trim_p_r[0] ),
    .I(net14),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[1].ntrimn  (.EN(\u_inj.trim_n_r[1] ),
    .I(net33),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[1].ntrimp  (.EN(\u_inj.trim_n_r[1] ),
    .I(net34),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[1].ptrimn  (.EN(\u_inj.trim_p_r[1] ),
    .I(net14),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[1].ptrimp  (.EN(\u_inj.trim_p_r[1] ),
    .I(net14),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[2].ntrimn  (.EN(\u_inj.trim_n_r[2] ),
    .I(net35),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[2].ntrimp  (.EN(\u_inj.trim_n_r[2] ),
    .I(net36),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[2].ptrimn  (.EN(\u_inj.trim_p_r[2] ),
    .I(net14),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[2].ptrimp  (.EN(\u_inj.trim_p_r[2] ),
    .I(net14),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[3].ntrimn  (.EN(\u_inj.trim_n_r[3] ),
    .I(net37),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[3].ntrimp  (.EN(\u_inj.trim_n_r[3] ),
    .I(net38),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[3].ptrimn  (.EN(\u_inj.trim_p_r[3] ),
    .I(net14),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__invz_1 \u_inj.gen_TRIM[3].ptrimp  (.EN(\u_inj.trim_p_r[3] ),
    .I(net14),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.nsijn  (.I(_001_),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.nsijp  (.I(net214),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.psijn  (.I(net215),
    .ZN(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \u_inj.psijp  (.I(_001_),
    .ZN(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \u_inj.siginv  (.I(net39),
    .ZN(\u_inj.signal_n ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(io_in[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(io_in[9]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 fanout11 (.I(net13),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 fanout12 (.I(net13),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout13 (.I(net14),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout14 (.I(_000_),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u_inj.gen_PD[0].pdn_15  (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__I (.I(\u_inj.outn ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__I (.I(\u_inj.outp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__030__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__035__D (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__036__D (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__037__D (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__038__D (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__039__D (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__040__D (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__040__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__039__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__038__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__037__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__036__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__035__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__034__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__033__CLK (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[8].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[7].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[6].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[5].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[4].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[2].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[1].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[18].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[17].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[16].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[15].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[14].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[13].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[12].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[10].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[0].pup_I  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[6].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[5].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[4].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[3].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[2].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[1].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[18].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[17].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[16].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[15].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[14].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[13].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[12].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[11].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[10].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_PU[0].pun_I  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[3].ptrimp_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[3].ptrimn_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[2].ptrimp_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[2].ptrimn_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout13_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[1].ptrimp_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[1].ptrimn_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[0].ptrimp_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_inj.gen_TRIM[0].ptrimn_I  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__031__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1577 ();
 assign io_oeb[0] = net143;
 assign io_oeb[10] = net153;
 assign io_oeb[11] = net154;
 assign io_oeb[12] = net155;
 assign io_oeb[13] = net156;
 assign io_oeb[14] = net157;
 assign io_oeb[15] = net158;
 assign io_oeb[16] = net159;
 assign io_oeb[17] = net160;
 assign io_oeb[18] = net161;
 assign io_oeb[19] = net162;
 assign io_oeb[1] = net144;
 assign io_oeb[20] = net163;
 assign io_oeb[21] = net164;
 assign io_oeb[22] = net165;
 assign io_oeb[23] = net166;
 assign io_oeb[24] = net167;
 assign io_oeb[25] = net168;
 assign io_oeb[26] = net169;
 assign io_oeb[27] = net170;
 assign io_oeb[28] = net171;
 assign io_oeb[29] = net172;
 assign io_oeb[2] = net145;
 assign io_oeb[30] = net173;
 assign io_oeb[31] = net174;
 assign io_oeb[32] = net175;
 assign io_oeb[33] = net176;
 assign io_oeb[34] = net177;
 assign io_oeb[35] = net178;
 assign io_oeb[36] = net179;
 assign io_oeb[37] = net180;
 assign io_oeb[3] = net146;
 assign io_oeb[4] = net147;
 assign io_oeb[5] = net148;
 assign io_oeb[6] = net149;
 assign io_oeb[7] = net150;
 assign io_oeb[8] = net151;
 assign io_oeb[9] = net152;
 assign io_out[0] = net105;
 assign io_out[10] = net115;
 assign io_out[11] = net116;
 assign io_out[12] = net117;
 assign io_out[13] = net118;
 assign io_out[14] = net119;
 assign io_out[15] = net120;
 assign io_out[16] = net121;
 assign io_out[17] = net122;
 assign io_out[18] = net123;
 assign io_out[19] = net124;
 assign io_out[1] = net106;
 assign io_out[20] = net125;
 assign io_out[21] = net126;
 assign io_out[22] = net127;
 assign io_out[23] = net128;
 assign io_out[24] = net129;
 assign io_out[25] = net130;
 assign io_out[26] = net131;
 assign io_out[27] = net132;
 assign io_out[28] = net133;
 assign io_out[29] = net134;
 assign io_out[2] = net107;
 assign io_out[30] = net135;
 assign io_out[31] = net136;
 assign io_out[32] = net137;
 assign io_out[33] = net138;
 assign io_out[34] = net139;
 assign io_out[35] = net140;
 assign io_out[36] = net141;
 assign io_out[37] = net142;
 assign io_out[3] = net108;
 assign io_out[4] = net109;
 assign io_out[5] = net110;
 assign io_out[6] = net111;
 assign io_out[7] = net112;
 assign io_out[8] = net113;
 assign io_out[9] = net114;
 assign irq[0] = net102;
 assign irq[1] = net103;
 assign irq[2] = net104;
 assign la_data_out[0] = net40;
 assign la_data_out[10] = net50;
 assign la_data_out[11] = net51;
 assign la_data_out[12] = net52;
 assign la_data_out[13] = net53;
 assign la_data_out[14] = net54;
 assign la_data_out[15] = net55;
 assign la_data_out[16] = net56;
 assign la_data_out[17] = net57;
 assign la_data_out[18] = net58;
 assign la_data_out[19] = net59;
 assign la_data_out[1] = net41;
 assign la_data_out[20] = net60;
 assign la_data_out[21] = net61;
 assign la_data_out[22] = net62;
 assign la_data_out[23] = net63;
 assign la_data_out[24] = net64;
 assign la_data_out[25] = net65;
 assign la_data_out[26] = net66;
 assign la_data_out[27] = net67;
 assign la_data_out[28] = net68;
 assign la_data_out[29] = net69;
 assign la_data_out[2] = net42;
 assign la_data_out[30] = net70;
 assign la_data_out[31] = net71;
 assign la_data_out[34] = net72;
 assign la_data_out[35] = net73;
 assign la_data_out[36] = net74;
 assign la_data_out[37] = net75;
 assign la_data_out[38] = net76;
 assign la_data_out[39] = net77;
 assign la_data_out[3] = net43;
 assign la_data_out[40] = net78;
 assign la_data_out[41] = net79;
 assign la_data_out[42] = net80;
 assign la_data_out[43] = net81;
 assign la_data_out[44] = net82;
 assign la_data_out[45] = net83;
 assign la_data_out[46] = net84;
 assign la_data_out[47] = net85;
 assign la_data_out[48] = net86;
 assign la_data_out[49] = net87;
 assign la_data_out[4] = net44;
 assign la_data_out[50] = net88;
 assign la_data_out[51] = net89;
 assign la_data_out[52] = net90;
 assign la_data_out[53] = net91;
 assign la_data_out[54] = net92;
 assign la_data_out[55] = net93;
 assign la_data_out[56] = net94;
 assign la_data_out[57] = net95;
 assign la_data_out[58] = net96;
 assign la_data_out[59] = net97;
 assign la_data_out[5] = net45;
 assign la_data_out[60] = net98;
 assign la_data_out[61] = net99;
 assign la_data_out[62] = net100;
 assign la_data_out[63] = net101;
 assign la_data_out[6] = net46;
 assign la_data_out[7] = net47;
 assign la_data_out[8] = net48;
 assign la_data_out[9] = net49;
 assign wbs_ack_o = net181;
 assign wbs_dat_o[0] = net182;
 assign wbs_dat_o[10] = net192;
 assign wbs_dat_o[11] = net193;
 assign wbs_dat_o[12] = net194;
 assign wbs_dat_o[13] = net195;
 assign wbs_dat_o[14] = net196;
 assign wbs_dat_o[15] = net197;
 assign wbs_dat_o[16] = net198;
 assign wbs_dat_o[17] = net199;
 assign wbs_dat_o[18] = net200;
 assign wbs_dat_o[19] = net201;
 assign wbs_dat_o[1] = net183;
 assign wbs_dat_o[20] = net202;
 assign wbs_dat_o[21] = net203;
 assign wbs_dat_o[22] = net204;
 assign wbs_dat_o[23] = net205;
 assign wbs_dat_o[24] = net206;
 assign wbs_dat_o[25] = net207;
 assign wbs_dat_o[26] = net208;
 assign wbs_dat_o[27] = net209;
 assign wbs_dat_o[28] = net210;
 assign wbs_dat_o[29] = net211;
 assign wbs_dat_o[2] = net184;
 assign wbs_dat_o[30] = net212;
 assign wbs_dat_o[31] = net213;
 assign wbs_dat_o[3] = net185;
 assign wbs_dat_o[4] = net186;
 assign wbs_dat_o[5] = net187;
 assign wbs_dat_o[6] = net188;
 assign wbs_dat_o[7] = net189;
 assign wbs_dat_o[8] = net190;
 assign wbs_dat_o[9] = net191;
endmodule

