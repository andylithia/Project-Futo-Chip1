magic
tech gf180mcuC
magscale 1 5
timestamp 1670013958
<< metal1 >>
rect 672 6285 6408 6302
rect 672 6259 2021 6285
rect 2047 6259 2073 6285
rect 2099 6259 2125 6285
rect 2151 6259 3435 6285
rect 3461 6259 3487 6285
rect 3513 6259 3539 6285
rect 3565 6259 4849 6285
rect 4875 6259 4901 6285
rect 4927 6259 4953 6285
rect 4979 6259 6263 6285
rect 6289 6259 6315 6285
rect 6341 6259 6367 6285
rect 6393 6259 6408 6285
rect 672 6242 6408 6259
rect 1807 6201 1833 6207
rect 1807 6169 1833 6175
rect 2927 6145 2953 6151
rect 2927 6113 2953 6119
rect 3655 6145 3681 6151
rect 3655 6113 3681 6119
rect 4271 6145 4297 6151
rect 4271 6113 4297 6119
rect 1135 6089 1161 6095
rect 1135 6057 1161 6063
rect 1415 6089 1441 6095
rect 1415 6057 1441 6063
rect 1751 6089 1777 6095
rect 1751 6057 1777 6063
rect 2087 6089 2113 6095
rect 2087 6057 2113 6063
rect 2423 6089 2449 6095
rect 2423 6057 2449 6063
rect 2479 6089 2505 6095
rect 2479 6057 2505 6063
rect 3263 6089 3289 6095
rect 3263 6057 3289 6063
rect 3599 6089 3625 6095
rect 3599 6057 3625 6063
rect 3935 6089 3961 6095
rect 3935 6057 3961 6063
rect 3991 6089 4017 6095
rect 3991 6057 4017 6063
rect 4327 6089 4353 6095
rect 4327 6057 4353 6063
rect 1079 5977 1105 5983
rect 1079 5945 1105 5951
rect 1471 5977 1497 5983
rect 1471 5945 1497 5951
rect 2143 5977 2169 5983
rect 2143 5945 2169 5951
rect 2983 5977 3009 5983
rect 2983 5945 3009 5951
rect 3319 5977 3345 5983
rect 3319 5945 3345 5951
rect 672 5893 6328 5910
rect 672 5867 1314 5893
rect 1340 5867 1366 5893
rect 1392 5867 1418 5893
rect 1444 5867 2728 5893
rect 2754 5867 2780 5893
rect 2806 5867 2832 5893
rect 2858 5867 4142 5893
rect 4168 5867 4194 5893
rect 4220 5867 4246 5893
rect 4272 5867 5556 5893
rect 5582 5867 5608 5893
rect 5634 5867 5660 5893
rect 5686 5867 6328 5893
rect 672 5850 6328 5867
rect 2423 5809 2449 5815
rect 2423 5777 2449 5783
rect 3039 5809 3065 5815
rect 3039 5777 3065 5783
rect 3375 5809 3401 5815
rect 3375 5777 3401 5783
rect 3935 5809 3961 5815
rect 3935 5777 3961 5783
rect 1079 5697 1105 5703
rect 1079 5665 1105 5671
rect 1807 5697 1833 5703
rect 1807 5665 1833 5671
rect 2143 5697 2169 5703
rect 2143 5665 2169 5671
rect 2479 5697 2505 5703
rect 2479 5665 2505 5671
rect 3095 5697 3121 5703
rect 3095 5665 3121 5671
rect 3431 5697 3457 5703
rect 3431 5665 3457 5671
rect 1471 5641 1497 5647
rect 1471 5609 1497 5615
rect 3991 5641 4017 5647
rect 3991 5609 4017 5615
rect 4271 5641 4297 5647
rect 4271 5609 4297 5615
rect 4327 5641 4353 5647
rect 4327 5609 4353 5615
rect 1135 5585 1161 5591
rect 1135 5553 1161 5559
rect 1415 5585 1441 5591
rect 1415 5553 1441 5559
rect 1751 5585 1777 5591
rect 1751 5553 1777 5559
rect 2087 5585 2113 5591
rect 2087 5553 2113 5559
rect 672 5501 6408 5518
rect 672 5475 2021 5501
rect 2047 5475 2073 5501
rect 2099 5475 2125 5501
rect 2151 5475 3435 5501
rect 3461 5475 3487 5501
rect 3513 5475 3539 5501
rect 3565 5475 4849 5501
rect 4875 5475 4901 5501
rect 4927 5475 4953 5501
rect 4979 5475 6263 5501
rect 6289 5475 6315 5501
rect 6341 5475 6367 5501
rect 6393 5475 6408 5501
rect 672 5458 6408 5475
rect 3879 5417 3905 5423
rect 3879 5385 3905 5391
rect 2479 5361 2505 5367
rect 2479 5329 2505 5335
rect 3543 5361 3569 5367
rect 3543 5329 3569 5335
rect 4215 5361 4241 5367
rect 4215 5329 4241 5335
rect 1135 5305 1161 5311
rect 1135 5273 1161 5279
rect 1471 5305 1497 5311
rect 1471 5273 1497 5279
rect 1527 5305 1553 5311
rect 1527 5273 1553 5279
rect 1807 5305 1833 5311
rect 1807 5273 1833 5279
rect 1863 5305 1889 5311
rect 1863 5273 1889 5279
rect 2143 5305 2169 5311
rect 2143 5273 2169 5279
rect 2815 5305 2841 5311
rect 2815 5273 2841 5279
rect 2871 5305 2897 5311
rect 2871 5273 2897 5279
rect 3151 5305 3177 5311
rect 3151 5273 3177 5279
rect 3207 5305 3233 5311
rect 3207 5273 3233 5279
rect 3487 5305 3513 5311
rect 3487 5273 3513 5279
rect 3823 5305 3849 5311
rect 3823 5273 3849 5279
rect 4159 5305 4185 5311
rect 4159 5273 4185 5279
rect 1191 5193 1217 5199
rect 1191 5161 1217 5167
rect 2199 5193 2225 5199
rect 2199 5161 2225 5167
rect 2535 5193 2561 5199
rect 2535 5161 2561 5167
rect 672 5109 6328 5126
rect 672 5083 1314 5109
rect 1340 5083 1366 5109
rect 1392 5083 1418 5109
rect 1444 5083 2728 5109
rect 2754 5083 2780 5109
rect 2806 5083 2832 5109
rect 2858 5083 4142 5109
rect 4168 5083 4194 5109
rect 4220 5083 4246 5109
rect 4272 5083 5556 5109
rect 5582 5083 5608 5109
rect 5634 5083 5660 5109
rect 5686 5083 6328 5109
rect 672 5066 6328 5083
rect 1415 5025 1441 5031
rect 1415 4993 1441 4999
rect 1751 5025 1777 5031
rect 1751 4993 1777 4999
rect 3095 5025 3121 5031
rect 3095 4993 3121 4999
rect 3431 5025 3457 5031
rect 3431 4993 3457 4999
rect 1079 4913 1105 4919
rect 1079 4881 1105 4887
rect 1807 4913 1833 4919
rect 1807 4881 1833 4887
rect 2087 4913 2113 4919
rect 2087 4881 2113 4887
rect 2423 4913 2449 4919
rect 2423 4881 2449 4887
rect 2479 4913 2505 4919
rect 2479 4881 2505 4887
rect 3151 4913 3177 4919
rect 3151 4881 3177 4887
rect 1471 4857 1497 4863
rect 1471 4825 1497 4831
rect 3487 4857 3513 4863
rect 3487 4825 3513 4831
rect 3823 4857 3849 4863
rect 3823 4825 3849 4831
rect 1135 4801 1161 4807
rect 1135 4769 1161 4775
rect 2143 4801 2169 4807
rect 2143 4769 2169 4775
rect 3767 4801 3793 4807
rect 3767 4769 3793 4775
rect 672 4717 6408 4734
rect 672 4691 2021 4717
rect 2047 4691 2073 4717
rect 2099 4691 2125 4717
rect 2151 4691 3435 4717
rect 3461 4691 3487 4717
rect 3513 4691 3539 4717
rect 3565 4691 4849 4717
rect 4875 4691 4901 4717
rect 4927 4691 4953 4717
rect 4979 4691 6263 4717
rect 6289 4691 6315 4717
rect 6341 4691 6367 4717
rect 6393 4691 6408 4717
rect 672 4674 6408 4691
rect 1191 4633 1217 4639
rect 1191 4601 1217 4607
rect 2871 4633 2897 4639
rect 2871 4601 2897 4607
rect 3207 4633 3233 4639
rect 3207 4601 3233 4607
rect 3543 4633 3569 4639
rect 3543 4601 3569 4607
rect 1527 4577 1553 4583
rect 1527 4545 1553 4551
rect 2143 4577 2169 4583
rect 2143 4545 2169 4551
rect 3151 4577 3177 4583
rect 3151 4545 3177 4551
rect 3487 4577 3513 4583
rect 3487 4545 3513 4551
rect 1135 4521 1161 4527
rect 1135 4489 1161 4495
rect 1471 4521 1497 4527
rect 1471 4489 1497 4495
rect 1807 4521 1833 4527
rect 1807 4489 1833 4495
rect 2479 4521 2505 4527
rect 2479 4489 2505 4495
rect 2815 4521 2841 4527
rect 2815 4489 2841 4495
rect 3879 4521 3905 4527
rect 3879 4489 3905 4495
rect 1863 4409 1889 4415
rect 1863 4377 1889 4383
rect 2199 4409 2225 4415
rect 2199 4377 2225 4383
rect 2535 4409 2561 4415
rect 2535 4377 2561 4383
rect 3823 4409 3849 4415
rect 3823 4377 3849 4383
rect 672 4325 6328 4342
rect 672 4299 1314 4325
rect 1340 4299 1366 4325
rect 1392 4299 1418 4325
rect 1444 4299 2728 4325
rect 2754 4299 2780 4325
rect 2806 4299 2832 4325
rect 2858 4299 4142 4325
rect 4168 4299 4194 4325
rect 4220 4299 4246 4325
rect 4272 4299 5556 4325
rect 5582 4299 5608 4325
rect 5634 4299 5660 4325
rect 5686 4299 6328 4325
rect 672 4282 6328 4299
rect 1527 4241 1553 4247
rect 1527 4209 1553 4215
rect 2311 4241 2337 4247
rect 2311 4209 2337 4215
rect 3095 4241 3121 4247
rect 3095 4209 3121 4215
rect 2031 4185 2057 4191
rect 2031 4153 2057 4159
rect 3431 4185 3457 4191
rect 3431 4153 3457 4159
rect 1583 4129 1609 4135
rect 1583 4097 1609 4103
rect 1975 4129 2001 4135
rect 1975 4097 2001 4103
rect 2367 4129 2393 4135
rect 2367 4097 2393 4103
rect 3151 4129 3177 4135
rect 3151 4097 3177 4103
rect 1079 4073 1105 4079
rect 1079 4041 1105 4047
rect 3487 4073 3513 4079
rect 3487 4041 3513 4047
rect 3767 4073 3793 4079
rect 3767 4041 3793 4047
rect 3823 4073 3849 4079
rect 3823 4041 3849 4047
rect 4103 4073 4129 4079
rect 4103 4041 4129 4047
rect 4159 4017 4185 4023
rect 4159 3985 4185 3991
rect 672 3933 6408 3950
rect 672 3907 2021 3933
rect 2047 3907 2073 3933
rect 2099 3907 2125 3933
rect 2151 3907 3435 3933
rect 3461 3907 3487 3933
rect 3513 3907 3539 3933
rect 3565 3907 4849 3933
rect 4875 3907 4901 3933
rect 4927 3907 4953 3933
rect 4979 3907 6263 3933
rect 6289 3907 6315 3933
rect 6341 3907 6367 3933
rect 6393 3907 6408 3933
rect 672 3890 6408 3907
rect 1359 3849 1385 3855
rect 1359 3817 1385 3823
rect 2703 3849 2729 3855
rect 2703 3817 2729 3823
rect 3039 3849 3065 3855
rect 3039 3817 3065 3823
rect 2367 3793 2393 3799
rect 2367 3761 2393 3767
rect 3375 3793 3401 3799
rect 3375 3761 3401 3767
rect 967 3737 993 3743
rect 967 3705 993 3711
rect 1303 3737 1329 3743
rect 1303 3705 1329 3711
rect 1639 3737 1665 3743
rect 1639 3705 1665 3711
rect 1975 3737 2001 3743
rect 1975 3705 2001 3711
rect 2311 3737 2337 3743
rect 2311 3705 2337 3711
rect 2647 3737 2673 3743
rect 2647 3705 2673 3711
rect 2983 3737 3009 3743
rect 2983 3705 3009 3711
rect 3319 3737 3345 3743
rect 3319 3705 3345 3711
rect 3711 3737 3737 3743
rect 3711 3705 3737 3711
rect 4047 3737 4073 3743
rect 4047 3705 4073 3711
rect 4327 3737 4353 3743
rect 4327 3705 4353 3711
rect 4383 3737 4409 3743
rect 4383 3705 4409 3711
rect 1023 3625 1049 3631
rect 1023 3593 1049 3599
rect 1695 3625 1721 3631
rect 1695 3593 1721 3599
rect 2031 3625 2057 3631
rect 2031 3593 2057 3599
rect 3655 3625 3681 3631
rect 3655 3593 3681 3599
rect 3991 3625 4017 3631
rect 3991 3593 4017 3599
rect 672 3541 6328 3558
rect 672 3515 1314 3541
rect 1340 3515 1366 3541
rect 1392 3515 1418 3541
rect 1444 3515 2728 3541
rect 2754 3515 2780 3541
rect 2806 3515 2832 3541
rect 2858 3515 4142 3541
rect 4168 3515 4194 3541
rect 4220 3515 4246 3541
rect 4272 3515 5556 3541
rect 5582 3515 5608 3541
rect 5634 3515 5660 3541
rect 5686 3515 6328 3541
rect 672 3498 6328 3515
rect 1415 3457 1441 3463
rect 1415 3425 1441 3431
rect 2983 3457 3009 3463
rect 2983 3425 3009 3431
rect 3375 3457 3401 3463
rect 3375 3425 3401 3431
rect 4327 3457 4353 3463
rect 4327 3425 4353 3431
rect 1135 3345 1161 3351
rect 1135 3313 1161 3319
rect 1807 3345 1833 3351
rect 1807 3313 1833 3319
rect 2199 3345 2225 3351
rect 2199 3313 2225 3319
rect 2255 3345 2281 3351
rect 2255 3313 2281 3319
rect 3039 3345 3065 3351
rect 3039 3313 3065 3319
rect 4383 3345 4409 3351
rect 4383 3313 4409 3319
rect 1471 3289 1497 3295
rect 1471 3257 1497 3263
rect 1751 3289 1777 3295
rect 1751 3257 1777 3263
rect 3319 3289 3345 3295
rect 3319 3257 3345 3263
rect 3711 3289 3737 3295
rect 3711 3257 3737 3263
rect 4047 3289 4073 3295
rect 4047 3257 4073 3263
rect 4663 3289 4689 3295
rect 4663 3257 4689 3263
rect 1079 3233 1105 3239
rect 1079 3201 1105 3207
rect 3655 3233 3681 3239
rect 3655 3201 3681 3207
rect 3991 3233 4017 3239
rect 3991 3201 4017 3207
rect 4719 3233 4745 3239
rect 4719 3201 4745 3207
rect 672 3149 6408 3166
rect 672 3123 2021 3149
rect 2047 3123 2073 3149
rect 2099 3123 2125 3149
rect 2151 3123 3435 3149
rect 3461 3123 3487 3149
rect 3513 3123 3539 3149
rect 3565 3123 4849 3149
rect 4875 3123 4901 3149
rect 4927 3123 4953 3149
rect 4979 3123 6263 3149
rect 6289 3123 6315 3149
rect 6341 3123 6367 3149
rect 6393 3123 6408 3149
rect 672 3106 6408 3123
rect 2311 3065 2337 3071
rect 2311 3033 2337 3039
rect 3151 3065 3177 3071
rect 3151 3033 3177 3039
rect 3487 3065 3513 3071
rect 3487 3033 3513 3039
rect 1023 3009 1049 3015
rect 1023 2977 1049 2983
rect 2759 3009 2785 3015
rect 2759 2977 2785 2983
rect 3095 3009 3121 3015
rect 3095 2977 3121 2983
rect 3767 3009 3793 3015
rect 3767 2977 3793 2983
rect 1303 2953 1329 2959
rect 1303 2921 1329 2927
rect 1639 2953 1665 2959
rect 1639 2921 1665 2927
rect 1695 2953 1721 2959
rect 1695 2921 1721 2927
rect 1975 2953 2001 2959
rect 1975 2921 2001 2927
rect 2031 2953 2057 2959
rect 2031 2921 2057 2927
rect 2367 2953 2393 2959
rect 2367 2921 2393 2927
rect 2815 2953 2841 2959
rect 2815 2921 2841 2927
rect 3431 2953 3457 2959
rect 3431 2921 3457 2927
rect 3823 2953 3849 2959
rect 3823 2921 3849 2927
rect 4103 2953 4129 2959
rect 4103 2921 4129 2927
rect 4159 2953 4185 2959
rect 4159 2921 4185 2927
rect 4439 2953 4465 2959
rect 4439 2921 4465 2927
rect 4887 2953 4913 2959
rect 4887 2921 4913 2927
rect 5223 2953 5249 2959
rect 5223 2921 5249 2927
rect 967 2841 993 2847
rect 967 2809 993 2815
rect 1359 2841 1385 2847
rect 1359 2809 1385 2815
rect 4495 2841 4521 2847
rect 4495 2809 4521 2815
rect 4943 2841 4969 2847
rect 4943 2809 4969 2815
rect 5279 2841 5305 2847
rect 5279 2809 5305 2815
rect 672 2757 6328 2774
rect 672 2731 1314 2757
rect 1340 2731 1366 2757
rect 1392 2731 1418 2757
rect 1444 2731 2728 2757
rect 2754 2731 2780 2757
rect 2806 2731 2832 2757
rect 2858 2731 4142 2757
rect 4168 2731 4194 2757
rect 4220 2731 4246 2757
rect 4272 2731 5556 2757
rect 5582 2731 5608 2757
rect 5634 2731 5660 2757
rect 5686 2731 6328 2757
rect 672 2714 6328 2731
rect 1527 2673 1553 2679
rect 1527 2641 1553 2647
rect 1863 2673 1889 2679
rect 1863 2641 1889 2647
rect 2423 2673 2449 2679
rect 2423 2641 2449 2647
rect 5223 2673 5249 2679
rect 5223 2641 5249 2647
rect 5895 2673 5921 2679
rect 5895 2641 5921 2647
rect 4215 2617 4241 2623
rect 4215 2585 4241 2591
rect 1023 2561 1049 2567
rect 1023 2529 1049 2535
rect 1919 2561 1945 2567
rect 1919 2529 1945 2535
rect 2367 2561 2393 2567
rect 2367 2529 2393 2535
rect 2871 2561 2897 2567
rect 2871 2529 2897 2535
rect 3207 2561 3233 2567
rect 3207 2529 3233 2535
rect 3263 2561 3289 2567
rect 3263 2529 3289 2535
rect 3543 2561 3569 2567
rect 3543 2529 3569 2535
rect 3599 2561 3625 2567
rect 3599 2529 3625 2535
rect 3935 2561 3961 2567
rect 3935 2529 3961 2535
rect 4271 2561 4297 2567
rect 4271 2529 4297 2535
rect 4887 2561 4913 2567
rect 4887 2529 4913 2535
rect 4943 2561 4969 2567
rect 4943 2529 4969 2535
rect 5279 2561 5305 2567
rect 5279 2529 5305 2535
rect 5559 2561 5585 2567
rect 5559 2529 5585 2535
rect 5951 2561 5977 2567
rect 5951 2529 5977 2535
rect 1583 2505 1609 2511
rect 1583 2473 1609 2479
rect 3879 2505 3905 2511
rect 3879 2473 3905 2479
rect 4607 2505 4633 2511
rect 4607 2473 4633 2479
rect 967 2449 993 2455
rect 967 2417 993 2423
rect 2927 2449 2953 2455
rect 2927 2417 2953 2423
rect 4551 2449 4577 2455
rect 4551 2417 4577 2423
rect 5615 2449 5641 2455
rect 5615 2417 5641 2423
rect 672 2365 6408 2382
rect 672 2339 2021 2365
rect 2047 2339 2073 2365
rect 2099 2339 2125 2365
rect 2151 2339 3435 2365
rect 3461 2339 3487 2365
rect 3513 2339 3539 2365
rect 3565 2339 4849 2365
rect 4875 2339 4901 2365
rect 4927 2339 4953 2365
rect 4979 2339 6263 2365
rect 6289 2339 6315 2365
rect 6341 2339 6367 2365
rect 6393 2339 6408 2365
rect 672 2322 6408 2339
rect 1191 2281 1217 2287
rect 1191 2249 1217 2255
rect 1527 2281 1553 2287
rect 1527 2249 1553 2255
rect 3039 2281 3065 2287
rect 3039 2249 3065 2255
rect 3935 2281 3961 2287
rect 3935 2249 3961 2255
rect 5223 2281 5249 2287
rect 5223 2249 5249 2255
rect 5895 2281 5921 2287
rect 5895 2249 5921 2255
rect 1471 2225 1497 2231
rect 1471 2193 1497 2199
rect 2367 2225 2393 2231
rect 2367 2193 2393 2199
rect 3375 2225 3401 2231
rect 3375 2193 3401 2199
rect 4943 2225 4969 2231
rect 4943 2193 4969 2199
rect 5559 2225 5585 2231
rect 5559 2193 5585 2199
rect 1135 2169 1161 2175
rect 1135 2137 1161 2143
rect 1975 2169 2001 2175
rect 1975 2137 2001 2143
rect 2311 2169 2337 2175
rect 2311 2137 2337 2143
rect 2647 2169 2673 2175
rect 2647 2137 2673 2143
rect 2703 2169 2729 2175
rect 2703 2137 2729 2143
rect 2983 2169 3009 2175
rect 2983 2137 3009 2143
rect 3319 2169 3345 2175
rect 3319 2137 3345 2143
rect 3991 2169 4017 2175
rect 3991 2137 4017 2143
rect 4271 2169 4297 2175
rect 4271 2137 4297 2143
rect 4327 2169 4353 2175
rect 4327 2137 4353 2143
rect 5279 2169 5305 2175
rect 5279 2137 5305 2143
rect 5615 2169 5641 2175
rect 5615 2137 5641 2143
rect 5951 2169 5977 2175
rect 5951 2137 5977 2143
rect 4887 2113 4913 2119
rect 4887 2081 4913 2087
rect 2031 2057 2057 2063
rect 2031 2025 2057 2031
rect 672 1973 6328 1990
rect 672 1947 1314 1973
rect 1340 1947 1366 1973
rect 1392 1947 1418 1973
rect 1444 1947 2728 1973
rect 2754 1947 2780 1973
rect 2806 1947 2832 1973
rect 2858 1947 4142 1973
rect 4168 1947 4194 1973
rect 4220 1947 4246 1973
rect 4272 1947 5556 1973
rect 5582 1947 5608 1973
rect 5634 1947 5660 1973
rect 5686 1947 6328 1973
rect 672 1930 6328 1947
rect 1751 1889 1777 1895
rect 1751 1857 1777 1863
rect 2031 1889 2057 1895
rect 2031 1857 2057 1863
rect 3879 1889 3905 1895
rect 3879 1857 3905 1863
rect 5223 1889 5249 1895
rect 5223 1857 5249 1863
rect 1079 1833 1105 1839
rect 1079 1801 1105 1807
rect 4831 1833 4857 1839
rect 4831 1801 4857 1807
rect 1023 1777 1049 1783
rect 1023 1745 1049 1751
rect 1359 1777 1385 1783
rect 1359 1745 1385 1751
rect 2423 1777 2449 1783
rect 2423 1745 2449 1751
rect 3151 1777 3177 1783
rect 3151 1745 3177 1751
rect 3543 1777 3569 1783
rect 3543 1745 3569 1751
rect 3823 1777 3849 1783
rect 3823 1745 3849 1751
rect 4159 1777 4185 1783
rect 4159 1745 4185 1751
rect 4215 1777 4241 1783
rect 4215 1745 4241 1751
rect 4887 1777 4913 1783
rect 4887 1745 4913 1751
rect 5167 1777 5193 1783
rect 5167 1745 5193 1751
rect 5503 1777 5529 1783
rect 5503 1745 5529 1751
rect 5895 1777 5921 1783
rect 5895 1745 5921 1751
rect 1415 1721 1441 1727
rect 1415 1689 1441 1695
rect 1695 1721 1721 1727
rect 1695 1689 1721 1695
rect 2087 1721 2113 1727
rect 2087 1689 2113 1695
rect 2367 1721 2393 1727
rect 2367 1689 2393 1695
rect 3207 1721 3233 1727
rect 3207 1689 3233 1695
rect 3487 1721 3513 1727
rect 3487 1689 3513 1695
rect 5559 1721 5585 1727
rect 5559 1689 5585 1695
rect 5839 1721 5865 1727
rect 5839 1689 5865 1695
rect 672 1581 6408 1598
rect 672 1555 2021 1581
rect 2047 1555 2073 1581
rect 2099 1555 2125 1581
rect 2151 1555 3435 1581
rect 3461 1555 3487 1581
rect 3513 1555 3539 1581
rect 3565 1555 4849 1581
rect 4875 1555 4901 1581
rect 4927 1555 4953 1581
rect 4979 1555 6263 1581
rect 6289 1555 6315 1581
rect 6341 1555 6367 1581
rect 6393 1555 6408 1581
rect 672 1538 6408 1555
<< via1 >>
rect 2021 6259 2047 6285
rect 2073 6259 2099 6285
rect 2125 6259 2151 6285
rect 3435 6259 3461 6285
rect 3487 6259 3513 6285
rect 3539 6259 3565 6285
rect 4849 6259 4875 6285
rect 4901 6259 4927 6285
rect 4953 6259 4979 6285
rect 6263 6259 6289 6285
rect 6315 6259 6341 6285
rect 6367 6259 6393 6285
rect 1807 6175 1833 6201
rect 2927 6119 2953 6145
rect 3655 6119 3681 6145
rect 4271 6119 4297 6145
rect 1135 6063 1161 6089
rect 1415 6063 1441 6089
rect 1751 6063 1777 6089
rect 2087 6063 2113 6089
rect 2423 6063 2449 6089
rect 2479 6063 2505 6089
rect 3263 6063 3289 6089
rect 3599 6063 3625 6089
rect 3935 6063 3961 6089
rect 3991 6063 4017 6089
rect 4327 6063 4353 6089
rect 1079 5951 1105 5977
rect 1471 5951 1497 5977
rect 2143 5951 2169 5977
rect 2983 5951 3009 5977
rect 3319 5951 3345 5977
rect 1314 5867 1340 5893
rect 1366 5867 1392 5893
rect 1418 5867 1444 5893
rect 2728 5867 2754 5893
rect 2780 5867 2806 5893
rect 2832 5867 2858 5893
rect 4142 5867 4168 5893
rect 4194 5867 4220 5893
rect 4246 5867 4272 5893
rect 5556 5867 5582 5893
rect 5608 5867 5634 5893
rect 5660 5867 5686 5893
rect 2423 5783 2449 5809
rect 3039 5783 3065 5809
rect 3375 5783 3401 5809
rect 3935 5783 3961 5809
rect 1079 5671 1105 5697
rect 1807 5671 1833 5697
rect 2143 5671 2169 5697
rect 2479 5671 2505 5697
rect 3095 5671 3121 5697
rect 3431 5671 3457 5697
rect 1471 5615 1497 5641
rect 3991 5615 4017 5641
rect 4271 5615 4297 5641
rect 4327 5615 4353 5641
rect 1135 5559 1161 5585
rect 1415 5559 1441 5585
rect 1751 5559 1777 5585
rect 2087 5559 2113 5585
rect 2021 5475 2047 5501
rect 2073 5475 2099 5501
rect 2125 5475 2151 5501
rect 3435 5475 3461 5501
rect 3487 5475 3513 5501
rect 3539 5475 3565 5501
rect 4849 5475 4875 5501
rect 4901 5475 4927 5501
rect 4953 5475 4979 5501
rect 6263 5475 6289 5501
rect 6315 5475 6341 5501
rect 6367 5475 6393 5501
rect 3879 5391 3905 5417
rect 2479 5335 2505 5361
rect 3543 5335 3569 5361
rect 4215 5335 4241 5361
rect 1135 5279 1161 5305
rect 1471 5279 1497 5305
rect 1527 5279 1553 5305
rect 1807 5279 1833 5305
rect 1863 5279 1889 5305
rect 2143 5279 2169 5305
rect 2815 5279 2841 5305
rect 2871 5279 2897 5305
rect 3151 5279 3177 5305
rect 3207 5279 3233 5305
rect 3487 5279 3513 5305
rect 3823 5279 3849 5305
rect 4159 5279 4185 5305
rect 1191 5167 1217 5193
rect 2199 5167 2225 5193
rect 2535 5167 2561 5193
rect 1314 5083 1340 5109
rect 1366 5083 1392 5109
rect 1418 5083 1444 5109
rect 2728 5083 2754 5109
rect 2780 5083 2806 5109
rect 2832 5083 2858 5109
rect 4142 5083 4168 5109
rect 4194 5083 4220 5109
rect 4246 5083 4272 5109
rect 5556 5083 5582 5109
rect 5608 5083 5634 5109
rect 5660 5083 5686 5109
rect 1415 4999 1441 5025
rect 1751 4999 1777 5025
rect 3095 4999 3121 5025
rect 3431 4999 3457 5025
rect 1079 4887 1105 4913
rect 1807 4887 1833 4913
rect 2087 4887 2113 4913
rect 2423 4887 2449 4913
rect 2479 4887 2505 4913
rect 3151 4887 3177 4913
rect 1471 4831 1497 4857
rect 3487 4831 3513 4857
rect 3823 4831 3849 4857
rect 1135 4775 1161 4801
rect 2143 4775 2169 4801
rect 3767 4775 3793 4801
rect 2021 4691 2047 4717
rect 2073 4691 2099 4717
rect 2125 4691 2151 4717
rect 3435 4691 3461 4717
rect 3487 4691 3513 4717
rect 3539 4691 3565 4717
rect 4849 4691 4875 4717
rect 4901 4691 4927 4717
rect 4953 4691 4979 4717
rect 6263 4691 6289 4717
rect 6315 4691 6341 4717
rect 6367 4691 6393 4717
rect 1191 4607 1217 4633
rect 2871 4607 2897 4633
rect 3207 4607 3233 4633
rect 3543 4607 3569 4633
rect 1527 4551 1553 4577
rect 2143 4551 2169 4577
rect 3151 4551 3177 4577
rect 3487 4551 3513 4577
rect 1135 4495 1161 4521
rect 1471 4495 1497 4521
rect 1807 4495 1833 4521
rect 2479 4495 2505 4521
rect 2815 4495 2841 4521
rect 3879 4495 3905 4521
rect 1863 4383 1889 4409
rect 2199 4383 2225 4409
rect 2535 4383 2561 4409
rect 3823 4383 3849 4409
rect 1314 4299 1340 4325
rect 1366 4299 1392 4325
rect 1418 4299 1444 4325
rect 2728 4299 2754 4325
rect 2780 4299 2806 4325
rect 2832 4299 2858 4325
rect 4142 4299 4168 4325
rect 4194 4299 4220 4325
rect 4246 4299 4272 4325
rect 5556 4299 5582 4325
rect 5608 4299 5634 4325
rect 5660 4299 5686 4325
rect 1527 4215 1553 4241
rect 2311 4215 2337 4241
rect 3095 4215 3121 4241
rect 2031 4159 2057 4185
rect 3431 4159 3457 4185
rect 1583 4103 1609 4129
rect 1975 4103 2001 4129
rect 2367 4103 2393 4129
rect 3151 4103 3177 4129
rect 1079 4047 1105 4073
rect 3487 4047 3513 4073
rect 3767 4047 3793 4073
rect 3823 4047 3849 4073
rect 4103 4047 4129 4073
rect 4159 3991 4185 4017
rect 2021 3907 2047 3933
rect 2073 3907 2099 3933
rect 2125 3907 2151 3933
rect 3435 3907 3461 3933
rect 3487 3907 3513 3933
rect 3539 3907 3565 3933
rect 4849 3907 4875 3933
rect 4901 3907 4927 3933
rect 4953 3907 4979 3933
rect 6263 3907 6289 3933
rect 6315 3907 6341 3933
rect 6367 3907 6393 3933
rect 1359 3823 1385 3849
rect 2703 3823 2729 3849
rect 3039 3823 3065 3849
rect 2367 3767 2393 3793
rect 3375 3767 3401 3793
rect 967 3711 993 3737
rect 1303 3711 1329 3737
rect 1639 3711 1665 3737
rect 1975 3711 2001 3737
rect 2311 3711 2337 3737
rect 2647 3711 2673 3737
rect 2983 3711 3009 3737
rect 3319 3711 3345 3737
rect 3711 3711 3737 3737
rect 4047 3711 4073 3737
rect 4327 3711 4353 3737
rect 4383 3711 4409 3737
rect 1023 3599 1049 3625
rect 1695 3599 1721 3625
rect 2031 3599 2057 3625
rect 3655 3599 3681 3625
rect 3991 3599 4017 3625
rect 1314 3515 1340 3541
rect 1366 3515 1392 3541
rect 1418 3515 1444 3541
rect 2728 3515 2754 3541
rect 2780 3515 2806 3541
rect 2832 3515 2858 3541
rect 4142 3515 4168 3541
rect 4194 3515 4220 3541
rect 4246 3515 4272 3541
rect 5556 3515 5582 3541
rect 5608 3515 5634 3541
rect 5660 3515 5686 3541
rect 1415 3431 1441 3457
rect 2983 3431 3009 3457
rect 3375 3431 3401 3457
rect 4327 3431 4353 3457
rect 1135 3319 1161 3345
rect 1807 3319 1833 3345
rect 2199 3319 2225 3345
rect 2255 3319 2281 3345
rect 3039 3319 3065 3345
rect 4383 3319 4409 3345
rect 1471 3263 1497 3289
rect 1751 3263 1777 3289
rect 3319 3263 3345 3289
rect 3711 3263 3737 3289
rect 4047 3263 4073 3289
rect 4663 3263 4689 3289
rect 1079 3207 1105 3233
rect 3655 3207 3681 3233
rect 3991 3207 4017 3233
rect 4719 3207 4745 3233
rect 2021 3123 2047 3149
rect 2073 3123 2099 3149
rect 2125 3123 2151 3149
rect 3435 3123 3461 3149
rect 3487 3123 3513 3149
rect 3539 3123 3565 3149
rect 4849 3123 4875 3149
rect 4901 3123 4927 3149
rect 4953 3123 4979 3149
rect 6263 3123 6289 3149
rect 6315 3123 6341 3149
rect 6367 3123 6393 3149
rect 2311 3039 2337 3065
rect 3151 3039 3177 3065
rect 3487 3039 3513 3065
rect 1023 2983 1049 3009
rect 2759 2983 2785 3009
rect 3095 2983 3121 3009
rect 3767 2983 3793 3009
rect 1303 2927 1329 2953
rect 1639 2927 1665 2953
rect 1695 2927 1721 2953
rect 1975 2927 2001 2953
rect 2031 2927 2057 2953
rect 2367 2927 2393 2953
rect 2815 2927 2841 2953
rect 3431 2927 3457 2953
rect 3823 2927 3849 2953
rect 4103 2927 4129 2953
rect 4159 2927 4185 2953
rect 4439 2927 4465 2953
rect 4887 2927 4913 2953
rect 5223 2927 5249 2953
rect 967 2815 993 2841
rect 1359 2815 1385 2841
rect 4495 2815 4521 2841
rect 4943 2815 4969 2841
rect 5279 2815 5305 2841
rect 1314 2731 1340 2757
rect 1366 2731 1392 2757
rect 1418 2731 1444 2757
rect 2728 2731 2754 2757
rect 2780 2731 2806 2757
rect 2832 2731 2858 2757
rect 4142 2731 4168 2757
rect 4194 2731 4220 2757
rect 4246 2731 4272 2757
rect 5556 2731 5582 2757
rect 5608 2731 5634 2757
rect 5660 2731 5686 2757
rect 1527 2647 1553 2673
rect 1863 2647 1889 2673
rect 2423 2647 2449 2673
rect 5223 2647 5249 2673
rect 5895 2647 5921 2673
rect 4215 2591 4241 2617
rect 1023 2535 1049 2561
rect 1919 2535 1945 2561
rect 2367 2535 2393 2561
rect 2871 2535 2897 2561
rect 3207 2535 3233 2561
rect 3263 2535 3289 2561
rect 3543 2535 3569 2561
rect 3599 2535 3625 2561
rect 3935 2535 3961 2561
rect 4271 2535 4297 2561
rect 4887 2535 4913 2561
rect 4943 2535 4969 2561
rect 5279 2535 5305 2561
rect 5559 2535 5585 2561
rect 5951 2535 5977 2561
rect 1583 2479 1609 2505
rect 3879 2479 3905 2505
rect 4607 2479 4633 2505
rect 967 2423 993 2449
rect 2927 2423 2953 2449
rect 4551 2423 4577 2449
rect 5615 2423 5641 2449
rect 2021 2339 2047 2365
rect 2073 2339 2099 2365
rect 2125 2339 2151 2365
rect 3435 2339 3461 2365
rect 3487 2339 3513 2365
rect 3539 2339 3565 2365
rect 4849 2339 4875 2365
rect 4901 2339 4927 2365
rect 4953 2339 4979 2365
rect 6263 2339 6289 2365
rect 6315 2339 6341 2365
rect 6367 2339 6393 2365
rect 1191 2255 1217 2281
rect 1527 2255 1553 2281
rect 3039 2255 3065 2281
rect 3935 2255 3961 2281
rect 5223 2255 5249 2281
rect 5895 2255 5921 2281
rect 1471 2199 1497 2225
rect 2367 2199 2393 2225
rect 3375 2199 3401 2225
rect 4943 2199 4969 2225
rect 5559 2199 5585 2225
rect 1135 2143 1161 2169
rect 1975 2143 2001 2169
rect 2311 2143 2337 2169
rect 2647 2143 2673 2169
rect 2703 2143 2729 2169
rect 2983 2143 3009 2169
rect 3319 2143 3345 2169
rect 3991 2143 4017 2169
rect 4271 2143 4297 2169
rect 4327 2143 4353 2169
rect 5279 2143 5305 2169
rect 5615 2143 5641 2169
rect 5951 2143 5977 2169
rect 4887 2087 4913 2113
rect 2031 2031 2057 2057
rect 1314 1947 1340 1973
rect 1366 1947 1392 1973
rect 1418 1947 1444 1973
rect 2728 1947 2754 1973
rect 2780 1947 2806 1973
rect 2832 1947 2858 1973
rect 4142 1947 4168 1973
rect 4194 1947 4220 1973
rect 4246 1947 4272 1973
rect 5556 1947 5582 1973
rect 5608 1947 5634 1973
rect 5660 1947 5686 1973
rect 1751 1863 1777 1889
rect 2031 1863 2057 1889
rect 3879 1863 3905 1889
rect 5223 1863 5249 1889
rect 1079 1807 1105 1833
rect 4831 1807 4857 1833
rect 1023 1751 1049 1777
rect 1359 1751 1385 1777
rect 2423 1751 2449 1777
rect 3151 1751 3177 1777
rect 3543 1751 3569 1777
rect 3823 1751 3849 1777
rect 4159 1751 4185 1777
rect 4215 1751 4241 1777
rect 4887 1751 4913 1777
rect 5167 1751 5193 1777
rect 5503 1751 5529 1777
rect 5895 1751 5921 1777
rect 1415 1695 1441 1721
rect 1695 1695 1721 1721
rect 2087 1695 2113 1721
rect 2367 1695 2393 1721
rect 3207 1695 3233 1721
rect 3487 1695 3513 1721
rect 5559 1695 5585 1721
rect 5839 1695 5865 1721
rect 2021 1555 2047 1581
rect 2073 1555 2099 1581
rect 2125 1555 2151 1581
rect 3435 1555 3461 1581
rect 3487 1555 3513 1581
rect 3539 1555 3565 1581
rect 4849 1555 4875 1581
rect 4901 1555 4927 1581
rect 4953 1555 4979 1581
rect 6263 1555 6289 1581
rect 6315 1555 6341 1581
rect 6367 1555 6393 1581
<< metal2 >>
rect 2020 6286 2152 6291
rect 2048 6258 2072 6286
rect 2100 6258 2124 6286
rect 2020 6253 2152 6258
rect 3434 6286 3566 6291
rect 3462 6258 3486 6286
rect 3514 6258 3538 6286
rect 3434 6253 3566 6258
rect 4848 6286 4980 6291
rect 4876 6258 4900 6286
rect 4928 6258 4952 6286
rect 4848 6253 4980 6258
rect 6262 6286 6394 6291
rect 6290 6258 6314 6286
rect 6342 6258 6366 6286
rect 6262 6253 6394 6258
rect 1806 6202 1834 6207
rect 1806 6201 2002 6202
rect 1806 6175 1807 6201
rect 1833 6175 2002 6201
rect 1806 6174 2002 6175
rect 1806 6169 1834 6174
rect 1134 6090 1162 6095
rect 1134 6043 1162 6062
rect 1414 6090 1442 6095
rect 1694 6090 1722 6095
rect 1414 6089 1554 6090
rect 1414 6063 1415 6089
rect 1441 6063 1554 6089
rect 1414 6062 1554 6063
rect 1414 6057 1442 6062
rect 1078 5977 1106 5983
rect 1078 5951 1079 5977
rect 1105 5951 1106 5977
rect 1078 5697 1106 5951
rect 1470 5978 1498 5997
rect 1470 5945 1498 5950
rect 1526 5922 1554 6062
rect 1313 5894 1445 5899
rect 1341 5866 1365 5894
rect 1393 5866 1417 5894
rect 1526 5889 1554 5894
rect 1313 5861 1445 5866
rect 1078 5671 1079 5697
rect 1105 5671 1106 5697
rect 1078 5665 1106 5671
rect 1470 5641 1498 5647
rect 1470 5615 1471 5641
rect 1497 5615 1498 5641
rect 1134 5586 1162 5591
rect 1414 5586 1442 5591
rect 1022 5585 1162 5586
rect 1022 5559 1135 5585
rect 1161 5559 1162 5585
rect 1022 5558 1162 5559
rect 1022 4578 1050 5558
rect 1134 5553 1162 5558
rect 1190 5585 1442 5586
rect 1190 5559 1415 5585
rect 1441 5559 1442 5585
rect 1190 5558 1442 5559
rect 1190 5418 1218 5558
rect 1414 5553 1442 5558
rect 1470 5418 1498 5615
rect 1694 5586 1722 6062
rect 1750 6090 1778 6095
rect 1750 6089 1890 6090
rect 1750 6063 1751 6089
rect 1777 6063 1890 6089
rect 1750 6062 1890 6063
rect 1750 6057 1778 6062
rect 1750 5978 1778 5983
rect 1750 5698 1778 5950
rect 1862 5810 1890 6062
rect 1974 5978 2002 6174
rect 2926 6146 2954 6151
rect 2926 6099 2954 6118
rect 3374 6146 3402 6151
rect 2086 6090 2114 6095
rect 2422 6090 2450 6095
rect 2086 6089 2450 6090
rect 2086 6063 2087 6089
rect 2113 6063 2423 6089
rect 2449 6063 2450 6089
rect 2086 6062 2450 6063
rect 2086 6057 2114 6062
rect 2422 6057 2450 6062
rect 2478 6090 2506 6095
rect 2478 6043 2506 6062
rect 2870 6090 2898 6095
rect 2142 5978 2170 5983
rect 2870 5978 2898 6062
rect 3262 6090 3290 6095
rect 3262 6043 3290 6062
rect 2982 5978 3010 5983
rect 1974 5950 2114 5978
rect 1862 5777 1890 5782
rect 2030 5866 2058 5871
rect 1806 5698 1834 5703
rect 1750 5697 1834 5698
rect 1750 5671 1807 5697
rect 1833 5671 1834 5697
rect 1750 5670 1834 5671
rect 1806 5665 1834 5670
rect 1750 5586 1778 5591
rect 1694 5585 1778 5586
rect 1694 5559 1751 5585
rect 1777 5559 1778 5585
rect 1694 5558 1778 5559
rect 2030 5586 2058 5838
rect 2086 5698 2114 5950
rect 2142 5977 2506 5978
rect 2142 5951 2143 5977
rect 2169 5951 2506 5977
rect 2142 5950 2506 5951
rect 2870 5950 2954 5978
rect 2142 5945 2170 5950
rect 2422 5810 2450 5815
rect 2422 5763 2450 5782
rect 2142 5698 2170 5703
rect 2086 5697 2170 5698
rect 2086 5671 2143 5697
rect 2169 5671 2170 5697
rect 2086 5670 2170 5671
rect 2142 5665 2170 5670
rect 2478 5697 2506 5950
rect 2727 5894 2859 5899
rect 2755 5866 2779 5894
rect 2807 5866 2831 5894
rect 2727 5861 2859 5866
rect 2926 5866 2954 5950
rect 2982 5977 3122 5978
rect 2982 5951 2983 5977
rect 3009 5951 3122 5977
rect 2982 5950 3122 5951
rect 2982 5945 3010 5950
rect 2926 5838 3066 5866
rect 3038 5809 3066 5838
rect 3038 5783 3039 5809
rect 3065 5783 3066 5809
rect 3038 5777 3066 5783
rect 2478 5671 2479 5697
rect 2505 5671 2506 5697
rect 2478 5665 2506 5671
rect 3094 5697 3122 5950
rect 3094 5671 3095 5697
rect 3121 5671 3122 5697
rect 3094 5665 3122 5671
rect 3318 5977 3346 5983
rect 3318 5951 3319 5977
rect 3345 5951 3346 5977
rect 3318 5698 3346 5951
rect 3374 5809 3402 6118
rect 3654 6146 3682 6151
rect 3654 6099 3682 6118
rect 4270 6146 4298 6151
rect 4270 6099 4298 6118
rect 3598 6090 3626 6095
rect 3598 6043 3626 6062
rect 3934 6089 3962 6095
rect 3934 6063 3935 6089
rect 3961 6063 3962 6089
rect 3374 5783 3375 5809
rect 3401 5783 3402 5809
rect 3374 5777 3402 5783
rect 3934 5809 3962 6063
rect 3990 6090 4018 6095
rect 3990 6043 4018 6062
rect 4326 6090 4354 6095
rect 4326 6043 4354 6062
rect 4141 5894 4273 5899
rect 4169 5866 4193 5894
rect 4221 5866 4245 5894
rect 4141 5861 4273 5866
rect 5555 5894 5687 5899
rect 5583 5866 5607 5894
rect 5635 5866 5659 5894
rect 5555 5861 5687 5866
rect 3934 5783 3935 5809
rect 3961 5783 3962 5809
rect 3934 5777 3962 5783
rect 3430 5698 3458 5703
rect 3318 5697 3458 5698
rect 3318 5671 3431 5697
rect 3457 5671 3458 5697
rect 3318 5670 3458 5671
rect 3430 5665 3458 5670
rect 3990 5642 4018 5647
rect 3990 5595 4018 5614
rect 4270 5642 4298 5647
rect 4270 5595 4298 5614
rect 4326 5641 4354 5647
rect 4326 5615 4327 5641
rect 4353 5615 4354 5641
rect 2086 5586 2114 5591
rect 2030 5585 2114 5586
rect 2030 5559 2087 5585
rect 2113 5559 2114 5585
rect 2030 5558 2114 5559
rect 1750 5553 1778 5558
rect 2086 5553 2114 5558
rect 2020 5502 2152 5507
rect 2048 5474 2072 5502
rect 2100 5474 2124 5502
rect 2020 5469 2152 5474
rect 3434 5502 3566 5507
rect 3462 5474 3486 5502
rect 3514 5474 3538 5502
rect 3434 5469 3566 5474
rect 1078 5390 1218 5418
rect 1246 5390 1498 5418
rect 3878 5418 3906 5423
rect 1078 4913 1106 5390
rect 1134 5305 1162 5311
rect 1134 5279 1135 5305
rect 1161 5279 1162 5305
rect 1134 5026 1162 5279
rect 1134 4993 1162 4998
rect 1190 5193 1218 5199
rect 1190 5167 1191 5193
rect 1217 5167 1218 5193
rect 1078 4887 1079 4913
rect 1105 4887 1106 4913
rect 1078 4881 1106 4887
rect 1190 4914 1218 5167
rect 1190 4881 1218 4886
rect 1134 4802 1162 4807
rect 1022 4545 1050 4550
rect 1078 4801 1162 4802
rect 1078 4775 1135 4801
rect 1161 4775 1162 4801
rect 1078 4774 1162 4775
rect 1078 4214 1106 4774
rect 1134 4769 1162 4774
rect 1190 4634 1218 4639
rect 1246 4634 1274 5390
rect 3878 5371 3906 5390
rect 4326 5418 4354 5615
rect 4848 5502 4980 5507
rect 4876 5474 4900 5502
rect 4928 5474 4952 5502
rect 4848 5469 4980 5474
rect 6262 5502 6394 5507
rect 6290 5474 6314 5502
rect 6342 5474 6366 5502
rect 6262 5469 6394 5474
rect 4326 5385 4354 5390
rect 2478 5362 2506 5367
rect 2478 5315 2506 5334
rect 3430 5362 3458 5367
rect 1470 5305 1498 5311
rect 1470 5279 1471 5305
rect 1497 5279 1498 5305
rect 1470 5194 1498 5279
rect 1526 5306 1554 5311
rect 1526 5259 1554 5278
rect 1806 5306 1834 5311
rect 1806 5259 1834 5278
rect 1862 5306 1890 5311
rect 2142 5306 2170 5311
rect 1862 5305 2170 5306
rect 1862 5279 1863 5305
rect 1889 5279 2143 5305
rect 2169 5279 2170 5305
rect 1862 5278 2170 5279
rect 1862 5273 1890 5278
rect 2142 5273 2170 5278
rect 2814 5305 2842 5311
rect 2814 5279 2815 5305
rect 2841 5279 2842 5305
rect 2198 5194 2226 5199
rect 2534 5194 2562 5199
rect 2814 5194 2842 5279
rect 2870 5306 2898 5311
rect 3150 5306 3178 5311
rect 2870 5305 3178 5306
rect 2870 5279 2871 5305
rect 2897 5279 3151 5305
rect 3177 5279 3178 5305
rect 2870 5278 3178 5279
rect 2870 5273 2898 5278
rect 3150 5273 3178 5278
rect 3206 5306 3234 5311
rect 3206 5259 3234 5278
rect 1470 5166 1666 5194
rect 1313 5110 1445 5115
rect 1341 5082 1365 5110
rect 1393 5082 1417 5110
rect 1313 5077 1445 5082
rect 1414 5026 1442 5031
rect 1638 5026 1666 5166
rect 2198 5193 2506 5194
rect 2198 5167 2199 5193
rect 2225 5167 2506 5193
rect 2198 5166 2506 5167
rect 2198 5161 2226 5166
rect 1750 5026 1778 5031
rect 1638 5025 1778 5026
rect 1638 4999 1751 5025
rect 1777 4999 1778 5025
rect 1638 4998 1778 4999
rect 1414 4979 1442 4998
rect 1750 4993 1778 4998
rect 1806 4914 1834 4919
rect 1806 4867 1834 4886
rect 2086 4914 2114 4919
rect 2422 4914 2450 4919
rect 2086 4913 2450 4914
rect 2086 4887 2087 4913
rect 2113 4887 2423 4913
rect 2449 4887 2450 4913
rect 2086 4886 2450 4887
rect 2086 4881 2114 4886
rect 2422 4881 2450 4886
rect 2478 4913 2506 5166
rect 2534 5193 2674 5194
rect 2534 5167 2535 5193
rect 2561 5167 2674 5193
rect 2534 5166 2674 5167
rect 2814 5166 3122 5194
rect 2534 5161 2562 5166
rect 2646 4970 2674 5166
rect 2727 5110 2859 5115
rect 2755 5082 2779 5110
rect 2807 5082 2831 5110
rect 2727 5077 2859 5082
rect 3094 5025 3122 5166
rect 3094 4999 3095 5025
rect 3121 4999 3122 5025
rect 3094 4993 3122 4999
rect 3430 5025 3458 5334
rect 3542 5362 3570 5367
rect 3542 5315 3570 5334
rect 4214 5362 4242 5367
rect 4214 5315 4242 5334
rect 3486 5306 3514 5311
rect 3486 5259 3514 5278
rect 3822 5306 3850 5311
rect 4158 5306 4186 5311
rect 3822 5305 4186 5306
rect 3822 5279 3823 5305
rect 3849 5279 4159 5305
rect 4185 5279 4186 5305
rect 3822 5278 4186 5279
rect 3822 5273 3850 5278
rect 4158 5273 4186 5278
rect 4141 5110 4273 5115
rect 4169 5082 4193 5110
rect 4221 5082 4245 5110
rect 4141 5077 4273 5082
rect 5555 5110 5687 5115
rect 5583 5082 5607 5110
rect 5635 5082 5659 5110
rect 5555 5077 5687 5082
rect 3430 4999 3431 5025
rect 3457 4999 3458 5025
rect 3430 4993 3458 4999
rect 2646 4942 3066 4970
rect 2478 4887 2479 4913
rect 2505 4887 2506 4913
rect 2478 4881 2506 4887
rect 3038 4914 3066 4942
rect 3150 4914 3178 4919
rect 3038 4913 3178 4914
rect 3038 4887 3151 4913
rect 3177 4887 3178 4913
rect 3038 4886 3178 4887
rect 3150 4881 3178 4886
rect 1470 4858 1498 4863
rect 3206 4858 3234 4863
rect 1470 4857 1610 4858
rect 1470 4831 1471 4857
rect 1497 4831 1610 4857
rect 1470 4830 1610 4831
rect 1470 4825 1498 4830
rect 1190 4633 1274 4634
rect 1190 4607 1191 4633
rect 1217 4607 1274 4633
rect 1190 4606 1274 4607
rect 1190 4601 1218 4606
rect 1526 4578 1554 4583
rect 1526 4531 1554 4550
rect 1134 4522 1162 4527
rect 1470 4522 1498 4527
rect 1134 4521 1498 4522
rect 1134 4495 1135 4521
rect 1161 4495 1471 4521
rect 1497 4495 1498 4521
rect 1134 4494 1498 4495
rect 1134 4489 1162 4494
rect 1470 4489 1498 4494
rect 1313 4326 1445 4331
rect 1341 4298 1365 4326
rect 1393 4298 1417 4326
rect 1313 4293 1445 4298
rect 1526 4242 1554 4247
rect 1582 4242 1610 4830
rect 2142 4802 2170 4807
rect 3150 4802 3178 4807
rect 2142 4801 2226 4802
rect 2142 4775 2143 4801
rect 2169 4775 2226 4801
rect 2142 4774 2226 4775
rect 2142 4769 2170 4774
rect 2020 4718 2152 4723
rect 2048 4690 2072 4718
rect 2100 4690 2124 4718
rect 2020 4685 2152 4690
rect 2142 4578 2170 4583
rect 2198 4578 2226 4774
rect 2870 4634 2898 4639
rect 2870 4587 2898 4606
rect 2142 4577 2226 4578
rect 2142 4551 2143 4577
rect 2169 4551 2226 4577
rect 2142 4550 2226 4551
rect 3150 4577 3178 4774
rect 3206 4633 3234 4830
rect 3486 4858 3514 4863
rect 3486 4811 3514 4830
rect 3822 4857 3850 4863
rect 3822 4831 3823 4857
rect 3849 4831 3850 4857
rect 3766 4802 3794 4807
rect 3766 4755 3794 4774
rect 3434 4718 3566 4723
rect 3462 4690 3486 4718
rect 3514 4690 3538 4718
rect 3822 4690 3850 4831
rect 3434 4685 3566 4690
rect 3598 4662 3850 4690
rect 4848 4718 4980 4723
rect 4876 4690 4900 4718
rect 4928 4690 4952 4718
rect 4848 4685 4980 4690
rect 6262 4718 6394 4723
rect 6290 4690 6314 4718
rect 6342 4690 6366 4718
rect 6262 4685 6394 4690
rect 3206 4607 3207 4633
rect 3233 4607 3234 4633
rect 3206 4601 3234 4607
rect 3486 4634 3514 4639
rect 3150 4551 3151 4577
rect 3177 4551 3178 4577
rect 2142 4545 2170 4550
rect 3150 4545 3178 4551
rect 3486 4577 3514 4606
rect 3542 4634 3570 4639
rect 3598 4634 3626 4662
rect 3542 4633 3626 4634
rect 3542 4607 3543 4633
rect 3569 4607 3626 4633
rect 3542 4606 3626 4607
rect 3542 4601 3570 4606
rect 3486 4551 3487 4577
rect 3513 4551 3514 4577
rect 3486 4545 3514 4551
rect 1806 4522 1834 4527
rect 2478 4522 2506 4527
rect 1806 4521 2114 4522
rect 1806 4495 1807 4521
rect 1833 4495 2114 4521
rect 1806 4494 2114 4495
rect 1806 4489 1834 4494
rect 1526 4241 1610 4242
rect 1526 4215 1527 4241
rect 1553 4215 1610 4241
rect 1526 4214 1610 4215
rect 1862 4409 1890 4415
rect 1862 4383 1863 4409
rect 1889 4383 1890 4409
rect 1078 4186 1498 4214
rect 1526 4209 1554 4214
rect 1470 4130 1498 4186
rect 1582 4130 1610 4135
rect 1470 4129 1610 4130
rect 1470 4103 1583 4129
rect 1609 4103 1610 4129
rect 1470 4102 1610 4103
rect 1862 4130 1890 4383
rect 2030 4242 2058 4247
rect 2086 4242 2114 4494
rect 2478 4475 2506 4494
rect 2814 4522 2842 4527
rect 3430 4522 3458 4527
rect 2814 4521 3122 4522
rect 2814 4495 2815 4521
rect 2841 4495 3122 4521
rect 2814 4494 3122 4495
rect 2814 4489 2842 4494
rect 2198 4410 2226 4415
rect 2422 4410 2450 4415
rect 2198 4409 2394 4410
rect 2198 4383 2199 4409
rect 2225 4383 2394 4409
rect 2198 4382 2394 4383
rect 2198 4377 2226 4382
rect 2310 4242 2338 4247
rect 2086 4241 2338 4242
rect 2086 4215 2311 4241
rect 2337 4215 2338 4241
rect 2086 4214 2338 4215
rect 2030 4185 2058 4214
rect 2310 4209 2338 4214
rect 2030 4159 2031 4185
rect 2057 4159 2058 4185
rect 2030 4153 2058 4159
rect 1974 4130 2002 4135
rect 1862 4129 2002 4130
rect 1862 4103 1975 4129
rect 2001 4103 2002 4129
rect 1862 4102 2002 4103
rect 1582 4097 1610 4102
rect 1974 4097 2002 4102
rect 2366 4129 2394 4382
rect 2366 4103 2367 4129
rect 2393 4103 2394 4129
rect 2366 4097 2394 4103
rect 1078 4074 1106 4079
rect 1078 4027 1106 4046
rect 910 4018 938 4023
rect 910 2450 938 3990
rect 2020 3934 2152 3939
rect 2048 3906 2072 3934
rect 2100 3906 2124 3934
rect 2020 3901 2152 3906
rect 1358 3850 1386 3855
rect 1358 3849 1610 3850
rect 1358 3823 1359 3849
rect 1385 3823 1610 3849
rect 1358 3822 1610 3823
rect 1358 3817 1386 3822
rect 966 3738 994 3743
rect 1302 3738 1330 3743
rect 966 3737 1274 3738
rect 966 3711 967 3737
rect 993 3711 1274 3737
rect 966 3710 1274 3711
rect 966 3705 994 3710
rect 1022 3626 1050 3631
rect 1190 3626 1218 3631
rect 1022 3625 1162 3626
rect 1022 3599 1023 3625
rect 1049 3599 1162 3625
rect 1022 3598 1162 3599
rect 1022 3593 1050 3598
rect 1134 3345 1162 3598
rect 1134 3319 1135 3345
rect 1161 3319 1162 3345
rect 1134 3313 1162 3319
rect 1078 3233 1106 3239
rect 1078 3207 1079 3233
rect 1105 3207 1106 3233
rect 1022 3010 1050 3015
rect 1078 3010 1106 3207
rect 1022 3009 1106 3010
rect 1022 2983 1023 3009
rect 1049 2983 1106 3009
rect 1022 2982 1106 2983
rect 1022 2977 1050 2982
rect 966 2841 994 2847
rect 966 2815 967 2841
rect 993 2815 994 2841
rect 966 2562 994 2815
rect 1190 2674 1218 3598
rect 1246 3458 1274 3710
rect 1302 3737 1554 3738
rect 1302 3711 1303 3737
rect 1329 3711 1554 3737
rect 1302 3710 1554 3711
rect 1302 3705 1330 3710
rect 1313 3542 1445 3547
rect 1341 3514 1365 3542
rect 1393 3514 1417 3542
rect 1313 3509 1445 3514
rect 1414 3458 1442 3463
rect 1246 3457 1442 3458
rect 1246 3431 1415 3457
rect 1441 3431 1442 3457
rect 1246 3430 1442 3431
rect 1414 3425 1442 3430
rect 1470 3290 1498 3295
rect 1470 3243 1498 3262
rect 1526 3066 1554 3710
rect 1526 3033 1554 3038
rect 1302 2954 1330 2959
rect 1302 2953 1554 2954
rect 1302 2927 1303 2953
rect 1329 2927 1554 2953
rect 1302 2926 1554 2927
rect 1302 2921 1330 2926
rect 1358 2842 1386 2861
rect 1358 2809 1386 2814
rect 1313 2758 1445 2763
rect 1341 2730 1365 2758
rect 1393 2730 1417 2758
rect 1313 2725 1445 2730
rect 1190 2646 1498 2674
rect 1022 2562 1050 2567
rect 966 2561 1050 2562
rect 966 2535 1023 2561
rect 1049 2535 1050 2561
rect 966 2534 1050 2535
rect 1022 2529 1050 2534
rect 1190 2506 1218 2511
rect 966 2450 994 2455
rect 910 2449 994 2450
rect 910 2423 967 2449
rect 993 2423 994 2449
rect 910 2422 994 2423
rect 966 2417 994 2422
rect 1190 2281 1218 2478
rect 1190 2255 1191 2281
rect 1217 2255 1218 2281
rect 1190 2249 1218 2255
rect 1022 2226 1050 2231
rect 1022 1777 1050 2198
rect 1470 2225 1498 2646
rect 1526 2673 1554 2926
rect 1526 2647 1527 2673
rect 1553 2647 1554 2673
rect 1526 2641 1554 2647
rect 1582 2618 1610 3822
rect 2366 3794 2394 3799
rect 2422 3794 2450 4382
rect 2534 4409 2562 4415
rect 2534 4383 2535 4409
rect 2561 4383 2562 4409
rect 2534 4214 2562 4383
rect 2727 4326 2859 4331
rect 2755 4298 2779 4326
rect 2807 4298 2831 4326
rect 2727 4293 2859 4298
rect 3094 4241 3122 4494
rect 3094 4215 3095 4241
rect 3121 4215 3122 4241
rect 2534 4186 3066 4214
rect 3094 4209 3122 4215
rect 3038 4130 3066 4186
rect 3430 4185 3458 4494
rect 3878 4521 3906 4527
rect 3878 4495 3879 4521
rect 3905 4495 3906 4521
rect 3822 4410 3850 4415
rect 3822 4363 3850 4382
rect 3878 4242 3906 4495
rect 4141 4326 4273 4331
rect 4169 4298 4193 4326
rect 4221 4298 4245 4326
rect 4141 4293 4273 4298
rect 5555 4326 5687 4331
rect 5583 4298 5607 4326
rect 5635 4298 5659 4326
rect 5555 4293 5687 4298
rect 3878 4209 3906 4214
rect 3430 4159 3431 4185
rect 3457 4159 3458 4185
rect 3430 4153 3458 4159
rect 3150 4130 3178 4135
rect 3038 4129 3178 4130
rect 3038 4103 3151 4129
rect 3177 4103 3178 4129
rect 3038 4102 3178 4103
rect 3150 4097 3178 4102
rect 3486 4073 3514 4079
rect 3486 4047 3487 4073
rect 3513 4047 3514 4073
rect 3038 4018 3066 4023
rect 2702 3850 2730 3855
rect 2702 3803 2730 3822
rect 3038 3849 3066 3990
rect 3486 4018 3514 4047
rect 3766 4074 3794 4079
rect 3766 4027 3794 4046
rect 3822 4074 3850 4079
rect 4102 4074 4130 4079
rect 3822 4073 4130 4074
rect 3822 4047 3823 4073
rect 3849 4047 4103 4073
rect 4129 4047 4130 4073
rect 3822 4046 4130 4047
rect 3822 4041 3850 4046
rect 4102 4041 4130 4046
rect 3486 3985 3514 3990
rect 4158 4017 4186 4023
rect 4158 3991 4159 4017
rect 4185 3991 4186 4017
rect 3434 3934 3566 3939
rect 3462 3906 3486 3934
rect 3514 3906 3538 3934
rect 3434 3901 3566 3906
rect 3038 3823 3039 3849
rect 3065 3823 3066 3849
rect 3038 3817 3066 3823
rect 3374 3850 3402 3855
rect 2366 3793 2450 3794
rect 2366 3767 2367 3793
rect 2393 3767 2450 3793
rect 2366 3766 2450 3767
rect 3374 3793 3402 3822
rect 3374 3767 3375 3793
rect 3401 3767 3402 3793
rect 2366 3761 2394 3766
rect 3374 3761 3402 3767
rect 1638 3737 1666 3743
rect 1638 3711 1639 3737
rect 1665 3711 1666 3737
rect 1638 3346 1666 3711
rect 1974 3738 2002 3743
rect 2310 3738 2338 3743
rect 1974 3737 2338 3738
rect 1974 3711 1975 3737
rect 2001 3711 2311 3737
rect 2337 3711 2338 3737
rect 1974 3710 2338 3711
rect 1974 3705 2002 3710
rect 2310 3705 2338 3710
rect 2646 3738 2674 3743
rect 2982 3738 3010 3743
rect 3318 3738 3346 3743
rect 3710 3738 3738 3743
rect 2646 3737 2954 3738
rect 2646 3711 2647 3737
rect 2673 3711 2954 3737
rect 2646 3710 2954 3711
rect 2646 3705 2674 3710
rect 1694 3626 1722 3631
rect 2030 3626 2058 3631
rect 1694 3625 1834 3626
rect 1694 3599 1695 3625
rect 1721 3599 1834 3625
rect 1694 3598 1834 3599
rect 1694 3593 1722 3598
rect 1638 3313 1666 3318
rect 1806 3345 1834 3598
rect 2030 3625 2282 3626
rect 2030 3599 2031 3625
rect 2057 3599 2282 3625
rect 2030 3598 2282 3599
rect 2030 3593 2058 3598
rect 1806 3319 1807 3345
rect 1833 3319 1834 3345
rect 1806 3313 1834 3319
rect 2198 3346 2226 3351
rect 2198 3299 2226 3318
rect 2254 3345 2282 3598
rect 2727 3542 2859 3547
rect 2755 3514 2779 3542
rect 2807 3514 2831 3542
rect 2727 3509 2859 3514
rect 2926 3458 2954 3710
rect 2982 3737 3346 3738
rect 2982 3711 2983 3737
rect 3009 3711 3319 3737
rect 3345 3711 3346 3737
rect 2982 3710 3346 3711
rect 2982 3705 3010 3710
rect 3318 3705 3346 3710
rect 3430 3737 3738 3738
rect 3430 3711 3711 3737
rect 3737 3711 3738 3737
rect 3430 3710 3738 3711
rect 2982 3458 3010 3463
rect 2926 3457 3010 3458
rect 2926 3431 2983 3457
rect 3009 3431 3010 3457
rect 2926 3430 3010 3431
rect 2982 3425 3010 3430
rect 3374 3458 3402 3463
rect 3430 3458 3458 3710
rect 3710 3705 3738 3710
rect 4046 3738 4074 3743
rect 4046 3691 4074 3710
rect 3374 3457 3458 3458
rect 3374 3431 3375 3457
rect 3401 3431 3458 3457
rect 3374 3430 3458 3431
rect 3654 3625 3682 3631
rect 3654 3599 3655 3625
rect 3681 3599 3682 3625
rect 3374 3425 3402 3430
rect 2254 3319 2255 3345
rect 2281 3319 2282 3345
rect 2254 3313 2282 3319
rect 3038 3402 3066 3407
rect 3038 3345 3066 3374
rect 3654 3402 3682 3599
rect 3990 3626 4018 3631
rect 4158 3626 4186 3991
rect 4848 3934 4980 3939
rect 4876 3906 4900 3934
rect 4928 3906 4952 3934
rect 4848 3901 4980 3906
rect 6262 3934 6394 3939
rect 6290 3906 6314 3934
rect 6342 3906 6366 3934
rect 6262 3901 6394 3906
rect 4326 3738 4354 3743
rect 4326 3691 4354 3710
rect 4382 3737 4410 3743
rect 4382 3711 4383 3737
rect 4409 3711 4410 3737
rect 3990 3579 4018 3598
rect 4046 3598 4186 3626
rect 4046 3402 4074 3598
rect 4141 3542 4273 3547
rect 4169 3514 4193 3542
rect 4221 3514 4245 3542
rect 4141 3509 4273 3514
rect 4326 3458 4354 3463
rect 4382 3458 4410 3711
rect 5555 3542 5687 3547
rect 5583 3514 5607 3542
rect 5635 3514 5659 3542
rect 5555 3509 5687 3514
rect 4326 3457 4410 3458
rect 4326 3431 4327 3457
rect 4353 3431 4410 3457
rect 4326 3430 4410 3431
rect 4326 3425 4354 3430
rect 4046 3374 4130 3402
rect 3654 3369 3682 3374
rect 3038 3319 3039 3345
rect 3065 3319 3066 3345
rect 3038 3313 3066 3319
rect 4102 3346 4130 3374
rect 4102 3313 4130 3318
rect 4382 3346 4410 3351
rect 4382 3299 4410 3318
rect 1750 3290 1778 3295
rect 1750 3243 1778 3262
rect 2422 3290 2450 3295
rect 3318 3290 3346 3295
rect 2020 3150 2152 3155
rect 2048 3122 2072 3150
rect 2100 3122 2124 3150
rect 2020 3117 2152 3122
rect 2310 3066 2338 3071
rect 2310 3019 2338 3038
rect 1638 2953 1666 2959
rect 1638 2927 1639 2953
rect 1665 2927 1666 2953
rect 1638 2674 1666 2927
rect 1694 2954 1722 2959
rect 1974 2954 2002 2959
rect 1694 2953 2002 2954
rect 1694 2927 1695 2953
rect 1721 2927 1975 2953
rect 2001 2927 2002 2953
rect 1694 2926 2002 2927
rect 1694 2921 1722 2926
rect 1974 2921 2002 2926
rect 2030 2954 2058 2959
rect 2366 2954 2394 2959
rect 2030 2953 2394 2954
rect 2030 2927 2031 2953
rect 2057 2927 2367 2953
rect 2393 2927 2394 2953
rect 2030 2926 2394 2927
rect 2030 2921 2058 2926
rect 2366 2921 2394 2926
rect 1918 2842 1946 2847
rect 1638 2641 1666 2646
rect 1862 2674 1890 2679
rect 1862 2627 1890 2646
rect 1582 2585 1610 2590
rect 1918 2561 1946 2814
rect 2422 2673 2450 3262
rect 3150 3289 3346 3290
rect 3150 3263 3319 3289
rect 3345 3263 3346 3289
rect 3150 3262 3346 3263
rect 3094 3234 3122 3239
rect 2758 3010 2786 3015
rect 2758 2963 2786 2982
rect 3094 3009 3122 3206
rect 3150 3065 3178 3262
rect 3318 3257 3346 3262
rect 3710 3289 3738 3295
rect 3710 3263 3711 3289
rect 3737 3263 3738 3289
rect 3654 3234 3682 3239
rect 3654 3187 3682 3206
rect 3434 3150 3566 3155
rect 3462 3122 3486 3150
rect 3514 3122 3538 3150
rect 3434 3117 3566 3122
rect 3150 3039 3151 3065
rect 3177 3039 3178 3065
rect 3150 3033 3178 3039
rect 3486 3066 3514 3071
rect 3710 3066 3738 3263
rect 4046 3290 4074 3295
rect 4046 3243 4074 3262
rect 4662 3290 4690 3295
rect 4662 3243 4690 3262
rect 6006 3290 6034 3295
rect 3486 3065 3738 3066
rect 3486 3039 3487 3065
rect 3513 3039 3738 3065
rect 3486 3038 3738 3039
rect 3990 3233 4018 3239
rect 3990 3207 3991 3233
rect 4017 3207 4018 3233
rect 3486 3033 3514 3038
rect 3094 2983 3095 3009
rect 3121 2983 3122 3009
rect 3094 2977 3122 2983
rect 3766 3010 3794 3015
rect 3766 2963 3794 2982
rect 2814 2954 2842 2959
rect 2814 2907 2842 2926
rect 3430 2954 3458 2959
rect 3430 2907 3458 2926
rect 3822 2953 3850 2959
rect 3822 2927 3823 2953
rect 3849 2927 3850 2953
rect 2727 2758 2859 2763
rect 2755 2730 2779 2758
rect 2807 2730 2831 2758
rect 2727 2725 2859 2730
rect 2422 2647 2423 2673
rect 2449 2647 2450 2673
rect 2422 2641 2450 2647
rect 3318 2674 3346 2679
rect 1918 2535 1919 2561
rect 1945 2535 1946 2561
rect 1918 2529 1946 2535
rect 2366 2618 2394 2623
rect 2366 2561 2394 2590
rect 2366 2535 2367 2561
rect 2393 2535 2394 2561
rect 2366 2529 2394 2535
rect 2870 2562 2898 2567
rect 3206 2562 3234 2567
rect 2870 2561 3234 2562
rect 2870 2535 2871 2561
rect 2897 2535 3207 2561
rect 3233 2535 3234 2561
rect 2870 2534 3234 2535
rect 2870 2529 2898 2534
rect 3206 2529 3234 2534
rect 3262 2562 3290 2567
rect 3262 2515 3290 2534
rect 1582 2505 1610 2511
rect 1582 2479 1583 2505
rect 1609 2479 1610 2505
rect 1526 2282 1554 2287
rect 1582 2282 1610 2479
rect 2926 2450 2954 2455
rect 3318 2450 3346 2646
rect 3822 2674 3850 2927
rect 3822 2641 3850 2646
rect 3598 2618 3626 2623
rect 3542 2562 3570 2567
rect 3542 2515 3570 2534
rect 3598 2561 3626 2590
rect 3598 2535 3599 2561
rect 3625 2535 3626 2561
rect 3598 2529 3626 2535
rect 3934 2562 3962 2567
rect 3934 2515 3962 2534
rect 3878 2505 3906 2511
rect 3878 2479 3879 2505
rect 3905 2479 3906 2505
rect 2926 2403 2954 2422
rect 3038 2422 3346 2450
rect 3374 2450 3402 2455
rect 2020 2366 2152 2371
rect 2048 2338 2072 2366
rect 2100 2338 2124 2366
rect 2020 2333 2152 2338
rect 1526 2281 1610 2282
rect 1526 2255 1527 2281
rect 1553 2255 1610 2281
rect 1526 2254 1610 2255
rect 2366 2282 2394 2287
rect 1526 2249 1554 2254
rect 1470 2199 1471 2225
rect 1497 2199 1498 2225
rect 1470 2193 1498 2199
rect 2366 2225 2394 2254
rect 3038 2281 3066 2422
rect 3038 2255 3039 2281
rect 3065 2255 3066 2281
rect 3038 2249 3066 2255
rect 2366 2199 2367 2225
rect 2393 2199 2394 2225
rect 2366 2193 2394 2199
rect 3374 2225 3402 2422
rect 3598 2450 3626 2455
rect 3434 2366 3566 2371
rect 3462 2338 3486 2366
rect 3514 2338 3538 2366
rect 3434 2333 3566 2338
rect 3374 2199 3375 2225
rect 3401 2199 3402 2225
rect 3374 2193 3402 2199
rect 1134 2169 1162 2175
rect 1134 2143 1135 2169
rect 1161 2143 1162 2169
rect 1134 1890 1162 2143
rect 1974 2170 2002 2175
rect 2310 2170 2338 2175
rect 1974 2169 2338 2170
rect 1974 2143 1975 2169
rect 2001 2143 2311 2169
rect 2337 2143 2338 2169
rect 1974 2142 2338 2143
rect 1974 2137 2002 2142
rect 2310 2137 2338 2142
rect 2646 2170 2674 2175
rect 2646 2123 2674 2142
rect 2702 2170 2730 2175
rect 2982 2170 3010 2175
rect 2702 2169 3010 2170
rect 2702 2143 2703 2169
rect 2729 2143 2983 2169
rect 3009 2143 3010 2169
rect 2702 2142 3010 2143
rect 2702 2137 2730 2142
rect 2982 2137 3010 2142
rect 3318 2170 3346 2175
rect 3318 2123 3346 2142
rect 1526 2114 1554 2119
rect 1313 1974 1445 1979
rect 1341 1946 1365 1974
rect 1393 1946 1417 1974
rect 1313 1941 1445 1946
rect 1526 1890 1554 2086
rect 1134 1857 1162 1862
rect 1358 1862 1554 1890
rect 1750 2058 1778 2063
rect 1750 1889 1778 2030
rect 2030 2058 2058 2063
rect 2030 2057 2450 2058
rect 2030 2031 2031 2057
rect 2057 2031 2450 2057
rect 2030 2030 2450 2031
rect 2030 2025 2058 2030
rect 1750 1863 1751 1889
rect 1777 1863 1778 1889
rect 1078 1834 1106 1839
rect 1078 1787 1106 1806
rect 1022 1751 1023 1777
rect 1049 1751 1050 1777
rect 1022 1745 1050 1751
rect 1358 1777 1386 1862
rect 1750 1857 1778 1863
rect 2030 1890 2058 1895
rect 2030 1843 2058 1862
rect 1358 1751 1359 1777
rect 1385 1751 1386 1777
rect 1358 1745 1386 1751
rect 2422 1777 2450 2030
rect 2727 1974 2859 1979
rect 2755 1946 2779 1974
rect 2807 1946 2831 1974
rect 2727 1941 2859 1946
rect 3598 1890 3626 2422
rect 3878 2282 3906 2479
rect 3934 2282 3962 2287
rect 3878 2281 3962 2282
rect 3878 2255 3935 2281
rect 3961 2255 3962 2281
rect 3878 2254 3962 2255
rect 3934 2249 3962 2254
rect 3990 2282 4018 3207
rect 4718 3234 4746 3239
rect 4718 3187 4746 3206
rect 5950 3234 5978 3239
rect 4848 3150 4980 3155
rect 4876 3122 4900 3150
rect 4928 3122 4952 3150
rect 4848 3117 4980 3122
rect 4102 2954 4130 2959
rect 4046 2953 4130 2954
rect 4046 2927 4103 2953
rect 4129 2927 4130 2953
rect 4046 2926 4130 2927
rect 4046 2506 4074 2926
rect 4102 2921 4130 2926
rect 4158 2954 4186 2959
rect 4158 2907 4186 2926
rect 4438 2954 4466 2959
rect 4438 2907 4466 2926
rect 4886 2954 4914 2959
rect 4886 2907 4914 2926
rect 5166 2954 5194 2959
rect 4494 2842 4522 2847
rect 4942 2842 4970 2847
rect 4494 2841 4914 2842
rect 4494 2815 4495 2841
rect 4521 2815 4914 2841
rect 4494 2814 4914 2815
rect 4494 2809 4522 2814
rect 4141 2758 4273 2763
rect 4169 2730 4193 2758
rect 4221 2730 4245 2758
rect 4141 2725 4273 2730
rect 4214 2618 4242 2623
rect 4214 2571 4242 2590
rect 4270 2562 4298 2567
rect 4270 2515 4298 2534
rect 4886 2561 4914 2814
rect 4942 2841 5026 2842
rect 4942 2815 4943 2841
rect 4969 2815 5026 2841
rect 4942 2814 5026 2815
rect 4942 2809 4970 2814
rect 4886 2535 4887 2561
rect 4913 2535 4914 2561
rect 4886 2529 4914 2535
rect 4942 2562 4970 2567
rect 4942 2515 4970 2534
rect 4046 2473 4074 2478
rect 4606 2505 4634 2511
rect 4606 2479 4607 2505
rect 4633 2479 4634 2505
rect 3990 2249 4018 2254
rect 4550 2449 4578 2455
rect 4550 2423 4551 2449
rect 4577 2423 4578 2449
rect 4550 2226 4578 2423
rect 4606 2282 4634 2479
rect 4774 2450 4802 2455
rect 4774 2282 4802 2422
rect 4998 2450 5026 2814
rect 5166 2674 5194 2926
rect 5222 2953 5250 2959
rect 5222 2927 5223 2953
rect 5249 2927 5250 2953
rect 5222 2842 5250 2927
rect 5222 2809 5250 2814
rect 5278 2842 5306 2847
rect 5894 2842 5922 2847
rect 5278 2841 5474 2842
rect 5278 2815 5279 2841
rect 5305 2815 5474 2841
rect 5278 2814 5474 2815
rect 5278 2809 5306 2814
rect 5222 2674 5250 2679
rect 5166 2673 5250 2674
rect 5166 2647 5223 2673
rect 5249 2647 5250 2673
rect 5166 2646 5250 2647
rect 5446 2674 5474 2814
rect 5555 2758 5687 2763
rect 5583 2730 5607 2758
rect 5635 2730 5659 2758
rect 5555 2725 5687 2730
rect 5446 2646 5586 2674
rect 5222 2641 5250 2646
rect 5278 2562 5306 2567
rect 5278 2515 5306 2534
rect 5558 2561 5586 2646
rect 5894 2673 5922 2814
rect 5894 2647 5895 2673
rect 5921 2647 5922 2673
rect 5894 2641 5922 2647
rect 5558 2535 5559 2561
rect 5585 2535 5586 2561
rect 5558 2529 5586 2535
rect 5950 2561 5978 3206
rect 5950 2535 5951 2561
rect 5977 2535 5978 2561
rect 5950 2529 5978 2535
rect 4998 2417 5026 2422
rect 5558 2450 5586 2455
rect 4848 2366 4980 2371
rect 4876 2338 4900 2366
rect 4928 2338 4952 2366
rect 4848 2333 4980 2338
rect 5222 2282 5250 2287
rect 4774 2254 4970 2282
rect 4606 2249 4634 2254
rect 4550 2193 4578 2198
rect 4942 2225 4970 2254
rect 5222 2235 5250 2254
rect 4942 2199 4943 2225
rect 4969 2199 4970 2225
rect 4942 2193 4970 2199
rect 5558 2225 5586 2422
rect 5614 2450 5642 2455
rect 5614 2449 5866 2450
rect 5614 2423 5615 2449
rect 5641 2423 5866 2449
rect 5614 2422 5866 2423
rect 5614 2417 5642 2422
rect 5558 2199 5559 2225
rect 5585 2199 5586 2225
rect 5558 2193 5586 2199
rect 3990 2170 4018 2175
rect 3990 2123 4018 2142
rect 4270 2170 4298 2175
rect 4270 2123 4298 2142
rect 4326 2169 4354 2175
rect 4326 2143 4327 2169
rect 4353 2143 4354 2169
rect 4141 1974 4273 1979
rect 4169 1946 4193 1974
rect 4221 1946 4245 1974
rect 4141 1941 4273 1946
rect 3598 1857 3626 1862
rect 3878 1890 3906 1895
rect 3878 1843 3906 1862
rect 4326 1890 4354 2143
rect 5278 2169 5306 2175
rect 5278 2143 5279 2169
rect 5305 2143 5306 2169
rect 4886 2114 4914 2119
rect 4886 2067 4914 2086
rect 4326 1857 4354 1862
rect 4886 2002 4914 2007
rect 2422 1751 2423 1777
rect 2449 1751 2450 1777
rect 2422 1745 2450 1751
rect 3150 1834 3178 1839
rect 3150 1777 3178 1806
rect 4830 1834 4858 1839
rect 4830 1787 4858 1806
rect 3150 1751 3151 1777
rect 3177 1751 3178 1777
rect 3150 1745 3178 1751
rect 3542 1778 3570 1783
rect 3542 1731 3570 1750
rect 3822 1778 3850 1783
rect 4158 1778 4186 1783
rect 3822 1777 4186 1778
rect 3822 1751 3823 1777
rect 3849 1751 4159 1777
rect 4185 1751 4186 1777
rect 3822 1750 4186 1751
rect 3822 1745 3850 1750
rect 4158 1745 4186 1750
rect 4214 1778 4242 1783
rect 4214 1731 4242 1750
rect 4886 1777 4914 1974
rect 5222 1890 5250 1895
rect 5278 1890 5306 2143
rect 5614 2170 5642 2175
rect 5614 2123 5642 2142
rect 5555 1974 5687 1979
rect 5583 1946 5607 1974
rect 5635 1946 5659 1974
rect 5555 1941 5687 1946
rect 5838 1946 5866 2422
rect 5894 2282 5922 2287
rect 6006 2282 6034 3262
rect 6262 3150 6394 3155
rect 6290 3122 6314 3150
rect 6342 3122 6366 3150
rect 6262 3117 6394 3122
rect 6262 2366 6394 2371
rect 6290 2338 6314 2366
rect 6342 2338 6366 2366
rect 6262 2333 6394 2338
rect 5894 2281 6034 2282
rect 5894 2255 5895 2281
rect 5921 2255 6034 2281
rect 5894 2254 6034 2255
rect 5894 2249 5922 2254
rect 5950 2170 5978 2175
rect 5950 2123 5978 2142
rect 5838 1918 5922 1946
rect 5222 1889 5306 1890
rect 5222 1863 5223 1889
rect 5249 1863 5306 1889
rect 5222 1862 5306 1863
rect 5222 1857 5250 1862
rect 4886 1751 4887 1777
rect 4913 1751 4914 1777
rect 4886 1745 4914 1751
rect 5166 1778 5194 1783
rect 5502 1778 5530 1783
rect 5166 1777 5530 1778
rect 5166 1751 5167 1777
rect 5193 1751 5503 1777
rect 5529 1751 5530 1777
rect 5166 1750 5530 1751
rect 5166 1745 5194 1750
rect 5502 1745 5530 1750
rect 5894 1777 5922 1918
rect 5894 1751 5895 1777
rect 5921 1751 5922 1777
rect 5894 1745 5922 1751
rect 1414 1722 1442 1727
rect 1414 1675 1442 1694
rect 1694 1722 1722 1727
rect 1694 1675 1722 1694
rect 2086 1722 2114 1727
rect 2366 1722 2394 1727
rect 2086 1721 2394 1722
rect 2086 1695 2087 1721
rect 2113 1695 2367 1721
rect 2393 1695 2394 1721
rect 2086 1694 2394 1695
rect 2086 1689 2114 1694
rect 2366 1689 2394 1694
rect 3206 1722 3234 1727
rect 3206 1675 3234 1694
rect 3486 1722 3514 1727
rect 3486 1675 3514 1694
rect 5558 1722 5586 1727
rect 5838 1722 5866 1727
rect 5558 1721 5866 1722
rect 5558 1695 5559 1721
rect 5585 1695 5839 1721
rect 5865 1695 5866 1721
rect 5558 1694 5866 1695
rect 5558 1689 5586 1694
rect 5838 1689 5866 1694
rect 2020 1582 2152 1587
rect 2048 1554 2072 1582
rect 2100 1554 2124 1582
rect 2020 1549 2152 1554
rect 3434 1582 3566 1587
rect 3462 1554 3486 1582
rect 3514 1554 3538 1582
rect 3434 1549 3566 1554
rect 4848 1582 4980 1587
rect 4876 1554 4900 1582
rect 4928 1554 4952 1582
rect 4848 1549 4980 1554
rect 6262 1582 6394 1587
rect 6290 1554 6314 1582
rect 6342 1554 6366 1582
rect 6262 1549 6394 1554
<< via2 >>
rect 2020 6285 2048 6286
rect 2020 6259 2021 6285
rect 2021 6259 2047 6285
rect 2047 6259 2048 6285
rect 2020 6258 2048 6259
rect 2072 6285 2100 6286
rect 2072 6259 2073 6285
rect 2073 6259 2099 6285
rect 2099 6259 2100 6285
rect 2072 6258 2100 6259
rect 2124 6285 2152 6286
rect 2124 6259 2125 6285
rect 2125 6259 2151 6285
rect 2151 6259 2152 6285
rect 2124 6258 2152 6259
rect 3434 6285 3462 6286
rect 3434 6259 3435 6285
rect 3435 6259 3461 6285
rect 3461 6259 3462 6285
rect 3434 6258 3462 6259
rect 3486 6285 3514 6286
rect 3486 6259 3487 6285
rect 3487 6259 3513 6285
rect 3513 6259 3514 6285
rect 3486 6258 3514 6259
rect 3538 6285 3566 6286
rect 3538 6259 3539 6285
rect 3539 6259 3565 6285
rect 3565 6259 3566 6285
rect 3538 6258 3566 6259
rect 4848 6285 4876 6286
rect 4848 6259 4849 6285
rect 4849 6259 4875 6285
rect 4875 6259 4876 6285
rect 4848 6258 4876 6259
rect 4900 6285 4928 6286
rect 4900 6259 4901 6285
rect 4901 6259 4927 6285
rect 4927 6259 4928 6285
rect 4900 6258 4928 6259
rect 4952 6285 4980 6286
rect 4952 6259 4953 6285
rect 4953 6259 4979 6285
rect 4979 6259 4980 6285
rect 4952 6258 4980 6259
rect 6262 6285 6290 6286
rect 6262 6259 6263 6285
rect 6263 6259 6289 6285
rect 6289 6259 6290 6285
rect 6262 6258 6290 6259
rect 6314 6285 6342 6286
rect 6314 6259 6315 6285
rect 6315 6259 6341 6285
rect 6341 6259 6342 6285
rect 6314 6258 6342 6259
rect 6366 6285 6394 6286
rect 6366 6259 6367 6285
rect 6367 6259 6393 6285
rect 6393 6259 6394 6285
rect 6366 6258 6394 6259
rect 1134 6089 1162 6090
rect 1134 6063 1135 6089
rect 1135 6063 1161 6089
rect 1161 6063 1162 6089
rect 1134 6062 1162 6063
rect 1470 5977 1498 5978
rect 1470 5951 1471 5977
rect 1471 5951 1497 5977
rect 1497 5951 1498 5977
rect 1470 5950 1498 5951
rect 1313 5893 1341 5894
rect 1313 5867 1314 5893
rect 1314 5867 1340 5893
rect 1340 5867 1341 5893
rect 1313 5866 1341 5867
rect 1365 5893 1393 5894
rect 1365 5867 1366 5893
rect 1366 5867 1392 5893
rect 1392 5867 1393 5893
rect 1365 5866 1393 5867
rect 1417 5893 1445 5894
rect 1417 5867 1418 5893
rect 1418 5867 1444 5893
rect 1444 5867 1445 5893
rect 1526 5894 1554 5922
rect 1694 6062 1722 6090
rect 1417 5866 1445 5867
rect 1750 5950 1778 5978
rect 2926 6145 2954 6146
rect 2926 6119 2927 6145
rect 2927 6119 2953 6145
rect 2953 6119 2954 6145
rect 2926 6118 2954 6119
rect 3374 6118 3402 6146
rect 2478 6089 2506 6090
rect 2478 6063 2479 6089
rect 2479 6063 2505 6089
rect 2505 6063 2506 6089
rect 2478 6062 2506 6063
rect 2870 6062 2898 6090
rect 3262 6089 3290 6090
rect 3262 6063 3263 6089
rect 3263 6063 3289 6089
rect 3289 6063 3290 6089
rect 3262 6062 3290 6063
rect 1862 5782 1890 5810
rect 2030 5838 2058 5866
rect 2422 5809 2450 5810
rect 2422 5783 2423 5809
rect 2423 5783 2449 5809
rect 2449 5783 2450 5809
rect 2422 5782 2450 5783
rect 2727 5893 2755 5894
rect 2727 5867 2728 5893
rect 2728 5867 2754 5893
rect 2754 5867 2755 5893
rect 2727 5866 2755 5867
rect 2779 5893 2807 5894
rect 2779 5867 2780 5893
rect 2780 5867 2806 5893
rect 2806 5867 2807 5893
rect 2779 5866 2807 5867
rect 2831 5893 2859 5894
rect 2831 5867 2832 5893
rect 2832 5867 2858 5893
rect 2858 5867 2859 5893
rect 2831 5866 2859 5867
rect 3654 6145 3682 6146
rect 3654 6119 3655 6145
rect 3655 6119 3681 6145
rect 3681 6119 3682 6145
rect 3654 6118 3682 6119
rect 4270 6145 4298 6146
rect 4270 6119 4271 6145
rect 4271 6119 4297 6145
rect 4297 6119 4298 6145
rect 4270 6118 4298 6119
rect 3598 6089 3626 6090
rect 3598 6063 3599 6089
rect 3599 6063 3625 6089
rect 3625 6063 3626 6089
rect 3598 6062 3626 6063
rect 3990 6089 4018 6090
rect 3990 6063 3991 6089
rect 3991 6063 4017 6089
rect 4017 6063 4018 6089
rect 3990 6062 4018 6063
rect 4326 6089 4354 6090
rect 4326 6063 4327 6089
rect 4327 6063 4353 6089
rect 4353 6063 4354 6089
rect 4326 6062 4354 6063
rect 4141 5893 4169 5894
rect 4141 5867 4142 5893
rect 4142 5867 4168 5893
rect 4168 5867 4169 5893
rect 4141 5866 4169 5867
rect 4193 5893 4221 5894
rect 4193 5867 4194 5893
rect 4194 5867 4220 5893
rect 4220 5867 4221 5893
rect 4193 5866 4221 5867
rect 4245 5893 4273 5894
rect 4245 5867 4246 5893
rect 4246 5867 4272 5893
rect 4272 5867 4273 5893
rect 4245 5866 4273 5867
rect 5555 5893 5583 5894
rect 5555 5867 5556 5893
rect 5556 5867 5582 5893
rect 5582 5867 5583 5893
rect 5555 5866 5583 5867
rect 5607 5893 5635 5894
rect 5607 5867 5608 5893
rect 5608 5867 5634 5893
rect 5634 5867 5635 5893
rect 5607 5866 5635 5867
rect 5659 5893 5687 5894
rect 5659 5867 5660 5893
rect 5660 5867 5686 5893
rect 5686 5867 5687 5893
rect 5659 5866 5687 5867
rect 3990 5641 4018 5642
rect 3990 5615 3991 5641
rect 3991 5615 4017 5641
rect 4017 5615 4018 5641
rect 3990 5614 4018 5615
rect 4270 5641 4298 5642
rect 4270 5615 4271 5641
rect 4271 5615 4297 5641
rect 4297 5615 4298 5641
rect 4270 5614 4298 5615
rect 2020 5501 2048 5502
rect 2020 5475 2021 5501
rect 2021 5475 2047 5501
rect 2047 5475 2048 5501
rect 2020 5474 2048 5475
rect 2072 5501 2100 5502
rect 2072 5475 2073 5501
rect 2073 5475 2099 5501
rect 2099 5475 2100 5501
rect 2072 5474 2100 5475
rect 2124 5501 2152 5502
rect 2124 5475 2125 5501
rect 2125 5475 2151 5501
rect 2151 5475 2152 5501
rect 2124 5474 2152 5475
rect 3434 5501 3462 5502
rect 3434 5475 3435 5501
rect 3435 5475 3461 5501
rect 3461 5475 3462 5501
rect 3434 5474 3462 5475
rect 3486 5501 3514 5502
rect 3486 5475 3487 5501
rect 3487 5475 3513 5501
rect 3513 5475 3514 5501
rect 3486 5474 3514 5475
rect 3538 5501 3566 5502
rect 3538 5475 3539 5501
rect 3539 5475 3565 5501
rect 3565 5475 3566 5501
rect 3538 5474 3566 5475
rect 3878 5417 3906 5418
rect 3878 5391 3879 5417
rect 3879 5391 3905 5417
rect 3905 5391 3906 5417
rect 3878 5390 3906 5391
rect 1134 4998 1162 5026
rect 1190 4886 1218 4914
rect 1022 4550 1050 4578
rect 4848 5501 4876 5502
rect 4848 5475 4849 5501
rect 4849 5475 4875 5501
rect 4875 5475 4876 5501
rect 4848 5474 4876 5475
rect 4900 5501 4928 5502
rect 4900 5475 4901 5501
rect 4901 5475 4927 5501
rect 4927 5475 4928 5501
rect 4900 5474 4928 5475
rect 4952 5501 4980 5502
rect 4952 5475 4953 5501
rect 4953 5475 4979 5501
rect 4979 5475 4980 5501
rect 4952 5474 4980 5475
rect 6262 5501 6290 5502
rect 6262 5475 6263 5501
rect 6263 5475 6289 5501
rect 6289 5475 6290 5501
rect 6262 5474 6290 5475
rect 6314 5501 6342 5502
rect 6314 5475 6315 5501
rect 6315 5475 6341 5501
rect 6341 5475 6342 5501
rect 6314 5474 6342 5475
rect 6366 5501 6394 5502
rect 6366 5475 6367 5501
rect 6367 5475 6393 5501
rect 6393 5475 6394 5501
rect 6366 5474 6394 5475
rect 4326 5390 4354 5418
rect 2478 5361 2506 5362
rect 2478 5335 2479 5361
rect 2479 5335 2505 5361
rect 2505 5335 2506 5361
rect 2478 5334 2506 5335
rect 3430 5334 3458 5362
rect 1526 5305 1554 5306
rect 1526 5279 1527 5305
rect 1527 5279 1553 5305
rect 1553 5279 1554 5305
rect 1526 5278 1554 5279
rect 1806 5305 1834 5306
rect 1806 5279 1807 5305
rect 1807 5279 1833 5305
rect 1833 5279 1834 5305
rect 1806 5278 1834 5279
rect 3206 5305 3234 5306
rect 3206 5279 3207 5305
rect 3207 5279 3233 5305
rect 3233 5279 3234 5305
rect 3206 5278 3234 5279
rect 1313 5109 1341 5110
rect 1313 5083 1314 5109
rect 1314 5083 1340 5109
rect 1340 5083 1341 5109
rect 1313 5082 1341 5083
rect 1365 5109 1393 5110
rect 1365 5083 1366 5109
rect 1366 5083 1392 5109
rect 1392 5083 1393 5109
rect 1365 5082 1393 5083
rect 1417 5109 1445 5110
rect 1417 5083 1418 5109
rect 1418 5083 1444 5109
rect 1444 5083 1445 5109
rect 1417 5082 1445 5083
rect 1414 5025 1442 5026
rect 1414 4999 1415 5025
rect 1415 4999 1441 5025
rect 1441 4999 1442 5025
rect 1414 4998 1442 4999
rect 1806 4913 1834 4914
rect 1806 4887 1807 4913
rect 1807 4887 1833 4913
rect 1833 4887 1834 4913
rect 1806 4886 1834 4887
rect 2727 5109 2755 5110
rect 2727 5083 2728 5109
rect 2728 5083 2754 5109
rect 2754 5083 2755 5109
rect 2727 5082 2755 5083
rect 2779 5109 2807 5110
rect 2779 5083 2780 5109
rect 2780 5083 2806 5109
rect 2806 5083 2807 5109
rect 2779 5082 2807 5083
rect 2831 5109 2859 5110
rect 2831 5083 2832 5109
rect 2832 5083 2858 5109
rect 2858 5083 2859 5109
rect 2831 5082 2859 5083
rect 3542 5361 3570 5362
rect 3542 5335 3543 5361
rect 3543 5335 3569 5361
rect 3569 5335 3570 5361
rect 3542 5334 3570 5335
rect 4214 5361 4242 5362
rect 4214 5335 4215 5361
rect 4215 5335 4241 5361
rect 4241 5335 4242 5361
rect 4214 5334 4242 5335
rect 3486 5305 3514 5306
rect 3486 5279 3487 5305
rect 3487 5279 3513 5305
rect 3513 5279 3514 5305
rect 3486 5278 3514 5279
rect 4141 5109 4169 5110
rect 4141 5083 4142 5109
rect 4142 5083 4168 5109
rect 4168 5083 4169 5109
rect 4141 5082 4169 5083
rect 4193 5109 4221 5110
rect 4193 5083 4194 5109
rect 4194 5083 4220 5109
rect 4220 5083 4221 5109
rect 4193 5082 4221 5083
rect 4245 5109 4273 5110
rect 4245 5083 4246 5109
rect 4246 5083 4272 5109
rect 4272 5083 4273 5109
rect 4245 5082 4273 5083
rect 5555 5109 5583 5110
rect 5555 5083 5556 5109
rect 5556 5083 5582 5109
rect 5582 5083 5583 5109
rect 5555 5082 5583 5083
rect 5607 5109 5635 5110
rect 5607 5083 5608 5109
rect 5608 5083 5634 5109
rect 5634 5083 5635 5109
rect 5607 5082 5635 5083
rect 5659 5109 5687 5110
rect 5659 5083 5660 5109
rect 5660 5083 5686 5109
rect 5686 5083 5687 5109
rect 5659 5082 5687 5083
rect 1526 4577 1554 4578
rect 1526 4551 1527 4577
rect 1527 4551 1553 4577
rect 1553 4551 1554 4577
rect 1526 4550 1554 4551
rect 1313 4325 1341 4326
rect 1313 4299 1314 4325
rect 1314 4299 1340 4325
rect 1340 4299 1341 4325
rect 1313 4298 1341 4299
rect 1365 4325 1393 4326
rect 1365 4299 1366 4325
rect 1366 4299 1392 4325
rect 1392 4299 1393 4325
rect 1365 4298 1393 4299
rect 1417 4325 1445 4326
rect 1417 4299 1418 4325
rect 1418 4299 1444 4325
rect 1444 4299 1445 4325
rect 1417 4298 1445 4299
rect 3206 4830 3234 4858
rect 2020 4717 2048 4718
rect 2020 4691 2021 4717
rect 2021 4691 2047 4717
rect 2047 4691 2048 4717
rect 2020 4690 2048 4691
rect 2072 4717 2100 4718
rect 2072 4691 2073 4717
rect 2073 4691 2099 4717
rect 2099 4691 2100 4717
rect 2072 4690 2100 4691
rect 2124 4717 2152 4718
rect 2124 4691 2125 4717
rect 2125 4691 2151 4717
rect 2151 4691 2152 4717
rect 2124 4690 2152 4691
rect 3150 4774 3178 4802
rect 2870 4633 2898 4634
rect 2870 4607 2871 4633
rect 2871 4607 2897 4633
rect 2897 4607 2898 4633
rect 2870 4606 2898 4607
rect 3486 4857 3514 4858
rect 3486 4831 3487 4857
rect 3487 4831 3513 4857
rect 3513 4831 3514 4857
rect 3486 4830 3514 4831
rect 3766 4801 3794 4802
rect 3766 4775 3767 4801
rect 3767 4775 3793 4801
rect 3793 4775 3794 4801
rect 3766 4774 3794 4775
rect 3434 4717 3462 4718
rect 3434 4691 3435 4717
rect 3435 4691 3461 4717
rect 3461 4691 3462 4717
rect 3434 4690 3462 4691
rect 3486 4717 3514 4718
rect 3486 4691 3487 4717
rect 3487 4691 3513 4717
rect 3513 4691 3514 4717
rect 3486 4690 3514 4691
rect 3538 4717 3566 4718
rect 3538 4691 3539 4717
rect 3539 4691 3565 4717
rect 3565 4691 3566 4717
rect 3538 4690 3566 4691
rect 4848 4717 4876 4718
rect 4848 4691 4849 4717
rect 4849 4691 4875 4717
rect 4875 4691 4876 4717
rect 4848 4690 4876 4691
rect 4900 4717 4928 4718
rect 4900 4691 4901 4717
rect 4901 4691 4927 4717
rect 4927 4691 4928 4717
rect 4900 4690 4928 4691
rect 4952 4717 4980 4718
rect 4952 4691 4953 4717
rect 4953 4691 4979 4717
rect 4979 4691 4980 4717
rect 4952 4690 4980 4691
rect 6262 4717 6290 4718
rect 6262 4691 6263 4717
rect 6263 4691 6289 4717
rect 6289 4691 6290 4717
rect 6262 4690 6290 4691
rect 6314 4717 6342 4718
rect 6314 4691 6315 4717
rect 6315 4691 6341 4717
rect 6341 4691 6342 4717
rect 6314 4690 6342 4691
rect 6366 4717 6394 4718
rect 6366 4691 6367 4717
rect 6367 4691 6393 4717
rect 6393 4691 6394 4717
rect 6366 4690 6394 4691
rect 3486 4606 3514 4634
rect 2030 4214 2058 4242
rect 2478 4521 2506 4522
rect 2478 4495 2479 4521
rect 2479 4495 2505 4521
rect 2505 4495 2506 4521
rect 2478 4494 2506 4495
rect 2422 4382 2450 4410
rect 1078 4073 1106 4074
rect 1078 4047 1079 4073
rect 1079 4047 1105 4073
rect 1105 4047 1106 4073
rect 1078 4046 1106 4047
rect 910 3990 938 4018
rect 2020 3933 2048 3934
rect 2020 3907 2021 3933
rect 2021 3907 2047 3933
rect 2047 3907 2048 3933
rect 2020 3906 2048 3907
rect 2072 3933 2100 3934
rect 2072 3907 2073 3933
rect 2073 3907 2099 3933
rect 2099 3907 2100 3933
rect 2072 3906 2100 3907
rect 2124 3933 2152 3934
rect 2124 3907 2125 3933
rect 2125 3907 2151 3933
rect 2151 3907 2152 3933
rect 2124 3906 2152 3907
rect 1190 3598 1218 3626
rect 1313 3541 1341 3542
rect 1313 3515 1314 3541
rect 1314 3515 1340 3541
rect 1340 3515 1341 3541
rect 1313 3514 1341 3515
rect 1365 3541 1393 3542
rect 1365 3515 1366 3541
rect 1366 3515 1392 3541
rect 1392 3515 1393 3541
rect 1365 3514 1393 3515
rect 1417 3541 1445 3542
rect 1417 3515 1418 3541
rect 1418 3515 1444 3541
rect 1444 3515 1445 3541
rect 1417 3514 1445 3515
rect 1470 3289 1498 3290
rect 1470 3263 1471 3289
rect 1471 3263 1497 3289
rect 1497 3263 1498 3289
rect 1470 3262 1498 3263
rect 1526 3038 1554 3066
rect 1358 2841 1386 2842
rect 1358 2815 1359 2841
rect 1359 2815 1385 2841
rect 1385 2815 1386 2841
rect 1358 2814 1386 2815
rect 1313 2757 1341 2758
rect 1313 2731 1314 2757
rect 1314 2731 1340 2757
rect 1340 2731 1341 2757
rect 1313 2730 1341 2731
rect 1365 2757 1393 2758
rect 1365 2731 1366 2757
rect 1366 2731 1392 2757
rect 1392 2731 1393 2757
rect 1365 2730 1393 2731
rect 1417 2757 1445 2758
rect 1417 2731 1418 2757
rect 1418 2731 1444 2757
rect 1444 2731 1445 2757
rect 1417 2730 1445 2731
rect 1190 2478 1218 2506
rect 1022 2198 1050 2226
rect 2727 4325 2755 4326
rect 2727 4299 2728 4325
rect 2728 4299 2754 4325
rect 2754 4299 2755 4325
rect 2727 4298 2755 4299
rect 2779 4325 2807 4326
rect 2779 4299 2780 4325
rect 2780 4299 2806 4325
rect 2806 4299 2807 4325
rect 2779 4298 2807 4299
rect 2831 4325 2859 4326
rect 2831 4299 2832 4325
rect 2832 4299 2858 4325
rect 2858 4299 2859 4325
rect 2831 4298 2859 4299
rect 3430 4494 3458 4522
rect 3822 4409 3850 4410
rect 3822 4383 3823 4409
rect 3823 4383 3849 4409
rect 3849 4383 3850 4409
rect 3822 4382 3850 4383
rect 4141 4325 4169 4326
rect 4141 4299 4142 4325
rect 4142 4299 4168 4325
rect 4168 4299 4169 4325
rect 4141 4298 4169 4299
rect 4193 4325 4221 4326
rect 4193 4299 4194 4325
rect 4194 4299 4220 4325
rect 4220 4299 4221 4325
rect 4193 4298 4221 4299
rect 4245 4325 4273 4326
rect 4245 4299 4246 4325
rect 4246 4299 4272 4325
rect 4272 4299 4273 4325
rect 4245 4298 4273 4299
rect 5555 4325 5583 4326
rect 5555 4299 5556 4325
rect 5556 4299 5582 4325
rect 5582 4299 5583 4325
rect 5555 4298 5583 4299
rect 5607 4325 5635 4326
rect 5607 4299 5608 4325
rect 5608 4299 5634 4325
rect 5634 4299 5635 4325
rect 5607 4298 5635 4299
rect 5659 4325 5687 4326
rect 5659 4299 5660 4325
rect 5660 4299 5686 4325
rect 5686 4299 5687 4325
rect 5659 4298 5687 4299
rect 3878 4214 3906 4242
rect 3038 3990 3066 4018
rect 2702 3849 2730 3850
rect 2702 3823 2703 3849
rect 2703 3823 2729 3849
rect 2729 3823 2730 3849
rect 2702 3822 2730 3823
rect 3766 4073 3794 4074
rect 3766 4047 3767 4073
rect 3767 4047 3793 4073
rect 3793 4047 3794 4073
rect 3766 4046 3794 4047
rect 3486 3990 3514 4018
rect 3434 3933 3462 3934
rect 3434 3907 3435 3933
rect 3435 3907 3461 3933
rect 3461 3907 3462 3933
rect 3434 3906 3462 3907
rect 3486 3933 3514 3934
rect 3486 3907 3487 3933
rect 3487 3907 3513 3933
rect 3513 3907 3514 3933
rect 3486 3906 3514 3907
rect 3538 3933 3566 3934
rect 3538 3907 3539 3933
rect 3539 3907 3565 3933
rect 3565 3907 3566 3933
rect 3538 3906 3566 3907
rect 3374 3822 3402 3850
rect 1638 3318 1666 3346
rect 2198 3345 2226 3346
rect 2198 3319 2199 3345
rect 2199 3319 2225 3345
rect 2225 3319 2226 3345
rect 2198 3318 2226 3319
rect 2727 3541 2755 3542
rect 2727 3515 2728 3541
rect 2728 3515 2754 3541
rect 2754 3515 2755 3541
rect 2727 3514 2755 3515
rect 2779 3541 2807 3542
rect 2779 3515 2780 3541
rect 2780 3515 2806 3541
rect 2806 3515 2807 3541
rect 2779 3514 2807 3515
rect 2831 3541 2859 3542
rect 2831 3515 2832 3541
rect 2832 3515 2858 3541
rect 2858 3515 2859 3541
rect 2831 3514 2859 3515
rect 4046 3737 4074 3738
rect 4046 3711 4047 3737
rect 4047 3711 4073 3737
rect 4073 3711 4074 3737
rect 4046 3710 4074 3711
rect 3038 3374 3066 3402
rect 4848 3933 4876 3934
rect 4848 3907 4849 3933
rect 4849 3907 4875 3933
rect 4875 3907 4876 3933
rect 4848 3906 4876 3907
rect 4900 3933 4928 3934
rect 4900 3907 4901 3933
rect 4901 3907 4927 3933
rect 4927 3907 4928 3933
rect 4900 3906 4928 3907
rect 4952 3933 4980 3934
rect 4952 3907 4953 3933
rect 4953 3907 4979 3933
rect 4979 3907 4980 3933
rect 4952 3906 4980 3907
rect 6262 3933 6290 3934
rect 6262 3907 6263 3933
rect 6263 3907 6289 3933
rect 6289 3907 6290 3933
rect 6262 3906 6290 3907
rect 6314 3933 6342 3934
rect 6314 3907 6315 3933
rect 6315 3907 6341 3933
rect 6341 3907 6342 3933
rect 6314 3906 6342 3907
rect 6366 3933 6394 3934
rect 6366 3907 6367 3933
rect 6367 3907 6393 3933
rect 6393 3907 6394 3933
rect 6366 3906 6394 3907
rect 4326 3737 4354 3738
rect 4326 3711 4327 3737
rect 4327 3711 4353 3737
rect 4353 3711 4354 3737
rect 4326 3710 4354 3711
rect 3990 3625 4018 3626
rect 3990 3599 3991 3625
rect 3991 3599 4017 3625
rect 4017 3599 4018 3625
rect 3990 3598 4018 3599
rect 3654 3374 3682 3402
rect 4141 3541 4169 3542
rect 4141 3515 4142 3541
rect 4142 3515 4168 3541
rect 4168 3515 4169 3541
rect 4141 3514 4169 3515
rect 4193 3541 4221 3542
rect 4193 3515 4194 3541
rect 4194 3515 4220 3541
rect 4220 3515 4221 3541
rect 4193 3514 4221 3515
rect 4245 3541 4273 3542
rect 4245 3515 4246 3541
rect 4246 3515 4272 3541
rect 4272 3515 4273 3541
rect 4245 3514 4273 3515
rect 5555 3541 5583 3542
rect 5555 3515 5556 3541
rect 5556 3515 5582 3541
rect 5582 3515 5583 3541
rect 5555 3514 5583 3515
rect 5607 3541 5635 3542
rect 5607 3515 5608 3541
rect 5608 3515 5634 3541
rect 5634 3515 5635 3541
rect 5607 3514 5635 3515
rect 5659 3541 5687 3542
rect 5659 3515 5660 3541
rect 5660 3515 5686 3541
rect 5686 3515 5687 3541
rect 5659 3514 5687 3515
rect 4102 3318 4130 3346
rect 4382 3345 4410 3346
rect 4382 3319 4383 3345
rect 4383 3319 4409 3345
rect 4409 3319 4410 3345
rect 4382 3318 4410 3319
rect 1750 3289 1778 3290
rect 1750 3263 1751 3289
rect 1751 3263 1777 3289
rect 1777 3263 1778 3289
rect 1750 3262 1778 3263
rect 2422 3262 2450 3290
rect 2020 3149 2048 3150
rect 2020 3123 2021 3149
rect 2021 3123 2047 3149
rect 2047 3123 2048 3149
rect 2020 3122 2048 3123
rect 2072 3149 2100 3150
rect 2072 3123 2073 3149
rect 2073 3123 2099 3149
rect 2099 3123 2100 3149
rect 2072 3122 2100 3123
rect 2124 3149 2152 3150
rect 2124 3123 2125 3149
rect 2125 3123 2151 3149
rect 2151 3123 2152 3149
rect 2124 3122 2152 3123
rect 2310 3065 2338 3066
rect 2310 3039 2311 3065
rect 2311 3039 2337 3065
rect 2337 3039 2338 3065
rect 2310 3038 2338 3039
rect 1918 2814 1946 2842
rect 1638 2646 1666 2674
rect 1862 2673 1890 2674
rect 1862 2647 1863 2673
rect 1863 2647 1889 2673
rect 1889 2647 1890 2673
rect 1862 2646 1890 2647
rect 1582 2590 1610 2618
rect 3094 3206 3122 3234
rect 2758 3009 2786 3010
rect 2758 2983 2759 3009
rect 2759 2983 2785 3009
rect 2785 2983 2786 3009
rect 2758 2982 2786 2983
rect 3654 3233 3682 3234
rect 3654 3207 3655 3233
rect 3655 3207 3681 3233
rect 3681 3207 3682 3233
rect 3654 3206 3682 3207
rect 3434 3149 3462 3150
rect 3434 3123 3435 3149
rect 3435 3123 3461 3149
rect 3461 3123 3462 3149
rect 3434 3122 3462 3123
rect 3486 3149 3514 3150
rect 3486 3123 3487 3149
rect 3487 3123 3513 3149
rect 3513 3123 3514 3149
rect 3486 3122 3514 3123
rect 3538 3149 3566 3150
rect 3538 3123 3539 3149
rect 3539 3123 3565 3149
rect 3565 3123 3566 3149
rect 3538 3122 3566 3123
rect 4046 3289 4074 3290
rect 4046 3263 4047 3289
rect 4047 3263 4073 3289
rect 4073 3263 4074 3289
rect 4046 3262 4074 3263
rect 4662 3289 4690 3290
rect 4662 3263 4663 3289
rect 4663 3263 4689 3289
rect 4689 3263 4690 3289
rect 4662 3262 4690 3263
rect 6006 3262 6034 3290
rect 3766 3009 3794 3010
rect 3766 2983 3767 3009
rect 3767 2983 3793 3009
rect 3793 2983 3794 3009
rect 3766 2982 3794 2983
rect 2814 2953 2842 2954
rect 2814 2927 2815 2953
rect 2815 2927 2841 2953
rect 2841 2927 2842 2953
rect 2814 2926 2842 2927
rect 3430 2953 3458 2954
rect 3430 2927 3431 2953
rect 3431 2927 3457 2953
rect 3457 2927 3458 2953
rect 3430 2926 3458 2927
rect 2727 2757 2755 2758
rect 2727 2731 2728 2757
rect 2728 2731 2754 2757
rect 2754 2731 2755 2757
rect 2727 2730 2755 2731
rect 2779 2757 2807 2758
rect 2779 2731 2780 2757
rect 2780 2731 2806 2757
rect 2806 2731 2807 2757
rect 2779 2730 2807 2731
rect 2831 2757 2859 2758
rect 2831 2731 2832 2757
rect 2832 2731 2858 2757
rect 2858 2731 2859 2757
rect 2831 2730 2859 2731
rect 3318 2646 3346 2674
rect 2366 2590 2394 2618
rect 3262 2561 3290 2562
rect 3262 2535 3263 2561
rect 3263 2535 3289 2561
rect 3289 2535 3290 2561
rect 3262 2534 3290 2535
rect 3822 2646 3850 2674
rect 3598 2590 3626 2618
rect 3542 2561 3570 2562
rect 3542 2535 3543 2561
rect 3543 2535 3569 2561
rect 3569 2535 3570 2561
rect 3542 2534 3570 2535
rect 3934 2561 3962 2562
rect 3934 2535 3935 2561
rect 3935 2535 3961 2561
rect 3961 2535 3962 2561
rect 3934 2534 3962 2535
rect 2926 2449 2954 2450
rect 2926 2423 2927 2449
rect 2927 2423 2953 2449
rect 2953 2423 2954 2449
rect 2926 2422 2954 2423
rect 3374 2422 3402 2450
rect 2020 2365 2048 2366
rect 2020 2339 2021 2365
rect 2021 2339 2047 2365
rect 2047 2339 2048 2365
rect 2020 2338 2048 2339
rect 2072 2365 2100 2366
rect 2072 2339 2073 2365
rect 2073 2339 2099 2365
rect 2099 2339 2100 2365
rect 2072 2338 2100 2339
rect 2124 2365 2152 2366
rect 2124 2339 2125 2365
rect 2125 2339 2151 2365
rect 2151 2339 2152 2365
rect 2124 2338 2152 2339
rect 2366 2254 2394 2282
rect 3598 2422 3626 2450
rect 3434 2365 3462 2366
rect 3434 2339 3435 2365
rect 3435 2339 3461 2365
rect 3461 2339 3462 2365
rect 3434 2338 3462 2339
rect 3486 2365 3514 2366
rect 3486 2339 3487 2365
rect 3487 2339 3513 2365
rect 3513 2339 3514 2365
rect 3486 2338 3514 2339
rect 3538 2365 3566 2366
rect 3538 2339 3539 2365
rect 3539 2339 3565 2365
rect 3565 2339 3566 2365
rect 3538 2338 3566 2339
rect 2646 2169 2674 2170
rect 2646 2143 2647 2169
rect 2647 2143 2673 2169
rect 2673 2143 2674 2169
rect 2646 2142 2674 2143
rect 3318 2169 3346 2170
rect 3318 2143 3319 2169
rect 3319 2143 3345 2169
rect 3345 2143 3346 2169
rect 3318 2142 3346 2143
rect 1526 2086 1554 2114
rect 1313 1973 1341 1974
rect 1313 1947 1314 1973
rect 1314 1947 1340 1973
rect 1340 1947 1341 1973
rect 1313 1946 1341 1947
rect 1365 1973 1393 1974
rect 1365 1947 1366 1973
rect 1366 1947 1392 1973
rect 1392 1947 1393 1973
rect 1365 1946 1393 1947
rect 1417 1973 1445 1974
rect 1417 1947 1418 1973
rect 1418 1947 1444 1973
rect 1444 1947 1445 1973
rect 1417 1946 1445 1947
rect 1134 1862 1162 1890
rect 1750 2030 1778 2058
rect 1078 1833 1106 1834
rect 1078 1807 1079 1833
rect 1079 1807 1105 1833
rect 1105 1807 1106 1833
rect 1078 1806 1106 1807
rect 2030 1889 2058 1890
rect 2030 1863 2031 1889
rect 2031 1863 2057 1889
rect 2057 1863 2058 1889
rect 2030 1862 2058 1863
rect 2727 1973 2755 1974
rect 2727 1947 2728 1973
rect 2728 1947 2754 1973
rect 2754 1947 2755 1973
rect 2727 1946 2755 1947
rect 2779 1973 2807 1974
rect 2779 1947 2780 1973
rect 2780 1947 2806 1973
rect 2806 1947 2807 1973
rect 2779 1946 2807 1947
rect 2831 1973 2859 1974
rect 2831 1947 2832 1973
rect 2832 1947 2858 1973
rect 2858 1947 2859 1973
rect 2831 1946 2859 1947
rect 4718 3233 4746 3234
rect 4718 3207 4719 3233
rect 4719 3207 4745 3233
rect 4745 3207 4746 3233
rect 4718 3206 4746 3207
rect 5950 3206 5978 3234
rect 4848 3149 4876 3150
rect 4848 3123 4849 3149
rect 4849 3123 4875 3149
rect 4875 3123 4876 3149
rect 4848 3122 4876 3123
rect 4900 3149 4928 3150
rect 4900 3123 4901 3149
rect 4901 3123 4927 3149
rect 4927 3123 4928 3149
rect 4900 3122 4928 3123
rect 4952 3149 4980 3150
rect 4952 3123 4953 3149
rect 4953 3123 4979 3149
rect 4979 3123 4980 3149
rect 4952 3122 4980 3123
rect 4158 2953 4186 2954
rect 4158 2927 4159 2953
rect 4159 2927 4185 2953
rect 4185 2927 4186 2953
rect 4158 2926 4186 2927
rect 4438 2953 4466 2954
rect 4438 2927 4439 2953
rect 4439 2927 4465 2953
rect 4465 2927 4466 2953
rect 4438 2926 4466 2927
rect 4886 2953 4914 2954
rect 4886 2927 4887 2953
rect 4887 2927 4913 2953
rect 4913 2927 4914 2953
rect 4886 2926 4914 2927
rect 5166 2926 5194 2954
rect 4141 2757 4169 2758
rect 4141 2731 4142 2757
rect 4142 2731 4168 2757
rect 4168 2731 4169 2757
rect 4141 2730 4169 2731
rect 4193 2757 4221 2758
rect 4193 2731 4194 2757
rect 4194 2731 4220 2757
rect 4220 2731 4221 2757
rect 4193 2730 4221 2731
rect 4245 2757 4273 2758
rect 4245 2731 4246 2757
rect 4246 2731 4272 2757
rect 4272 2731 4273 2757
rect 4245 2730 4273 2731
rect 4214 2617 4242 2618
rect 4214 2591 4215 2617
rect 4215 2591 4241 2617
rect 4241 2591 4242 2617
rect 4214 2590 4242 2591
rect 4270 2561 4298 2562
rect 4270 2535 4271 2561
rect 4271 2535 4297 2561
rect 4297 2535 4298 2561
rect 4270 2534 4298 2535
rect 4942 2561 4970 2562
rect 4942 2535 4943 2561
rect 4943 2535 4969 2561
rect 4969 2535 4970 2561
rect 4942 2534 4970 2535
rect 4046 2478 4074 2506
rect 3990 2254 4018 2282
rect 4606 2254 4634 2282
rect 4774 2422 4802 2450
rect 5222 2814 5250 2842
rect 5894 2814 5922 2842
rect 5555 2757 5583 2758
rect 5555 2731 5556 2757
rect 5556 2731 5582 2757
rect 5582 2731 5583 2757
rect 5555 2730 5583 2731
rect 5607 2757 5635 2758
rect 5607 2731 5608 2757
rect 5608 2731 5634 2757
rect 5634 2731 5635 2757
rect 5607 2730 5635 2731
rect 5659 2757 5687 2758
rect 5659 2731 5660 2757
rect 5660 2731 5686 2757
rect 5686 2731 5687 2757
rect 5659 2730 5687 2731
rect 5278 2561 5306 2562
rect 5278 2535 5279 2561
rect 5279 2535 5305 2561
rect 5305 2535 5306 2561
rect 5278 2534 5306 2535
rect 4998 2422 5026 2450
rect 5558 2422 5586 2450
rect 4848 2365 4876 2366
rect 4848 2339 4849 2365
rect 4849 2339 4875 2365
rect 4875 2339 4876 2365
rect 4848 2338 4876 2339
rect 4900 2365 4928 2366
rect 4900 2339 4901 2365
rect 4901 2339 4927 2365
rect 4927 2339 4928 2365
rect 4900 2338 4928 2339
rect 4952 2365 4980 2366
rect 4952 2339 4953 2365
rect 4953 2339 4979 2365
rect 4979 2339 4980 2365
rect 4952 2338 4980 2339
rect 4550 2198 4578 2226
rect 5222 2281 5250 2282
rect 5222 2255 5223 2281
rect 5223 2255 5249 2281
rect 5249 2255 5250 2281
rect 5222 2254 5250 2255
rect 3990 2169 4018 2170
rect 3990 2143 3991 2169
rect 3991 2143 4017 2169
rect 4017 2143 4018 2169
rect 3990 2142 4018 2143
rect 4270 2169 4298 2170
rect 4270 2143 4271 2169
rect 4271 2143 4297 2169
rect 4297 2143 4298 2169
rect 4270 2142 4298 2143
rect 4141 1973 4169 1974
rect 4141 1947 4142 1973
rect 4142 1947 4168 1973
rect 4168 1947 4169 1973
rect 4141 1946 4169 1947
rect 4193 1973 4221 1974
rect 4193 1947 4194 1973
rect 4194 1947 4220 1973
rect 4220 1947 4221 1973
rect 4193 1946 4221 1947
rect 4245 1973 4273 1974
rect 4245 1947 4246 1973
rect 4246 1947 4272 1973
rect 4272 1947 4273 1973
rect 4245 1946 4273 1947
rect 3598 1862 3626 1890
rect 3878 1889 3906 1890
rect 3878 1863 3879 1889
rect 3879 1863 3905 1889
rect 3905 1863 3906 1889
rect 3878 1862 3906 1863
rect 4886 2113 4914 2114
rect 4886 2087 4887 2113
rect 4887 2087 4913 2113
rect 4913 2087 4914 2113
rect 4886 2086 4914 2087
rect 4326 1862 4354 1890
rect 4886 1974 4914 2002
rect 3150 1806 3178 1834
rect 4830 1833 4858 1834
rect 4830 1807 4831 1833
rect 4831 1807 4857 1833
rect 4857 1807 4858 1833
rect 4830 1806 4858 1807
rect 3542 1777 3570 1778
rect 3542 1751 3543 1777
rect 3543 1751 3569 1777
rect 3569 1751 3570 1777
rect 3542 1750 3570 1751
rect 4214 1777 4242 1778
rect 4214 1751 4215 1777
rect 4215 1751 4241 1777
rect 4241 1751 4242 1777
rect 4214 1750 4242 1751
rect 5614 2169 5642 2170
rect 5614 2143 5615 2169
rect 5615 2143 5641 2169
rect 5641 2143 5642 2169
rect 5614 2142 5642 2143
rect 5555 1973 5583 1974
rect 5555 1947 5556 1973
rect 5556 1947 5582 1973
rect 5582 1947 5583 1973
rect 5555 1946 5583 1947
rect 5607 1973 5635 1974
rect 5607 1947 5608 1973
rect 5608 1947 5634 1973
rect 5634 1947 5635 1973
rect 5607 1946 5635 1947
rect 5659 1973 5687 1974
rect 5659 1947 5660 1973
rect 5660 1947 5686 1973
rect 5686 1947 5687 1973
rect 5659 1946 5687 1947
rect 6262 3149 6290 3150
rect 6262 3123 6263 3149
rect 6263 3123 6289 3149
rect 6289 3123 6290 3149
rect 6262 3122 6290 3123
rect 6314 3149 6342 3150
rect 6314 3123 6315 3149
rect 6315 3123 6341 3149
rect 6341 3123 6342 3149
rect 6314 3122 6342 3123
rect 6366 3149 6394 3150
rect 6366 3123 6367 3149
rect 6367 3123 6393 3149
rect 6393 3123 6394 3149
rect 6366 3122 6394 3123
rect 6262 2365 6290 2366
rect 6262 2339 6263 2365
rect 6263 2339 6289 2365
rect 6289 2339 6290 2365
rect 6262 2338 6290 2339
rect 6314 2365 6342 2366
rect 6314 2339 6315 2365
rect 6315 2339 6341 2365
rect 6341 2339 6342 2365
rect 6314 2338 6342 2339
rect 6366 2365 6394 2366
rect 6366 2339 6367 2365
rect 6367 2339 6393 2365
rect 6393 2339 6394 2365
rect 6366 2338 6394 2339
rect 5950 2169 5978 2170
rect 5950 2143 5951 2169
rect 5951 2143 5977 2169
rect 5977 2143 5978 2169
rect 5950 2142 5978 2143
rect 1414 1721 1442 1722
rect 1414 1695 1415 1721
rect 1415 1695 1441 1721
rect 1441 1695 1442 1721
rect 1414 1694 1442 1695
rect 1694 1721 1722 1722
rect 1694 1695 1695 1721
rect 1695 1695 1721 1721
rect 1721 1695 1722 1721
rect 1694 1694 1722 1695
rect 3206 1721 3234 1722
rect 3206 1695 3207 1721
rect 3207 1695 3233 1721
rect 3233 1695 3234 1721
rect 3206 1694 3234 1695
rect 3486 1721 3514 1722
rect 3486 1695 3487 1721
rect 3487 1695 3513 1721
rect 3513 1695 3514 1721
rect 3486 1694 3514 1695
rect 2020 1581 2048 1582
rect 2020 1555 2021 1581
rect 2021 1555 2047 1581
rect 2047 1555 2048 1581
rect 2020 1554 2048 1555
rect 2072 1581 2100 1582
rect 2072 1555 2073 1581
rect 2073 1555 2099 1581
rect 2099 1555 2100 1581
rect 2072 1554 2100 1555
rect 2124 1581 2152 1582
rect 2124 1555 2125 1581
rect 2125 1555 2151 1581
rect 2151 1555 2152 1581
rect 2124 1554 2152 1555
rect 3434 1581 3462 1582
rect 3434 1555 3435 1581
rect 3435 1555 3461 1581
rect 3461 1555 3462 1581
rect 3434 1554 3462 1555
rect 3486 1581 3514 1582
rect 3486 1555 3487 1581
rect 3487 1555 3513 1581
rect 3513 1555 3514 1581
rect 3486 1554 3514 1555
rect 3538 1581 3566 1582
rect 3538 1555 3539 1581
rect 3539 1555 3565 1581
rect 3565 1555 3566 1581
rect 3538 1554 3566 1555
rect 4848 1581 4876 1582
rect 4848 1555 4849 1581
rect 4849 1555 4875 1581
rect 4875 1555 4876 1581
rect 4848 1554 4876 1555
rect 4900 1581 4928 1582
rect 4900 1555 4901 1581
rect 4901 1555 4927 1581
rect 4927 1555 4928 1581
rect 4900 1554 4928 1555
rect 4952 1581 4980 1582
rect 4952 1555 4953 1581
rect 4953 1555 4979 1581
rect 4979 1555 4980 1581
rect 4952 1554 4980 1555
rect 6262 1581 6290 1582
rect 6262 1555 6263 1581
rect 6263 1555 6289 1581
rect 6289 1555 6290 1581
rect 6262 1554 6290 1555
rect 6314 1581 6342 1582
rect 6314 1555 6315 1581
rect 6315 1555 6341 1581
rect 6341 1555 6342 1581
rect 6314 1554 6342 1555
rect 6366 1581 6394 1582
rect 6366 1555 6367 1581
rect 6367 1555 6393 1581
rect 6393 1555 6394 1581
rect 6366 1554 6394 1555
<< metal3 >>
rect 2015 6258 2020 6286
rect 2048 6258 2072 6286
rect 2100 6258 2124 6286
rect 2152 6258 2157 6286
rect 3429 6258 3434 6286
rect 3462 6258 3486 6286
rect 3514 6258 3538 6286
rect 3566 6258 3571 6286
rect 4843 6258 4848 6286
rect 4876 6258 4900 6286
rect 4928 6258 4952 6286
rect 4980 6258 4985 6286
rect 6257 6258 6262 6286
rect 6290 6258 6314 6286
rect 6342 6258 6366 6286
rect 6394 6258 6399 6286
rect 2921 6118 2926 6146
rect 2954 6118 3374 6146
rect 3402 6118 3407 6146
rect 3649 6118 3654 6146
rect 3682 6118 4270 6146
rect 4298 6118 4303 6146
rect 1129 6062 1134 6090
rect 1162 6062 1694 6090
rect 1722 6062 1727 6090
rect 2473 6062 2478 6090
rect 2506 6062 2870 6090
rect 2898 6062 2903 6090
rect 3257 6062 3262 6090
rect 3290 6062 3598 6090
rect 3626 6062 3631 6090
rect 3985 6062 3990 6090
rect 4018 6062 4326 6090
rect 4354 6062 4359 6090
rect 1465 5950 1470 5978
rect 1498 5950 1750 5978
rect 1778 5950 1783 5978
rect 1521 5894 1526 5922
rect 1554 5894 2058 5922
rect 1308 5866 1313 5894
rect 1341 5866 1365 5894
rect 1393 5866 1417 5894
rect 1445 5866 1450 5894
rect 2030 5866 2058 5894
rect 2722 5866 2727 5894
rect 2755 5866 2779 5894
rect 2807 5866 2831 5894
rect 2859 5866 2864 5894
rect 4136 5866 4141 5894
rect 4169 5866 4193 5894
rect 4221 5866 4245 5894
rect 4273 5866 4278 5894
rect 5550 5866 5555 5894
rect 5583 5866 5607 5894
rect 5635 5866 5659 5894
rect 5687 5866 5692 5894
rect 2025 5838 2030 5866
rect 2058 5838 2063 5866
rect 1857 5782 1862 5810
rect 1890 5782 2422 5810
rect 2450 5782 2455 5810
rect 3985 5614 3990 5642
rect 4018 5614 4270 5642
rect 4298 5614 4303 5642
rect 2015 5474 2020 5502
rect 2048 5474 2072 5502
rect 2100 5474 2124 5502
rect 2152 5474 2157 5502
rect 3429 5474 3434 5502
rect 3462 5474 3486 5502
rect 3514 5474 3538 5502
rect 3566 5474 3571 5502
rect 4843 5474 4848 5502
rect 4876 5474 4900 5502
rect 4928 5474 4952 5502
rect 4980 5474 4985 5502
rect 6257 5474 6262 5502
rect 6290 5474 6314 5502
rect 6342 5474 6366 5502
rect 6394 5474 6399 5502
rect 3873 5390 3878 5418
rect 3906 5390 4326 5418
rect 4354 5390 4359 5418
rect 2473 5334 2478 5362
rect 2506 5334 3430 5362
rect 3458 5334 3463 5362
rect 3537 5334 3542 5362
rect 3570 5334 4214 5362
rect 4242 5334 4247 5362
rect 1521 5278 1526 5306
rect 1554 5278 1806 5306
rect 1834 5278 1839 5306
rect 3201 5278 3206 5306
rect 3234 5278 3486 5306
rect 3514 5278 3519 5306
rect 1308 5082 1313 5110
rect 1341 5082 1365 5110
rect 1393 5082 1417 5110
rect 1445 5082 1450 5110
rect 2722 5082 2727 5110
rect 2755 5082 2779 5110
rect 2807 5082 2831 5110
rect 2859 5082 2864 5110
rect 4136 5082 4141 5110
rect 4169 5082 4193 5110
rect 4221 5082 4245 5110
rect 4273 5082 4278 5110
rect 5550 5082 5555 5110
rect 5583 5082 5607 5110
rect 5635 5082 5659 5110
rect 5687 5082 5692 5110
rect 1129 4998 1134 5026
rect 1162 4998 1414 5026
rect 1442 4998 1447 5026
rect 1185 4886 1190 4914
rect 1218 4886 1806 4914
rect 1834 4886 1839 4914
rect 3201 4830 3206 4858
rect 3234 4830 3486 4858
rect 3514 4830 3519 4858
rect 3145 4774 3150 4802
rect 3178 4774 3766 4802
rect 3794 4774 3799 4802
rect 2015 4690 2020 4718
rect 2048 4690 2072 4718
rect 2100 4690 2124 4718
rect 2152 4690 2157 4718
rect 3429 4690 3434 4718
rect 3462 4690 3486 4718
rect 3514 4690 3538 4718
rect 3566 4690 3571 4718
rect 4843 4690 4848 4718
rect 4876 4690 4900 4718
rect 4928 4690 4952 4718
rect 4980 4690 4985 4718
rect 6257 4690 6262 4718
rect 6290 4690 6314 4718
rect 6342 4690 6366 4718
rect 6394 4690 6399 4718
rect 2865 4606 2870 4634
rect 2898 4606 3486 4634
rect 3514 4606 3519 4634
rect 1017 4550 1022 4578
rect 1050 4550 1526 4578
rect 1554 4550 1559 4578
rect 2473 4494 2478 4522
rect 2506 4494 3430 4522
rect 3458 4494 3463 4522
rect 2417 4382 2422 4410
rect 2450 4382 3822 4410
rect 3850 4382 3855 4410
rect 1308 4298 1313 4326
rect 1341 4298 1365 4326
rect 1393 4298 1417 4326
rect 1445 4298 1450 4326
rect 2722 4298 2727 4326
rect 2755 4298 2779 4326
rect 2807 4298 2831 4326
rect 2859 4298 2864 4326
rect 4136 4298 4141 4326
rect 4169 4298 4193 4326
rect 4221 4298 4245 4326
rect 4273 4298 4278 4326
rect 5550 4298 5555 4326
rect 5583 4298 5607 4326
rect 5635 4298 5659 4326
rect 5687 4298 5692 4326
rect 2025 4214 2030 4242
rect 2058 4214 3878 4242
rect 3906 4214 3911 4242
rect 1073 4046 1078 4074
rect 1106 4046 3766 4074
rect 3794 4046 3799 4074
rect 0 4018 400 4032
rect 1078 4018 1106 4046
rect 0 3990 910 4018
rect 938 3990 1106 4018
rect 3033 3990 3038 4018
rect 3066 3990 3486 4018
rect 3514 3990 3519 4018
rect 0 3976 400 3990
rect 2015 3906 2020 3934
rect 2048 3906 2072 3934
rect 2100 3906 2124 3934
rect 2152 3906 2157 3934
rect 3429 3906 3434 3934
rect 3462 3906 3486 3934
rect 3514 3906 3538 3934
rect 3566 3906 3571 3934
rect 4843 3906 4848 3934
rect 4876 3906 4900 3934
rect 4928 3906 4952 3934
rect 4980 3906 4985 3934
rect 6257 3906 6262 3934
rect 6290 3906 6314 3934
rect 6342 3906 6366 3934
rect 6394 3906 6399 3934
rect 2697 3822 2702 3850
rect 2730 3822 3374 3850
rect 3402 3822 3407 3850
rect 4041 3710 4046 3738
rect 4074 3710 4326 3738
rect 4354 3710 4359 3738
rect 1185 3598 1190 3626
rect 1218 3598 3990 3626
rect 4018 3598 4023 3626
rect 1308 3514 1313 3542
rect 1341 3514 1365 3542
rect 1393 3514 1417 3542
rect 1445 3514 1450 3542
rect 2722 3514 2727 3542
rect 2755 3514 2779 3542
rect 2807 3514 2831 3542
rect 2859 3514 2864 3542
rect 4136 3514 4141 3542
rect 4169 3514 4193 3542
rect 4221 3514 4245 3542
rect 4273 3514 4278 3542
rect 5550 3514 5555 3542
rect 5583 3514 5607 3542
rect 5635 3514 5659 3542
rect 5687 3514 5692 3542
rect 3033 3374 3038 3402
rect 3066 3374 3654 3402
rect 3682 3374 3687 3402
rect 1633 3318 1638 3346
rect 1666 3318 2198 3346
rect 2226 3318 2231 3346
rect 4097 3318 4102 3346
rect 4130 3318 4382 3346
rect 4410 3318 4415 3346
rect 1465 3262 1470 3290
rect 1498 3262 1750 3290
rect 1778 3262 1783 3290
rect 2417 3262 2422 3290
rect 2450 3262 4046 3290
rect 4074 3262 4079 3290
rect 4657 3262 4662 3290
rect 4690 3262 6006 3290
rect 6034 3262 6039 3290
rect 3089 3206 3094 3234
rect 3122 3206 3654 3234
rect 3682 3206 3687 3234
rect 4713 3206 4718 3234
rect 4746 3206 5950 3234
rect 5978 3206 5983 3234
rect 2015 3122 2020 3150
rect 2048 3122 2072 3150
rect 2100 3122 2124 3150
rect 2152 3122 2157 3150
rect 3429 3122 3434 3150
rect 3462 3122 3486 3150
rect 3514 3122 3538 3150
rect 3566 3122 3571 3150
rect 4843 3122 4848 3150
rect 4876 3122 4900 3150
rect 4928 3122 4952 3150
rect 4980 3122 4985 3150
rect 6257 3122 6262 3150
rect 6290 3122 6314 3150
rect 6342 3122 6366 3150
rect 6394 3122 6399 3150
rect 1521 3038 1526 3066
rect 1554 3038 2310 3066
rect 2338 3038 2343 3066
rect 2753 2982 2758 3010
rect 2786 2982 3766 3010
rect 3794 2982 3799 3010
rect 2809 2926 2814 2954
rect 2842 2926 3430 2954
rect 3458 2926 3463 2954
rect 4153 2926 4158 2954
rect 4186 2926 4438 2954
rect 4466 2926 4471 2954
rect 4881 2926 4886 2954
rect 4914 2926 5166 2954
rect 5194 2926 5199 2954
rect 1353 2814 1358 2842
rect 1386 2814 1918 2842
rect 1946 2814 1951 2842
rect 5217 2814 5222 2842
rect 5250 2814 5894 2842
rect 5922 2814 5927 2842
rect 1308 2730 1313 2758
rect 1341 2730 1365 2758
rect 1393 2730 1417 2758
rect 1445 2730 1450 2758
rect 2722 2730 2727 2758
rect 2755 2730 2779 2758
rect 2807 2730 2831 2758
rect 2859 2730 2864 2758
rect 4136 2730 4141 2758
rect 4169 2730 4193 2758
rect 4221 2730 4245 2758
rect 4273 2730 4278 2758
rect 5550 2730 5555 2758
rect 5583 2730 5607 2758
rect 5635 2730 5659 2758
rect 5687 2730 5692 2758
rect 1633 2646 1638 2674
rect 1666 2646 1862 2674
rect 1890 2646 1895 2674
rect 3313 2646 3318 2674
rect 3346 2646 3822 2674
rect 3850 2646 3855 2674
rect 1577 2590 1582 2618
rect 1610 2590 2366 2618
rect 2394 2590 2399 2618
rect 3593 2590 3598 2618
rect 3626 2590 4214 2618
rect 4242 2590 4247 2618
rect 3257 2534 3262 2562
rect 3290 2534 3542 2562
rect 3570 2534 3575 2562
rect 3929 2534 3934 2562
rect 3962 2534 4270 2562
rect 4298 2534 4303 2562
rect 4937 2534 4942 2562
rect 4970 2534 5278 2562
rect 5306 2534 5311 2562
rect 1185 2478 1190 2506
rect 1218 2478 4046 2506
rect 4074 2478 4079 2506
rect 2921 2422 2926 2450
rect 2954 2422 3374 2450
rect 3402 2422 3407 2450
rect 3593 2422 3598 2450
rect 3626 2422 4774 2450
rect 4802 2422 4807 2450
rect 4993 2422 4998 2450
rect 5026 2422 5558 2450
rect 5586 2422 5591 2450
rect 2015 2338 2020 2366
rect 2048 2338 2072 2366
rect 2100 2338 2124 2366
rect 2152 2338 2157 2366
rect 3429 2338 3434 2366
rect 3462 2338 3486 2366
rect 3514 2338 3538 2366
rect 3566 2338 3571 2366
rect 4843 2338 4848 2366
rect 4876 2338 4900 2366
rect 4928 2338 4952 2366
rect 4980 2338 4985 2366
rect 6257 2338 6262 2366
rect 6290 2338 6314 2366
rect 6342 2338 6366 2366
rect 6394 2338 6399 2366
rect 2361 2254 2366 2282
rect 2394 2254 3990 2282
rect 4018 2254 4023 2282
rect 4601 2254 4606 2282
rect 4634 2254 5222 2282
rect 5250 2254 5255 2282
rect 1017 2198 1022 2226
rect 1050 2198 4550 2226
rect 4578 2198 4583 2226
rect 2641 2142 2646 2170
rect 2674 2142 3318 2170
rect 3346 2142 3351 2170
rect 3985 2142 3990 2170
rect 4018 2142 4270 2170
rect 4298 2142 4303 2170
rect 5609 2142 5614 2170
rect 5642 2142 5950 2170
rect 5978 2142 5983 2170
rect 1521 2086 1526 2114
rect 1554 2086 4886 2114
rect 4914 2086 4919 2114
rect 1745 2030 1750 2058
rect 1778 2030 4914 2058
rect 4886 2002 4914 2030
rect 4881 1974 4886 2002
rect 4914 1974 4919 2002
rect 1308 1946 1313 1974
rect 1341 1946 1365 1974
rect 1393 1946 1417 1974
rect 1445 1946 1450 1974
rect 2722 1946 2727 1974
rect 2755 1946 2779 1974
rect 2807 1946 2831 1974
rect 2859 1946 2864 1974
rect 4136 1946 4141 1974
rect 4169 1946 4193 1974
rect 4221 1946 4245 1974
rect 4273 1946 4278 1974
rect 5550 1946 5555 1974
rect 5583 1946 5607 1974
rect 5635 1946 5659 1974
rect 5687 1946 5692 1974
rect 1129 1862 1134 1890
rect 1162 1862 2030 1890
rect 2058 1862 2063 1890
rect 2646 1862 3598 1890
rect 3626 1862 3631 1890
rect 3873 1862 3878 1890
rect 3906 1862 4326 1890
rect 4354 1862 4359 1890
rect 2646 1834 2674 1862
rect 1073 1806 1078 1834
rect 1106 1806 2674 1834
rect 3145 1806 3150 1834
rect 3178 1806 4830 1834
rect 4858 1806 4863 1834
rect 3537 1750 3542 1778
rect 3570 1750 4214 1778
rect 4242 1750 4247 1778
rect 1409 1694 1414 1722
rect 1442 1694 1694 1722
rect 1722 1694 1727 1722
rect 3201 1694 3206 1722
rect 3234 1694 3486 1722
rect 3514 1694 3519 1722
rect 2015 1554 2020 1582
rect 2048 1554 2072 1582
rect 2100 1554 2124 1582
rect 2152 1554 2157 1582
rect 3429 1554 3434 1582
rect 3462 1554 3486 1582
rect 3514 1554 3538 1582
rect 3566 1554 3571 1582
rect 4843 1554 4848 1582
rect 4876 1554 4900 1582
rect 4928 1554 4952 1582
rect 4980 1554 4985 1582
rect 6257 1554 6262 1582
rect 6290 1554 6314 1582
rect 6342 1554 6366 1582
rect 6394 1554 6399 1582
<< via3 >>
rect 2020 6258 2048 6286
rect 2072 6258 2100 6286
rect 2124 6258 2152 6286
rect 3434 6258 3462 6286
rect 3486 6258 3514 6286
rect 3538 6258 3566 6286
rect 4848 6258 4876 6286
rect 4900 6258 4928 6286
rect 4952 6258 4980 6286
rect 6262 6258 6290 6286
rect 6314 6258 6342 6286
rect 6366 6258 6394 6286
rect 1313 5866 1341 5894
rect 1365 5866 1393 5894
rect 1417 5866 1445 5894
rect 2727 5866 2755 5894
rect 2779 5866 2807 5894
rect 2831 5866 2859 5894
rect 4141 5866 4169 5894
rect 4193 5866 4221 5894
rect 4245 5866 4273 5894
rect 5555 5866 5583 5894
rect 5607 5866 5635 5894
rect 5659 5866 5687 5894
rect 2020 5474 2048 5502
rect 2072 5474 2100 5502
rect 2124 5474 2152 5502
rect 3434 5474 3462 5502
rect 3486 5474 3514 5502
rect 3538 5474 3566 5502
rect 4848 5474 4876 5502
rect 4900 5474 4928 5502
rect 4952 5474 4980 5502
rect 6262 5474 6290 5502
rect 6314 5474 6342 5502
rect 6366 5474 6394 5502
rect 1313 5082 1341 5110
rect 1365 5082 1393 5110
rect 1417 5082 1445 5110
rect 2727 5082 2755 5110
rect 2779 5082 2807 5110
rect 2831 5082 2859 5110
rect 4141 5082 4169 5110
rect 4193 5082 4221 5110
rect 4245 5082 4273 5110
rect 5555 5082 5583 5110
rect 5607 5082 5635 5110
rect 5659 5082 5687 5110
rect 2020 4690 2048 4718
rect 2072 4690 2100 4718
rect 2124 4690 2152 4718
rect 3434 4690 3462 4718
rect 3486 4690 3514 4718
rect 3538 4690 3566 4718
rect 4848 4690 4876 4718
rect 4900 4690 4928 4718
rect 4952 4690 4980 4718
rect 6262 4690 6290 4718
rect 6314 4690 6342 4718
rect 6366 4690 6394 4718
rect 1313 4298 1341 4326
rect 1365 4298 1393 4326
rect 1417 4298 1445 4326
rect 2727 4298 2755 4326
rect 2779 4298 2807 4326
rect 2831 4298 2859 4326
rect 4141 4298 4169 4326
rect 4193 4298 4221 4326
rect 4245 4298 4273 4326
rect 5555 4298 5583 4326
rect 5607 4298 5635 4326
rect 5659 4298 5687 4326
rect 2020 3906 2048 3934
rect 2072 3906 2100 3934
rect 2124 3906 2152 3934
rect 3434 3906 3462 3934
rect 3486 3906 3514 3934
rect 3538 3906 3566 3934
rect 4848 3906 4876 3934
rect 4900 3906 4928 3934
rect 4952 3906 4980 3934
rect 6262 3906 6290 3934
rect 6314 3906 6342 3934
rect 6366 3906 6394 3934
rect 1313 3514 1341 3542
rect 1365 3514 1393 3542
rect 1417 3514 1445 3542
rect 2727 3514 2755 3542
rect 2779 3514 2807 3542
rect 2831 3514 2859 3542
rect 4141 3514 4169 3542
rect 4193 3514 4221 3542
rect 4245 3514 4273 3542
rect 5555 3514 5583 3542
rect 5607 3514 5635 3542
rect 5659 3514 5687 3542
rect 2020 3122 2048 3150
rect 2072 3122 2100 3150
rect 2124 3122 2152 3150
rect 3434 3122 3462 3150
rect 3486 3122 3514 3150
rect 3538 3122 3566 3150
rect 4848 3122 4876 3150
rect 4900 3122 4928 3150
rect 4952 3122 4980 3150
rect 6262 3122 6290 3150
rect 6314 3122 6342 3150
rect 6366 3122 6394 3150
rect 1313 2730 1341 2758
rect 1365 2730 1393 2758
rect 1417 2730 1445 2758
rect 2727 2730 2755 2758
rect 2779 2730 2807 2758
rect 2831 2730 2859 2758
rect 4141 2730 4169 2758
rect 4193 2730 4221 2758
rect 4245 2730 4273 2758
rect 5555 2730 5583 2758
rect 5607 2730 5635 2758
rect 5659 2730 5687 2758
rect 2020 2338 2048 2366
rect 2072 2338 2100 2366
rect 2124 2338 2152 2366
rect 3434 2338 3462 2366
rect 3486 2338 3514 2366
rect 3538 2338 3566 2366
rect 4848 2338 4876 2366
rect 4900 2338 4928 2366
rect 4952 2338 4980 2366
rect 6262 2338 6290 2366
rect 6314 2338 6342 2366
rect 6366 2338 6394 2366
rect 1313 1946 1341 1974
rect 1365 1946 1393 1974
rect 1417 1946 1445 1974
rect 2727 1946 2755 1974
rect 2779 1946 2807 1974
rect 2831 1946 2859 1974
rect 4141 1946 4169 1974
rect 4193 1946 4221 1974
rect 4245 1946 4273 1974
rect 5555 1946 5583 1974
rect 5607 1946 5635 1974
rect 5659 1946 5687 1974
rect 2020 1554 2048 1582
rect 2072 1554 2100 1582
rect 2124 1554 2152 1582
rect 3434 1554 3462 1582
rect 3486 1554 3514 1582
rect 3538 1554 3566 1582
rect 4848 1554 4876 1582
rect 4900 1554 4928 1582
rect 4952 1554 4980 1582
rect 6262 1554 6290 1582
rect 6314 1554 6342 1582
rect 6366 1554 6394 1582
<< metal4 >>
rect 1299 5894 1459 6302
rect 1299 5866 1313 5894
rect 1341 5866 1365 5894
rect 1393 5866 1417 5894
rect 1445 5866 1459 5894
rect 1299 5110 1459 5866
rect 1299 5082 1313 5110
rect 1341 5082 1365 5110
rect 1393 5082 1417 5110
rect 1445 5082 1459 5110
rect 1299 4326 1459 5082
rect 1299 4298 1313 4326
rect 1341 4298 1365 4326
rect 1393 4298 1417 4326
rect 1445 4298 1459 4326
rect 1299 3542 1459 4298
rect 1299 3514 1313 3542
rect 1341 3514 1365 3542
rect 1393 3514 1417 3542
rect 1445 3514 1459 3542
rect 1299 2758 1459 3514
rect 1299 2730 1313 2758
rect 1341 2730 1365 2758
rect 1393 2730 1417 2758
rect 1445 2730 1459 2758
rect 1299 1974 1459 2730
rect 1299 1946 1313 1974
rect 1341 1946 1365 1974
rect 1393 1946 1417 1974
rect 1445 1946 1459 1974
rect 1299 1538 1459 1946
rect 2006 6286 2166 6302
rect 2006 6258 2020 6286
rect 2048 6258 2072 6286
rect 2100 6258 2124 6286
rect 2152 6258 2166 6286
rect 2006 5502 2166 6258
rect 2006 5474 2020 5502
rect 2048 5474 2072 5502
rect 2100 5474 2124 5502
rect 2152 5474 2166 5502
rect 2006 4718 2166 5474
rect 2006 4690 2020 4718
rect 2048 4690 2072 4718
rect 2100 4690 2124 4718
rect 2152 4690 2166 4718
rect 2006 3934 2166 4690
rect 2006 3906 2020 3934
rect 2048 3906 2072 3934
rect 2100 3906 2124 3934
rect 2152 3906 2166 3934
rect 2006 3150 2166 3906
rect 2006 3122 2020 3150
rect 2048 3122 2072 3150
rect 2100 3122 2124 3150
rect 2152 3122 2166 3150
rect 2006 2366 2166 3122
rect 2006 2338 2020 2366
rect 2048 2338 2072 2366
rect 2100 2338 2124 2366
rect 2152 2338 2166 2366
rect 2006 1582 2166 2338
rect 2006 1554 2020 1582
rect 2048 1554 2072 1582
rect 2100 1554 2124 1582
rect 2152 1554 2166 1582
rect 2006 1538 2166 1554
rect 2713 5894 2873 6302
rect 2713 5866 2727 5894
rect 2755 5866 2779 5894
rect 2807 5866 2831 5894
rect 2859 5866 2873 5894
rect 2713 5110 2873 5866
rect 2713 5082 2727 5110
rect 2755 5082 2779 5110
rect 2807 5082 2831 5110
rect 2859 5082 2873 5110
rect 2713 4326 2873 5082
rect 2713 4298 2727 4326
rect 2755 4298 2779 4326
rect 2807 4298 2831 4326
rect 2859 4298 2873 4326
rect 2713 3542 2873 4298
rect 2713 3514 2727 3542
rect 2755 3514 2779 3542
rect 2807 3514 2831 3542
rect 2859 3514 2873 3542
rect 2713 2758 2873 3514
rect 2713 2730 2727 2758
rect 2755 2730 2779 2758
rect 2807 2730 2831 2758
rect 2859 2730 2873 2758
rect 2713 1974 2873 2730
rect 2713 1946 2727 1974
rect 2755 1946 2779 1974
rect 2807 1946 2831 1974
rect 2859 1946 2873 1974
rect 2713 1538 2873 1946
rect 3420 6286 3580 6302
rect 3420 6258 3434 6286
rect 3462 6258 3486 6286
rect 3514 6258 3538 6286
rect 3566 6258 3580 6286
rect 3420 5502 3580 6258
rect 3420 5474 3434 5502
rect 3462 5474 3486 5502
rect 3514 5474 3538 5502
rect 3566 5474 3580 5502
rect 3420 4718 3580 5474
rect 3420 4690 3434 4718
rect 3462 4690 3486 4718
rect 3514 4690 3538 4718
rect 3566 4690 3580 4718
rect 3420 3934 3580 4690
rect 3420 3906 3434 3934
rect 3462 3906 3486 3934
rect 3514 3906 3538 3934
rect 3566 3906 3580 3934
rect 3420 3150 3580 3906
rect 3420 3122 3434 3150
rect 3462 3122 3486 3150
rect 3514 3122 3538 3150
rect 3566 3122 3580 3150
rect 3420 2366 3580 3122
rect 3420 2338 3434 2366
rect 3462 2338 3486 2366
rect 3514 2338 3538 2366
rect 3566 2338 3580 2366
rect 3420 1582 3580 2338
rect 3420 1554 3434 1582
rect 3462 1554 3486 1582
rect 3514 1554 3538 1582
rect 3566 1554 3580 1582
rect 3420 1538 3580 1554
rect 4127 5894 4287 6302
rect 4127 5866 4141 5894
rect 4169 5866 4193 5894
rect 4221 5866 4245 5894
rect 4273 5866 4287 5894
rect 4127 5110 4287 5866
rect 4127 5082 4141 5110
rect 4169 5082 4193 5110
rect 4221 5082 4245 5110
rect 4273 5082 4287 5110
rect 4127 4326 4287 5082
rect 4127 4298 4141 4326
rect 4169 4298 4193 4326
rect 4221 4298 4245 4326
rect 4273 4298 4287 4326
rect 4127 3542 4287 4298
rect 4127 3514 4141 3542
rect 4169 3514 4193 3542
rect 4221 3514 4245 3542
rect 4273 3514 4287 3542
rect 4127 2758 4287 3514
rect 4127 2730 4141 2758
rect 4169 2730 4193 2758
rect 4221 2730 4245 2758
rect 4273 2730 4287 2758
rect 4127 1974 4287 2730
rect 4127 1946 4141 1974
rect 4169 1946 4193 1974
rect 4221 1946 4245 1974
rect 4273 1946 4287 1974
rect 4127 1538 4287 1946
rect 4834 6286 4994 6302
rect 4834 6258 4848 6286
rect 4876 6258 4900 6286
rect 4928 6258 4952 6286
rect 4980 6258 4994 6286
rect 4834 5502 4994 6258
rect 4834 5474 4848 5502
rect 4876 5474 4900 5502
rect 4928 5474 4952 5502
rect 4980 5474 4994 5502
rect 4834 4718 4994 5474
rect 4834 4690 4848 4718
rect 4876 4690 4900 4718
rect 4928 4690 4952 4718
rect 4980 4690 4994 4718
rect 4834 3934 4994 4690
rect 4834 3906 4848 3934
rect 4876 3906 4900 3934
rect 4928 3906 4952 3934
rect 4980 3906 4994 3934
rect 4834 3150 4994 3906
rect 4834 3122 4848 3150
rect 4876 3122 4900 3150
rect 4928 3122 4952 3150
rect 4980 3122 4994 3150
rect 4834 2366 4994 3122
rect 4834 2338 4848 2366
rect 4876 2338 4900 2366
rect 4928 2338 4952 2366
rect 4980 2338 4994 2366
rect 4834 1582 4994 2338
rect 4834 1554 4848 1582
rect 4876 1554 4900 1582
rect 4928 1554 4952 1582
rect 4980 1554 4994 1582
rect 4834 1538 4994 1554
rect 5541 5894 5701 6302
rect 5541 5866 5555 5894
rect 5583 5866 5607 5894
rect 5635 5866 5659 5894
rect 5687 5866 5701 5894
rect 5541 5110 5701 5866
rect 5541 5082 5555 5110
rect 5583 5082 5607 5110
rect 5635 5082 5659 5110
rect 5687 5082 5701 5110
rect 5541 4326 5701 5082
rect 5541 4298 5555 4326
rect 5583 4298 5607 4326
rect 5635 4298 5659 4326
rect 5687 4298 5701 4326
rect 5541 3542 5701 4298
rect 5541 3514 5555 3542
rect 5583 3514 5607 3542
rect 5635 3514 5659 3542
rect 5687 3514 5701 3542
rect 5541 2758 5701 3514
rect 5541 2730 5555 2758
rect 5583 2730 5607 2758
rect 5635 2730 5659 2758
rect 5687 2730 5701 2758
rect 5541 1974 5701 2730
rect 5541 1946 5555 1974
rect 5583 1946 5607 1974
rect 5635 1946 5659 1974
rect 5687 1946 5701 1974
rect 5541 1538 5701 1946
rect 6248 6286 6408 6302
rect 6248 6258 6262 6286
rect 6290 6258 6314 6286
rect 6342 6258 6366 6286
rect 6394 6258 6408 6286
rect 6248 5502 6408 6258
rect 6248 5474 6262 5502
rect 6290 5474 6314 5502
rect 6342 5474 6366 5502
rect 6394 5474 6408 5502
rect 6248 4718 6408 5474
rect 6248 4690 6262 4718
rect 6290 4690 6314 4718
rect 6342 4690 6366 4718
rect 6394 4690 6408 4718
rect 6248 3934 6408 4690
rect 6248 3906 6262 3934
rect 6290 3906 6314 3934
rect 6342 3906 6366 3934
rect 6394 3906 6408 3934
rect 6248 3150 6408 3906
rect 6248 3122 6262 3150
rect 6290 3122 6314 3150
rect 6342 3122 6366 3150
rect 6394 3122 6408 3150
rect 6248 2366 6408 3122
rect 6248 2338 6262 2366
rect 6290 2338 6314 2366
rect 6342 2338 6366 2366
rect 6394 2338 6408 2366
rect 6248 1582 6408 2338
rect 6248 1554 6262 1582
rect 6290 1554 6314 1582
rect 6342 1554 6366 1582
rect 6394 1554 6408 1582
rect 6248 1538 6408 1554
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 896 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9
timestamp 1667941163
transform 1 0 1176 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15
timestamp 1667941163
transform 1 0 1512 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21
timestamp 1667941163
transform 1 0 1848 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27
timestamp 1667941163
transform 1 0 2184 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33
timestamp 1667941163
transform 1 0 2520 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2744 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41
timestamp 1667941163
transform 1 0 2968 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47
timestamp 1667941163
transform 1 0 3304 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53
timestamp 1667941163
transform 1 0 3640 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59
timestamp 1667941163
transform 1 0 3976 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65
timestamp 1667941163
transform 1 0 4312 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 4536 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77
timestamp 1667941163
transform 1 0 4984 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83
timestamp 1667941163
transform 1 0 5320 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89
timestamp 1667941163
transform 1 0 5656 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95
timestamp 1667941163
transform 1 0 5992 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1667941163
transform 1 0 784 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_6
timestamp 1667941163
transform 1 0 1008 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_11
timestamp 1667941163
transform 1 0 1288 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_17
timestamp 1667941163
transform 1 0 1624 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_21
timestamp 1667941163
transform 1 0 1848 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_26
timestamp 1667941163
transform 1 0 2128 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_32
timestamp 1667941163
transform 1 0 2464 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_38
timestamp 1667941163
transform 1 0 2800 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_44
timestamp 1667941163
transform 1 0 3136 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_50
timestamp 1667941163
transform 1 0 3472 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 3696 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_56
timestamp 1667941163
transform 1 0 3808 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_61
timestamp 1667941163
transform 1 0 4088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_67
timestamp 1667941163
transform 1 0 4424 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_78
timestamp 1667941163
transform 1 0 5040 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_84
timestamp 1667941163
transform 1 0 5376 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_90
timestamp 1667941163
transform 1 0 5712 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_96
timestamp 1667941163
transform 1 0 6048 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_98
timestamp 1667941163
transform 1 0 6160 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_8
timestamp 1667941163
transform 1 0 1120 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_12
timestamp 1667941163
transform 1 0 1344 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_18
timestamp 1667941163
transform 1 0 1680 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_24
timestamp 1667941163
transform 1 0 2016 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_28
timestamp 1667941163
transform 1 0 2240 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1667941163
transform 1 0 2520 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_42
timestamp 1667941163
transform 1 0 3024 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_48
timestamp 1667941163
transform 1 0 3360 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_54
timestamp 1667941163
transform 1 0 3696 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_60
timestamp 1667941163
transform 1 0 4032 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_66
timestamp 1667941163
transform 1 0 4368 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_72
timestamp 1667941163
transform 1 0 4704 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_78
timestamp 1667941163
transform 1 0 5040 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_84
timestamp 1667941163
transform 1 0 5376 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_90
timestamp 1667941163
transform 1 0 5712 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_96
timestamp 1667941163
transform 1 0 6048 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_98
timestamp 1667941163
transform 1 0 6160 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_8
timestamp 1667941163
transform 1 0 1120 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_14
timestamp 1667941163
transform 1 0 1456 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_20
timestamp 1667941163
transform 1 0 1792 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_26
timestamp 1667941163
transform 1 0 2128 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_32
timestamp 1667941163
transform 1 0 2464 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_40
timestamp 1667941163
transform 1 0 2912 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_46
timestamp 1667941163
transform 1 0 3248 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_52
timestamp 1667941163
transform 1 0 3584 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_58
timestamp 1667941163
transform 1 0 3920 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_64
timestamp 1667941163
transform 1 0 4256 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_78
timestamp 1667941163
transform 1 0 5040 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_84 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 5376 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_92
timestamp 1667941163
transform 1 0 5824 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_96
timestamp 1667941163
transform 1 0 6048 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_98
timestamp 1667941163
transform 1 0 6160 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_10
timestamp 1667941163
transform 1 0 1232 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_16
timestamp 1667941163
transform 1 0 1568 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_22
timestamp 1667941163
transform 1 0 1904 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_30
timestamp 1667941163
transform 1 0 2352 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_39
timestamp 1667941163
transform 1 0 2856 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_44
timestamp 1667941163
transform 1 0 3136 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_50
timestamp 1667941163
transform 1 0 3472 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_56
timestamp 1667941163
transform 1 0 3808 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_62
timestamp 1667941163
transform 1 0 4144 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_68
timestamp 1667941163
transform 1 0 4480 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_74 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 4816 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_90
timestamp 1667941163
transform 1 0 5712 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_98
timestamp 1667941163
transform 1 0 6160 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_8
timestamp 1667941163
transform 1 0 1120 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_14
timestamp 1667941163
transform 1 0 1456 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_20
timestamp 1667941163
transform 1 0 1792 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_26
timestamp 1667941163
transform 1 0 2128 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_32
timestamp 1667941163
transform 1 0 2464 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_38
timestamp 1667941163
transform 1 0 2800 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_44
timestamp 1667941163
transform 1 0 3136 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_50
timestamp 1667941163
transform 1 0 3472 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_56
timestamp 1667941163
transform 1 0 3808 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_62
timestamp 1667941163
transform 1 0 4144 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_68
timestamp 1667941163
transform 1 0 4480 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_89
timestamp 1667941163
transform 1 0 5656 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_97
timestamp 1667941163
transform 1 0 6104 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_9
timestamp 1667941163
transform 1 0 1176 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_13
timestamp 1667941163
transform 1 0 1400 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_18
timestamp 1667941163
transform 1 0 1680 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 2128 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_32
timestamp 1667941163
transform 1 0 2464 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_41
timestamp 1667941163
transform 1 0 2968 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_46
timestamp 1667941163
transform 1 0 3248 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_52
timestamp 1667941163
transform 1 0 3584 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_58
timestamp 1667941163
transform 1 0 3920 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_64 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 4256 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_96
timestamp 1667941163
transform 1 0 6048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_98
timestamp 1667941163
transform 1 0 6160 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_2
timestamp 1667941163
transform 1 0 784 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_6
timestamp 1667941163
transform 1 0 1008 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_11
timestamp 1667941163
transform 1 0 1288 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_17
timestamp 1667941163
transform 1 0 1624 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_23
timestamp 1667941163
transform 1 0 1960 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_29
timestamp 1667941163
transform 1 0 2296 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_35
timestamp 1667941163
transform 1 0 2632 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_41
timestamp 1667941163
transform 1 0 2968 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_47
timestamp 1667941163
transform 1 0 3304 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_53
timestamp 1667941163
transform 1 0 3640 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_59
timestamp 1667941163
transform 1 0 3976 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_67
timestamp 1667941163
transform 1 0 4424 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1667941163
transform 1 0 4760 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_89
timestamp 1667941163
transform 1 0 5656 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_97
timestamp 1667941163
transform 1 0 6104 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_2
timestamp 1667941163
transform 1 0 784 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_10
timestamp 1667941163
transform 1 0 1232 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_16
timestamp 1667941163
transform 1 0 1568 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_22
timestamp 1667941163
transform 1 0 1904 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_28
timestamp 1667941163
transform 1 0 2240 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_37
timestamp 1667941163
transform 1 0 2744 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_41
timestamp 1667941163
transform 1 0 2968 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_46
timestamp 1667941163
transform 1 0 3248 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_52
timestamp 1667941163
transform 1 0 3584 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_58
timestamp 1667941163
transform 1 0 3920 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_90
timestamp 1667941163
transform 1 0 5712 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_98
timestamp 1667941163
transform 1 0 6160 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_2
timestamp 1667941163
transform 1 0 784 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_6
timestamp 1667941163
transform 1 0 1008 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_11
timestamp 1667941163
transform 1 0 1288 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_17
timestamp 1667941163
transform 1 0 1624 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_23
timestamp 1667941163
transform 1 0 1960 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_29
timestamp 1667941163
transform 1 0 2296 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_35
timestamp 1667941163
transform 1 0 2632 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_41
timestamp 1667941163
transform 1 0 2968 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_47
timestamp 1667941163
transform 1 0 3304 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_53
timestamp 1667941163
transform 1 0 3640 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_59
timestamp 1667941163
transform 1 0 3976 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_65
timestamp 1667941163
transform 1 0 4312 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_69
timestamp 1667941163
transform 1 0 4536 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_73
timestamp 1667941163
transform 1 0 4760 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_89
timestamp 1667941163
transform 1 0 5656 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_97
timestamp 1667941163
transform 1 0 6104 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_2
timestamp 1667941163
transform 1 0 784 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_10
timestamp 1667941163
transform 1 0 1232 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_16
timestamp 1667941163
transform 1 0 1568 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_22
timestamp 1667941163
transform 1 0 1904 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_28
timestamp 1667941163
transform 1 0 2240 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 2576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_37
timestamp 1667941163
transform 1 0 2744 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_45
timestamp 1667941163
transform 1 0 3192 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_51
timestamp 1667941163
transform 1 0 3528 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_55
timestamp 1667941163
transform 1 0 3752 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_61
timestamp 1667941163
transform 1 0 4088 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_67
timestamp 1667941163
transform 1 0 4424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1667941163
transform 1 0 784 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_10
timestamp 1667941163
transform 1 0 1232 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_16
timestamp 1667941163
transform 1 0 1568 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_22
timestamp 1667941163
transform 1 0 1904 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_28
timestamp 1667941163
transform 1 0 2240 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_34
timestamp 1667941163
transform 1 0 2576 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_37
timestamp 1667941163
transform 1 0 2744 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_43
timestamp 1667941163
transform 1 0 3080 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_49
timestamp 1667941163
transform 1 0 3416 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_55
timestamp 1667941163
transform 1 0 3752 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_61
timestamp 1667941163
transform 1 0 4088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_67
timestamp 1667941163
transform 1 0 4424 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1667941163
transform 1 0 4536 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_72
timestamp 1667941163
transform 1 0 4704 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_88
timestamp 1667941163
transform 1 0 5600 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_96
timestamp 1667941163
transform 1 0 6048 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_98
timestamp 1667941163
transform 1 0 6160 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 6328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 6328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 6328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 6328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 6328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 6328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 6328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 6328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 6328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 6328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 6328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 6328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1667941163
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1667941163
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1667941163
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1667941163
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1667941163
transform 1 0 2632 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1667941163
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0_ pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 1176 0 1 3920
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[0\].u_uinv pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 4480 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[1\].u_uinv
timestamp 1667941163
transform -1 0 4480 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[2\].u_uinv
timestamp 1667941163
transform -1 0 4144 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[3\].u_uinv
timestamp 1667941163
transform 1 0 1400 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[4\].u_uinv
timestamp 1667941163
transform -1 0 1680 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[5\].u_uinv
timestamp 1667941163
transform 1 0 1232 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[6\].u_uinv
timestamp 1667941163
transform -1 0 2016 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[7\].u_uinv
timestamp 1667941163
transform 1 0 1568 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[8\].u_uinv
timestamp 1667941163
transform 1 0 1904 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[9\].u_uinv
timestamp 1667941163
transform -1 0 2464 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[10\].u_uinv
timestamp 1667941163
transform 1 0 1232 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[11\].u_uinv
timestamp 1667941163
transform 1 0 2296 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[12\].u_uinv
timestamp 1667941163
transform -1 0 4144 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[13\].u_uinv
timestamp 1667941163
transform -1 0 2464 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[14\].u_uinv
timestamp 1667941163
transform 1 0 1904 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[15\].u_uinv
timestamp 1667941163
transform -1 0 2520 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[16\].u_uinv
timestamp 1667941163
transform -1 0 2184 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[17\].u_uinv
timestamp 1667941163
transform 1 0 1064 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[18\].u_uinv
timestamp 1667941163
transform 1 0 4032 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[19\].u_uinv
timestamp 1667941163
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[20\].u_uinv
timestamp 1667941163
transform 1 0 4816 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[21\].u_uinv
timestamp 1667941163
transform -1 0 5376 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[22\].u_uinv
timestamp 1667941163
transform 1 0 4816 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[23\].u_uinv
timestamp 1667941163
transform 1 0 5488 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[24\].u_uinv
timestamp 1667941163
transform -1 0 6048 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[25\].u_uinv
timestamp 1667941163
transform 1 0 4592 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[26\].u_uinv
timestamp 1667941163
transform -1 0 6048 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[27\].u_uinv
timestamp 1667941163
transform 1 0 5152 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[28\].u_uinv
timestamp 1667941163
transform 1 0 5488 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[29\].u_uinv
timestamp 1667941163
transform -1 0 5992 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[30\].u_uinv
timestamp 1667941163
transform -1 0 5656 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[31\].u_uinv
timestamp 1667941163
transform 1 0 5096 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[32\].u_uinv
timestamp 1667941163
transform -1 0 5376 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[33\].u_uinv
timestamp 1667941163
transform -1 0 4704 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[34\].u_uinv
timestamp 1667941163
transform 1 0 952 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[35\].u_uinv
timestamp 1667941163
transform -1 0 5040 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[36\].u_uinv
timestamp 1667941163
transform 1 0 1288 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[37\].u_uinv
timestamp 1667941163
transform 1 0 1624 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[38\].u_uinv
timestamp 1667941163
transform -1 0 4984 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[39\].u_uinv
timestamp 1667941163
transform 1 0 3080 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[40\].u_uinv
timestamp 1667941163
transform 1 0 3416 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[41\].u_uinv
timestamp 1667941163
transform -1 0 4312 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[42\].u_uinv
timestamp 1667941163
transform 1 0 3752 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[43\].u_uinv
timestamp 1667941163
transform -1 0 4424 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[44\].u_uinv
timestamp 1667941163
transform -1 0 4088 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[45\].u_uinv
timestamp 1667941163
transform 1 0 3808 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[46\].u_uinv
timestamp 1667941163
transform -1 0 4368 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[47\].u_uinv
timestamp 1667941163
transform -1 0 3696 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[48\].u_uinv
timestamp 1667941163
transform -1 0 3360 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[49\].u_uinv
timestamp 1667941163
transform 1 0 2800 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[50\].u_uinv
timestamp 1667941163
transform -1 0 3472 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[51\].u_uinv
timestamp 1667941163
transform 1 0 2576 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[52\].u_uinv
timestamp 1667941163
transform 1 0 2912 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[53\].u_uinv
timestamp 1667941163
transform -1 0 3920 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[54\].u_uinv
timestamp 1667941163
transform 1 0 2688 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[55\].u_uinv
timestamp 1667941163
transform 1 0 3360 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[56\].u_uinv
timestamp 1667941163
transform -1 0 3808 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[57\].u_uinv
timestamp 1667941163
transform 1 0 3024 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[58\].u_uinv
timestamp 1667941163
transform 1 0 3248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[59\].u_uinv
timestamp 1667941163
transform -1 0 3808 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[60\].u_uinv
timestamp 1667941163
transform -1 0 3136 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[61\].u_uinv
timestamp 1667941163
transform 1 0 2576 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[62\].u_uinv
timestamp 1667941163
transform -1 0 3472 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[63\].u_uinv
timestamp 1667941163
transform 1 0 2912 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[64\].u_uinv
timestamp 1667941163
transform -1 0 3584 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[65\].u_uinv
timestamp 1667941163
transform 1 0 2408 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[66\].u_uinv
timestamp 1667941163
transform -1 0 3248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[67\].u_uinv
timestamp 1667941163
transform 1 0 2744 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[68\].u_uinv
timestamp 1667941163
transform 1 0 3416 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[69\].u_uinv
timestamp 1667941163
transform -1 0 3920 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[70\].u_uinv
timestamp 1667941163
transform 1 0 3080 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[71\].u_uinv
timestamp 1667941163
transform -1 0 3584 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[72\].u_uinv
timestamp 1667941163
transform 1 0 2408 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[73\].u_uinv
timestamp 1667941163
transform -1 0 3248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[74\].u_uinv
timestamp 1667941163
transform 1 0 2744 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[75\].u_uinv
timestamp 1667941163
transform 1 0 3080 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[76\].u_uinv
timestamp 1667941163
transform 1 0 3416 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[77\].u_uinv
timestamp 1667941163
transform -1 0 4312 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[78\].u_uinv
timestamp 1667941163
transform 1 0 3752 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[79\].u_uinv
timestamp 1667941163
transform -1 0 4424 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[80\].u_uinv
timestamp 1667941163
transform -1 0 4088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[81\].u_uinv
timestamp 1667941163
transform 1 0 3864 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[82\].u_uinv
timestamp 1667941163
transform -1 0 4424 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[83\].u_uinv
timestamp 1667941163
transform -1 0 3752 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[84\].u_uinv
timestamp 1667941163
transform 1 0 3192 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[85\].u_uinv
timestamp 1667941163
transform -1 0 3528 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[86\].u_uinv
timestamp 1667941163
transform 1 0 2856 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[87\].u_uinv
timestamp 1667941163
transform -1 0 3192 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[88\].u_uinv
timestamp 1667941163
transform -1 0 2576 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[89\].u_uinv
timestamp 1667941163
transform 1 0 2016 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[90\].u_uinv
timestamp 1667941163
transform -1 0 2576 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[91\].u_uinv
timestamp 1667941163
transform 1 0 1680 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[92\].u_uinv
timestamp 1667941163
transform -1 0 2240 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[93\].u_uinv
timestamp 1667941163
transform 1 0 1344 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[94\].u_uinv
timestamp 1667941163
transform -1 0 1904 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[95\].u_uinv
timestamp 1667941163
transform -1 0 1232 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[96\].u_uinv
timestamp 1667941163
transform 1 0 1008 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[97\].u_uinv
timestamp 1667941163
transform -1 0 1624 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[98\].u_uinv
timestamp 1667941163
transform 1 0 1064 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[99\].u_uinv
timestamp 1667941163
transform -1 0 1568 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[100\].u_uinv
timestamp 1667941163
transform 1 0 1008 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[101\].u_uinv
timestamp 1667941163
transform -1 0 1680 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[102\].u_uinv
timestamp 1667941163
transform -1 0 1568 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[103\].u_uinv
timestamp 1667941163
transform 1 0 1064 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[104\].u_uinv
timestamp 1667941163
transform -1 0 1904 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[105\].u_uinv
timestamp 1667941163
transform 1 0 1400 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[106\].u_uinv
timestamp 1667941163
transform 1 0 1736 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[107\].u_uinv
timestamp 1667941163
transform 1 0 2072 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[108\].u_uinv
timestamp 1667941163
transform -1 0 2576 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[109\].u_uinv
timestamp 1667941163
transform 1 0 2016 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[110\].u_uinv
timestamp 1667941163
transform 1 0 2072 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[111\].u_uinv
timestamp 1667941163
transform -1 0 2464 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[112\].u_uinv
timestamp 1667941163
transform 1 0 1736 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[113\].u_uinv
timestamp 1667941163
transform 1 0 1904 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[114\].u_uinv
timestamp 1667941163
transform -1 0 3976 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[115\].u_uinv
timestamp 1667941163
transform -1 0 2464 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[116\].u_uinv
timestamp 1667941163
transform 1 0 1904 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[117\].u_uinv
timestamp 1667941163
transform -1 0 2352 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[118\].u_uinv
timestamp 1667941163
transform 1 0 1568 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[119\].u_uinv
timestamp 1667941163
transform -1 0 1904 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[120\].u_uinv
timestamp 1667941163
transform -1 0 1568 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[121\].u_uinv
timestamp 1667941163
transform 1 0 896 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[122\].u_uinv
timestamp 1667941163
transform -1 0 1232 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[123\].u_uinv
timestamp 1667941163
transform -1 0 1120 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[124\].u_uinv
timestamp 1667941163
transform -1 0 1120 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gen_ring\[125\].u_uinv
timestamp 1667941163
transform 1 0 3696 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_uinv_init
timestamp 1667941163
transform 1 0 4032 0 1 3920
box -43 -43 267 435
<< labels >>
flabel metal3 s 0 3976 400 4032 0 FreeSans 224 0 0 0 Y
port 0 nsew signal tristate
flabel metal4 s 1299 1538 1459 6302 0 FreeSans 640 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 2713 1538 2873 6302 0 FreeSans 640 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 4127 1538 4287 6302 0 FreeSans 640 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 5541 1538 5701 6302 0 FreeSans 640 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 2006 1538 2166 6302 0 FreeSans 640 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 3420 1538 3580 6302 0 FreeSans 640 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 4834 1538 4994 6302 0 FreeSans 640 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 6248 1538 6408 6302 0 FreeSans 640 90 0 0 vss
port 2 nsew ground bidirectional
rlabel metal1 3500 5880 3500 5880 0 vdd
rlabel via1 3540 6272 3540 6272 0 vss
rlabel metal3 2436 4060 2436 4060 0 Y
rlabel metal2 4116 3360 4116 3360 0 con\[0\]
rlabel metal2 1092 5152 1092 5152 0 con\[100\]
rlabel metal2 1540 4116 1540 4116 0 con\[101\]
rlabel metal2 1568 4228 1568 4228 0 con\[102\]
rlabel metal3 1288 5012 1288 5012 0 con\[103\]
rlabel metal3 1512 4900 1512 4900 0 con\[104\]
rlabel metal2 1708 5012 1708 5012 0 con\[105\]
rlabel metal3 1680 5292 1680 5292 0 con\[106\]
rlabel metal2 2016 5292 2016 5292 0 con\[107\]
rlabel metal2 2492 5040 2492 5040 0 con\[108\]
rlabel metal2 2268 4900 2268 4900 0 con\[109\]
rlabel metal3 1932 3052 1932 3052 0 con\[10\]
rlabel metal2 2184 4564 2184 4564 0 con\[110\]
rlabel metal2 2296 4396 2296 4396 0 con\[111\]
rlabel metal2 2212 4228 2212 4228 0 con\[112\]
rlabel metal2 1932 4116 1932 4116 0 con\[113\]
rlabel metal3 2968 4228 2968 4228 0 con\[114\]
rlabel metal2 2408 3780 2408 3780 0 con\[115\]
rlabel metal2 2156 3724 2156 3724 0 con\[116\]
rlabel metal2 2268 3472 2268 3472 0 con\[117\]
rlabel metal3 1932 3332 1932 3332 0 con\[118\]
rlabel metal2 1820 3472 1820 3472 0 con\[119\]
rlabel metal2 2380 2576 2380 2576 0 con\[11\]
rlabel metal3 1624 3276 1624 3276 0 con\[120\]
rlabel metal2 1344 3444 1344 3444 0 con\[121\]
rlabel metal2 1148 3472 1148 3472 0 con\[122\]
rlabel metal2 1064 2996 1064 2996 0 con\[123\]
rlabel metal2 1008 2548 1008 2548 0 con\[124\]
rlabel metal2 3976 4060 3976 4060 0 con\[126\]
rlabel metal2 2436 2968 2436 2968 0 con\[12\]
rlabel metal2 2380 2240 2380 2240 0 con\[13\]
rlabel metal2 2156 2156 2156 2156 0 con\[14\]
rlabel metal2 2436 1904 2436 1904 0 con\[15\]
rlabel metal2 2240 1708 2240 1708 0 con\[16\]
rlabel metal3 1596 1876 1596 1876 0 con\[17\]
rlabel metal2 1204 2380 1204 2380 0 con\[18\]
rlabel metal3 4312 2940 4312 2940 0 con\[19\]
rlabel metal2 4368 3444 4368 3444 0 con\[1\]
rlabel metal2 4900 2688 4900 2688 0 con\[20\]
rlabel metal3 5124 2548 5124 2548 0 con\[21\]
rlabel metal2 5208 2660 5208 2660 0 con\[22\]
rlabel metal2 5572 2324 5572 2324 0 con\[23\]
rlabel metal3 5796 2156 5796 2156 0 con\[24\]
rlabel metal2 5964 2268 5964 2268 0 con\[25\]
rlabel metal2 5964 2884 5964 2884 0 con\[26\]
rlabel metal2 5908 2744 5908 2744 0 con\[27\]
rlabel metal2 5572 2604 5572 2604 0 con\[28\]
rlabel metal2 5908 1848 5908 1848 0 con\[29\]
rlabel metal3 4200 3724 4200 3724 0 con\[2\]
rlabel metal2 5712 1708 5712 1708 0 con\[30\]
rlabel metal2 5348 1764 5348 1764 0 con\[31\]
rlabel metal2 5264 1876 5264 1876 0 con\[32\]
rlabel metal3 4928 2268 4928 2268 0 con\[33\]
rlabel metal2 1036 1988 1036 1988 0 con\[34\]
rlabel metal3 1876 1820 1876 1820 0 con\[35\]
rlabel metal2 1372 1820 1372 1820 0 con\[36\]
rlabel metal3 1568 1708 1568 1708 0 con\[37\]
rlabel metal2 1764 1960 1764 1960 0 con\[38\]
rlabel metal2 3164 1792 3164 1792 0 con\[39\]
rlabel metal2 1484 2436 1484 2436 0 con\[3\]
rlabel metal3 3360 1708 3360 1708 0 con\[40\]
rlabel metal3 3892 1764 3892 1764 0 con\[41\]
rlabel metal2 4004 1764 4004 1764 0 con\[42\]
rlabel metal2 4340 2016 4340 2016 0 con\[43\]
rlabel metal3 4144 2156 4144 2156 0 con\[44\]
rlabel metal2 3920 2268 3920 2268 0 con\[45\]
rlabel metal3 4116 2548 4116 2548 0 con\[46\]
rlabel metal2 3612 2576 3612 2576 0 con\[47\]
rlabel metal3 3416 2548 3416 2548 0 con\[48\]
rlabel metal2 3052 2548 3052 2548 0 con\[49\]
rlabel metal2 1568 2268 1568 2268 0 con\[4\]
rlabel metal2 3388 2324 3388 2324 0 con\[50\]
rlabel metal3 2996 2156 2996 2156 0 con\[51\]
rlabel metal2 2856 2156 2856 2156 0 con\[52\]
rlabel metal2 3052 2352 3052 2352 0 con\[53\]
rlabel metal3 3276 2996 3276 2996 0 con\[54\]
rlabel metal3 3136 2940 3136 2940 0 con\[55\]
rlabel metal2 3612 3052 3612 3052 0 con\[56\]
rlabel metal2 3108 3108 3108 3108 0 con\[57\]
rlabel metal2 3164 3164 3164 3164 0 con\[58\]
rlabel metal2 3416 3444 3416 3444 0 con\[59\]
rlabel metal2 1540 2800 1540 2800 0 con\[5\]
rlabel metal2 3052 3360 3052 3360 0 con\[60\]
rlabel metal2 2968 3444 2968 3444 0 con\[61\]
rlabel metal2 3388 3808 3388 3808 0 con\[62\]
rlabel metal2 3164 3724 3164 3724 0 con\[63\]
rlabel metal2 3052 3920 3052 3920 0 con\[64\]
rlabel metal3 2968 4508 2968 4508 0 con\[65\]
rlabel metal2 3108 4116 3108 4116 0 con\[66\]
rlabel metal2 3108 4368 3108 4368 0 con\[67\]
rlabel metal2 3500 4592 3500 4592 0 con\[68\]
rlabel metal2 3584 4620 3584 4620 0 con\[69\]
rlabel metal2 1932 2688 1932 2688 0 con\[6\]
rlabel metal2 3164 4676 3164 4676 0 con\[70\]
rlabel metal2 3220 4732 3220 4732 0 con\[71\]
rlabel metal2 3444 5180 3444 5180 0 con\[72\]
rlabel metal2 3108 4900 3108 4900 0 con\[73\]
rlabel metal2 3108 5096 3108 5096 0 con\[74\]
rlabel metal2 3024 5292 3024 5292 0 con\[75\]
rlabel metal3 3360 5292 3360 5292 0 con\[76\]
rlabel metal3 3892 5348 3892 5348 0 con\[77\]
rlabel metal2 4004 5292 4004 5292 0 con\[78\]
rlabel metal2 4340 5516 4340 5516 0 con\[79\]
rlabel metal3 1764 2660 1764 2660 0 con\[7\]
rlabel metal3 4144 5628 4144 5628 0 con\[80\]
rlabel metal2 3948 5936 3948 5936 0 con\[81\]
rlabel metal3 4172 6076 4172 6076 0 con\[82\]
rlabel metal3 3976 6132 3976 6132 0 con\[83\]
rlabel metal3 3444 6076 3444 6076 0 con\[84\]
rlabel metal2 3388 5684 3388 5684 0 con\[85\]
rlabel metal2 3388 5964 3388 5964 0 con\[86\]
rlabel metal2 3108 5824 3108 5824 0 con\[87\]
rlabel metal2 3052 5824 3052 5824 0 con\[88\]
rlabel metal2 2268 6076 2268 6076 0 con\[89\]
rlabel metal2 1848 2940 1848 2940 0 con\[8\]
rlabel metal2 2492 5824 2492 5824 0 con\[90\]
rlabel metal3 2156 5796 2156 5796 0 con\[91\]
rlabel metal2 2128 5684 2128 5684 0 con\[92\]
rlabel metal2 2072 5572 2072 5572 0 con\[93\]
rlabel metal2 1792 5684 1792 5684 0 con\[94\]
rlabel metal2 1736 5572 1736 5572 0 con\[95\]
rlabel metal2 1092 5824 1092 5824 0 con\[96\]
rlabel metal3 1288 4564 1288 4564 0 con\[97\]
rlabel metal2 1316 4508 1316 4508 0 con\[98\]
rlabel metal2 1232 4620 1232 4620 0 con\[99\]
rlabel metal2 2212 2940 2212 2940 0 con\[9\]
<< properties >>
string FIXED_BBOX 0 0 7000 8000
<< end >>
