// This is the unpowered netlist.
module shiftreg (latch,
    sclk,
    sdin,
    sr_out,
    tune_s1_series_gy,
    tune_s1_series_gygy,
    tune_s1_shunt,
    tune_s1_shunt_gy,
    tune_s2_series_gy,
    tune_s2_series_gygy,
    tune_s2_shunt,
    tune_s2_shunt_gy);
 input latch;
 input sclk;
 input sdin;
 output sr_out;
 output [5:0] tune_s1_series_gy;
 output [5:0] tune_s1_series_gygy;
 output [7:0] tune_s1_shunt;
 output [6:0] tune_s1_shunt_gy;
 output [7:0] tune_s2_series_gy;
 output [7:0] tune_s2_series_gygy;
 output [10:0] tune_s2_shunt;
 output [4:0] tune_s2_shunt_gy;

 wire \sr[0] ;
 wire \sr[10] ;
 wire \sr[11] ;
 wire \sr[12] ;
 wire \sr[13] ;
 wire \sr[14] ;
 wire \sr[15] ;
 wire \sr[16] ;
 wire \sr[17] ;
 wire \sr[18] ;
 wire \sr[19] ;
 wire \sr[1] ;
 wire \sr[20] ;
 wire \sr[21] ;
 wire \sr[22] ;
 wire \sr[23] ;
 wire \sr[24] ;
 wire \sr[25] ;
 wire \sr[26] ;
 wire \sr[27] ;
 wire \sr[28] ;
 wire \sr[29] ;
 wire \sr[2] ;
 wire \sr[30] ;
 wire \sr[31] ;
 wire \sr[32] ;
 wire \sr[33] ;
 wire \sr[34] ;
 wire \sr[35] ;
 wire \sr[36] ;
 wire \sr[37] ;
 wire \sr[38] ;
 wire \sr[39] ;
 wire \sr[3] ;
 wire \sr[40] ;
 wire \sr[41] ;
 wire \sr[42] ;
 wire \sr[43] ;
 wire \sr[44] ;
 wire \sr[45] ;
 wire \sr[46] ;
 wire \sr[47] ;
 wire \sr[48] ;
 wire \sr[49] ;
 wire \sr[4] ;
 wire \sr[50] ;
 wire \sr[51] ;
 wire \sr[52] ;
 wire \sr[53] ;
 wire \sr[54] ;
 wire \sr[55] ;
 wire \sr[56] ;
 wire \sr[57] ;
 wire \sr[5] ;
 wire \sr[6] ;
 wire \sr[7] ;
 wire \sr[8] ;
 wire \sr[9] ;
 wire clknet_0_sclk;
 wire clknet_3_0__leaf_sclk;
 wire clknet_3_1__leaf_sclk;
 wire clknet_3_2__leaf_sclk;
 wire clknet_3_3__leaf_sclk;
 wire clknet_3_4__leaf_sclk;
 wire clknet_3_5__leaf_sclk;
 wire clknet_3_6__leaf_sclk;
 wire clknet_3_7__leaf_sclk;

 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _000_ (.D(\sr[18] ),
    .CLK(latch),
    .Q(tune_s1_series_gy[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _001_ (.D(\sr[19] ),
    .CLK(latch),
    .Q(tune_s1_series_gy[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _002_ (.D(\sr[20] ),
    .CLK(latch),
    .Q(tune_s1_series_gy[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _003_ (.D(\sr[21] ),
    .CLK(latch),
    .Q(tune_s1_series_gygy[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _004_ (.D(\sr[22] ),
    .CLK(latch),
    .Q(tune_s1_series_gygy[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _005_ (.D(\sr[23] ),
    .CLK(latch),
    .Q(tune_s1_series_gygy[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _006_ (.D(\sr[24] ),
    .CLK(latch),
    .Q(tune_s1_series_gygy[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _007_ (.D(\sr[25] ),
    .CLK(latch),
    .Q(tune_s1_series_gygy[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _008_ (.D(\sr[26] ),
    .CLK(latch),
    .Q(tune_s1_series_gygy[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _009_ (.D(\sr[27] ),
    .CLK(latch),
    .Q(tune_s2_shunt[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _010_ (.D(\sr[28] ),
    .CLK(latch),
    .Q(tune_s2_shunt[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _011_ (.D(\sr[29] ),
    .CLK(latch),
    .Q(tune_s2_shunt[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _012_ (.D(\sr[30] ),
    .CLK(latch),
    .Q(tune_s2_shunt[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _013_ (.D(\sr[31] ),
    .CLK(latch),
    .Q(tune_s2_shunt[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _014_ (.D(\sr[32] ),
    .CLK(latch),
    .Q(tune_s2_shunt[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _015_ (.D(\sr[33] ),
    .CLK(latch),
    .Q(tune_s2_shunt[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _016_ (.D(\sr[34] ),
    .CLK(latch),
    .Q(tune_s2_shunt[7]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _017_ (.D(\sr[35] ),
    .CLK(latch),
    .Q(tune_s2_shunt[8]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _018_ (.D(\sr[36] ),
    .CLK(latch),
    .Q(tune_s2_shunt[9]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _019_ (.D(\sr[37] ),
    .CLK(latch),
    .Q(tune_s2_shunt[10]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _020_ (.D(\sr[38] ),
    .CLK(latch),
    .Q(tune_s2_shunt_gy[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _021_ (.D(\sr[39] ),
    .CLK(latch),
    .Q(tune_s2_shunt_gy[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _022_ (.D(\sr[40] ),
    .CLK(latch),
    .Q(tune_s2_shunt_gy[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _023_ (.D(\sr[41] ),
    .CLK(latch),
    .Q(tune_s2_shunt_gy[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _024_ (.D(\sr[42] ),
    .CLK(latch),
    .Q(tune_s2_shunt_gy[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _025_ (.D(\sr[43] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _026_ (.D(\sr[44] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _027_ (.D(\sr[45] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _028_ (.D(\sr[46] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _029_ (.D(\sr[47] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _030_ (.D(\sr[48] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _031_ (.D(\sr[49] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _032_ (.D(\sr[50] ),
    .CLK(latch),
    .Q(tune_s2_series_gy[7]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _033_ (.D(\sr[51] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _034_ (.D(\sr[52] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _035_ (.D(\sr[53] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _036_ (.D(\sr[54] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _037_ (.D(\sr[55] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _038_ (.D(\sr[56] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _039_ (.D(\sr[57] ),
    .CLK(latch),
    .Q(tune_s2_series_gygy[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _040_ (.D(sr_out),
    .CLK(latch),
    .Q(tune_s2_series_gygy[7]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _041_ (.D(sdin),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _042_ (.D(\sr[0] ),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _043_ (.D(\sr[1] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _044_ (.D(\sr[2] ),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _045_ (.D(\sr[3] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _046_ (.D(\sr[4] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _047_ (.D(\sr[5] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _048_ (.D(\sr[6] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _049_ (.D(\sr[7] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _050_ (.D(\sr[8] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _051_ (.D(\sr[9] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _052_ (.D(\sr[10] ),
    .CLK(clknet_3_1__leaf_sclk),
    .Q(\sr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _053_ (.D(\sr[11] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _054_ (.D(\sr[12] ),
    .CLK(clknet_3_1__leaf_sclk),
    .Q(\sr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _055_ (.D(\sr[13] ),
    .CLK(clknet_3_1__leaf_sclk),
    .Q(\sr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _056_ (.D(\sr[14] ),
    .CLK(clknet_3_1__leaf_sclk),
    .Q(\sr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _057_ (.D(\sr[15] ),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _058_ (.D(\sr[16] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _059_ (.D(\sr[17] ),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _060_ (.D(\sr[18] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _061_ (.D(\sr[19] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _062_ (.D(\sr[20] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _063_ (.D(\sr[21] ),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _064_ (.D(\sr[22] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _065_ (.D(\sr[23] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _066_ (.D(\sr[24] ),
    .CLK(clknet_3_0__leaf_sclk),
    .Q(\sr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _067_ (.D(\sr[25] ),
    .CLK(clknet_3_2__leaf_sclk),
    .Q(\sr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _068_ (.D(\sr[26] ),
    .CLK(clknet_3_3__leaf_sclk),
    .Q(\sr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _069_ (.D(\sr[27] ),
    .CLK(clknet_3_1__leaf_sclk),
    .Q(\sr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _070_ (.D(\sr[28] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _071_ (.D(\sr[29] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _072_ (.D(\sr[30] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _073_ (.D(\sr[31] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _074_ (.D(\sr[32] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _075_ (.D(\sr[33] ),
    .CLK(clknet_3_4__leaf_sclk),
    .Q(\sr[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _076_ (.D(\sr[34] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _077_ (.D(\sr[35] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _078_ (.D(\sr[36] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _079_ (.D(\sr[37] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _080_ (.D(\sr[38] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _081_ (.D(\sr[39] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _082_ (.D(\sr[40] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _083_ (.D(\sr[41] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _084_ (.D(\sr[42] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _085_ (.D(\sr[43] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _086_ (.D(\sr[44] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _087_ (.D(\sr[45] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _088_ (.D(\sr[46] ),
    .CLK(clknet_3_4__leaf_sclk),
    .Q(\sr[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _089_ (.D(\sr[47] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _090_ (.D(\sr[48] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _091_ (.D(\sr[49] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _092_ (.D(\sr[50] ),
    .CLK(clknet_3_4__leaf_sclk),
    .Q(\sr[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _093_ (.D(\sr[51] ),
    .CLK(clknet_3_4__leaf_sclk),
    .Q(\sr[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _094_ (.D(\sr[52] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(\sr[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _095_ (.D(\sr[53] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _096_ (.D(\sr[54] ),
    .CLK(clknet_3_4__leaf_sclk),
    .Q(\sr[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _097_ (.D(\sr[55] ),
    .CLK(clknet_3_6__leaf_sclk),
    .Q(\sr[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _098_ (.D(\sr[56] ),
    .CLK(clknet_3_5__leaf_sclk),
    .Q(\sr[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _099_ (.D(\sr[57] ),
    .CLK(clknet_3_7__leaf_sclk),
    .Q(sr_out));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _100_ (.D(\sr[0] ),
    .CLK(latch),
    .Q(tune_s1_shunt[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _101_ (.D(\sr[1] ),
    .CLK(latch),
    .Q(tune_s1_shunt[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _102_ (.D(\sr[2] ),
    .CLK(latch),
    .Q(tune_s1_shunt[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _103_ (.D(\sr[3] ),
    .CLK(latch),
    .Q(tune_s1_shunt[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _104_ (.D(\sr[4] ),
    .CLK(latch),
    .Q(tune_s1_shunt[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _105_ (.D(\sr[5] ),
    .CLK(latch),
    .Q(tune_s1_shunt[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _106_ (.D(\sr[6] ),
    .CLK(latch),
    .Q(tune_s1_shunt[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _107_ (.D(\sr[7] ),
    .CLK(latch),
    .Q(tune_s1_shunt[7]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _108_ (.D(\sr[8] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _109_ (.D(\sr[9] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _110_ (.D(\sr[10] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[2]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _111_ (.D(\sr[11] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[3]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _112_ (.D(\sr[12] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[4]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _113_ (.D(\sr[13] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[5]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _114_ (.D(\sr[14] ),
    .CLK(latch),
    .Q(tune_s1_shunt_gy[6]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _115_ (.D(\sr[15] ),
    .CLK(latch),
    .Q(tune_s1_series_gy[0]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _116_ (.D(\sr[16] ),
    .CLK(latch),
    .Q(tune_s1_series_gy[1]));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _117_ (.D(\sr[17] ),
    .CLK(latch),
    .Q(tune_s1_series_gy[2]));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_17 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_18 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_19 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_20 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_21 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_22 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_23 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_24 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_25 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_26 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_27 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_28 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_29 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_30 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_sclk (.I(sclk),
    .Z(clknet_0_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_0__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_1__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_2__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_3__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_4__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_5__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_6__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_sclk (.I(clknet_0_sclk),
    .Z(clknet_3_7__leaf_sclk));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1399 ();
endmodule

