* NGSPICE file created from caparray_s1.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

.subckt caparray_s1 cap_series_gygyn cap_series_gygyp cap_series_gyn cap_series_gyp
+ cap_shunt_gyn cap_shunt_gyp cap_shunt_n cap_shunt_p tune_series_gy[0] tune_series_gy[1]
+ tune_series_gy[2] tune_series_gy[3] tune_series_gy[4] tune_series_gy[5] tune_series_gygy[0]
+ tune_series_gygy[1] tune_series_gygy[2] tune_series_gygy[3] tune_series_gygy[4]
+ tune_series_gygy[5] tune_shunt[0] tune_shunt[1] tune_shunt[2] tune_shunt[3] tune_shunt[4]
+ tune_shunt[5] tune_shunt[6] tune_shunt[7] tune_shunt_gy[0] tune_shunt_gy[1] tune_shunt_gy[2]
+ tune_shunt_gy[3] tune_shunt_gy[4] tune_shunt_gy[5] tune_shunt_gy[6] vdd vss
XFILLER_39_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[12\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[12\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[72\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[72\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g3\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[117\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[117\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[7\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[7\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[61\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[61\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g8\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[0] gen_shunt_g8\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[3\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[3\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[11\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[11\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[88\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[88\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g2\[3\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[3\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[114\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[114\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[37\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[37\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g1\[20\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[20\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[71\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[71\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g3\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[116\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[116\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[39\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[39\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[60\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[60\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[87\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[87\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g1\[3\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[3\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[113\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[113\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[36\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[36\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[70\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[70\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gygy_g1\[5\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[5\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[89\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[89\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[115\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[115\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[38\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[38\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[86\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[86\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[112\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[112\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[35\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[35\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[3\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[3\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[88\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[88\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[114\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[114\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[37\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[37\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[85\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[85\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[111\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[111\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[18\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[18\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[34\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[34\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[87\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[87\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[113\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[113\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g3\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[36\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[36\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g1\[5\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[5\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[84\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[84\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_66_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[26\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[26\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[110\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[110\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[33\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[33\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[86\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[86\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[112\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[112\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[35\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[35\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[83\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[83\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_66_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[32\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[32\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[13\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[13\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g3\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[3]
+ gen_shunt_gygy_g3\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[85\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[85\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[18\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[18\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[111\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[111\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[6\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[6\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[34\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[34\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g11\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[12\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[12\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[82\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[82\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g3\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[127\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[127\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[21\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[21\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[84\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[84\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g3\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g2\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[26\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[26\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[110\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[110\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[33\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[33\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[39\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[39\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[81\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[81\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[126\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[126\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[49\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[49\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[83\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[83\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[32\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[32\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[38\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[38\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[6\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[6\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[13\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[13\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g3\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[3]
+ gen_shunt_gygy_g3\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[80\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[80\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[99\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[99\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[6\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[6\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g7\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[1] gen_shunt_g7\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[125\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[125\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[48\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[48\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_series_gy_g11\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[12\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[12\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[82\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[82\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[37\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[37\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[127\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[127\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[21\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[21\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[6\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[6\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[98\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[98\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g3\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[39\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[39\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g7\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[1] gen_shunt_g7\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[124\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[124\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_53_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[47\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[47\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gygy_g2\[2\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[2\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[81\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[81\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[36\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[36\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[126\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[126\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_58_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[49\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[49\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g2\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[97\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[97\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[38\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[38\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[123\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[123\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[6\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[6\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[46\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[46\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g3\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_79_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[80\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[80\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[2\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[2\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[99\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[99\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g7\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[1] gen_shunt_g7\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[35\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[35\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[125\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[125\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[48\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[48\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[96\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[96\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[37\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[37\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_3_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[122\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[122\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[45\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[45\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[6\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[6\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g4\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[98\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[98\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g7\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[1] gen_shunt_g7\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g1\[19\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[19\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[34\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[34\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[124\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[124\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g1\[2\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[2\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[47\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[47\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g3\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[2] gen_shunt_gy_g3\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[2\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[2\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[2]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[95\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[95\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g3\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[36\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[36\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_80_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[121\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[121\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[44\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[44\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g4\[0\].u_shunt_n cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[0] gen_shunt_gy_g4\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[97\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[97\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[27\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[27\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[33\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[33\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[123\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[123\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[46\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[46\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g4\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[2\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[2\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g3\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[1] gen_shunt_gy_g3\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[94\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[94\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[35\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[35\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp2 cap_series_gygyp cap_series_gygyp tune_series_gygy[1]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[120\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[120\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[4\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[4\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[43\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[43\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[96\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[96\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[32\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[32\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[122\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[122\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[45\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[45\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[14\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[14\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[93\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[93\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g3\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[19\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[19\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[34\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[34\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[7\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[7\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[2\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[2\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g3\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[2] gen_shunt_gy_g3\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[42\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[42\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g6\[0\].u_shunt_gyp3 cap_series_gygyp cap_series_gygyp tune_series_gygy[0]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyp3/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[2]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[13\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[13\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g4\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[95\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[95\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g3\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g3\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_series_gy_g11\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[121\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[121\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[44\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[44\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[22\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[22\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g4\[0\].u_shunt_p cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[0] gen_shunt_gy_g4\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_80_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[92\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[92\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[27\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[27\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[33\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[33\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[41\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[41\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g3\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[1] gen_shunt_gy_g3\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[94\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[94\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn2 cap_series_gygyn cap_series_gygyn tune_series_gygy[1]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn2/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g2\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g2\[3\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[3\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g1\[4\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[4\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[120\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[120\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[43\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[43\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[49\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[49\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[30\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[30\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[91\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[91\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[32\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[32\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[14\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[14\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[40\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[40\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[2\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[2\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[59\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[59\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[93\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[93\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[21\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[21\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[7\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[7\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[42\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[42\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[48\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[48\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g6\[0\].u_shunt_gyn3 cap_series_gygyn cap_series_gygyn tune_series_gygy[0]
+ gen_shunt_gygy_g6\[0\].u_shunt_gyn3/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g2\[3\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[3\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g11\[13\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[13\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[90\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[90\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[22\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[22\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[58\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[58\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[92\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[92\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[20\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[20\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[41\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[41\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[47\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[47\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g6\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g2\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[3\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[3\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[49\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[49\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[30\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[30\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[57\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[57\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g1\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[91\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[91\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g5\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[0]
+ gen_series_gy_g5\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[40\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[40\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[46\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[46\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[2\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[2\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[59\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[59\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g6\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[48\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[48\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[56\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[56\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g2\[3\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[3\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[90\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[90\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[5\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[5\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[45\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[45\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[58\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[58\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[47\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[47\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[55\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[55\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[8\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[8\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[44\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[44\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[57\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[57\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[5\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[5\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g2\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[2] gen_shunt_g6\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g5\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[0]
+ gen_series_gy_g5\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[28\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[28\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g2\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[46\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[46\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[54\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[54\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g6\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[43\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[43\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[56\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[56\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[5\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[5\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[45\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[45\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_29_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[15\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[15\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[7\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[7\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[53\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[53\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[8\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[8\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[42\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[42\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_46_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[55\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[55\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g11\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[14\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[14\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[31\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[31\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[8\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[8\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[44\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[44\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g2\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[23\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[23\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[5\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[5\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[52\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[52\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g6\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[2] gen_shunt_g6\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[28\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[28\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g3\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[2] gen_shunt_gy_g3\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[41\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[41\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[54\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[54\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[30\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[30\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[43\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[43\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[31\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[31\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[51\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[51\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[10\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[10\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g2\[40\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[40\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[15\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[15\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[3\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[3\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gygy_g1\[7\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[7\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[53\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[53\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g2\[59\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[59\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gy_g3\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[1] gen_shunt_gy_g3\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g4\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[1]
+ gen_series_gy_g4\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[3\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[3\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g1\[8\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[8\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[42\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[42\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[50\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[50\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[14\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[14\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[69\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[69\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g3\[31\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[31\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_80_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[23\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[23\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[52\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[52\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[58\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[58\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g3\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[2] gen_shunt_gy_g3\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[41\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[41\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[68\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[68\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[30\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[5] gen_shunt_g3\[30\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[31\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[31\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[51\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[51\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[57\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[57\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g5\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[10\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[10\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g2\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[40\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[40\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[3\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[3\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[59\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[59\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_gy_g3\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[1] gen_shunt_gy_g3\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g4\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[1]
+ gen_series_gy_g4\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[67\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[67\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[2\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[2\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[3\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[3\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[50\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[50\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[56\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[56\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[69\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[69\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_52_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g2\[58\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[58\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[66\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[66\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gy_g2\[2\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[2\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[55\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[55\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g5\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[68\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[68\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_37_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[9\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[9\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[57\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[57\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g5\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[65\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[65\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g2\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_series_gy_g1\[29\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[29\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[54\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[54\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g5\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[67\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[67\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g2\[2\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[2\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[56\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[56\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g5\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[64\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[64\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[109\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[109\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[16\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[16\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[53\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[53\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_80_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g5\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[66\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[66\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[9\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[9\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[2\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[2\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g3\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g2\[55\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[55\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g5\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[63\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[63\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[4\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[15\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[15\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g11\[9\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[9\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[108\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[108\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_51_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_series_gy_g1\[24\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[24\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[52\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[52\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g5\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[65\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[65\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[29\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[29\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[54\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[54\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[62\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[62\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gy_g1\[4\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[4\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_g1\[107\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[107\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_28_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[51\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[51\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[3] gen_shunt_g5\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[64\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[64\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[11\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[11\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[0\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[0\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[109\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[109\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_24_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[16\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[16\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[4\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[4\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[53\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[53\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g5\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[61\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[61\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g4\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[1]
+ gen_series_gy_g4\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[9\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[9\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g11\[10\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[10\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[106\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[106\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_series_gy_g3\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g11\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[50\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[50\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[63\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[63\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[4\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g11\[15\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[15\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g1\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[108\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[108\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g1\[6\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[6\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[0\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[0\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[24\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[24\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[52\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[52\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[60\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[60\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_58_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[79\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[79\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[105\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[105\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[62\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[62\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[3\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[3\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_17_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[4\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[4\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[107\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[107\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[51\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[51\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g5\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[3] gen_shunt_g5\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_gy_g1\[0\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[0\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g1\[11\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[11\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_gygy_g2\[0\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[4]
+ gen_shunt_gygy_g2\[0\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[78\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[78\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[19\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[19\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_79_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g4\[9\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[9\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[104\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[104\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[27\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[27\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g1\[4\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[4\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_61_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[61\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[61\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_series_gy_g4\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[1]
+ gen_series_gy_g4\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[10\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[10\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[2\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[2\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_55_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[16\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[16\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[10\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[10\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[106\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[106\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_4_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[29\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[29\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[50\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[50\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[77\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[77\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[18\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[18\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_gygy_g1\[6\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[6\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[0\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[0\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_g4\[8\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[8\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[103\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[103\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[26\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[26\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[60\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[60\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_79_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g1\[2\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[5]
+ gen_shunt_gygy_g1\[2\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[79\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[79\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[1\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[1\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[15\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[15\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[105\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[105\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[28\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[28\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[76\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[76\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[17\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[17\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g2\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[3]
+ gen_series_gy_g2\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[7\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[7\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[102\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[102\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[25\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[25\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g1\[0\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[5] gen_shunt_gy_g1\[0\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_series_gy_g2\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[78\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[78\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[0\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[0\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g2\[14\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[14\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[104\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[104\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g4\[9\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[9\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[27\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[27\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_30_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gygy_g3\[1\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[3]
+ gen_shunt_gygy_g3\[1\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_80_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[75\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[75\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[16\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[16\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[101\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[101\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[6\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[6\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[24\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[24\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xgen_shunt_g1\[77\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[77\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g2\[13\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[13\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[103\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[103\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[8\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[8\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[26\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[26\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_series_gy_g1\[17\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[17\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_21_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g2\[1\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[4] gen_shunt_gy_g2\[1\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xgen_shunt_gygy_g1\[2\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[5]
+ gen_shunt_gygy_g1\[2\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[74\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[74\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[15\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[15\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[100\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[100\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[5\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[5\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[23\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[23\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[119\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[119\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[1\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[2]
+ gen_series_gy_g3\[1\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g11\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[63\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[63\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xgen_shunt_g1\[76\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[76\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g2\[0\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[3]
+ gen_series_gy_g2\[0\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_63_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[12\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[12\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[102\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[102\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[7\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[7\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[25\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[25\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[25\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[25\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_45_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[73\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[73\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[7\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[7\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[14\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[14\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g2\[1\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[3] gen_shunt_gy_g2\[1\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_gygy_g3\[1\].u_shunt_gyn1 cap_series_gygyn cap_series_gygyn tune_series_gygy[3]
+ gen_shunt_gygy_g3\[1\].u_shunt_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[4\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[4\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[22\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[22\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_2_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[118\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[118\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[62\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[62\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g1\[75\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[75\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[11\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[11\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[101\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[101\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g4\[6\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[6\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[24\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[24\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g1\[12\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[12\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[72\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[72\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[13\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[13\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g3\[19\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[19\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[3\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[3\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[21\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[21\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_series_gy_g1\[17\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[17\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[117\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[117\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[7\].u_shunt_gyp2 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[5] gen_shunt_gy_g1\[7\].u_shunt_gyp2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_series_gy_g1\[5\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[5\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gy_g2\[1\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[4] gen_shunt_gy_g2\[1\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[61\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[61\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g8\[0\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[0] gen_shunt_g8\[0\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_80_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[0\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[0\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[74\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[74\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_series_gy_g11\[11\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[4]
+ gen_series_gy_g11\[11\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_75_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_gygy_g2\[3\].u_shunt_gyp1 cap_series_gygyp cap_series_gygyp tune_series_gygy[4]
+ gen_shunt_gygy_g2\[3\].u_shunt_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[10\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[10\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[100\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[100\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[5\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[5\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[23\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[23\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[29\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[29\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[119\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[119\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g3\[1\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[2]
+ gen_series_gy_g3\[1\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_series_gy_g11\[5\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[4]
+ gen_series_gy_g11\[5\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[63\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[63\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_series_gy_g1\[20\].u_series_gyp1 cap_series_gyp cap_series_gyp tune_series_gy[5]
+ gen_series_gy_g1\[20\].u_series_gyp1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xgen_shunt_g1\[71\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[71\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g3\[18\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[18\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[12\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[12\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g4\[2\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[2\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[20\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[20\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_series_gy_g1\[25\].u_series_gyn1 cap_series_gyn cap_series_gyn tune_series_gy[5]
+ gen_series_gy_g1\[25\].u_series_gyn1/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_33_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g1\[116\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[116\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[39\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[39\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g2\[60\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[60\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_10_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[73\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[73\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_gy_g1\[7\].u_shunt_gyn1 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[6] gen_shunt_gy_g1\[7\].u_shunt_gyn1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xgen_shunt_gy_g2\[1\].u_shunt_gyn2 cap_shunt_gyn cap_shunt_gyn tune_shunt_gy[3] gen_shunt_gy_g2\[1\].u_shunt_gyn2/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g4\[4\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[4] gen_shunt_g4\[4\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[28\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[6] gen_shunt_g2\[28\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[22\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[22\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g1\[118\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[7] gen_shunt_g1\[118\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_gy_g1\[3\].u_shunt_gyp1 cap_shunt_gyp cap_shunt_gyp tune_shunt_gy[6] gen_shunt_gy_g1\[3\].u_shunt_gyp1/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g2\[62\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[62\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xgen_shunt_g1\[70\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[70\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[89\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[89\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xgen_shunt_g3\[17\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[5] gen_shunt_g3\[17\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xgen_shunt_g2\[11\].u_shunt_p cap_shunt_p cap_shunt_p tune_shunt[6] gen_shunt_g2\[11\].u_shunt_p/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_16_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xgen_shunt_g4\[1\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[4] gen_shunt_g4\[1\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xgen_shunt_g1\[115\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[115\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xgen_shunt_g1\[38\].u_shunt_n cap_shunt_n cap_shunt_n tune_shunt[7] gen_shunt_g1\[38\].u_shunt_n/ZN
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_36_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

