magic
tech gf180mcuC
magscale 1 5
timestamp 1669699727
<< obsm1 >>
rect 672 1538 11392 8262
<< metal2 >>
rect 1064 0 1120 400
rect 3024 0 3080 400
rect 4984 0 5040 400
rect 6944 0 7000 400
rect 8904 0 8960 400
rect 10864 0 10920 400
<< obsm2 >>
rect 1022 430 11378 8251
rect 1022 400 1034 430
rect 1150 400 2994 430
rect 3110 400 4954 430
rect 5070 400 6914 430
rect 7030 400 8874 430
rect 8990 400 10834 430
rect 10950 400 11378 430
<< metal3 >>
rect 0 7448 400 7504
rect 11600 7448 12000 7504
rect 0 2464 400 2520
rect 11600 2464 12000 2520
<< obsm3 >>
rect 400 7534 11600 8246
rect 430 7418 11570 7534
rect 400 2550 11600 7418
rect 430 2434 11570 2550
rect 400 1554 11600 2434
<< metal4 >>
rect 1922 1538 2082 8262
rect 3252 1538 3412 8262
rect 4582 1538 4742 8262
rect 5912 1538 6072 8262
rect 7242 1538 7402 8262
rect 8572 1538 8732 8262
rect 9902 1538 10062 8262
rect 11232 1538 11392 8262
<< labels >>
rlabel metal3 s 0 7448 400 7504 6 nbusin_nshunt
port 1 nsew signal bidirectional
rlabel metal3 s 11600 7448 12000 7504 6 nbusout
port 2 nsew signal bidirectional
rlabel metal2 s 6944 0 7000 400 6 nseries_gy
port 3 nsew signal bidirectional
rlabel metal2 s 10864 0 10920 400 6 nseries_gygy
port 4 nsew signal bidirectional
rlabel metal2 s 3024 0 3080 400 6 nshunt_gy
port 5 nsew signal bidirectional
rlabel metal3 s 0 2464 400 2520 6 pbusin_pshunt
port 6 nsew signal bidirectional
rlabel metal3 s 11600 2464 12000 2520 6 pbusout
port 7 nsew signal bidirectional
rlabel metal2 s 4984 0 5040 400 6 pseries_gy
port 8 nsew signal bidirectional
rlabel metal2 s 8904 0 8960 400 6 pseries_gygy
port 9 nsew signal bidirectional
rlabel metal2 s 1064 0 1120 400 6 pshunt_gy
port 10 nsew signal bidirectional
rlabel metal4 s 1922 1538 2082 8262 6 vdd
port 11 nsew power bidirectional
rlabel metal4 s 4582 1538 4742 8262 6 vdd
port 11 nsew power bidirectional
rlabel metal4 s 7242 1538 7402 8262 6 vdd
port 11 nsew power bidirectional
rlabel metal4 s 9902 1538 10062 8262 6 vdd
port 11 nsew power bidirectional
rlabel metal4 s 3252 1538 3412 8262 6 vss
port 12 nsew ground bidirectional
rlabel metal4 s 5912 1538 6072 8262 6 vss
port 12 nsew ground bidirectional
rlabel metal4 s 8572 1538 8732 8262 6 vss
port 12 nsew ground bidirectional
rlabel metal4 s 11232 1538 11392 8262 6 vss
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 361376
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/dlc/runs/22_11_29_00_28/results/signoff/filterstage.magic.gds
string GDS_START 48204
<< end >>

