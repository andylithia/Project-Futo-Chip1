magic
tech gf180mcuC
magscale 1 10
timestamp 1670004454
<< deepnwell >>
rect 199000 199000 206000 206000
<< nwell >>
rect 200000 204000 205000 205200
rect 200000 201000 201000 204000
rect 204000 201000 205000 204000
rect 200000 199800 205000 201000
<< pwell >>
rect 194000 210000 211000 211000
rect 194000 195000 195000 210000
rect 210000 195000 211000 210000
rect 194000 194000 211000 195000
<< psubdiff >>
rect 194200 210700 210800 210800
rect 194200 210300 194800 210700
rect 210200 210300 210800 210700
rect 194200 210200 210800 210300
rect 194200 194800 194800 210200
rect 210200 194800 210800 210200
rect 194200 194700 210800 194800
rect 194200 194300 194800 194700
rect 210200 194300 210800 194700
rect 194200 194200 210800 194300
<< nsubdiff >>
rect 200200 204800 204800 205000
rect 200200 204400 200400 204800
rect 204600 204400 204800 204800
rect 200200 204200 204800 204400
rect 200200 200800 200800 204200
rect 204200 200800 204800 204200
rect 200200 200600 204800 200800
rect 200200 200200 200400 200600
rect 204600 200200 204800 200600
rect 200200 200000 204800 200200
<< psubdiffcont >>
rect 194800 210300 210200 210700
rect 194800 194300 210200 194700
<< nsubdiffcont >>
rect 200400 204400 204600 204800
rect 200400 200200 204600 200600
<< metal1 >>
rect 194200 210700 210800 210800
rect 194200 210300 194800 210700
rect 210200 210300 210800 210700
rect 194200 210200 210800 210300
rect 200200 204800 204800 205000
rect 200200 204400 200400 204800
rect 204600 204400 204800 204800
rect 200200 204200 204800 204400
rect 200200 200600 204800 200800
rect 200200 200200 200400 200600
rect 204600 200200 204800 200600
rect 200200 200000 204800 200200
rect 194200 194700 210800 194800
rect 194200 194300 194800 194700
rect 210200 194300 210800 194700
rect 194200 194200 210800 194300
<< metal2 >>
rect 10108 599564 11508 599620
rect 11592 599592 11816 600960
rect 33768 599592 33992 600960
rect 10108 596288 10164 599564
rect 11452 599508 11508 599564
rect 11564 599520 11816 599592
rect 33740 599520 33992 599592
rect 55468 599564 55860 599620
rect 55944 599592 56168 600960
rect 11564 599508 11620 599520
rect 11452 599452 11620 599508
rect 33740 596288 33796 599520
rect 55468 596288 55524 599564
rect 55804 599508 55860 599564
rect 55916 599520 56168 599592
rect 78120 599592 78344 600960
rect 100296 599592 100520 600960
rect 78120 599520 78372 599592
rect 100296 599520 100548 599592
rect 55916 599508 55972 599520
rect 55804 599452 55972 599508
rect 78316 596288 78372 599520
rect 100492 596288 100548 599520
rect 120988 599564 122388 599620
rect 122472 599592 122696 600960
rect 120988 596288 121044 599564
rect 122332 599508 122388 599564
rect 122444 599520 122696 599592
rect 144648 599592 144872 600960
rect 144648 599520 144900 599592
rect 122444 599508 122500 599520
rect 122332 599452 122500 599508
rect 144844 596288 144900 599520
rect 166348 599564 166740 599620
rect 166824 599592 167048 600960
rect 166348 596288 166404 599564
rect 166684 599508 166740 599564
rect 166796 599520 167048 599592
rect 189000 599592 189224 600960
rect 211176 599592 211400 600960
rect 233352 599592 233576 600960
rect 255528 599592 255752 600960
rect 277704 599592 277928 600960
rect 299880 599592 300104 600960
rect 189000 599520 189252 599592
rect 211176 599520 211428 599592
rect 166796 599508 166852 599520
rect 166684 599452 166852 599508
rect 188188 598164 188244 598174
rect 188188 596288 188244 598108
rect 189196 596288 189252 599520
rect 211372 596288 211428 599520
rect 233324 599520 233576 599592
rect 255500 599520 255752 599592
rect 277676 599520 277928 599592
rect 299852 599520 300104 599592
rect 320908 599564 321972 599620
rect 322056 599592 322280 600960
rect 233324 596288 233380 599520
rect 255500 596288 255556 599520
rect 277676 596288 277732 599520
rect 299852 596288 299908 599520
rect 320908 596288 320964 599564
rect 321916 599508 321972 599564
rect 322028 599520 322280 599592
rect 342748 599564 344148 599620
rect 344232 599592 344456 600960
rect 366408 599592 366632 600960
rect 322028 599508 322084 599520
rect 321916 599452 322084 599508
rect 342748 596288 342804 599564
rect 344092 599508 344148 599564
rect 344204 599520 344456 599592
rect 366380 599520 366632 599592
rect 388108 599564 388500 599620
rect 388584 599592 388808 600960
rect 344204 599508 344260 599520
rect 344092 599452 344260 599508
rect 366380 596288 366436 599520
rect 388108 596288 388164 599564
rect 388444 599508 388500 599564
rect 388556 599520 388808 599592
rect 409948 599564 410676 599620
rect 410760 599592 410984 600960
rect 388556 599508 388612 599520
rect 388444 599452 388612 599508
rect 409948 596288 410004 599564
rect 410620 599508 410676 599564
rect 410732 599520 410984 599592
rect 431788 599564 432852 599620
rect 432936 599592 433160 600960
rect 410732 599508 410788 599520
rect 410620 599452 410788 599508
rect 431788 596288 431844 599564
rect 432796 599508 432852 599564
rect 432908 599520 433160 599592
rect 453628 599564 455028 599620
rect 455112 599592 455336 600960
rect 477288 599592 477512 600960
rect 432908 599508 432964 599520
rect 432796 599452 432964 599508
rect 453628 596288 453684 599564
rect 454972 599508 455028 599564
rect 455084 599520 455336 599592
rect 477260 599520 477512 599592
rect 498988 599564 499380 599620
rect 499464 599592 499688 600960
rect 455084 599508 455140 599520
rect 454972 599452 455140 599508
rect 477260 596288 477316 599520
rect 498988 596288 499044 599564
rect 499324 599508 499380 599564
rect 499436 599520 499688 599592
rect 520828 599564 521556 599620
rect 521640 599592 521864 600960
rect 543816 599592 544040 600960
rect 499436 599508 499492 599520
rect 499324 599452 499492 599508
rect 520828 596288 520884 599564
rect 521500 599508 521556 599564
rect 521612 599520 521864 599592
rect 543788 599520 544040 599592
rect 564508 599564 565908 599620
rect 565992 599592 566216 600960
rect 588168 599592 588392 600960
rect 521612 599508 521668 599520
rect 521500 599452 521668 599508
rect 543788 596288 543844 599520
rect 564508 596288 564564 599564
rect 565852 599508 565908 599564
rect 565964 599520 566216 599592
rect 588140 599520 588392 599592
rect 565964 599508 566020 599520
rect 565852 599452 566020 599508
rect 588140 598164 588196 599520
rect 588140 598098 588196 598108
rect 598108 579796 598164 579806
rect 4172 534548 4228 534558
rect 4172 291956 4228 534492
rect 4396 477652 4452 477662
rect 4284 434980 4340 434990
rect 4284 304948 4340 434924
rect 4284 304882 4340 304892
rect 4172 291890 4228 291900
rect 4284 300804 4340 300814
rect 4172 130228 4228 130238
rect 4172 65380 4228 130172
rect 4284 79604 4340 300748
rect 4396 291844 4452 477596
rect 595756 406644 595812 406654
rect 4396 291778 4452 291788
rect 4620 363860 4676 363870
rect 4620 291732 4676 363804
rect 595644 312564 595700 312574
rect 595532 307524 595588 307534
rect 4620 291666 4676 291676
rect 4844 306964 4900 306974
rect 4844 291620 4900 306908
rect 4844 291554 4900 291564
rect 595532 126868 595588 307468
rect 595644 153524 595700 312508
rect 595756 306628 595812 406588
rect 595756 306562 595812 306572
rect 595868 315924 595924 315934
rect 595868 220052 595924 315868
rect 595980 314244 596036 314254
rect 595980 260148 596036 314188
rect 596092 313236 596148 313246
rect 596092 291508 596148 313180
rect 598108 303268 598164 579740
rect 598108 303202 598164 303212
rect 596092 291442 596148 291452
rect 595980 260082 596036 260092
rect 595868 219986 595924 219996
rect 595644 153458 595700 153468
rect 595532 126802 595588 126812
rect 595644 141988 595700 141998
rect 4284 79538 4340 79548
rect 4172 65314 4228 65324
rect 595644 33572 595700 141932
rect 595644 33506 595700 33516
rect 11788 420 11844 2326
rect 13132 480 13300 532
rect 15148 480 15204 2326
rect 17052 480 17108 2326
rect 13132 476 13496 480
rect 13132 420 13188 476
rect 11788 364 13188 420
rect 13244 392 13496 476
rect 15148 392 15400 480
rect 17052 392 17304 480
rect 13272 -960 13496 392
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18508 420 18564 2326
rect 18844 480 19012 532
rect 21084 480 21140 2326
rect 22988 480 23044 2326
rect 18844 476 19208 480
rect 18844 420 18900 476
rect 18508 364 18900 420
rect 18956 392 19208 476
rect 18984 -960 19208 392
rect 20888 392 21140 480
rect 22792 392 23044 480
rect 23548 420 23604 2326
rect 24556 480 24724 532
rect 24556 476 24920 480
rect 24556 420 24612 476
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 23548 364 24612 420
rect 24668 392 24920 476
rect 24696 -960 24920 392
rect 25228 420 25284 2326
rect 26460 480 26628 532
rect 28700 480 28756 2326
rect 30604 480 30660 2326
rect 26460 476 26824 480
rect 26460 420 26516 476
rect 25228 364 26516 420
rect 26572 392 26824 476
rect 26600 -960 26824 392
rect 28504 392 28756 480
rect 30408 392 30660 480
rect 31948 420 32004 2326
rect 32172 480 32340 532
rect 32172 476 32536 480
rect 32172 420 32228 476
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 31948 364 32228 420
rect 32284 392 32536 476
rect 32312 -960 32536 392
rect 33628 420 33684 2326
rect 34076 480 34244 532
rect 34076 476 34440 480
rect 34076 420 34132 476
rect 33628 364 34132 420
rect 34188 392 34440 476
rect 34216 -960 34440 392
rect 35308 420 35364 2326
rect 35980 480 36148 532
rect 35980 476 36344 480
rect 35980 420 36036 476
rect 35308 364 36036 420
rect 36092 392 36344 476
rect 36120 -960 36344 392
rect 36988 420 37044 2326
rect 37884 480 38052 532
rect 40124 480 40180 2326
rect 41916 480 41972 2326
rect 43932 480 43988 2326
rect 45836 480 45892 2326
rect 47740 480 47796 2326
rect 37884 476 38248 480
rect 37884 420 37940 476
rect 36988 364 37940 420
rect 37996 392 38248 476
rect 38024 -960 38248 392
rect 39928 392 40180 480
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 392 43988 480
rect 45640 392 45892 480
rect 47544 392 47796 480
rect 48748 420 48804 2326
rect 49308 480 49476 532
rect 49308 476 49672 480
rect 49308 420 49364 476
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 48748 364 49364 420
rect 49420 392 49672 476
rect 49448 -960 49672 392
rect 50428 420 50484 2326
rect 51212 480 51380 532
rect 53452 480 53508 2326
rect 51212 476 51576 480
rect 51212 420 51268 476
rect 50428 364 51268 420
rect 51324 392 51576 476
rect 51352 -960 51576 392
rect 53256 392 53508 480
rect 53788 420 53844 2326
rect 55020 480 55188 532
rect 57148 480 57204 2326
rect 59164 480 59220 2326
rect 55020 476 55384 480
rect 55020 420 55076 476
rect 53256 -960 53480 392
rect 53788 364 55076 420
rect 55132 392 55384 476
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58968 392 59220 480
rect 60508 420 60564 2326
rect 60732 480 60900 532
rect 62972 480 63028 2326
rect 64876 480 64932 2326
rect 60732 476 61096 480
rect 60732 420 60788 476
rect 58968 -960 59192 392
rect 60508 364 60788 420
rect 60844 392 61096 476
rect 60872 -960 61096 392
rect 62776 392 63028 480
rect 64680 392 64932 480
rect 65548 420 65604 2326
rect 66444 480 66612 532
rect 66444 476 66808 480
rect 66444 420 66500 476
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 65548 364 66500 420
rect 66556 392 66808 476
rect 66584 -960 66808 392
rect 67228 420 67284 2326
rect 68348 480 68516 532
rect 70476 480 70532 2326
rect 72268 480 72324 2326
rect 74172 480 74228 2326
rect 76300 480 76356 2326
rect 78204 480 78260 2326
rect 80108 480 80164 2326
rect 82012 480 82068 2326
rect 68348 476 68712 480
rect 68348 420 68404 476
rect 67228 364 68404 420
rect 68460 392 68712 476
rect 68488 -960 68712 392
rect 70392 -960 70616 480
rect 72268 392 72520 480
rect 74172 392 74424 480
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 392 76356 480
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 82348 420 82404 2326
rect 83580 480 83748 532
rect 85708 480 85764 2326
rect 87724 480 87780 2326
rect 89628 480 89684 2326
rect 91532 480 91588 2326
rect 83580 476 83944 480
rect 83580 420 83636 476
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 82348 364 83636 420
rect 83692 392 83944 476
rect 83720 -960 83944 392
rect 85624 -960 85848 480
rect 87528 392 87780 480
rect 89432 392 89684 480
rect 91336 392 91588 480
rect 92428 420 92484 2326
rect 93100 480 93268 532
rect 95340 480 95396 2326
rect 93100 476 93464 480
rect 93100 420 93156 476
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 92428 364 93156 420
rect 93212 392 93464 476
rect 93240 -960 93464 392
rect 95144 392 95396 480
rect 95788 420 95844 2326
rect 96908 480 97076 532
rect 99036 480 99092 2326
rect 101052 480 101108 2326
rect 96908 476 97272 480
rect 96908 420 96964 476
rect 95144 -960 95368 392
rect 95788 364 96964 420
rect 97020 392 97272 476
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102732 480 102788 2326
rect 102732 392 102984 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104188 420 104244 2326
rect 104524 480 104692 532
rect 104524 476 104888 480
rect 104524 420 104580 476
rect 104188 364 104580 420
rect 104636 392 104888 476
rect 104664 -960 104888 392
rect 105868 420 105924 2326
rect 106428 480 106596 532
rect 106428 476 106792 480
rect 106428 420 106484 476
rect 105868 364 106484 420
rect 106540 392 106792 476
rect 106568 -960 106792 392
rect 107548 420 107604 2326
rect 108332 480 108500 532
rect 108332 476 108696 480
rect 108332 420 108388 476
rect 107548 364 108388 420
rect 108444 392 108696 476
rect 108472 -960 108696 392
rect 109228 420 109284 2326
rect 110236 480 110404 532
rect 110236 476 110600 480
rect 110236 420 110292 476
rect 109228 364 110292 420
rect 110348 392 110600 476
rect 110376 -960 110600 392
rect 110908 420 110964 2326
rect 112140 480 112308 532
rect 114268 480 114324 2326
rect 116284 480 116340 2326
rect 118188 480 118244 2326
rect 119980 480 120036 2326
rect 112140 476 112504 480
rect 112140 420 112196 476
rect 110908 364 112196 420
rect 112252 392 112504 476
rect 112280 -960 112504 392
rect 114184 -960 114408 480
rect 116088 392 116340 480
rect 117992 392 118244 480
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 480
rect 120988 420 121044 2326
rect 121660 480 121828 532
rect 121660 476 122024 480
rect 121660 420 121716 476
rect 120988 364 121716 420
rect 121772 392 122024 476
rect 121800 -960 122024 392
rect 122668 420 122724 2326
rect 123564 480 123732 532
rect 123564 476 123928 480
rect 123564 420 123620 476
rect 122668 364 123620 420
rect 123676 392 123928 476
rect 123704 -960 123928 392
rect 124684 420 124740 2326
rect 125468 480 125636 532
rect 127596 480 127652 2326
rect 129500 480 129556 2326
rect 131516 480 131572 2326
rect 125468 476 125832 480
rect 125468 420 125524 476
rect 124684 364 125524 420
rect 125580 392 125832 476
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129416 -960 129640 480
rect 131320 392 131572 480
rect 133196 480 133252 2326
rect 135324 480 135380 2326
rect 137228 480 137284 2326
rect 139132 480 139188 2326
rect 133196 392 133448 480
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 392 135380 480
rect 137032 392 137284 480
rect 138936 392 139188 480
rect 139468 420 139524 2326
rect 140700 480 140868 532
rect 142828 480 142884 2326
rect 144844 480 144900 2326
rect 140700 476 141064 480
rect 140700 420 140756 476
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 139468 364 140756 420
rect 140812 392 141064 476
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144648 392 144900 480
rect 146188 420 146244 2326
rect 146412 480 146580 532
rect 148652 480 148708 2326
rect 146412 476 146776 480
rect 146412 420 146468 476
rect 144648 -960 144872 392
rect 146188 364 146468 420
rect 146524 392 146776 476
rect 146552 -960 146776 392
rect 148456 392 148708 480
rect 149548 420 149604 2326
rect 150220 480 150388 532
rect 150220 476 150584 480
rect 150220 420 150276 476
rect 148456 -960 148680 392
rect 149548 364 150276 420
rect 150332 392 150584 476
rect 150360 -960 150584 392
rect 151228 420 151284 2326
rect 152124 480 152292 532
rect 154364 480 154420 2326
rect 152124 476 152488 480
rect 152124 420 152180 476
rect 151228 364 152180 420
rect 152236 392 152488 476
rect 152264 -960 152488 392
rect 154168 392 154420 480
rect 154588 420 154644 2326
rect 155932 480 156100 532
rect 158172 480 158228 2326
rect 159964 480 160020 2326
rect 155932 476 156296 480
rect 155932 420 155988 476
rect 154168 -960 154392 392
rect 154588 364 155988 420
rect 156044 392 156296 476
rect 156072 -960 156296 392
rect 157976 392 158228 480
rect 157976 -960 158200 392
rect 159880 -960 160104 480
rect 161308 420 161364 2326
rect 161644 480 161812 532
rect 161644 476 162008 480
rect 161644 420 161700 476
rect 161308 364 161700 420
rect 161756 392 162008 476
rect 161784 -960 162008 392
rect 163324 420 163380 2326
rect 163548 480 163716 532
rect 163548 476 163912 480
rect 163548 420 163604 476
rect 163324 364 163604 420
rect 163660 392 163912 476
rect 163688 -960 163912 392
rect 164668 420 164724 2326
rect 165452 480 165620 532
rect 167692 480 167748 2326
rect 165452 476 165816 480
rect 165452 420 165508 476
rect 164668 364 165508 420
rect 165564 392 165816 476
rect 165592 -960 165816 392
rect 167496 392 167748 480
rect 168700 420 168756 2326
rect 169260 480 169428 532
rect 171388 480 171444 2326
rect 173180 480 173236 2326
rect 175084 480 175140 2326
rect 169260 476 169624 480
rect 169260 420 169316 476
rect 167496 -960 167720 392
rect 168700 364 169316 420
rect 169372 392 169624 476
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 176428 420 176484 2326
rect 176876 480 177044 532
rect 176876 476 177240 480
rect 176876 420 176932 476
rect 176428 364 176932 420
rect 176988 392 177240 476
rect 177016 -960 177240 392
rect 178220 420 178276 2326
rect 178780 480 178948 532
rect 180796 480 180852 2326
rect 182700 480 182756 2326
rect 178780 476 179144 480
rect 178780 420 178836 476
rect 178220 364 178836 420
rect 178892 392 179144 476
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 183260 420 183316 2326
rect 184492 480 184660 532
rect 186508 480 186564 2326
rect 188412 480 188468 2326
rect 190316 480 190372 2326
rect 192220 480 192276 2326
rect 194124 480 194180 2326
rect 184492 476 184856 480
rect 184492 420 184548 476
rect 183260 364 184548 420
rect 184604 392 184856 476
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 190316 392 190568 480
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 194908 420 194964 2326
rect 195916 480 196084 532
rect 197932 480 197988 2326
rect 200060 480 200116 2326
rect 195916 476 196280 480
rect 195916 420 195972 476
rect 194908 364 195972 420
rect 196028 392 196280 476
rect 197932 392 198184 480
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 392 200116 480
rect 201740 480 201796 2326
rect 203644 480 203700 2326
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 199864 -960 200088 392
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 204988 420 205044 2326
rect 205436 480 205604 532
rect 207452 480 207508 2326
rect 209356 480 209412 2326
rect 205436 476 205800 480
rect 205436 420 205492 476
rect 204988 364 205492 420
rect 205548 392 205800 476
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 210140 420 210196 2326
rect 211148 480 211316 532
rect 213164 480 213220 2326
rect 211148 476 211512 480
rect 211148 420 211204 476
rect 210140 364 211204 420
rect 211260 392 211512 476
rect 213164 392 213416 480
rect 211288 -960 211512 392
rect 213192 -960 213416 392
rect 214060 196 214116 2326
rect 215068 480 215124 2326
rect 217084 480 217140 2326
rect 215068 392 215320 480
rect 214060 130 214116 140
rect 215096 -960 215320 392
rect 217000 -960 217224 480
rect 218428 420 218484 2326
rect 218764 480 218932 532
rect 220780 480 220836 2326
rect 222684 480 222740 2326
rect 218764 476 219128 480
rect 218764 420 218820 476
rect 218428 364 218820 420
rect 218876 392 219128 476
rect 220780 392 221032 480
rect 222684 392 222936 480
rect 218904 -960 219128 392
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 223468 420 223524 2326
rect 224476 480 224644 532
rect 224476 476 224840 480
rect 224476 420 224532 476
rect 223468 364 224532 420
rect 224588 392 224840 476
rect 224616 -960 224840 392
rect 225260 420 225316 2326
rect 226380 480 226548 532
rect 228620 480 228676 2326
rect 226380 476 226744 480
rect 226380 420 226436 476
rect 225260 364 226436 420
rect 226492 392 226744 476
rect 226520 -960 226744 392
rect 228424 392 228676 480
rect 228424 -960 228648 392
rect 228844 84 228900 2326
rect 230300 480 230356 2326
rect 232204 480 232260 2326
rect 234108 480 234164 2326
rect 230300 392 230552 480
rect 232204 392 232456 480
rect 234108 392 234360 480
rect 228844 18 228900 28
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 234136 -960 234360 392
rect 235228 420 235284 2326
rect 235900 480 236068 532
rect 237916 480 237972 2326
rect 235900 476 236264 480
rect 235900 420 235956 476
rect 235228 364 235956 420
rect 236012 392 236264 476
rect 237916 392 238168 480
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 238588 420 238644 2326
rect 239708 480 239876 532
rect 239708 476 240072 480
rect 239708 420 239764 476
rect 238588 364 239764 420
rect 239820 392 240072 476
rect 239848 -960 240072 392
rect 240380 420 240436 2326
rect 241612 480 241780 532
rect 243628 480 243684 2326
rect 245532 480 245588 2326
rect 247436 480 247492 2326
rect 241612 476 241976 480
rect 241612 420 241668 476
rect 240380 364 241668 420
rect 241724 392 241976 476
rect 243628 392 243880 480
rect 245532 392 245784 480
rect 247436 392 247688 480
rect 241752 -960 241976 392
rect 243656 -960 243880 392
rect 245560 -960 245784 392
rect 247464 -960 247688 392
rect 248780 420 248836 2326
rect 249228 480 249396 532
rect 249228 476 249592 480
rect 249228 420 249284 476
rect 248780 364 249284 420
rect 249340 392 249592 476
rect 249368 -960 249592 392
rect 250348 420 250404 2326
rect 251132 480 251300 532
rect 253148 480 253204 2326
rect 255052 480 255108 2326
rect 257068 480 257124 2326
rect 258860 480 258916 2326
rect 260764 480 260820 2326
rect 251132 476 251496 480
rect 251132 420 251188 476
rect 250348 364 251188 420
rect 251244 392 251496 476
rect 253148 392 253400 480
rect 255052 392 255304 480
rect 251272 -960 251496 392
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262220 420 262276 2326
rect 262556 480 262724 532
rect 264572 480 264628 2326
rect 262556 476 262920 480
rect 262556 420 262612 476
rect 262220 364 262612 420
rect 262668 392 262920 476
rect 264572 392 264824 480
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 265468 420 265524 2326
rect 266364 480 266532 532
rect 266364 476 266728 480
rect 266364 420 266420 476
rect 265468 364 266420 420
rect 266476 392 266728 476
rect 266504 -960 266728 392
rect 267148 420 267204 2326
rect 268268 480 268436 532
rect 270284 480 270340 2326
rect 272188 480 272244 2326
rect 274092 480 274148 2326
rect 268268 476 268632 480
rect 268268 420 268324 476
rect 267148 364 268324 420
rect 268380 392 268632 476
rect 270284 392 270536 480
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 268408 -960 268632 392
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 275548 420 275604 2326
rect 275884 480 276052 532
rect 277900 480 277956 2326
rect 275884 476 276248 480
rect 275884 420 275940 476
rect 275548 364 275940 420
rect 275996 392 276248 476
rect 277900 392 278152 480
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279020 420 279076 2326
rect 279692 480 279860 532
rect 279692 476 280056 480
rect 279692 420 279748 476
rect 279020 364 279748 420
rect 279804 392 280056 476
rect 279832 -960 280056 392
rect 280588 420 280644 2326
rect 281596 480 281764 532
rect 281596 476 281960 480
rect 281596 420 281652 476
rect 280588 364 281652 420
rect 281708 392 281960 476
rect 281736 -960 281960 392
rect 282268 420 282324 2326
rect 283500 480 283668 532
rect 285740 480 285796 2326
rect 283500 476 283864 480
rect 283500 420 283556 476
rect 282268 364 283556 420
rect 283612 392 283864 476
rect 283640 -960 283864 392
rect 285544 392 285796 480
rect 287420 480 287476 2326
rect 289324 480 289380 2326
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 285544 -960 285768 392
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 290668 420 290724 2326
rect 291116 480 291284 532
rect 291116 476 291480 480
rect 291116 420 291172 476
rect 290668 364 291172 420
rect 291228 392 291480 476
rect 291256 -960 291480 392
rect 292348 420 292404 2326
rect 293020 480 293188 532
rect 293020 476 293384 480
rect 293020 420 293076 476
rect 292348 364 293076 420
rect 293132 392 293384 476
rect 293160 -960 293384 392
rect 294028 420 294084 2326
rect 294924 480 295092 532
rect 294924 476 295288 480
rect 294924 420 294980 476
rect 294028 364 294980 420
rect 295036 392 295288 476
rect 295064 -960 295288 392
rect 295708 420 295764 2326
rect 296828 480 296996 532
rect 296828 476 297192 480
rect 296828 420 296884 476
rect 295708 364 296884 420
rect 296940 392 297192 476
rect 296968 -960 297192 392
rect 297388 420 297444 2326
rect 298732 480 298900 532
rect 300748 480 300804 2326
rect 302652 480 302708 2326
rect 298732 476 299096 480
rect 298732 420 298788 476
rect 297388 364 298788 420
rect 298844 392 299096 476
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304108 420 304164 2326
rect 304444 480 304612 532
rect 304444 476 304808 480
rect 304444 420 304500 476
rect 304108 364 304500 420
rect 304556 392 304808 476
rect 304584 -960 304808 392
rect 305788 420 305844 2326
rect 306348 480 306516 532
rect 306348 476 306712 480
rect 306348 420 306404 476
rect 305788 364 306404 420
rect 306460 392 306712 476
rect 306488 -960 306712 392
rect 307468 420 307524 2326
rect 308252 480 308420 532
rect 308252 476 308616 480
rect 308252 420 308308 476
rect 307468 364 308308 420
rect 308364 392 308616 476
rect 308392 -960 308616 392
rect 309148 420 309204 2326
rect 310156 480 310324 532
rect 310156 476 310520 480
rect 310156 420 310212 476
rect 309148 364 310212 420
rect 310268 392 310520 476
rect 310296 -960 310520 392
rect 310828 420 310884 2326
rect 312060 480 312228 532
rect 314188 480 314244 2326
rect 315980 480 316036 2326
rect 312060 476 312424 480
rect 312060 420 312116 476
rect 310828 364 312116 420
rect 312172 392 312424 476
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 316008 -960 316232 392
rect 317548 420 317604 2326
rect 317772 480 317940 532
rect 319676 480 319844 532
rect 317772 476 318136 480
rect 317772 420 317828 476
rect 317548 364 317828 420
rect 317884 392 318136 476
rect 317912 -960 318136 392
rect 319676 476 320040 480
rect 319676 196 319732 476
rect 319788 392 320040 476
rect 319676 130 319732 140
rect 319816 -960 320040 392
rect 320908 420 320964 2326
rect 321580 480 321748 532
rect 321580 476 321944 480
rect 321580 420 321636 476
rect 320908 364 321636 420
rect 321692 392 321944 476
rect 321720 -960 321944 392
rect 322588 420 322644 2326
rect 323484 480 323652 532
rect 323484 476 323848 480
rect 323484 420 323540 476
rect 322588 364 323540 420
rect 323596 392 323848 476
rect 323624 -960 323848 392
rect 324268 420 324324 2326
rect 325388 480 325556 532
rect 325388 476 325752 480
rect 325388 420 325444 476
rect 324268 364 325444 420
rect 325500 392 325752 476
rect 325528 -960 325752 392
rect 325948 420 326004 2326
rect 327292 480 327460 532
rect 329308 480 329364 2326
rect 331212 480 331268 2326
rect 333116 480 333172 2326
rect 327292 476 327656 480
rect 327292 420 327348 476
rect 325948 364 327348 420
rect 327404 392 327656 476
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 334348 420 334404 2326
rect 334908 480 335076 532
rect 334908 476 335272 480
rect 334908 420 334964 476
rect 334348 364 334964 420
rect 335020 392 335272 476
rect 335048 -960 335272 392
rect 336028 420 336084 2326
rect 336812 480 336980 532
rect 336812 476 337176 480
rect 336812 420 336868 476
rect 336028 364 336868 420
rect 336924 392 337176 476
rect 336952 -960 337176 392
rect 337708 420 337764 2326
rect 338716 480 338884 532
rect 338716 476 339080 480
rect 338716 420 338772 476
rect 337708 364 338772 420
rect 338828 392 339080 476
rect 338856 -960 339080 392
rect 339388 420 339444 2326
rect 340620 480 340788 532
rect 342748 480 342804 2326
rect 344540 480 344596 2326
rect 340620 476 340984 480
rect 340620 420 340676 476
rect 339388 364 340676 420
rect 340732 392 340984 476
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 344568 -960 344792 392
rect 346108 420 346164 2326
rect 346332 480 346500 532
rect 346332 476 346696 480
rect 346332 420 346388 476
rect 346108 364 346388 420
rect 346444 392 346696 476
rect 346472 -960 346696 392
rect 347788 420 347844 2326
rect 348236 480 348404 532
rect 350252 480 350308 2326
rect 348236 476 348600 480
rect 348236 420 348292 476
rect 347788 364 348292 420
rect 348348 392 348600 476
rect 350252 392 350504 480
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 351148 420 351204 2326
rect 352044 480 352212 532
rect 352044 476 352408 480
rect 352044 420 352100 476
rect 351148 364 352100 420
rect 352156 392 352408 476
rect 352184 -960 352408 392
rect 352828 420 352884 2326
rect 353948 480 354116 532
rect 353948 476 354312 480
rect 353948 420 354004 476
rect 352828 364 354004 420
rect 354060 392 354312 476
rect 354088 -960 354312 392
rect 354508 420 354564 2326
rect 355852 480 356020 532
rect 357868 480 357924 2326
rect 359772 480 359828 2326
rect 361676 480 361732 2326
rect 355852 476 356216 480
rect 355852 420 355908 476
rect 354508 364 355908 420
rect 355964 392 356216 476
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 362908 420 362964 2326
rect 363468 480 363636 532
rect 365484 480 365540 2326
rect 367388 480 367444 2326
rect 369292 480 369348 2326
rect 371308 480 371364 2326
rect 373100 480 373156 2326
rect 374892 480 375060 532
rect 363468 476 363832 480
rect 363468 420 363524 476
rect 362908 364 363524 420
rect 363580 392 363832 476
rect 365484 392 365736 480
rect 367388 392 367640 480
rect 369292 392 369544 480
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373100 392 373352 480
rect 373128 -960 373352 392
rect 374892 476 375256 480
rect 374892 84 374948 476
rect 375004 392 375256 476
rect 374892 18 374948 28
rect 375032 -960 375256 392
rect 376348 420 376404 2326
rect 376796 480 376964 532
rect 376796 476 377160 480
rect 376796 420 376852 476
rect 376348 364 376852 420
rect 376908 392 377160 476
rect 376936 -960 377160 392
rect 378028 420 378084 2326
rect 378700 480 378868 532
rect 378700 476 379064 480
rect 378700 420 378756 476
rect 378028 364 378756 420
rect 378812 392 379064 476
rect 378840 -960 379064 392
rect 379708 420 379764 2326
rect 380604 480 380772 532
rect 380604 476 380968 480
rect 380604 420 380660 476
rect 379708 364 380660 420
rect 380716 392 380968 476
rect 380744 -960 380968 392
rect 381388 420 381444 2326
rect 382508 480 382676 532
rect 384524 480 384580 2326
rect 386428 480 386484 2326
rect 388332 480 388388 2326
rect 382508 476 382872 480
rect 382508 420 382564 476
rect 381388 364 382564 420
rect 382620 392 382872 476
rect 384524 392 384776 480
rect 386428 392 386680 480
rect 388332 392 388584 480
rect 382648 -960 382872 392
rect 384552 -960 384776 392
rect 386456 -960 386680 392
rect 388360 -960 388584 392
rect 389788 420 389844 2326
rect 390124 480 390292 532
rect 390124 476 390488 480
rect 390124 420 390180 476
rect 389788 364 390180 420
rect 390236 392 390488 476
rect 390264 -960 390488 392
rect 391468 420 391524 2326
rect 392028 480 392196 532
rect 392028 476 392392 480
rect 392028 420 392084 476
rect 391468 364 392084 420
rect 392140 392 392392 476
rect 392168 -960 392392 392
rect 393148 420 393204 2326
rect 393932 480 394100 532
rect 393932 476 394296 480
rect 393932 420 393988 476
rect 393148 364 393988 420
rect 394044 392 394296 476
rect 394072 -960 394296 392
rect 394828 420 394884 2326
rect 395836 480 396004 532
rect 395836 476 396200 480
rect 395836 420 395892 476
rect 394828 364 395892 420
rect 395948 392 396200 476
rect 395976 -960 396200 392
rect 396508 420 396564 2326
rect 397740 480 397908 532
rect 399868 480 399924 2326
rect 401660 480 401716 2326
rect 397740 476 398104 480
rect 397740 420 397796 476
rect 396508 364 397796 420
rect 397852 392 398104 476
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401660 392 401912 480
rect 401688 -960 401912 392
rect 403228 420 403284 2326
rect 403452 480 403620 532
rect 405468 480 405524 2326
rect 403452 476 403816 480
rect 403452 420 403508 476
rect 403228 364 403508 420
rect 403564 392 403816 476
rect 405468 392 405720 480
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 406588 420 406644 2326
rect 407260 480 407428 532
rect 407260 476 407624 480
rect 407260 420 407316 476
rect 406588 364 407316 420
rect 407372 392 407624 476
rect 407400 -960 407624 392
rect 408268 420 408324 2326
rect 409164 480 409332 532
rect 409164 476 409528 480
rect 409164 420 409220 476
rect 408268 364 409220 420
rect 409276 392 409528 476
rect 409304 -960 409528 392
rect 409948 420 410004 2326
rect 411068 480 411236 532
rect 411068 476 411432 480
rect 411068 420 411124 476
rect 409948 364 411124 420
rect 411180 392 411432 476
rect 411208 -960 411432 392
rect 411628 420 411684 2326
rect 412972 480 413140 532
rect 414988 480 415044 2326
rect 416892 480 416948 2326
rect 418796 480 418852 2326
rect 412972 476 413336 480
rect 412972 420 413028 476
rect 411628 364 413028 420
rect 413084 392 413336 476
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 418796 392 419048 480
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 -960 419048 392
rect 420028 420 420084 2326
rect 420588 480 420756 532
rect 420588 476 420952 480
rect 420588 420 420644 476
rect 420028 364 420644 420
rect 420700 392 420952 476
rect 420728 -960 420952 392
rect 421708 420 421764 2326
rect 422492 480 422660 532
rect 422492 476 422856 480
rect 422492 420 422548 476
rect 421708 364 422548 420
rect 422604 392 422856 476
rect 422632 -960 422856 392
rect 423388 420 423444 2326
rect 424396 480 424564 532
rect 424396 476 424760 480
rect 424396 420 424452 476
rect 423388 364 424452 420
rect 424508 392 424760 476
rect 424536 -960 424760 392
rect 425068 420 425124 2326
rect 426300 480 426468 532
rect 428428 480 428484 2326
rect 430220 480 430276 2326
rect 426300 476 426664 480
rect 426300 420 426356 476
rect 425068 364 426356 420
rect 426412 392 426664 476
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430220 392 430472 480
rect 430248 -960 430472 392
rect 431788 420 431844 2326
rect 432012 480 432180 532
rect 432012 476 432376 480
rect 432012 420 432068 476
rect 431788 364 432068 420
rect 432124 392 432376 476
rect 432152 -960 432376 392
rect 433468 420 433524 2326
rect 433916 480 434084 532
rect 435932 480 435988 2326
rect 433916 476 434280 480
rect 433916 420 433972 476
rect 433468 364 433972 420
rect 434028 392 434280 476
rect 435932 392 436184 480
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 436828 420 436884 2326
rect 437724 480 437892 532
rect 437724 476 438088 480
rect 437724 420 437780 476
rect 436828 364 437780 420
rect 437836 392 438088 476
rect 437864 -960 438088 392
rect 438508 420 438564 2326
rect 439628 480 439796 532
rect 441644 480 441700 2326
rect 443548 480 443604 2326
rect 445452 480 445508 2326
rect 439628 476 439992 480
rect 439628 420 439684 476
rect 438508 364 439684 420
rect 439740 392 439992 476
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 446908 420 446964 2326
rect 447244 480 447412 532
rect 447244 476 447608 480
rect 447244 420 447300 476
rect 446908 364 447300 420
rect 447356 392 447608 476
rect 447384 -960 447608 392
rect 448588 420 448644 2326
rect 449148 480 449316 532
rect 449148 476 449512 480
rect 449148 420 449204 476
rect 448588 364 449204 420
rect 449260 392 449512 476
rect 449288 -960 449512 392
rect 450268 420 450324 2326
rect 451052 480 451220 532
rect 451052 476 451416 480
rect 451052 420 451108 476
rect 450268 364 451108 420
rect 451164 392 451416 476
rect 451192 -960 451416 392
rect 451948 420 452004 2326
rect 452956 480 453124 532
rect 452956 476 453320 480
rect 452956 420 453012 476
rect 451948 364 453012 420
rect 453068 392 453320 476
rect 453096 -960 453320 392
rect 453628 420 453684 2326
rect 454860 480 455028 532
rect 456988 480 457044 2326
rect 458780 480 458836 2326
rect 454860 476 455224 480
rect 454860 420 454916 476
rect 453628 364 454916 420
rect 454972 392 455224 476
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 458808 -960 459032 392
rect 460348 420 460404 2326
rect 460572 480 460740 532
rect 460572 476 460936 480
rect 460572 420 460628 476
rect 460348 364 460628 420
rect 460684 392 460936 476
rect 460712 -960 460936 392
rect 462028 420 462084 2326
rect 462476 480 462644 532
rect 462476 476 462840 480
rect 462476 420 462532 476
rect 462028 364 462532 420
rect 462588 392 462840 476
rect 462616 -960 462840 392
rect 463708 420 463764 2326
rect 464380 480 464548 532
rect 464380 476 464744 480
rect 464380 420 464436 476
rect 463708 364 464436 420
rect 464492 392 464744 476
rect 464520 -960 464744 392
rect 465388 420 465444 2326
rect 466284 480 466452 532
rect 466284 476 466648 480
rect 466284 420 466340 476
rect 465388 364 466340 420
rect 466396 392 466648 476
rect 466424 -960 466648 392
rect 467068 420 467124 2326
rect 468188 480 468356 532
rect 468188 476 468552 480
rect 468188 420 468244 476
rect 467068 364 468244 420
rect 468300 392 468552 476
rect 468328 -960 468552 392
rect 468748 420 468804 2326
rect 470092 480 470260 532
rect 472108 480 472164 2326
rect 474012 480 474068 2326
rect 475916 480 475972 2326
rect 470092 476 470456 480
rect 470092 420 470148 476
rect 468748 364 470148 420
rect 470204 392 470456 476
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 475916 392 476168 480
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475944 -960 476168 392
rect 477148 420 477204 2326
rect 477708 480 477876 532
rect 477708 476 478072 480
rect 477708 420 477764 476
rect 477148 364 477764 420
rect 477820 392 478072 476
rect 477848 -960 478072 392
rect 478828 420 478884 2326
rect 479612 480 479780 532
rect 479612 476 479976 480
rect 479612 420 479668 476
rect 478828 364 479668 420
rect 479724 392 479976 476
rect 479752 -960 479976 392
rect 480508 420 480564 2326
rect 481516 480 481684 532
rect 481516 476 481880 480
rect 481516 420 481572 476
rect 480508 364 481572 420
rect 481628 392 481880 476
rect 481656 -960 481880 392
rect 482188 420 482244 2326
rect 483420 480 483588 532
rect 485548 480 485604 2326
rect 487340 480 487396 2326
rect 483420 476 483784 480
rect 483420 420 483476 476
rect 482188 364 483476 420
rect 483532 392 483784 476
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 487368 -960 487592 392
rect 488908 420 488964 2326
rect 489132 480 489300 532
rect 491148 480 491204 2326
rect 489132 476 489496 480
rect 489132 420 489188 476
rect 488908 364 489188 420
rect 489244 392 489496 476
rect 491148 392 491400 480
rect 489272 -960 489496 392
rect 491176 -960 491400 392
rect 492268 420 492324 2326
rect 492940 480 493108 532
rect 494956 480 495012 2326
rect 492940 476 493304 480
rect 492940 420 492996 476
rect 492268 364 492996 420
rect 493052 392 493304 476
rect 494956 392 495208 480
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 495628 420 495684 2326
rect 496748 480 496916 532
rect 496748 476 497112 480
rect 496748 420 496804 476
rect 495628 364 496804 420
rect 496860 392 497112 476
rect 496888 -960 497112 392
rect 497308 420 497364 2326
rect 498652 480 498820 532
rect 500668 480 500724 2326
rect 502572 480 502628 2326
rect 498652 476 499016 480
rect 498652 420 498708 476
rect 497308 364 498708 420
rect 498764 392 499016 476
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504028 420 504084 2326
rect 504364 480 504532 532
rect 504364 476 504728 480
rect 504364 420 504420 476
rect 504028 364 504420 420
rect 504476 392 504728 476
rect 504504 -960 504728 392
rect 505708 420 505764 2326
rect 506268 480 506436 532
rect 506268 476 506632 480
rect 506268 420 506324 476
rect 505708 364 506324 420
rect 506380 392 506632 476
rect 506408 -960 506632 392
rect 507388 420 507444 2326
rect 508172 480 508340 532
rect 510188 480 510244 2326
rect 508172 476 508536 480
rect 508172 420 508228 476
rect 507388 364 508228 420
rect 508284 392 508536 476
rect 510188 392 510440 480
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 510748 420 510804 2326
rect 511980 480 512148 532
rect 514108 480 514164 2326
rect 515900 480 515956 2326
rect 511980 476 512344 480
rect 511980 420 512036 476
rect 510748 364 512036 420
rect 512092 392 512344 476
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 515928 -960 516152 392
rect 517468 420 517524 2326
rect 517692 480 517860 532
rect 517692 476 518056 480
rect 517692 420 517748 476
rect 517468 364 517748 420
rect 517804 392 518056 476
rect 517832 -960 518056 392
rect 519148 420 519204 2326
rect 519596 480 519764 532
rect 519596 476 519960 480
rect 519596 420 519652 476
rect 519148 364 519652 420
rect 519708 392 519960 476
rect 519736 -960 519960 392
rect 520828 420 520884 2326
rect 521500 480 521668 532
rect 521500 476 521864 480
rect 521500 420 521556 476
rect 520828 364 521556 420
rect 521612 392 521864 476
rect 521640 -960 521864 392
rect 522508 420 522564 2326
rect 523404 480 523572 532
rect 523404 476 523768 480
rect 523404 420 523460 476
rect 522508 364 523460 420
rect 523516 392 523768 476
rect 523544 -960 523768 392
rect 524188 420 524244 2326
rect 525308 480 525476 532
rect 527324 480 527380 2326
rect 529228 480 529284 2326
rect 531132 480 531188 2326
rect 525308 476 525672 480
rect 525308 420 525364 476
rect 524188 364 525364 420
rect 525420 392 525672 476
rect 527324 392 527576 480
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 532588 420 532644 2326
rect 532924 480 533092 532
rect 532924 476 533288 480
rect 532924 420 532980 476
rect 532588 364 532980 420
rect 533036 392 533288 476
rect 533064 -960 533288 392
rect 534268 420 534324 2326
rect 534828 480 534996 532
rect 534828 476 535192 480
rect 534828 420 534884 476
rect 534268 364 534884 420
rect 534940 392 535192 476
rect 534968 -960 535192 392
rect 535948 420 536004 2326
rect 536732 480 536900 532
rect 536732 476 537096 480
rect 536732 420 536788 476
rect 535948 364 536788 420
rect 536844 392 537096 476
rect 536872 -960 537096 392
rect 537628 420 537684 2326
rect 538636 480 538804 532
rect 538636 476 539000 480
rect 538636 420 538692 476
rect 537628 364 538692 420
rect 538748 392 539000 476
rect 538776 -960 539000 392
rect 539308 420 539364 2326
rect 540540 480 540708 532
rect 542668 480 542724 2326
rect 544460 480 544516 2326
rect 540540 476 540904 480
rect 540540 420 540596 476
rect 539308 364 540596 420
rect 540652 392 540904 476
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 544488 -960 544712 392
rect 546028 420 546084 2326
rect 546252 480 546420 532
rect 548268 480 548324 2326
rect 546252 476 546616 480
rect 546252 420 546308 476
rect 546028 364 546308 420
rect 546364 392 546616 476
rect 548268 392 548520 480
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 549388 420 549444 2326
rect 550060 480 550228 532
rect 550060 476 550424 480
rect 550060 420 550116 476
rect 549388 364 550116 420
rect 550172 392 550424 476
rect 550200 -960 550424 392
rect 551068 420 551124 2326
rect 551964 480 552132 532
rect 551964 476 552328 480
rect 551964 420 552020 476
rect 551068 364 552020 420
rect 552076 392 552328 476
rect 552104 -960 552328 392
rect 552748 420 552804 2326
rect 553868 480 554036 532
rect 553868 476 554232 480
rect 553868 420 553924 476
rect 552748 364 553924 420
rect 553980 392 554232 476
rect 554008 -960 554232 392
rect 554428 420 554484 2326
rect 555772 480 555940 532
rect 557788 480 557844 2326
rect 559692 480 559748 2326
rect 561596 480 561652 2326
rect 563500 480 563556 2326
rect 555772 476 556136 480
rect 555772 420 555828 476
rect 554428 364 555828 420
rect 555884 392 556136 476
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 563500 392 563752 480
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 -960 563752 392
rect 564508 420 564564 2326
rect 565292 480 565460 532
rect 567308 480 567364 2326
rect 565292 476 565656 480
rect 565292 420 565348 476
rect 564508 364 565348 420
rect 565404 392 565656 476
rect 567308 392 567560 480
rect 565432 -960 565656 392
rect 567336 -960 567560 392
rect 567868 420 567924 2326
rect 569100 480 569268 532
rect 571228 480 571284 2326
rect 573020 480 573076 2326
rect 569100 476 569464 480
rect 569100 420 569156 476
rect 567868 364 569156 420
rect 569212 392 569464 476
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 573048 -960 573272 392
rect 574588 420 574644 2326
rect 574812 480 574980 532
rect 574812 476 575176 480
rect 574812 420 574868 476
rect 574588 364 574868 420
rect 574924 392 575176 476
rect 574952 -960 575176 392
rect 576268 420 576324 2326
rect 576716 480 576884 532
rect 576716 476 577080 480
rect 576716 420 576772 476
rect 576268 364 576772 420
rect 576828 392 577080 476
rect 576856 -960 577080 392
rect 577948 420 578004 2326
rect 578620 480 578788 532
rect 582540 480 582596 2326
rect 578620 476 578984 480
rect 578620 420 578676 476
rect 577948 364 578676 420
rect 578732 392 578984 476
rect 578760 -960 578984 392
rect 580664 -960 580888 480
rect 582540 392 582792 480
rect 582568 -960 582792 392
rect 582988 420 583044 2326
rect 584332 480 584500 532
rect 586348 480 586404 2326
rect 584332 476 584696 480
rect 584332 420 584388 476
rect 582988 364 584388 420
rect 584444 392 584696 476
rect 586348 392 586600 480
rect 584472 -960 584696 392
rect 586376 -960 586600 392
<< via2 >>
rect 188188 598108 188244 598164
rect 588140 598108 588196 598164
rect 598108 579740 598164 579796
rect 4172 534492 4228 534548
rect 4396 477596 4452 477652
rect 4284 434924 4340 434980
rect 4284 304892 4340 304948
rect 4172 291900 4228 291956
rect 4284 300748 4340 300804
rect 4172 130172 4228 130228
rect 595756 406588 595812 406644
rect 4396 291788 4452 291844
rect 4620 363804 4676 363860
rect 595644 312508 595700 312564
rect 595532 307468 595588 307524
rect 4620 291676 4676 291732
rect 4844 306908 4900 306964
rect 4844 291564 4900 291620
rect 595756 306572 595812 306628
rect 595868 315868 595924 315924
rect 595980 314188 596036 314244
rect 596092 313180 596148 313236
rect 598108 303212 598164 303268
rect 596092 291452 596148 291508
rect 595980 260092 596036 260148
rect 595868 219996 595924 220052
rect 595644 153468 595700 153524
rect 595532 126812 595588 126868
rect 595644 141932 595700 141988
rect 4284 79548 4340 79604
rect 4172 65324 4228 65380
rect 595644 33516 595700 33572
rect 214060 140 214116 196
rect 228844 28 228900 84
rect 319676 140 319732 196
rect 374892 28 374948 84
<< metal3 >>
rect 188178 598108 188188 598164
rect 188244 598108 588140 598164
rect 588196 598108 588206 598164
rect 599520 593124 600960 593320
rect 595211 593096 600960 593124
rect 595211 593068 599592 593096
rect -960 591444 480 591640
rect -960 591416 6134 591444
rect 392 591388 6134 591416
rect 599520 579796 600960 579992
rect 598098 579740 598108 579796
rect 598164 579768 600960 579796
rect 598164 579740 599592 579768
rect -960 577220 480 577416
rect -960 577192 532 577220
rect 392 577164 532 577192
rect 476 577108 532 577164
rect 364 577052 532 577108
rect 364 576324 420 577052
rect 364 576268 6134 576324
rect 599520 566468 600960 566664
rect 595211 566440 600960 566468
rect 595211 566412 599592 566440
rect -960 562996 480 563192
rect -960 562968 6134 562996
rect 392 562940 6134 562968
rect 599520 553140 600960 553336
rect 599452 553112 600960 553140
rect 599452 553084 599592 553112
rect 599452 553028 599508 553084
rect 599452 552972 599620 553028
rect 599564 552804 599620 552972
rect 595211 552748 599620 552804
rect -960 548772 480 548968
rect -960 548744 532 548772
rect 392 548716 532 548744
rect 476 548660 532 548716
rect 364 548604 532 548660
rect 364 547764 420 548604
rect 364 547708 6134 547764
rect 599520 539812 600960 540008
rect 599452 539784 600960 539812
rect 599452 539756 599592 539784
rect 599452 539700 599508 539756
rect 599452 539644 599620 539700
rect 599564 539364 599620 539644
rect 595211 539308 599620 539364
rect -960 534548 480 534744
rect -960 534520 4172 534548
rect 392 534492 4172 534520
rect 4228 534492 4238 534548
rect 599520 526484 600960 526680
rect 599452 526456 600960 526484
rect 599452 526428 599592 526456
rect 599452 526372 599508 526428
rect 599452 526316 599620 526372
rect 599564 525924 599620 526316
rect 595211 525868 599620 525924
rect -960 520324 480 520520
rect -960 520296 532 520324
rect 392 520268 532 520296
rect 476 520212 532 520268
rect 364 520156 532 520212
rect 364 519204 420 520156
rect 364 519148 6134 519204
rect 599520 513156 600960 513352
rect 599452 513128 600960 513156
rect 599452 513100 599592 513128
rect 599452 513044 599508 513100
rect 599452 512988 599620 513044
rect 599564 512484 599620 512988
rect 595211 512428 599620 512484
rect -960 506100 480 506296
rect -960 506072 532 506100
rect 392 506044 532 506072
rect 476 505988 532 506044
rect 364 505932 532 505988
rect 364 505764 420 505932
rect 364 505708 6134 505764
rect 599520 499828 600960 500024
rect 599452 499800 600960 499828
rect 599452 499772 599592 499800
rect 599452 499716 599508 499772
rect 599452 499660 599620 499716
rect 599564 499044 599620 499660
rect 595211 498988 599620 499044
rect -960 491876 480 492072
rect -960 491848 532 491876
rect 392 491820 532 491848
rect 476 491764 532 491820
rect 364 491708 532 491764
rect 364 490644 420 491708
rect 364 490588 6134 490644
rect 599520 486500 600960 486696
rect 599452 486472 600960 486500
rect 599452 486444 599592 486472
rect 599452 486388 599508 486444
rect 599452 486332 599620 486388
rect 599564 485604 599620 486332
rect 595211 485548 599620 485604
rect -960 477652 480 477848
rect -960 477624 4396 477652
rect 392 477596 4396 477624
rect 4452 477596 4462 477652
rect 599520 473172 600960 473368
rect 599452 473144 600960 473172
rect 599452 473116 599592 473144
rect 599452 473060 599508 473116
rect 599452 473004 599620 473060
rect 599564 472164 599620 473004
rect 595211 472108 599620 472164
rect -960 463428 480 463624
rect -960 463400 532 463428
rect 392 463372 532 463400
rect 476 463316 532 463372
rect 364 463260 532 463316
rect 364 462084 420 463260
rect 364 462028 6134 462084
rect 599520 459844 600960 460040
rect 599452 459816 600960 459844
rect 599452 459788 599592 459816
rect 599452 459732 599508 459788
rect 599452 459676 599620 459732
rect 599564 458724 599620 459676
rect 595211 458668 599620 458724
rect -960 449204 480 449400
rect -960 449176 532 449204
rect 392 449148 532 449176
rect 476 449092 532 449148
rect 364 449036 532 449092
rect 364 448644 420 449036
rect 364 448588 6134 448644
rect 599520 446516 600960 446712
rect 599452 446488 600960 446516
rect 599452 446460 599592 446488
rect 599452 446404 599508 446460
rect 599452 446348 599620 446404
rect 599564 445284 599620 446348
rect 595211 445228 599620 445284
rect -960 434980 480 435176
rect -960 434952 4284 434980
rect 392 434924 4284 434952
rect 4340 434924 4350 434980
rect 599520 433188 600960 433384
rect 599452 433160 600960 433188
rect 599452 433132 599592 433160
rect 599452 433076 599508 433132
rect 599452 433020 599620 433076
rect 599564 431844 599620 433020
rect 595211 431788 599620 431844
rect -960 420756 480 420952
rect -960 420728 532 420756
rect 392 420700 532 420728
rect 476 420644 532 420700
rect 364 420588 532 420644
rect 364 420084 420 420588
rect 364 420028 6134 420084
rect 599520 419860 600960 420056
rect 599452 419832 600960 419860
rect 599452 419804 599592 419832
rect 599452 419748 599508 419804
rect 599452 419692 599620 419748
rect 599564 418404 599620 419692
rect 595211 418348 599620 418404
rect -960 406644 480 406728
rect 599520 406644 600960 406728
rect -960 406588 6134 406644
rect 595746 406588 595756 406644
rect 595812 406588 600960 406644
rect -960 406504 480 406588
rect 599520 406504 600960 406588
rect 599520 393204 600960 393400
rect 595211 393176 600960 393204
rect 595211 393148 599592 393176
rect -960 392308 480 392504
rect -960 392280 532 392308
rect 392 392252 532 392280
rect 476 392196 532 392252
rect 364 392140 532 392196
rect 364 391524 420 392140
rect 364 391468 6134 391524
rect 599520 379876 600960 380072
rect 595211 379848 600960 379876
rect 595211 379820 599592 379848
rect -960 378084 480 378280
rect -960 378056 6134 378084
rect 392 378028 6134 378056
rect 599520 366548 600960 366744
rect 595211 366520 600960 366548
rect 595211 366492 599592 366520
rect -960 363860 480 364056
rect -960 363832 4620 363860
rect 392 363804 4620 363832
rect 4676 363804 4686 363860
rect 599520 353220 600960 353416
rect 599452 353192 600960 353220
rect 599452 353164 599592 353192
rect 599452 353108 599508 353164
rect 599452 353052 599620 353108
rect 599564 352884 599620 353052
rect 595211 352828 599620 352884
rect -960 349636 480 349832
rect -960 349608 6134 349636
rect 392 349580 6134 349608
rect 599520 339892 600960 340088
rect 599452 339864 600960 339892
rect 599452 339836 599592 339864
rect 599452 339780 599508 339836
rect 599452 339724 599620 339780
rect 599564 339444 599620 339724
rect 595211 339388 599620 339444
rect -960 335412 480 335608
rect -960 335384 532 335412
rect 392 335356 532 335384
rect 476 335300 532 335356
rect 364 335244 532 335300
rect 364 334404 420 335244
rect 364 334348 6134 334404
rect 599520 326564 600960 326760
rect 599452 326536 600960 326564
rect 599452 326508 599592 326536
rect 599452 326452 599508 326508
rect 599452 326396 599620 326452
rect 599564 326004 599620 326396
rect 595211 325948 599620 326004
rect -960 321188 480 321384
rect -960 321160 6134 321188
rect 392 321132 6134 321160
rect 595211 315868 595868 315924
rect 595924 315868 595934 315924
rect 595211 314188 595980 314244
rect 596036 314188 596046 314244
rect 599520 313236 600960 313432
rect 596082 313180 596092 313236
rect 596148 313208 600960 313236
rect 596148 313180 599592 313208
rect 595211 312508 595644 312564
rect 595700 312508 595710 312564
rect 595211 307468 595532 307524
rect 595588 307468 595598 307524
rect -960 306964 480 307160
rect -960 306936 4844 306964
rect 392 306908 4844 306936
rect 4900 306908 4910 306964
rect 595211 306572 595756 306628
rect 595812 306572 595822 306628
rect 4274 304892 4284 304948
rect 4340 304892 6134 304948
rect 595211 303212 598108 303268
rect 598164 303212 598174 303268
rect 4274 300748 4284 300804
rect 4340 300748 6134 300804
rect 599520 299908 600960 300104
rect 599452 299880 600960 299908
rect 599452 299852 599592 299880
rect 599452 299796 599508 299852
rect 599452 299740 599620 299796
rect 599564 299124 599620 299740
rect 595211 299068 599620 299124
rect -960 292740 480 292936
rect -960 292712 532 292740
rect 392 292684 532 292712
rect 476 292628 532 292684
rect 364 292572 532 292628
rect 364 292404 420 292572
rect 364 292348 6134 292404
rect 4162 291900 4172 291956
rect 4228 291900 6134 291956
rect 4386 291788 4396 291844
rect 4452 291788 6134 291844
rect 4610 291676 4620 291732
rect 4676 291676 6134 291732
rect 4834 291564 4844 291620
rect 4900 291564 6134 291620
rect 595211 291452 596092 291508
rect 596148 291452 596158 291508
rect 599520 286580 600960 286776
rect 595211 286552 600960 286580
rect 595211 286524 599592 286552
rect -960 278516 480 278712
rect -960 278488 532 278516
rect 392 278460 532 278488
rect 476 278404 532 278460
rect 364 278348 532 278404
rect 364 277284 420 278348
rect 364 277228 6134 277284
rect 599520 273252 600960 273448
rect 599452 273224 600960 273252
rect 599452 273196 599592 273224
rect 599452 273140 599508 273196
rect 599452 273084 599620 273140
rect 599564 272244 599620 273084
rect 595211 272188 599620 272244
rect -960 264292 480 264488
rect -960 264264 532 264292
rect 392 264236 532 264264
rect 476 264180 532 264236
rect 364 264124 532 264180
rect 364 263844 420 264124
rect 364 263788 6134 263844
rect 595970 260092 595980 260148
rect 596036 260120 599592 260148
rect 596036 260092 600960 260120
rect 599520 259896 600960 260092
rect -960 250068 480 250264
rect -960 250040 532 250068
rect 392 250012 532 250040
rect 476 249956 532 250012
rect 364 249900 532 249956
rect 364 248724 420 249900
rect 364 248668 6134 248724
rect 599520 246596 600960 246792
rect 599452 246568 600960 246596
rect 599452 246540 599592 246568
rect 599452 246484 599508 246540
rect 599452 246428 599620 246484
rect 599564 245364 599620 246428
rect 595211 245308 599620 245364
rect -960 235844 480 236040
rect -960 235816 532 235844
rect 392 235788 532 235816
rect 476 235732 532 235788
rect 364 235676 532 235732
rect 364 235284 420 235676
rect 364 235228 6134 235284
rect 599520 233268 600960 233464
rect 599452 233240 600960 233268
rect 599452 233212 599592 233240
rect 599452 233156 599508 233212
rect 599452 233100 599620 233156
rect 599564 231924 599620 233100
rect 595211 231868 599620 231924
rect -960 221732 480 221816
rect -960 221676 6134 221732
rect -960 221592 480 221676
rect 599520 220052 600960 220136
rect 595858 219996 595868 220052
rect 595924 219996 600960 220052
rect 599520 219912 600960 219996
rect -960 207396 480 207592
rect -960 207368 532 207396
rect 392 207340 532 207368
rect 476 207284 532 207340
rect 364 207228 532 207284
rect 364 206724 420 207228
rect 599520 206724 600960 206808
rect 364 206668 6134 206724
rect 595211 206668 600960 206724
rect 599520 206584 600960 206668
rect -960 193284 480 193368
rect 599520 193284 600960 193480
rect -960 193228 6134 193284
rect 595211 193256 600960 193284
rect 595211 193228 599592 193256
rect -960 193144 480 193228
rect 599520 179956 600960 180152
rect 595211 179928 600960 179956
rect 595211 179900 599592 179928
rect -960 178948 480 179144
rect -960 178920 532 178948
rect 392 178892 532 178920
rect 476 178836 532 178892
rect 364 178780 532 178836
rect 364 178164 420 178780
rect 364 178108 6134 178164
rect 599520 166628 600960 166824
rect 595211 166600 600960 166628
rect 595211 166572 599592 166600
rect -960 164724 480 164920
rect -960 164696 6134 164724
rect 392 164668 6134 164696
rect 595634 153468 595644 153524
rect 595700 153496 599592 153524
rect 595700 153468 600960 153496
rect 599520 153272 600960 153468
rect -960 150500 480 150696
rect -960 150472 532 150500
rect 392 150444 532 150472
rect 476 150388 532 150444
rect 364 150332 532 150388
rect 364 149604 420 150332
rect 364 149548 6134 149604
rect 595211 141932 595644 141988
rect 595700 141932 595710 141988
rect 599520 139972 600960 140168
rect 599452 139944 600960 139972
rect 599452 139916 599592 139944
rect 599452 139860 599508 139916
rect 599452 139804 599620 139860
rect 599564 139524 599620 139804
rect 595211 139468 599620 139524
rect -960 136276 480 136472
rect -960 136248 6134 136276
rect 392 136220 6134 136248
rect 4162 130172 4172 130228
rect 4228 130172 6134 130228
rect 595522 126812 595532 126868
rect 595588 126840 599592 126868
rect 595588 126812 600960 126840
rect 599520 126616 600960 126812
rect -960 122052 480 122248
rect -960 122024 532 122052
rect 392 121996 532 122024
rect 476 121940 532 121996
rect 364 121884 532 121940
rect 364 121044 420 121884
rect 364 120988 6134 121044
rect 599520 113316 600960 113512
rect 599452 113288 600960 113316
rect 599452 113260 599592 113288
rect 599452 113204 599508 113260
rect 599452 113148 599620 113204
rect 599564 112644 599620 113148
rect 595211 112588 599620 112644
rect -960 107828 480 108024
rect -960 107800 6134 107828
rect 392 107772 6134 107800
rect 599520 99988 600960 100184
rect 599452 99960 600960 99988
rect 599452 99932 599592 99960
rect 599452 99876 599508 99932
rect 599452 99820 599620 99876
rect 599564 99204 599620 99820
rect 595211 99148 599620 99204
rect -960 93604 480 93800
rect -960 93576 532 93604
rect 392 93548 532 93576
rect 476 93492 532 93548
rect 364 93436 532 93492
rect 364 92484 420 93436
rect 364 92428 6134 92484
rect 599520 86660 600960 86856
rect 599452 86632 600960 86660
rect 599452 86604 599592 86632
rect 599452 86548 599508 86604
rect 599452 86492 599620 86548
rect 599564 85764 599620 86492
rect 595211 85708 599620 85764
rect 392 79576 4284 79604
rect -960 79548 4284 79576
rect 4340 79548 4350 79604
rect -960 79352 480 79548
rect 599520 73332 600960 73528
rect 599452 73304 600960 73332
rect 599452 73276 599592 73304
rect 599452 73220 599508 73276
rect 599452 73164 599620 73220
rect 599564 72324 599620 73164
rect 595211 72268 599620 72324
rect 392 65352 4172 65380
rect -960 65324 4172 65352
rect 4228 65324 4238 65380
rect -960 65128 480 65324
rect 599520 60004 600960 60200
rect 599452 59976 600960 60004
rect 599452 59948 599592 59976
rect 599452 59892 599508 59948
rect 599452 59836 599620 59892
rect 599564 58884 599620 59836
rect 595211 58828 599620 58884
rect -960 50932 480 51128
rect -960 50904 532 50932
rect 392 50876 532 50904
rect 476 50820 532 50876
rect 364 50764 532 50820
rect 364 50484 420 50764
rect 364 50428 6134 50484
rect 595211 46872 599592 46900
rect 595211 46844 600960 46872
rect 599520 46648 600960 46844
rect -960 36708 480 36904
rect -960 36680 532 36708
rect 392 36652 532 36680
rect 476 36596 532 36652
rect 364 36540 532 36596
rect 364 35364 420 36540
rect 364 35308 6134 35364
rect 595634 33516 595644 33572
rect 595700 33544 599592 33572
rect 595700 33516 600960 33544
rect 599520 33320 600960 33516
rect -960 22484 480 22680
rect -960 22456 532 22484
rect 392 22428 532 22456
rect 476 22372 532 22428
rect 364 22316 532 22372
rect 364 21924 420 22316
rect 364 21868 6134 21924
rect 599520 20020 600960 20216
rect 599452 19992 600960 20020
rect 599452 19964 599592 19992
rect 599452 19908 599508 19964
rect 599452 19852 599620 19908
rect 599564 18564 599620 19852
rect 595211 18508 599620 18564
rect -960 8372 480 8456
rect -960 8316 6134 8372
rect -960 8232 480 8316
rect 595211 6888 599592 6916
rect 595211 6860 600960 6888
rect 599520 6664 600960 6860
rect 214050 140 214060 196
rect 214116 140 319676 196
rect 319732 140 319742 196
rect 228834 28 228844 84
rect 228900 28 374892 84
rect 374948 28 374958 84
<< metal4 >>
rect -12 599340 608 599436
rect -12 599284 84 599340
rect 140 599284 208 599340
rect 264 599284 332 599340
rect 388 599284 456 599340
rect 512 599284 608 599340
rect -12 599216 608 599284
rect -12 599160 84 599216
rect 140 599160 208 599216
rect 264 599160 332 599216
rect 388 599160 456 599216
rect 512 599160 608 599216
rect -12 599092 608 599160
rect -12 599036 84 599092
rect 140 599036 208 599092
rect 264 599036 332 599092
rect 388 599036 456 599092
rect 512 599036 608 599092
rect -12 598968 608 599036
rect -12 598912 84 598968
rect 140 598912 208 598968
rect 264 598912 332 598968
rect 388 598912 456 598968
rect 512 598912 608 598968
rect -12 587918 608 598912
rect -12 587862 84 587918
rect 140 587862 208 587918
rect 264 587862 332 587918
rect 388 587862 456 587918
rect 512 587862 608 587918
rect -12 587794 608 587862
rect -12 587738 84 587794
rect 140 587738 208 587794
rect 264 587738 332 587794
rect 388 587738 456 587794
rect 512 587738 608 587794
rect -12 587670 608 587738
rect -12 587614 84 587670
rect 140 587614 208 587670
rect 264 587614 332 587670
rect 388 587614 456 587670
rect 512 587614 608 587670
rect -12 587546 608 587614
rect -12 587490 84 587546
rect 140 587490 208 587546
rect 264 587490 332 587546
rect 388 587490 456 587546
rect 512 587490 608 587546
rect -12 569918 608 587490
rect -12 569862 84 569918
rect 140 569862 208 569918
rect 264 569862 332 569918
rect 388 569862 456 569918
rect 512 569862 608 569918
rect -12 569794 608 569862
rect -12 569738 84 569794
rect 140 569738 208 569794
rect 264 569738 332 569794
rect 388 569738 456 569794
rect 512 569738 608 569794
rect -12 569670 608 569738
rect -12 569614 84 569670
rect 140 569614 208 569670
rect 264 569614 332 569670
rect 388 569614 456 569670
rect 512 569614 608 569670
rect -12 569546 608 569614
rect -12 569490 84 569546
rect 140 569490 208 569546
rect 264 569490 332 569546
rect 388 569490 456 569546
rect 512 569490 608 569546
rect -12 551918 608 569490
rect -12 551862 84 551918
rect 140 551862 208 551918
rect 264 551862 332 551918
rect 388 551862 456 551918
rect 512 551862 608 551918
rect -12 551794 608 551862
rect -12 551738 84 551794
rect 140 551738 208 551794
rect 264 551738 332 551794
rect 388 551738 456 551794
rect 512 551738 608 551794
rect -12 551670 608 551738
rect -12 551614 84 551670
rect 140 551614 208 551670
rect 264 551614 332 551670
rect 388 551614 456 551670
rect 512 551614 608 551670
rect -12 551546 608 551614
rect -12 551490 84 551546
rect 140 551490 208 551546
rect 264 551490 332 551546
rect 388 551490 456 551546
rect 512 551490 608 551546
rect -12 533918 608 551490
rect -12 533862 84 533918
rect 140 533862 208 533918
rect 264 533862 332 533918
rect 388 533862 456 533918
rect 512 533862 608 533918
rect -12 533794 608 533862
rect -12 533738 84 533794
rect 140 533738 208 533794
rect 264 533738 332 533794
rect 388 533738 456 533794
rect 512 533738 608 533794
rect -12 533670 608 533738
rect -12 533614 84 533670
rect 140 533614 208 533670
rect 264 533614 332 533670
rect 388 533614 456 533670
rect 512 533614 608 533670
rect -12 533546 608 533614
rect -12 533490 84 533546
rect 140 533490 208 533546
rect 264 533490 332 533546
rect 388 533490 456 533546
rect 512 533490 608 533546
rect -12 515918 608 533490
rect -12 515862 84 515918
rect 140 515862 208 515918
rect 264 515862 332 515918
rect 388 515862 456 515918
rect 512 515862 608 515918
rect -12 515794 608 515862
rect -12 515738 84 515794
rect 140 515738 208 515794
rect 264 515738 332 515794
rect 388 515738 456 515794
rect 512 515738 608 515794
rect -12 515670 608 515738
rect -12 515614 84 515670
rect 140 515614 208 515670
rect 264 515614 332 515670
rect 388 515614 456 515670
rect 512 515614 608 515670
rect -12 515546 608 515614
rect -12 515490 84 515546
rect 140 515490 208 515546
rect 264 515490 332 515546
rect 388 515490 456 515546
rect 512 515490 608 515546
rect -12 497918 608 515490
rect -12 497862 84 497918
rect 140 497862 208 497918
rect 264 497862 332 497918
rect 388 497862 456 497918
rect 512 497862 608 497918
rect -12 497794 608 497862
rect -12 497738 84 497794
rect 140 497738 208 497794
rect 264 497738 332 497794
rect 388 497738 456 497794
rect 512 497738 608 497794
rect -12 497670 608 497738
rect -12 497614 84 497670
rect 140 497614 208 497670
rect 264 497614 332 497670
rect 388 497614 456 497670
rect 512 497614 608 497670
rect -12 497546 608 497614
rect -12 497490 84 497546
rect 140 497490 208 497546
rect 264 497490 332 497546
rect 388 497490 456 497546
rect 512 497490 608 497546
rect -12 479918 608 497490
rect -12 479862 84 479918
rect 140 479862 208 479918
rect 264 479862 332 479918
rect 388 479862 456 479918
rect 512 479862 608 479918
rect -12 479794 608 479862
rect -12 479738 84 479794
rect 140 479738 208 479794
rect 264 479738 332 479794
rect 388 479738 456 479794
rect 512 479738 608 479794
rect -12 479670 608 479738
rect -12 479614 84 479670
rect 140 479614 208 479670
rect 264 479614 332 479670
rect 388 479614 456 479670
rect 512 479614 608 479670
rect -12 479546 608 479614
rect -12 479490 84 479546
rect 140 479490 208 479546
rect 264 479490 332 479546
rect 388 479490 456 479546
rect 512 479490 608 479546
rect -12 461918 608 479490
rect -12 461862 84 461918
rect 140 461862 208 461918
rect 264 461862 332 461918
rect 388 461862 456 461918
rect 512 461862 608 461918
rect -12 461794 608 461862
rect -12 461738 84 461794
rect 140 461738 208 461794
rect 264 461738 332 461794
rect 388 461738 456 461794
rect 512 461738 608 461794
rect -12 461670 608 461738
rect -12 461614 84 461670
rect 140 461614 208 461670
rect 264 461614 332 461670
rect 388 461614 456 461670
rect 512 461614 608 461670
rect -12 461546 608 461614
rect -12 461490 84 461546
rect 140 461490 208 461546
rect 264 461490 332 461546
rect 388 461490 456 461546
rect 512 461490 608 461546
rect -12 443918 608 461490
rect -12 443862 84 443918
rect 140 443862 208 443918
rect 264 443862 332 443918
rect 388 443862 456 443918
rect 512 443862 608 443918
rect -12 443794 608 443862
rect -12 443738 84 443794
rect 140 443738 208 443794
rect 264 443738 332 443794
rect 388 443738 456 443794
rect 512 443738 608 443794
rect -12 443670 608 443738
rect -12 443614 84 443670
rect 140 443614 208 443670
rect 264 443614 332 443670
rect 388 443614 456 443670
rect 512 443614 608 443670
rect -12 443546 608 443614
rect -12 443490 84 443546
rect 140 443490 208 443546
rect 264 443490 332 443546
rect 388 443490 456 443546
rect 512 443490 608 443546
rect -12 425918 608 443490
rect -12 425862 84 425918
rect 140 425862 208 425918
rect 264 425862 332 425918
rect 388 425862 456 425918
rect 512 425862 608 425918
rect -12 425794 608 425862
rect -12 425738 84 425794
rect 140 425738 208 425794
rect 264 425738 332 425794
rect 388 425738 456 425794
rect 512 425738 608 425794
rect -12 425670 608 425738
rect -12 425614 84 425670
rect 140 425614 208 425670
rect 264 425614 332 425670
rect 388 425614 456 425670
rect 512 425614 608 425670
rect -12 425546 608 425614
rect -12 425490 84 425546
rect 140 425490 208 425546
rect 264 425490 332 425546
rect 388 425490 456 425546
rect 512 425490 608 425546
rect -12 407918 608 425490
rect -12 407862 84 407918
rect 140 407862 208 407918
rect 264 407862 332 407918
rect 388 407862 456 407918
rect 512 407862 608 407918
rect -12 407794 608 407862
rect -12 407738 84 407794
rect 140 407738 208 407794
rect 264 407738 332 407794
rect 388 407738 456 407794
rect 512 407738 608 407794
rect -12 407670 608 407738
rect -12 407614 84 407670
rect 140 407614 208 407670
rect 264 407614 332 407670
rect 388 407614 456 407670
rect 512 407614 608 407670
rect -12 407546 608 407614
rect -12 407490 84 407546
rect 140 407490 208 407546
rect 264 407490 332 407546
rect 388 407490 456 407546
rect 512 407490 608 407546
rect -12 389918 608 407490
rect -12 389862 84 389918
rect 140 389862 208 389918
rect 264 389862 332 389918
rect 388 389862 456 389918
rect 512 389862 608 389918
rect -12 389794 608 389862
rect -12 389738 84 389794
rect 140 389738 208 389794
rect 264 389738 332 389794
rect 388 389738 456 389794
rect 512 389738 608 389794
rect -12 389670 608 389738
rect -12 389614 84 389670
rect 140 389614 208 389670
rect 264 389614 332 389670
rect 388 389614 456 389670
rect 512 389614 608 389670
rect -12 389546 608 389614
rect -12 389490 84 389546
rect 140 389490 208 389546
rect 264 389490 332 389546
rect 388 389490 456 389546
rect 512 389490 608 389546
rect -12 371918 608 389490
rect -12 371862 84 371918
rect 140 371862 208 371918
rect 264 371862 332 371918
rect 388 371862 456 371918
rect 512 371862 608 371918
rect -12 371794 608 371862
rect -12 371738 84 371794
rect 140 371738 208 371794
rect 264 371738 332 371794
rect 388 371738 456 371794
rect 512 371738 608 371794
rect -12 371670 608 371738
rect -12 371614 84 371670
rect 140 371614 208 371670
rect 264 371614 332 371670
rect 388 371614 456 371670
rect 512 371614 608 371670
rect -12 371546 608 371614
rect -12 371490 84 371546
rect 140 371490 208 371546
rect 264 371490 332 371546
rect 388 371490 456 371546
rect 512 371490 608 371546
rect -12 353918 608 371490
rect -12 353862 84 353918
rect 140 353862 208 353918
rect 264 353862 332 353918
rect 388 353862 456 353918
rect 512 353862 608 353918
rect -12 353794 608 353862
rect -12 353738 84 353794
rect 140 353738 208 353794
rect 264 353738 332 353794
rect 388 353738 456 353794
rect 512 353738 608 353794
rect -12 353670 608 353738
rect -12 353614 84 353670
rect 140 353614 208 353670
rect 264 353614 332 353670
rect 388 353614 456 353670
rect 512 353614 608 353670
rect -12 353546 608 353614
rect -12 353490 84 353546
rect 140 353490 208 353546
rect 264 353490 332 353546
rect 388 353490 456 353546
rect 512 353490 608 353546
rect -12 335918 608 353490
rect -12 335862 84 335918
rect 140 335862 208 335918
rect 264 335862 332 335918
rect 388 335862 456 335918
rect 512 335862 608 335918
rect -12 335794 608 335862
rect -12 335738 84 335794
rect 140 335738 208 335794
rect 264 335738 332 335794
rect 388 335738 456 335794
rect 512 335738 608 335794
rect -12 335670 608 335738
rect -12 335614 84 335670
rect 140 335614 208 335670
rect 264 335614 332 335670
rect 388 335614 456 335670
rect 512 335614 608 335670
rect -12 335546 608 335614
rect -12 335490 84 335546
rect 140 335490 208 335546
rect 264 335490 332 335546
rect 388 335490 456 335546
rect 512 335490 608 335546
rect -12 317918 608 335490
rect -12 317862 84 317918
rect 140 317862 208 317918
rect 264 317862 332 317918
rect 388 317862 456 317918
rect 512 317862 608 317918
rect -12 317794 608 317862
rect -12 317738 84 317794
rect 140 317738 208 317794
rect 264 317738 332 317794
rect 388 317738 456 317794
rect 512 317738 608 317794
rect -12 317670 608 317738
rect -12 317614 84 317670
rect 140 317614 208 317670
rect 264 317614 332 317670
rect 388 317614 456 317670
rect 512 317614 608 317670
rect -12 317546 608 317614
rect -12 317490 84 317546
rect 140 317490 208 317546
rect 264 317490 332 317546
rect 388 317490 456 317546
rect 512 317490 608 317546
rect -12 299918 608 317490
rect -12 299862 84 299918
rect 140 299862 208 299918
rect 264 299862 332 299918
rect 388 299862 456 299918
rect 512 299862 608 299918
rect -12 299794 608 299862
rect -12 299738 84 299794
rect 140 299738 208 299794
rect 264 299738 332 299794
rect 388 299738 456 299794
rect 512 299738 608 299794
rect -12 299670 608 299738
rect -12 299614 84 299670
rect 140 299614 208 299670
rect 264 299614 332 299670
rect 388 299614 456 299670
rect 512 299614 608 299670
rect -12 299546 608 299614
rect -12 299490 84 299546
rect 140 299490 208 299546
rect 264 299490 332 299546
rect 388 299490 456 299546
rect 512 299490 608 299546
rect -12 281918 608 299490
rect -12 281862 84 281918
rect 140 281862 208 281918
rect 264 281862 332 281918
rect 388 281862 456 281918
rect 512 281862 608 281918
rect -12 281794 608 281862
rect -12 281738 84 281794
rect 140 281738 208 281794
rect 264 281738 332 281794
rect 388 281738 456 281794
rect 512 281738 608 281794
rect -12 281670 608 281738
rect -12 281614 84 281670
rect 140 281614 208 281670
rect 264 281614 332 281670
rect 388 281614 456 281670
rect 512 281614 608 281670
rect -12 281546 608 281614
rect -12 281490 84 281546
rect 140 281490 208 281546
rect 264 281490 332 281546
rect 388 281490 456 281546
rect 512 281490 608 281546
rect -12 263918 608 281490
rect -12 263862 84 263918
rect 140 263862 208 263918
rect 264 263862 332 263918
rect 388 263862 456 263918
rect 512 263862 608 263918
rect -12 263794 608 263862
rect -12 263738 84 263794
rect 140 263738 208 263794
rect 264 263738 332 263794
rect 388 263738 456 263794
rect 512 263738 608 263794
rect -12 263670 608 263738
rect -12 263614 84 263670
rect 140 263614 208 263670
rect 264 263614 332 263670
rect 388 263614 456 263670
rect 512 263614 608 263670
rect -12 263546 608 263614
rect -12 263490 84 263546
rect 140 263490 208 263546
rect 264 263490 332 263546
rect 388 263490 456 263546
rect 512 263490 608 263546
rect -12 245918 608 263490
rect -12 245862 84 245918
rect 140 245862 208 245918
rect 264 245862 332 245918
rect 388 245862 456 245918
rect 512 245862 608 245918
rect -12 245794 608 245862
rect -12 245738 84 245794
rect 140 245738 208 245794
rect 264 245738 332 245794
rect 388 245738 456 245794
rect 512 245738 608 245794
rect -12 245670 608 245738
rect -12 245614 84 245670
rect 140 245614 208 245670
rect 264 245614 332 245670
rect 388 245614 456 245670
rect 512 245614 608 245670
rect -12 245546 608 245614
rect -12 245490 84 245546
rect 140 245490 208 245546
rect 264 245490 332 245546
rect 388 245490 456 245546
rect 512 245490 608 245546
rect -12 227918 608 245490
rect -12 227862 84 227918
rect 140 227862 208 227918
rect 264 227862 332 227918
rect 388 227862 456 227918
rect 512 227862 608 227918
rect -12 227794 608 227862
rect -12 227738 84 227794
rect 140 227738 208 227794
rect 264 227738 332 227794
rect 388 227738 456 227794
rect 512 227738 608 227794
rect -12 227670 608 227738
rect -12 227614 84 227670
rect 140 227614 208 227670
rect 264 227614 332 227670
rect 388 227614 456 227670
rect 512 227614 608 227670
rect -12 227546 608 227614
rect -12 227490 84 227546
rect 140 227490 208 227546
rect 264 227490 332 227546
rect 388 227490 456 227546
rect 512 227490 608 227546
rect -12 209918 608 227490
rect -12 209862 84 209918
rect 140 209862 208 209918
rect 264 209862 332 209918
rect 388 209862 456 209918
rect 512 209862 608 209918
rect -12 209794 608 209862
rect -12 209738 84 209794
rect 140 209738 208 209794
rect 264 209738 332 209794
rect 388 209738 456 209794
rect 512 209738 608 209794
rect -12 209670 608 209738
rect -12 209614 84 209670
rect 140 209614 208 209670
rect 264 209614 332 209670
rect 388 209614 456 209670
rect 512 209614 608 209670
rect -12 209546 608 209614
rect -12 209490 84 209546
rect 140 209490 208 209546
rect 264 209490 332 209546
rect 388 209490 456 209546
rect 512 209490 608 209546
rect -12 191918 608 209490
rect -12 191862 84 191918
rect 140 191862 208 191918
rect 264 191862 332 191918
rect 388 191862 456 191918
rect 512 191862 608 191918
rect -12 191794 608 191862
rect -12 191738 84 191794
rect 140 191738 208 191794
rect 264 191738 332 191794
rect 388 191738 456 191794
rect 512 191738 608 191794
rect -12 191670 608 191738
rect -12 191614 84 191670
rect 140 191614 208 191670
rect 264 191614 332 191670
rect 388 191614 456 191670
rect 512 191614 608 191670
rect -12 191546 608 191614
rect -12 191490 84 191546
rect 140 191490 208 191546
rect 264 191490 332 191546
rect 388 191490 456 191546
rect 512 191490 608 191546
rect -12 173918 608 191490
rect -12 173862 84 173918
rect 140 173862 208 173918
rect 264 173862 332 173918
rect 388 173862 456 173918
rect 512 173862 608 173918
rect -12 173794 608 173862
rect -12 173738 84 173794
rect 140 173738 208 173794
rect 264 173738 332 173794
rect 388 173738 456 173794
rect 512 173738 608 173794
rect -12 173670 608 173738
rect -12 173614 84 173670
rect 140 173614 208 173670
rect 264 173614 332 173670
rect 388 173614 456 173670
rect 512 173614 608 173670
rect -12 173546 608 173614
rect -12 173490 84 173546
rect 140 173490 208 173546
rect 264 173490 332 173546
rect 388 173490 456 173546
rect 512 173490 608 173546
rect -12 155918 608 173490
rect -12 155862 84 155918
rect 140 155862 208 155918
rect 264 155862 332 155918
rect 388 155862 456 155918
rect 512 155862 608 155918
rect -12 155794 608 155862
rect -12 155738 84 155794
rect 140 155738 208 155794
rect 264 155738 332 155794
rect 388 155738 456 155794
rect 512 155738 608 155794
rect -12 155670 608 155738
rect -12 155614 84 155670
rect 140 155614 208 155670
rect 264 155614 332 155670
rect 388 155614 456 155670
rect 512 155614 608 155670
rect -12 155546 608 155614
rect -12 155490 84 155546
rect 140 155490 208 155546
rect 264 155490 332 155546
rect 388 155490 456 155546
rect 512 155490 608 155546
rect -12 137918 608 155490
rect -12 137862 84 137918
rect 140 137862 208 137918
rect 264 137862 332 137918
rect 388 137862 456 137918
rect 512 137862 608 137918
rect -12 137794 608 137862
rect -12 137738 84 137794
rect 140 137738 208 137794
rect 264 137738 332 137794
rect 388 137738 456 137794
rect 512 137738 608 137794
rect -12 137670 608 137738
rect -12 137614 84 137670
rect 140 137614 208 137670
rect 264 137614 332 137670
rect 388 137614 456 137670
rect 512 137614 608 137670
rect -12 137546 608 137614
rect -12 137490 84 137546
rect 140 137490 208 137546
rect 264 137490 332 137546
rect 388 137490 456 137546
rect 512 137490 608 137546
rect -12 119918 608 137490
rect -12 119862 84 119918
rect 140 119862 208 119918
rect 264 119862 332 119918
rect 388 119862 456 119918
rect 512 119862 608 119918
rect -12 119794 608 119862
rect -12 119738 84 119794
rect 140 119738 208 119794
rect 264 119738 332 119794
rect 388 119738 456 119794
rect 512 119738 608 119794
rect -12 119670 608 119738
rect -12 119614 84 119670
rect 140 119614 208 119670
rect 264 119614 332 119670
rect 388 119614 456 119670
rect 512 119614 608 119670
rect -12 119546 608 119614
rect -12 119490 84 119546
rect 140 119490 208 119546
rect 264 119490 332 119546
rect 388 119490 456 119546
rect 512 119490 608 119546
rect -12 101918 608 119490
rect -12 101862 84 101918
rect 140 101862 208 101918
rect 264 101862 332 101918
rect 388 101862 456 101918
rect 512 101862 608 101918
rect -12 101794 608 101862
rect -12 101738 84 101794
rect 140 101738 208 101794
rect 264 101738 332 101794
rect 388 101738 456 101794
rect 512 101738 608 101794
rect -12 101670 608 101738
rect -12 101614 84 101670
rect 140 101614 208 101670
rect 264 101614 332 101670
rect 388 101614 456 101670
rect 512 101614 608 101670
rect -12 101546 608 101614
rect -12 101490 84 101546
rect 140 101490 208 101546
rect 264 101490 332 101546
rect 388 101490 456 101546
rect 512 101490 608 101546
rect -12 83918 608 101490
rect -12 83862 84 83918
rect 140 83862 208 83918
rect 264 83862 332 83918
rect 388 83862 456 83918
rect 512 83862 608 83918
rect -12 83794 608 83862
rect -12 83738 84 83794
rect 140 83738 208 83794
rect 264 83738 332 83794
rect 388 83738 456 83794
rect 512 83738 608 83794
rect -12 83670 608 83738
rect -12 83614 84 83670
rect 140 83614 208 83670
rect 264 83614 332 83670
rect 388 83614 456 83670
rect 512 83614 608 83670
rect -12 83546 608 83614
rect -12 83490 84 83546
rect 140 83490 208 83546
rect 264 83490 332 83546
rect 388 83490 456 83546
rect 512 83490 608 83546
rect -12 65918 608 83490
rect -12 65862 84 65918
rect 140 65862 208 65918
rect 264 65862 332 65918
rect 388 65862 456 65918
rect 512 65862 608 65918
rect -12 65794 608 65862
rect -12 65738 84 65794
rect 140 65738 208 65794
rect 264 65738 332 65794
rect 388 65738 456 65794
rect 512 65738 608 65794
rect -12 65670 608 65738
rect -12 65614 84 65670
rect 140 65614 208 65670
rect 264 65614 332 65670
rect 388 65614 456 65670
rect 512 65614 608 65670
rect -12 65546 608 65614
rect -12 65490 84 65546
rect 140 65490 208 65546
rect 264 65490 332 65546
rect 388 65490 456 65546
rect 512 65490 608 65546
rect -12 47918 608 65490
rect -12 47862 84 47918
rect 140 47862 208 47918
rect 264 47862 332 47918
rect 388 47862 456 47918
rect 512 47862 608 47918
rect -12 47794 608 47862
rect -12 47738 84 47794
rect 140 47738 208 47794
rect 264 47738 332 47794
rect 388 47738 456 47794
rect 512 47738 608 47794
rect -12 47670 608 47738
rect -12 47614 84 47670
rect 140 47614 208 47670
rect 264 47614 332 47670
rect 388 47614 456 47670
rect 512 47614 608 47670
rect -12 47546 608 47614
rect -12 47490 84 47546
rect 140 47490 208 47546
rect 264 47490 332 47546
rect 388 47490 456 47546
rect 512 47490 608 47546
rect -12 29918 608 47490
rect -12 29862 84 29918
rect 140 29862 208 29918
rect 264 29862 332 29918
rect 388 29862 456 29918
rect 512 29862 608 29918
rect -12 29794 608 29862
rect -12 29738 84 29794
rect 140 29738 208 29794
rect 264 29738 332 29794
rect 388 29738 456 29794
rect 512 29738 608 29794
rect -12 29670 608 29738
rect -12 29614 84 29670
rect 140 29614 208 29670
rect 264 29614 332 29670
rect 388 29614 456 29670
rect 512 29614 608 29670
rect -12 29546 608 29614
rect -12 29490 84 29546
rect 140 29490 208 29546
rect 264 29490 332 29546
rect 388 29490 456 29546
rect 512 29490 608 29546
rect -12 11918 608 29490
rect -12 11862 84 11918
rect 140 11862 208 11918
rect 264 11862 332 11918
rect 388 11862 456 11918
rect 512 11862 608 11918
rect -12 11794 608 11862
rect -12 11738 84 11794
rect 140 11738 208 11794
rect 264 11738 332 11794
rect 388 11738 456 11794
rect 512 11738 608 11794
rect -12 11670 608 11738
rect -12 11614 84 11670
rect 140 11614 208 11670
rect 264 11614 332 11670
rect 388 11614 456 11670
rect 512 11614 608 11670
rect -12 11546 608 11614
rect -12 11490 84 11546
rect 140 11490 208 11546
rect 264 11490 332 11546
rect 388 11490 456 11546
rect 512 11490 608 11546
rect -12 848 608 11490
rect 948 598380 1568 598476
rect 948 598324 1044 598380
rect 1100 598324 1168 598380
rect 1224 598324 1292 598380
rect 1348 598324 1416 598380
rect 1472 598324 1568 598380
rect 948 598256 1568 598324
rect 948 598200 1044 598256
rect 1100 598200 1168 598256
rect 1224 598200 1292 598256
rect 1348 598200 1416 598256
rect 1472 598200 1568 598256
rect 948 598132 1568 598200
rect 948 598076 1044 598132
rect 1100 598076 1168 598132
rect 1224 598076 1292 598132
rect 1348 598076 1416 598132
rect 1472 598076 1568 598132
rect 948 598008 1568 598076
rect 948 597952 1044 598008
rect 1100 597952 1168 598008
rect 1224 597952 1292 598008
rect 1348 597952 1416 598008
rect 1472 597952 1568 598008
rect 948 581918 1568 597952
rect 948 581862 1044 581918
rect 1100 581862 1168 581918
rect 1224 581862 1292 581918
rect 1348 581862 1416 581918
rect 1472 581862 1568 581918
rect 948 581794 1568 581862
rect 948 581738 1044 581794
rect 1100 581738 1168 581794
rect 1224 581738 1292 581794
rect 1348 581738 1416 581794
rect 1472 581738 1568 581794
rect 948 581670 1568 581738
rect 948 581614 1044 581670
rect 1100 581614 1168 581670
rect 1224 581614 1292 581670
rect 1348 581614 1416 581670
rect 1472 581614 1568 581670
rect 948 581546 1568 581614
rect 948 581490 1044 581546
rect 1100 581490 1168 581546
rect 1224 581490 1292 581546
rect 1348 581490 1416 581546
rect 1472 581490 1568 581546
rect 948 563918 1568 581490
rect 948 563862 1044 563918
rect 1100 563862 1168 563918
rect 1224 563862 1292 563918
rect 1348 563862 1416 563918
rect 1472 563862 1568 563918
rect 948 563794 1568 563862
rect 948 563738 1044 563794
rect 1100 563738 1168 563794
rect 1224 563738 1292 563794
rect 1348 563738 1416 563794
rect 1472 563738 1568 563794
rect 948 563670 1568 563738
rect 948 563614 1044 563670
rect 1100 563614 1168 563670
rect 1224 563614 1292 563670
rect 1348 563614 1416 563670
rect 1472 563614 1568 563670
rect 948 563546 1568 563614
rect 948 563490 1044 563546
rect 1100 563490 1168 563546
rect 1224 563490 1292 563546
rect 1348 563490 1416 563546
rect 1472 563490 1568 563546
rect 948 545918 1568 563490
rect 948 545862 1044 545918
rect 1100 545862 1168 545918
rect 1224 545862 1292 545918
rect 1348 545862 1416 545918
rect 1472 545862 1568 545918
rect 948 545794 1568 545862
rect 948 545738 1044 545794
rect 1100 545738 1168 545794
rect 1224 545738 1292 545794
rect 1348 545738 1416 545794
rect 1472 545738 1568 545794
rect 948 545670 1568 545738
rect 948 545614 1044 545670
rect 1100 545614 1168 545670
rect 1224 545614 1292 545670
rect 1348 545614 1416 545670
rect 1472 545614 1568 545670
rect 948 545546 1568 545614
rect 948 545490 1044 545546
rect 1100 545490 1168 545546
rect 1224 545490 1292 545546
rect 1348 545490 1416 545546
rect 1472 545490 1568 545546
rect 948 527918 1568 545490
rect 948 527862 1044 527918
rect 1100 527862 1168 527918
rect 1224 527862 1292 527918
rect 1348 527862 1416 527918
rect 1472 527862 1568 527918
rect 948 527794 1568 527862
rect 948 527738 1044 527794
rect 1100 527738 1168 527794
rect 1224 527738 1292 527794
rect 1348 527738 1416 527794
rect 1472 527738 1568 527794
rect 948 527670 1568 527738
rect 948 527614 1044 527670
rect 1100 527614 1168 527670
rect 1224 527614 1292 527670
rect 1348 527614 1416 527670
rect 1472 527614 1568 527670
rect 948 527546 1568 527614
rect 948 527490 1044 527546
rect 1100 527490 1168 527546
rect 1224 527490 1292 527546
rect 1348 527490 1416 527546
rect 1472 527490 1568 527546
rect 948 509918 1568 527490
rect 948 509862 1044 509918
rect 1100 509862 1168 509918
rect 1224 509862 1292 509918
rect 1348 509862 1416 509918
rect 1472 509862 1568 509918
rect 948 509794 1568 509862
rect 948 509738 1044 509794
rect 1100 509738 1168 509794
rect 1224 509738 1292 509794
rect 1348 509738 1416 509794
rect 1472 509738 1568 509794
rect 948 509670 1568 509738
rect 948 509614 1044 509670
rect 1100 509614 1168 509670
rect 1224 509614 1292 509670
rect 1348 509614 1416 509670
rect 1472 509614 1568 509670
rect 948 509546 1568 509614
rect 948 509490 1044 509546
rect 1100 509490 1168 509546
rect 1224 509490 1292 509546
rect 1348 509490 1416 509546
rect 1472 509490 1568 509546
rect 948 491918 1568 509490
rect 948 491862 1044 491918
rect 1100 491862 1168 491918
rect 1224 491862 1292 491918
rect 1348 491862 1416 491918
rect 1472 491862 1568 491918
rect 948 491794 1568 491862
rect 948 491738 1044 491794
rect 1100 491738 1168 491794
rect 1224 491738 1292 491794
rect 1348 491738 1416 491794
rect 1472 491738 1568 491794
rect 948 491670 1568 491738
rect 948 491614 1044 491670
rect 1100 491614 1168 491670
rect 1224 491614 1292 491670
rect 1348 491614 1416 491670
rect 1472 491614 1568 491670
rect 948 491546 1568 491614
rect 948 491490 1044 491546
rect 1100 491490 1168 491546
rect 1224 491490 1292 491546
rect 1348 491490 1416 491546
rect 1472 491490 1568 491546
rect 948 473918 1568 491490
rect 948 473862 1044 473918
rect 1100 473862 1168 473918
rect 1224 473862 1292 473918
rect 1348 473862 1416 473918
rect 1472 473862 1568 473918
rect 948 473794 1568 473862
rect 948 473738 1044 473794
rect 1100 473738 1168 473794
rect 1224 473738 1292 473794
rect 1348 473738 1416 473794
rect 1472 473738 1568 473794
rect 948 473670 1568 473738
rect 948 473614 1044 473670
rect 1100 473614 1168 473670
rect 1224 473614 1292 473670
rect 1348 473614 1416 473670
rect 1472 473614 1568 473670
rect 948 473546 1568 473614
rect 948 473490 1044 473546
rect 1100 473490 1168 473546
rect 1224 473490 1292 473546
rect 1348 473490 1416 473546
rect 1472 473490 1568 473546
rect 948 455918 1568 473490
rect 948 455862 1044 455918
rect 1100 455862 1168 455918
rect 1224 455862 1292 455918
rect 1348 455862 1416 455918
rect 1472 455862 1568 455918
rect 948 455794 1568 455862
rect 948 455738 1044 455794
rect 1100 455738 1168 455794
rect 1224 455738 1292 455794
rect 1348 455738 1416 455794
rect 1472 455738 1568 455794
rect 948 455670 1568 455738
rect 948 455614 1044 455670
rect 1100 455614 1168 455670
rect 1224 455614 1292 455670
rect 1348 455614 1416 455670
rect 1472 455614 1568 455670
rect 948 455546 1568 455614
rect 948 455490 1044 455546
rect 1100 455490 1168 455546
rect 1224 455490 1292 455546
rect 1348 455490 1416 455546
rect 1472 455490 1568 455546
rect 948 437918 1568 455490
rect 948 437862 1044 437918
rect 1100 437862 1168 437918
rect 1224 437862 1292 437918
rect 1348 437862 1416 437918
rect 1472 437862 1568 437918
rect 948 437794 1568 437862
rect 948 437738 1044 437794
rect 1100 437738 1168 437794
rect 1224 437738 1292 437794
rect 1348 437738 1416 437794
rect 1472 437738 1568 437794
rect 948 437670 1568 437738
rect 948 437614 1044 437670
rect 1100 437614 1168 437670
rect 1224 437614 1292 437670
rect 1348 437614 1416 437670
rect 1472 437614 1568 437670
rect 948 437546 1568 437614
rect 948 437490 1044 437546
rect 1100 437490 1168 437546
rect 1224 437490 1292 437546
rect 1348 437490 1416 437546
rect 1472 437490 1568 437546
rect 948 419918 1568 437490
rect 948 419862 1044 419918
rect 1100 419862 1168 419918
rect 1224 419862 1292 419918
rect 1348 419862 1416 419918
rect 1472 419862 1568 419918
rect 948 419794 1568 419862
rect 948 419738 1044 419794
rect 1100 419738 1168 419794
rect 1224 419738 1292 419794
rect 1348 419738 1416 419794
rect 1472 419738 1568 419794
rect 948 419670 1568 419738
rect 948 419614 1044 419670
rect 1100 419614 1168 419670
rect 1224 419614 1292 419670
rect 1348 419614 1416 419670
rect 1472 419614 1568 419670
rect 948 419546 1568 419614
rect 948 419490 1044 419546
rect 1100 419490 1168 419546
rect 1224 419490 1292 419546
rect 1348 419490 1416 419546
rect 1472 419490 1568 419546
rect 948 401918 1568 419490
rect 948 401862 1044 401918
rect 1100 401862 1168 401918
rect 1224 401862 1292 401918
rect 1348 401862 1416 401918
rect 1472 401862 1568 401918
rect 948 401794 1568 401862
rect 948 401738 1044 401794
rect 1100 401738 1168 401794
rect 1224 401738 1292 401794
rect 1348 401738 1416 401794
rect 1472 401738 1568 401794
rect 948 401670 1568 401738
rect 948 401614 1044 401670
rect 1100 401614 1168 401670
rect 1224 401614 1292 401670
rect 1348 401614 1416 401670
rect 1472 401614 1568 401670
rect 948 401546 1568 401614
rect 948 401490 1044 401546
rect 1100 401490 1168 401546
rect 1224 401490 1292 401546
rect 1348 401490 1416 401546
rect 1472 401490 1568 401546
rect 948 383918 1568 401490
rect 948 383862 1044 383918
rect 1100 383862 1168 383918
rect 1224 383862 1292 383918
rect 1348 383862 1416 383918
rect 1472 383862 1568 383918
rect 948 383794 1568 383862
rect 948 383738 1044 383794
rect 1100 383738 1168 383794
rect 1224 383738 1292 383794
rect 1348 383738 1416 383794
rect 1472 383738 1568 383794
rect 948 383670 1568 383738
rect 948 383614 1044 383670
rect 1100 383614 1168 383670
rect 1224 383614 1292 383670
rect 1348 383614 1416 383670
rect 1472 383614 1568 383670
rect 948 383546 1568 383614
rect 948 383490 1044 383546
rect 1100 383490 1168 383546
rect 1224 383490 1292 383546
rect 1348 383490 1416 383546
rect 1472 383490 1568 383546
rect 948 365918 1568 383490
rect 948 365862 1044 365918
rect 1100 365862 1168 365918
rect 1224 365862 1292 365918
rect 1348 365862 1416 365918
rect 1472 365862 1568 365918
rect 948 365794 1568 365862
rect 948 365738 1044 365794
rect 1100 365738 1168 365794
rect 1224 365738 1292 365794
rect 1348 365738 1416 365794
rect 1472 365738 1568 365794
rect 948 365670 1568 365738
rect 948 365614 1044 365670
rect 1100 365614 1168 365670
rect 1224 365614 1292 365670
rect 1348 365614 1416 365670
rect 1472 365614 1568 365670
rect 948 365546 1568 365614
rect 948 365490 1044 365546
rect 1100 365490 1168 365546
rect 1224 365490 1292 365546
rect 1348 365490 1416 365546
rect 1472 365490 1568 365546
rect 948 347918 1568 365490
rect 948 347862 1044 347918
rect 1100 347862 1168 347918
rect 1224 347862 1292 347918
rect 1348 347862 1416 347918
rect 1472 347862 1568 347918
rect 948 347794 1568 347862
rect 948 347738 1044 347794
rect 1100 347738 1168 347794
rect 1224 347738 1292 347794
rect 1348 347738 1416 347794
rect 1472 347738 1568 347794
rect 948 347670 1568 347738
rect 948 347614 1044 347670
rect 1100 347614 1168 347670
rect 1224 347614 1292 347670
rect 1348 347614 1416 347670
rect 1472 347614 1568 347670
rect 948 347546 1568 347614
rect 948 347490 1044 347546
rect 1100 347490 1168 347546
rect 1224 347490 1292 347546
rect 1348 347490 1416 347546
rect 1472 347490 1568 347546
rect 948 329918 1568 347490
rect 948 329862 1044 329918
rect 1100 329862 1168 329918
rect 1224 329862 1292 329918
rect 1348 329862 1416 329918
rect 1472 329862 1568 329918
rect 948 329794 1568 329862
rect 948 329738 1044 329794
rect 1100 329738 1168 329794
rect 1224 329738 1292 329794
rect 1348 329738 1416 329794
rect 1472 329738 1568 329794
rect 948 329670 1568 329738
rect 948 329614 1044 329670
rect 1100 329614 1168 329670
rect 1224 329614 1292 329670
rect 1348 329614 1416 329670
rect 1472 329614 1568 329670
rect 948 329546 1568 329614
rect 948 329490 1044 329546
rect 1100 329490 1168 329546
rect 1224 329490 1292 329546
rect 1348 329490 1416 329546
rect 1472 329490 1568 329546
rect 948 311918 1568 329490
rect 948 311862 1044 311918
rect 1100 311862 1168 311918
rect 1224 311862 1292 311918
rect 1348 311862 1416 311918
rect 1472 311862 1568 311918
rect 948 311794 1568 311862
rect 948 311738 1044 311794
rect 1100 311738 1168 311794
rect 1224 311738 1292 311794
rect 1348 311738 1416 311794
rect 1472 311738 1568 311794
rect 948 311670 1568 311738
rect 948 311614 1044 311670
rect 1100 311614 1168 311670
rect 1224 311614 1292 311670
rect 1348 311614 1416 311670
rect 1472 311614 1568 311670
rect 948 311546 1568 311614
rect 948 311490 1044 311546
rect 1100 311490 1168 311546
rect 1224 311490 1292 311546
rect 1348 311490 1416 311546
rect 1472 311490 1568 311546
rect 948 293918 1568 311490
rect 948 293862 1044 293918
rect 1100 293862 1168 293918
rect 1224 293862 1292 293918
rect 1348 293862 1416 293918
rect 1472 293862 1568 293918
rect 948 293794 1568 293862
rect 948 293738 1044 293794
rect 1100 293738 1168 293794
rect 1224 293738 1292 293794
rect 1348 293738 1416 293794
rect 1472 293738 1568 293794
rect 948 293670 1568 293738
rect 948 293614 1044 293670
rect 1100 293614 1168 293670
rect 1224 293614 1292 293670
rect 1348 293614 1416 293670
rect 1472 293614 1568 293670
rect 948 293546 1568 293614
rect 948 293490 1044 293546
rect 1100 293490 1168 293546
rect 1224 293490 1292 293546
rect 1348 293490 1416 293546
rect 1472 293490 1568 293546
rect 948 275918 1568 293490
rect 948 275862 1044 275918
rect 1100 275862 1168 275918
rect 1224 275862 1292 275918
rect 1348 275862 1416 275918
rect 1472 275862 1568 275918
rect 948 275794 1568 275862
rect 948 275738 1044 275794
rect 1100 275738 1168 275794
rect 1224 275738 1292 275794
rect 1348 275738 1416 275794
rect 1472 275738 1568 275794
rect 948 275670 1568 275738
rect 948 275614 1044 275670
rect 1100 275614 1168 275670
rect 1224 275614 1292 275670
rect 1348 275614 1416 275670
rect 1472 275614 1568 275670
rect 948 275546 1568 275614
rect 948 275490 1044 275546
rect 1100 275490 1168 275546
rect 1224 275490 1292 275546
rect 1348 275490 1416 275546
rect 1472 275490 1568 275546
rect 948 257918 1568 275490
rect 948 257862 1044 257918
rect 1100 257862 1168 257918
rect 1224 257862 1292 257918
rect 1348 257862 1416 257918
rect 1472 257862 1568 257918
rect 948 257794 1568 257862
rect 948 257738 1044 257794
rect 1100 257738 1168 257794
rect 1224 257738 1292 257794
rect 1348 257738 1416 257794
rect 1472 257738 1568 257794
rect 948 257670 1568 257738
rect 948 257614 1044 257670
rect 1100 257614 1168 257670
rect 1224 257614 1292 257670
rect 1348 257614 1416 257670
rect 1472 257614 1568 257670
rect 948 257546 1568 257614
rect 948 257490 1044 257546
rect 1100 257490 1168 257546
rect 1224 257490 1292 257546
rect 1348 257490 1416 257546
rect 1472 257490 1568 257546
rect 948 239918 1568 257490
rect 948 239862 1044 239918
rect 1100 239862 1168 239918
rect 1224 239862 1292 239918
rect 1348 239862 1416 239918
rect 1472 239862 1568 239918
rect 948 239794 1568 239862
rect 948 239738 1044 239794
rect 1100 239738 1168 239794
rect 1224 239738 1292 239794
rect 1348 239738 1416 239794
rect 1472 239738 1568 239794
rect 948 239670 1568 239738
rect 948 239614 1044 239670
rect 1100 239614 1168 239670
rect 1224 239614 1292 239670
rect 1348 239614 1416 239670
rect 1472 239614 1568 239670
rect 948 239546 1568 239614
rect 948 239490 1044 239546
rect 1100 239490 1168 239546
rect 1224 239490 1292 239546
rect 1348 239490 1416 239546
rect 1472 239490 1568 239546
rect 948 221918 1568 239490
rect 948 221862 1044 221918
rect 1100 221862 1168 221918
rect 1224 221862 1292 221918
rect 1348 221862 1416 221918
rect 1472 221862 1568 221918
rect 948 221794 1568 221862
rect 948 221738 1044 221794
rect 1100 221738 1168 221794
rect 1224 221738 1292 221794
rect 1348 221738 1416 221794
rect 1472 221738 1568 221794
rect 948 221670 1568 221738
rect 948 221614 1044 221670
rect 1100 221614 1168 221670
rect 1224 221614 1292 221670
rect 1348 221614 1416 221670
rect 1472 221614 1568 221670
rect 948 221546 1568 221614
rect 948 221490 1044 221546
rect 1100 221490 1168 221546
rect 1224 221490 1292 221546
rect 1348 221490 1416 221546
rect 1472 221490 1568 221546
rect 948 203918 1568 221490
rect 948 203862 1044 203918
rect 1100 203862 1168 203918
rect 1224 203862 1292 203918
rect 1348 203862 1416 203918
rect 1472 203862 1568 203918
rect 948 203794 1568 203862
rect 948 203738 1044 203794
rect 1100 203738 1168 203794
rect 1224 203738 1292 203794
rect 1348 203738 1416 203794
rect 1472 203738 1568 203794
rect 948 203670 1568 203738
rect 948 203614 1044 203670
rect 1100 203614 1168 203670
rect 1224 203614 1292 203670
rect 1348 203614 1416 203670
rect 1472 203614 1568 203670
rect 948 203546 1568 203614
rect 948 203490 1044 203546
rect 1100 203490 1168 203546
rect 1224 203490 1292 203546
rect 1348 203490 1416 203546
rect 1472 203490 1568 203546
rect 948 185918 1568 203490
rect 948 185862 1044 185918
rect 1100 185862 1168 185918
rect 1224 185862 1292 185918
rect 1348 185862 1416 185918
rect 1472 185862 1568 185918
rect 948 185794 1568 185862
rect 948 185738 1044 185794
rect 1100 185738 1168 185794
rect 1224 185738 1292 185794
rect 1348 185738 1416 185794
rect 1472 185738 1568 185794
rect 948 185670 1568 185738
rect 948 185614 1044 185670
rect 1100 185614 1168 185670
rect 1224 185614 1292 185670
rect 1348 185614 1416 185670
rect 1472 185614 1568 185670
rect 948 185546 1568 185614
rect 948 185490 1044 185546
rect 1100 185490 1168 185546
rect 1224 185490 1292 185546
rect 1348 185490 1416 185546
rect 1472 185490 1568 185546
rect 948 167918 1568 185490
rect 948 167862 1044 167918
rect 1100 167862 1168 167918
rect 1224 167862 1292 167918
rect 1348 167862 1416 167918
rect 1472 167862 1568 167918
rect 948 167794 1568 167862
rect 948 167738 1044 167794
rect 1100 167738 1168 167794
rect 1224 167738 1292 167794
rect 1348 167738 1416 167794
rect 1472 167738 1568 167794
rect 948 167670 1568 167738
rect 948 167614 1044 167670
rect 1100 167614 1168 167670
rect 1224 167614 1292 167670
rect 1348 167614 1416 167670
rect 1472 167614 1568 167670
rect 948 167546 1568 167614
rect 948 167490 1044 167546
rect 1100 167490 1168 167546
rect 1224 167490 1292 167546
rect 1348 167490 1416 167546
rect 1472 167490 1568 167546
rect 948 149918 1568 167490
rect 948 149862 1044 149918
rect 1100 149862 1168 149918
rect 1224 149862 1292 149918
rect 1348 149862 1416 149918
rect 1472 149862 1568 149918
rect 948 149794 1568 149862
rect 948 149738 1044 149794
rect 1100 149738 1168 149794
rect 1224 149738 1292 149794
rect 1348 149738 1416 149794
rect 1472 149738 1568 149794
rect 948 149670 1568 149738
rect 948 149614 1044 149670
rect 1100 149614 1168 149670
rect 1224 149614 1292 149670
rect 1348 149614 1416 149670
rect 1472 149614 1568 149670
rect 948 149546 1568 149614
rect 948 149490 1044 149546
rect 1100 149490 1168 149546
rect 1224 149490 1292 149546
rect 1348 149490 1416 149546
rect 1472 149490 1568 149546
rect 948 131918 1568 149490
rect 948 131862 1044 131918
rect 1100 131862 1168 131918
rect 1224 131862 1292 131918
rect 1348 131862 1416 131918
rect 1472 131862 1568 131918
rect 948 131794 1568 131862
rect 948 131738 1044 131794
rect 1100 131738 1168 131794
rect 1224 131738 1292 131794
rect 1348 131738 1416 131794
rect 1472 131738 1568 131794
rect 948 131670 1568 131738
rect 948 131614 1044 131670
rect 1100 131614 1168 131670
rect 1224 131614 1292 131670
rect 1348 131614 1416 131670
rect 1472 131614 1568 131670
rect 948 131546 1568 131614
rect 948 131490 1044 131546
rect 1100 131490 1168 131546
rect 1224 131490 1292 131546
rect 1348 131490 1416 131546
rect 1472 131490 1568 131546
rect 948 113918 1568 131490
rect 948 113862 1044 113918
rect 1100 113862 1168 113918
rect 1224 113862 1292 113918
rect 1348 113862 1416 113918
rect 1472 113862 1568 113918
rect 948 113794 1568 113862
rect 948 113738 1044 113794
rect 1100 113738 1168 113794
rect 1224 113738 1292 113794
rect 1348 113738 1416 113794
rect 1472 113738 1568 113794
rect 948 113670 1568 113738
rect 948 113614 1044 113670
rect 1100 113614 1168 113670
rect 1224 113614 1292 113670
rect 1348 113614 1416 113670
rect 1472 113614 1568 113670
rect 948 113546 1568 113614
rect 948 113490 1044 113546
rect 1100 113490 1168 113546
rect 1224 113490 1292 113546
rect 1348 113490 1416 113546
rect 1472 113490 1568 113546
rect 948 95918 1568 113490
rect 948 95862 1044 95918
rect 1100 95862 1168 95918
rect 1224 95862 1292 95918
rect 1348 95862 1416 95918
rect 1472 95862 1568 95918
rect 948 95794 1568 95862
rect 948 95738 1044 95794
rect 1100 95738 1168 95794
rect 1224 95738 1292 95794
rect 1348 95738 1416 95794
rect 1472 95738 1568 95794
rect 948 95670 1568 95738
rect 948 95614 1044 95670
rect 1100 95614 1168 95670
rect 1224 95614 1292 95670
rect 1348 95614 1416 95670
rect 1472 95614 1568 95670
rect 948 95546 1568 95614
rect 948 95490 1044 95546
rect 1100 95490 1168 95546
rect 1224 95490 1292 95546
rect 1348 95490 1416 95546
rect 1472 95490 1568 95546
rect 948 77918 1568 95490
rect 948 77862 1044 77918
rect 1100 77862 1168 77918
rect 1224 77862 1292 77918
rect 1348 77862 1416 77918
rect 1472 77862 1568 77918
rect 948 77794 1568 77862
rect 948 77738 1044 77794
rect 1100 77738 1168 77794
rect 1224 77738 1292 77794
rect 1348 77738 1416 77794
rect 1472 77738 1568 77794
rect 948 77670 1568 77738
rect 948 77614 1044 77670
rect 1100 77614 1168 77670
rect 1224 77614 1292 77670
rect 1348 77614 1416 77670
rect 1472 77614 1568 77670
rect 948 77546 1568 77614
rect 948 77490 1044 77546
rect 1100 77490 1168 77546
rect 1224 77490 1292 77546
rect 1348 77490 1416 77546
rect 1472 77490 1568 77546
rect 948 59918 1568 77490
rect 948 59862 1044 59918
rect 1100 59862 1168 59918
rect 1224 59862 1292 59918
rect 1348 59862 1416 59918
rect 1472 59862 1568 59918
rect 948 59794 1568 59862
rect 948 59738 1044 59794
rect 1100 59738 1168 59794
rect 1224 59738 1292 59794
rect 1348 59738 1416 59794
rect 1472 59738 1568 59794
rect 948 59670 1568 59738
rect 948 59614 1044 59670
rect 1100 59614 1168 59670
rect 1224 59614 1292 59670
rect 1348 59614 1416 59670
rect 1472 59614 1568 59670
rect 948 59546 1568 59614
rect 948 59490 1044 59546
rect 1100 59490 1168 59546
rect 1224 59490 1292 59546
rect 1348 59490 1416 59546
rect 1472 59490 1568 59546
rect 948 41918 1568 59490
rect 948 41862 1044 41918
rect 1100 41862 1168 41918
rect 1224 41862 1292 41918
rect 1348 41862 1416 41918
rect 1472 41862 1568 41918
rect 948 41794 1568 41862
rect 948 41738 1044 41794
rect 1100 41738 1168 41794
rect 1224 41738 1292 41794
rect 1348 41738 1416 41794
rect 1472 41738 1568 41794
rect 948 41670 1568 41738
rect 948 41614 1044 41670
rect 1100 41614 1168 41670
rect 1224 41614 1292 41670
rect 1348 41614 1416 41670
rect 1472 41614 1568 41670
rect 948 41546 1568 41614
rect 948 41490 1044 41546
rect 1100 41490 1168 41546
rect 1224 41490 1292 41546
rect 1348 41490 1416 41546
rect 1472 41490 1568 41546
rect 948 23918 1568 41490
rect 948 23862 1044 23918
rect 1100 23862 1168 23918
rect 1224 23862 1292 23918
rect 1348 23862 1416 23918
rect 1472 23862 1568 23918
rect 948 23794 1568 23862
rect 948 23738 1044 23794
rect 1100 23738 1168 23794
rect 1224 23738 1292 23794
rect 1348 23738 1416 23794
rect 1472 23738 1568 23794
rect 948 23670 1568 23738
rect 948 23614 1044 23670
rect 1100 23614 1168 23670
rect 1224 23614 1292 23670
rect 1348 23614 1416 23670
rect 1472 23614 1568 23670
rect 948 23546 1568 23614
rect 948 23490 1044 23546
rect 1100 23490 1168 23546
rect 1224 23490 1292 23546
rect 1348 23490 1416 23546
rect 1472 23490 1568 23546
rect 948 5918 1568 23490
rect 948 5862 1044 5918
rect 1100 5862 1168 5918
rect 1224 5862 1292 5918
rect 1348 5862 1416 5918
rect 1472 5862 1568 5918
rect 948 5794 1568 5862
rect 948 5738 1044 5794
rect 1100 5738 1168 5794
rect 1224 5738 1292 5794
rect 1348 5738 1416 5794
rect 1472 5738 1568 5794
rect 948 5670 1568 5738
rect 948 5614 1044 5670
rect 1100 5614 1168 5670
rect 1224 5614 1292 5670
rect 1348 5614 1416 5670
rect 1472 5614 1568 5670
rect 948 5546 1568 5614
rect 948 5490 1044 5546
rect 1100 5490 1168 5546
rect 1224 5490 1292 5546
rect 1348 5490 1416 5546
rect 1472 5490 1568 5546
rect 948 1808 1568 5490
rect 948 1752 1044 1808
rect 1100 1752 1168 1808
rect 1224 1752 1292 1808
rect 1348 1752 1416 1808
rect 1472 1752 1568 1808
rect 948 1684 1568 1752
rect 948 1628 1044 1684
rect 1100 1628 1168 1684
rect 1224 1628 1292 1684
rect 1348 1628 1416 1684
rect 1472 1628 1568 1684
rect 948 1560 1568 1628
rect 948 1504 1044 1560
rect 1100 1504 1168 1560
rect 1224 1504 1292 1560
rect 1348 1504 1416 1560
rect 1472 1504 1568 1560
rect 948 1436 1568 1504
rect 948 1380 1044 1436
rect 1100 1380 1168 1436
rect 1224 1380 1292 1436
rect 1348 1380 1416 1436
rect 1472 1380 1568 1436
rect 948 1284 1568 1380
rect 5058 598380 5678 599436
rect 5058 598324 5154 598380
rect 5210 598324 5278 598380
rect 5334 598324 5402 598380
rect 5458 598324 5526 598380
rect 5582 598324 5678 598380
rect 5058 598256 5678 598324
rect 5058 598200 5154 598256
rect 5210 598200 5278 598256
rect 5334 598200 5402 598256
rect 5458 598200 5526 598256
rect 5582 598200 5678 598256
rect 5058 598132 5678 598200
rect 5058 598076 5154 598132
rect 5210 598076 5278 598132
rect 5334 598076 5402 598132
rect 5458 598076 5526 598132
rect 5582 598076 5678 598132
rect 5058 598008 5678 598076
rect 5058 597952 5154 598008
rect 5210 597952 5278 598008
rect 5334 597952 5402 598008
rect 5458 597952 5526 598008
rect 5582 597952 5678 598008
rect 5058 581918 5678 597952
rect 8778 599340 9398 599436
rect 8778 599284 8874 599340
rect 8930 599284 8998 599340
rect 9054 599284 9122 599340
rect 9178 599284 9246 599340
rect 9302 599284 9398 599340
rect 8778 599216 9398 599284
rect 8778 599160 8874 599216
rect 8930 599160 8998 599216
rect 9054 599160 9122 599216
rect 9178 599160 9246 599216
rect 9302 599160 9398 599216
rect 8778 599092 9398 599160
rect 8778 599036 8874 599092
rect 8930 599036 8998 599092
rect 9054 599036 9122 599092
rect 9178 599036 9246 599092
rect 9302 599036 9398 599092
rect 8778 598968 9398 599036
rect 8778 598912 8874 598968
rect 8930 598912 8998 598968
rect 9054 598912 9122 598968
rect 9178 598912 9246 598968
rect 9302 598912 9398 598968
rect 8778 596288 9398 598912
rect 23058 598380 23678 599436
rect 23058 598324 23154 598380
rect 23210 598324 23278 598380
rect 23334 598324 23402 598380
rect 23458 598324 23526 598380
rect 23582 598324 23678 598380
rect 23058 598256 23678 598324
rect 23058 598200 23154 598256
rect 23210 598200 23278 598256
rect 23334 598200 23402 598256
rect 23458 598200 23526 598256
rect 23582 598200 23678 598256
rect 23058 598132 23678 598200
rect 23058 598076 23154 598132
rect 23210 598076 23278 598132
rect 23334 598076 23402 598132
rect 23458 598076 23526 598132
rect 23582 598076 23678 598132
rect 23058 598008 23678 598076
rect 23058 597952 23154 598008
rect 23210 597952 23278 598008
rect 23334 597952 23402 598008
rect 23458 597952 23526 598008
rect 23582 597952 23678 598008
rect 23058 596288 23678 597952
rect 26778 599340 27398 599436
rect 26778 599284 26874 599340
rect 26930 599284 26998 599340
rect 27054 599284 27122 599340
rect 27178 599284 27246 599340
rect 27302 599284 27398 599340
rect 26778 599216 27398 599284
rect 26778 599160 26874 599216
rect 26930 599160 26998 599216
rect 27054 599160 27122 599216
rect 27178 599160 27246 599216
rect 27302 599160 27398 599216
rect 26778 599092 27398 599160
rect 26778 599036 26874 599092
rect 26930 599036 26998 599092
rect 27054 599036 27122 599092
rect 27178 599036 27246 599092
rect 27302 599036 27398 599092
rect 26778 598968 27398 599036
rect 26778 598912 26874 598968
rect 26930 598912 26998 598968
rect 27054 598912 27122 598968
rect 27178 598912 27246 598968
rect 27302 598912 27398 598968
rect 26778 596288 27398 598912
rect 41058 598380 41678 599436
rect 41058 598324 41154 598380
rect 41210 598324 41278 598380
rect 41334 598324 41402 598380
rect 41458 598324 41526 598380
rect 41582 598324 41678 598380
rect 41058 598256 41678 598324
rect 41058 598200 41154 598256
rect 41210 598200 41278 598256
rect 41334 598200 41402 598256
rect 41458 598200 41526 598256
rect 41582 598200 41678 598256
rect 41058 598132 41678 598200
rect 41058 598076 41154 598132
rect 41210 598076 41278 598132
rect 41334 598076 41402 598132
rect 41458 598076 41526 598132
rect 41582 598076 41678 598132
rect 41058 598008 41678 598076
rect 41058 597952 41154 598008
rect 41210 597952 41278 598008
rect 41334 597952 41402 598008
rect 41458 597952 41526 598008
rect 41582 597952 41678 598008
rect 41058 596288 41678 597952
rect 44778 599340 45398 599436
rect 44778 599284 44874 599340
rect 44930 599284 44998 599340
rect 45054 599284 45122 599340
rect 45178 599284 45246 599340
rect 45302 599284 45398 599340
rect 44778 599216 45398 599284
rect 44778 599160 44874 599216
rect 44930 599160 44998 599216
rect 45054 599160 45122 599216
rect 45178 599160 45246 599216
rect 45302 599160 45398 599216
rect 44778 599092 45398 599160
rect 44778 599036 44874 599092
rect 44930 599036 44998 599092
rect 45054 599036 45122 599092
rect 45178 599036 45246 599092
rect 45302 599036 45398 599092
rect 44778 598968 45398 599036
rect 44778 598912 44874 598968
rect 44930 598912 44998 598968
rect 45054 598912 45122 598968
rect 45178 598912 45246 598968
rect 45302 598912 45398 598968
rect 44778 596288 45398 598912
rect 59058 598380 59678 599436
rect 59058 598324 59154 598380
rect 59210 598324 59278 598380
rect 59334 598324 59402 598380
rect 59458 598324 59526 598380
rect 59582 598324 59678 598380
rect 59058 598256 59678 598324
rect 59058 598200 59154 598256
rect 59210 598200 59278 598256
rect 59334 598200 59402 598256
rect 59458 598200 59526 598256
rect 59582 598200 59678 598256
rect 59058 598132 59678 598200
rect 59058 598076 59154 598132
rect 59210 598076 59278 598132
rect 59334 598076 59402 598132
rect 59458 598076 59526 598132
rect 59582 598076 59678 598132
rect 59058 598008 59678 598076
rect 59058 597952 59154 598008
rect 59210 597952 59278 598008
rect 59334 597952 59402 598008
rect 59458 597952 59526 598008
rect 59582 597952 59678 598008
rect 59058 596288 59678 597952
rect 62778 599340 63398 599436
rect 62778 599284 62874 599340
rect 62930 599284 62998 599340
rect 63054 599284 63122 599340
rect 63178 599284 63246 599340
rect 63302 599284 63398 599340
rect 62778 599216 63398 599284
rect 62778 599160 62874 599216
rect 62930 599160 62998 599216
rect 63054 599160 63122 599216
rect 63178 599160 63246 599216
rect 63302 599160 63398 599216
rect 62778 599092 63398 599160
rect 62778 599036 62874 599092
rect 62930 599036 62998 599092
rect 63054 599036 63122 599092
rect 63178 599036 63246 599092
rect 63302 599036 63398 599092
rect 62778 598968 63398 599036
rect 62778 598912 62874 598968
rect 62930 598912 62998 598968
rect 63054 598912 63122 598968
rect 63178 598912 63246 598968
rect 63302 598912 63398 598968
rect 62778 596288 63398 598912
rect 77058 598380 77678 599436
rect 77058 598324 77154 598380
rect 77210 598324 77278 598380
rect 77334 598324 77402 598380
rect 77458 598324 77526 598380
rect 77582 598324 77678 598380
rect 77058 598256 77678 598324
rect 77058 598200 77154 598256
rect 77210 598200 77278 598256
rect 77334 598200 77402 598256
rect 77458 598200 77526 598256
rect 77582 598200 77678 598256
rect 77058 598132 77678 598200
rect 77058 598076 77154 598132
rect 77210 598076 77278 598132
rect 77334 598076 77402 598132
rect 77458 598076 77526 598132
rect 77582 598076 77678 598132
rect 77058 598008 77678 598076
rect 77058 597952 77154 598008
rect 77210 597952 77278 598008
rect 77334 597952 77402 598008
rect 77458 597952 77526 598008
rect 77582 597952 77678 598008
rect 77058 596288 77678 597952
rect 80778 599340 81398 599436
rect 80778 599284 80874 599340
rect 80930 599284 80998 599340
rect 81054 599284 81122 599340
rect 81178 599284 81246 599340
rect 81302 599284 81398 599340
rect 80778 599216 81398 599284
rect 80778 599160 80874 599216
rect 80930 599160 80998 599216
rect 81054 599160 81122 599216
rect 81178 599160 81246 599216
rect 81302 599160 81398 599216
rect 80778 599092 81398 599160
rect 80778 599036 80874 599092
rect 80930 599036 80998 599092
rect 81054 599036 81122 599092
rect 81178 599036 81246 599092
rect 81302 599036 81398 599092
rect 80778 598968 81398 599036
rect 80778 598912 80874 598968
rect 80930 598912 80998 598968
rect 81054 598912 81122 598968
rect 81178 598912 81246 598968
rect 81302 598912 81398 598968
rect 80778 596288 81398 598912
rect 95058 598380 95678 599436
rect 95058 598324 95154 598380
rect 95210 598324 95278 598380
rect 95334 598324 95402 598380
rect 95458 598324 95526 598380
rect 95582 598324 95678 598380
rect 95058 598256 95678 598324
rect 95058 598200 95154 598256
rect 95210 598200 95278 598256
rect 95334 598200 95402 598256
rect 95458 598200 95526 598256
rect 95582 598200 95678 598256
rect 95058 598132 95678 598200
rect 95058 598076 95154 598132
rect 95210 598076 95278 598132
rect 95334 598076 95402 598132
rect 95458 598076 95526 598132
rect 95582 598076 95678 598132
rect 95058 598008 95678 598076
rect 95058 597952 95154 598008
rect 95210 597952 95278 598008
rect 95334 597952 95402 598008
rect 95458 597952 95526 598008
rect 95582 597952 95678 598008
rect 95058 596288 95678 597952
rect 98778 599340 99398 599436
rect 98778 599284 98874 599340
rect 98930 599284 98998 599340
rect 99054 599284 99122 599340
rect 99178 599284 99246 599340
rect 99302 599284 99398 599340
rect 98778 599216 99398 599284
rect 98778 599160 98874 599216
rect 98930 599160 98998 599216
rect 99054 599160 99122 599216
rect 99178 599160 99246 599216
rect 99302 599160 99398 599216
rect 98778 599092 99398 599160
rect 98778 599036 98874 599092
rect 98930 599036 98998 599092
rect 99054 599036 99122 599092
rect 99178 599036 99246 599092
rect 99302 599036 99398 599092
rect 98778 598968 99398 599036
rect 98778 598912 98874 598968
rect 98930 598912 98998 598968
rect 99054 598912 99122 598968
rect 99178 598912 99246 598968
rect 99302 598912 99398 598968
rect 98778 596288 99398 598912
rect 113058 598380 113678 599436
rect 113058 598324 113154 598380
rect 113210 598324 113278 598380
rect 113334 598324 113402 598380
rect 113458 598324 113526 598380
rect 113582 598324 113678 598380
rect 113058 598256 113678 598324
rect 113058 598200 113154 598256
rect 113210 598200 113278 598256
rect 113334 598200 113402 598256
rect 113458 598200 113526 598256
rect 113582 598200 113678 598256
rect 113058 598132 113678 598200
rect 113058 598076 113154 598132
rect 113210 598076 113278 598132
rect 113334 598076 113402 598132
rect 113458 598076 113526 598132
rect 113582 598076 113678 598132
rect 113058 598008 113678 598076
rect 113058 597952 113154 598008
rect 113210 597952 113278 598008
rect 113334 597952 113402 598008
rect 113458 597952 113526 598008
rect 113582 597952 113678 598008
rect 113058 596288 113678 597952
rect 116778 599340 117398 599436
rect 116778 599284 116874 599340
rect 116930 599284 116998 599340
rect 117054 599284 117122 599340
rect 117178 599284 117246 599340
rect 117302 599284 117398 599340
rect 116778 599216 117398 599284
rect 116778 599160 116874 599216
rect 116930 599160 116998 599216
rect 117054 599160 117122 599216
rect 117178 599160 117246 599216
rect 117302 599160 117398 599216
rect 116778 599092 117398 599160
rect 116778 599036 116874 599092
rect 116930 599036 116998 599092
rect 117054 599036 117122 599092
rect 117178 599036 117246 599092
rect 117302 599036 117398 599092
rect 116778 598968 117398 599036
rect 116778 598912 116874 598968
rect 116930 598912 116998 598968
rect 117054 598912 117122 598968
rect 117178 598912 117246 598968
rect 117302 598912 117398 598968
rect 116778 596288 117398 598912
rect 131058 598380 131678 599436
rect 131058 598324 131154 598380
rect 131210 598324 131278 598380
rect 131334 598324 131402 598380
rect 131458 598324 131526 598380
rect 131582 598324 131678 598380
rect 131058 598256 131678 598324
rect 131058 598200 131154 598256
rect 131210 598200 131278 598256
rect 131334 598200 131402 598256
rect 131458 598200 131526 598256
rect 131582 598200 131678 598256
rect 131058 598132 131678 598200
rect 131058 598076 131154 598132
rect 131210 598076 131278 598132
rect 131334 598076 131402 598132
rect 131458 598076 131526 598132
rect 131582 598076 131678 598132
rect 131058 598008 131678 598076
rect 131058 597952 131154 598008
rect 131210 597952 131278 598008
rect 131334 597952 131402 598008
rect 131458 597952 131526 598008
rect 131582 597952 131678 598008
rect 131058 596288 131678 597952
rect 134778 599340 135398 599436
rect 134778 599284 134874 599340
rect 134930 599284 134998 599340
rect 135054 599284 135122 599340
rect 135178 599284 135246 599340
rect 135302 599284 135398 599340
rect 134778 599216 135398 599284
rect 134778 599160 134874 599216
rect 134930 599160 134998 599216
rect 135054 599160 135122 599216
rect 135178 599160 135246 599216
rect 135302 599160 135398 599216
rect 134778 599092 135398 599160
rect 134778 599036 134874 599092
rect 134930 599036 134998 599092
rect 135054 599036 135122 599092
rect 135178 599036 135246 599092
rect 135302 599036 135398 599092
rect 134778 598968 135398 599036
rect 134778 598912 134874 598968
rect 134930 598912 134998 598968
rect 135054 598912 135122 598968
rect 135178 598912 135246 598968
rect 135302 598912 135398 598968
rect 134778 596288 135398 598912
rect 149058 598380 149678 599436
rect 149058 598324 149154 598380
rect 149210 598324 149278 598380
rect 149334 598324 149402 598380
rect 149458 598324 149526 598380
rect 149582 598324 149678 598380
rect 149058 598256 149678 598324
rect 149058 598200 149154 598256
rect 149210 598200 149278 598256
rect 149334 598200 149402 598256
rect 149458 598200 149526 598256
rect 149582 598200 149678 598256
rect 149058 598132 149678 598200
rect 149058 598076 149154 598132
rect 149210 598076 149278 598132
rect 149334 598076 149402 598132
rect 149458 598076 149526 598132
rect 149582 598076 149678 598132
rect 149058 598008 149678 598076
rect 149058 597952 149154 598008
rect 149210 597952 149278 598008
rect 149334 597952 149402 598008
rect 149458 597952 149526 598008
rect 149582 597952 149678 598008
rect 149058 596288 149678 597952
rect 152778 599340 153398 599436
rect 152778 599284 152874 599340
rect 152930 599284 152998 599340
rect 153054 599284 153122 599340
rect 153178 599284 153246 599340
rect 153302 599284 153398 599340
rect 152778 599216 153398 599284
rect 152778 599160 152874 599216
rect 152930 599160 152998 599216
rect 153054 599160 153122 599216
rect 153178 599160 153246 599216
rect 153302 599160 153398 599216
rect 152778 599092 153398 599160
rect 152778 599036 152874 599092
rect 152930 599036 152998 599092
rect 153054 599036 153122 599092
rect 153178 599036 153246 599092
rect 153302 599036 153398 599092
rect 152778 598968 153398 599036
rect 152778 598912 152874 598968
rect 152930 598912 152998 598968
rect 153054 598912 153122 598968
rect 153178 598912 153246 598968
rect 153302 598912 153398 598968
rect 152778 596288 153398 598912
rect 167058 598380 167678 599436
rect 167058 598324 167154 598380
rect 167210 598324 167278 598380
rect 167334 598324 167402 598380
rect 167458 598324 167526 598380
rect 167582 598324 167678 598380
rect 167058 598256 167678 598324
rect 167058 598200 167154 598256
rect 167210 598200 167278 598256
rect 167334 598200 167402 598256
rect 167458 598200 167526 598256
rect 167582 598200 167678 598256
rect 167058 598132 167678 598200
rect 167058 598076 167154 598132
rect 167210 598076 167278 598132
rect 167334 598076 167402 598132
rect 167458 598076 167526 598132
rect 167582 598076 167678 598132
rect 167058 598008 167678 598076
rect 167058 597952 167154 598008
rect 167210 597952 167278 598008
rect 167334 597952 167402 598008
rect 167458 597952 167526 598008
rect 167582 597952 167678 598008
rect 167058 596288 167678 597952
rect 170778 599340 171398 599436
rect 170778 599284 170874 599340
rect 170930 599284 170998 599340
rect 171054 599284 171122 599340
rect 171178 599284 171246 599340
rect 171302 599284 171398 599340
rect 170778 599216 171398 599284
rect 170778 599160 170874 599216
rect 170930 599160 170998 599216
rect 171054 599160 171122 599216
rect 171178 599160 171246 599216
rect 171302 599160 171398 599216
rect 170778 599092 171398 599160
rect 170778 599036 170874 599092
rect 170930 599036 170998 599092
rect 171054 599036 171122 599092
rect 171178 599036 171246 599092
rect 171302 599036 171398 599092
rect 170778 598968 171398 599036
rect 170778 598912 170874 598968
rect 170930 598912 170998 598968
rect 171054 598912 171122 598968
rect 171178 598912 171246 598968
rect 171302 598912 171398 598968
rect 170778 596288 171398 598912
rect 185058 598380 185678 599436
rect 185058 598324 185154 598380
rect 185210 598324 185278 598380
rect 185334 598324 185402 598380
rect 185458 598324 185526 598380
rect 185582 598324 185678 598380
rect 185058 598256 185678 598324
rect 185058 598200 185154 598256
rect 185210 598200 185278 598256
rect 185334 598200 185402 598256
rect 185458 598200 185526 598256
rect 185582 598200 185678 598256
rect 185058 598132 185678 598200
rect 185058 598076 185154 598132
rect 185210 598076 185278 598132
rect 185334 598076 185402 598132
rect 185458 598076 185526 598132
rect 185582 598076 185678 598132
rect 185058 598008 185678 598076
rect 185058 597952 185154 598008
rect 185210 597952 185278 598008
rect 185334 597952 185402 598008
rect 185458 597952 185526 598008
rect 185582 597952 185678 598008
rect 185058 596288 185678 597952
rect 188778 599340 189398 599436
rect 188778 599284 188874 599340
rect 188930 599284 188998 599340
rect 189054 599284 189122 599340
rect 189178 599284 189246 599340
rect 189302 599284 189398 599340
rect 188778 599216 189398 599284
rect 188778 599160 188874 599216
rect 188930 599160 188998 599216
rect 189054 599160 189122 599216
rect 189178 599160 189246 599216
rect 189302 599160 189398 599216
rect 188778 599092 189398 599160
rect 188778 599036 188874 599092
rect 188930 599036 188998 599092
rect 189054 599036 189122 599092
rect 189178 599036 189246 599092
rect 189302 599036 189398 599092
rect 188778 598968 189398 599036
rect 188778 598912 188874 598968
rect 188930 598912 188998 598968
rect 189054 598912 189122 598968
rect 189178 598912 189246 598968
rect 189302 598912 189398 598968
rect 188778 596288 189398 598912
rect 203058 598380 203678 599436
rect 203058 598324 203154 598380
rect 203210 598324 203278 598380
rect 203334 598324 203402 598380
rect 203458 598324 203526 598380
rect 203582 598324 203678 598380
rect 203058 598256 203678 598324
rect 203058 598200 203154 598256
rect 203210 598200 203278 598256
rect 203334 598200 203402 598256
rect 203458 598200 203526 598256
rect 203582 598200 203678 598256
rect 203058 598132 203678 598200
rect 203058 598076 203154 598132
rect 203210 598076 203278 598132
rect 203334 598076 203402 598132
rect 203458 598076 203526 598132
rect 203582 598076 203678 598132
rect 203058 598008 203678 598076
rect 203058 597952 203154 598008
rect 203210 597952 203278 598008
rect 203334 597952 203402 598008
rect 203458 597952 203526 598008
rect 203582 597952 203678 598008
rect 203058 596288 203678 597952
rect 206778 599340 207398 599436
rect 206778 599284 206874 599340
rect 206930 599284 206998 599340
rect 207054 599284 207122 599340
rect 207178 599284 207246 599340
rect 207302 599284 207398 599340
rect 206778 599216 207398 599284
rect 206778 599160 206874 599216
rect 206930 599160 206998 599216
rect 207054 599160 207122 599216
rect 207178 599160 207246 599216
rect 207302 599160 207398 599216
rect 206778 599092 207398 599160
rect 206778 599036 206874 599092
rect 206930 599036 206998 599092
rect 207054 599036 207122 599092
rect 207178 599036 207246 599092
rect 207302 599036 207398 599092
rect 206778 598968 207398 599036
rect 206778 598912 206874 598968
rect 206930 598912 206998 598968
rect 207054 598912 207122 598968
rect 207178 598912 207246 598968
rect 207302 598912 207398 598968
rect 206778 596288 207398 598912
rect 221058 598380 221678 599436
rect 221058 598324 221154 598380
rect 221210 598324 221278 598380
rect 221334 598324 221402 598380
rect 221458 598324 221526 598380
rect 221582 598324 221678 598380
rect 221058 598256 221678 598324
rect 221058 598200 221154 598256
rect 221210 598200 221278 598256
rect 221334 598200 221402 598256
rect 221458 598200 221526 598256
rect 221582 598200 221678 598256
rect 221058 598132 221678 598200
rect 221058 598076 221154 598132
rect 221210 598076 221278 598132
rect 221334 598076 221402 598132
rect 221458 598076 221526 598132
rect 221582 598076 221678 598132
rect 221058 598008 221678 598076
rect 221058 597952 221154 598008
rect 221210 597952 221278 598008
rect 221334 597952 221402 598008
rect 221458 597952 221526 598008
rect 221582 597952 221678 598008
rect 221058 596288 221678 597952
rect 224778 599340 225398 599436
rect 224778 599284 224874 599340
rect 224930 599284 224998 599340
rect 225054 599284 225122 599340
rect 225178 599284 225246 599340
rect 225302 599284 225398 599340
rect 224778 599216 225398 599284
rect 224778 599160 224874 599216
rect 224930 599160 224998 599216
rect 225054 599160 225122 599216
rect 225178 599160 225246 599216
rect 225302 599160 225398 599216
rect 224778 599092 225398 599160
rect 224778 599036 224874 599092
rect 224930 599036 224998 599092
rect 225054 599036 225122 599092
rect 225178 599036 225246 599092
rect 225302 599036 225398 599092
rect 224778 598968 225398 599036
rect 224778 598912 224874 598968
rect 224930 598912 224998 598968
rect 225054 598912 225122 598968
rect 225178 598912 225246 598968
rect 225302 598912 225398 598968
rect 224778 596288 225398 598912
rect 239058 598380 239678 599436
rect 239058 598324 239154 598380
rect 239210 598324 239278 598380
rect 239334 598324 239402 598380
rect 239458 598324 239526 598380
rect 239582 598324 239678 598380
rect 239058 598256 239678 598324
rect 239058 598200 239154 598256
rect 239210 598200 239278 598256
rect 239334 598200 239402 598256
rect 239458 598200 239526 598256
rect 239582 598200 239678 598256
rect 239058 598132 239678 598200
rect 239058 598076 239154 598132
rect 239210 598076 239278 598132
rect 239334 598076 239402 598132
rect 239458 598076 239526 598132
rect 239582 598076 239678 598132
rect 239058 598008 239678 598076
rect 239058 597952 239154 598008
rect 239210 597952 239278 598008
rect 239334 597952 239402 598008
rect 239458 597952 239526 598008
rect 239582 597952 239678 598008
rect 239058 596288 239678 597952
rect 242778 599340 243398 599436
rect 242778 599284 242874 599340
rect 242930 599284 242998 599340
rect 243054 599284 243122 599340
rect 243178 599284 243246 599340
rect 243302 599284 243398 599340
rect 242778 599216 243398 599284
rect 242778 599160 242874 599216
rect 242930 599160 242998 599216
rect 243054 599160 243122 599216
rect 243178 599160 243246 599216
rect 243302 599160 243398 599216
rect 242778 599092 243398 599160
rect 242778 599036 242874 599092
rect 242930 599036 242998 599092
rect 243054 599036 243122 599092
rect 243178 599036 243246 599092
rect 243302 599036 243398 599092
rect 242778 598968 243398 599036
rect 242778 598912 242874 598968
rect 242930 598912 242998 598968
rect 243054 598912 243122 598968
rect 243178 598912 243246 598968
rect 243302 598912 243398 598968
rect 242778 596288 243398 598912
rect 257058 598380 257678 599436
rect 257058 598324 257154 598380
rect 257210 598324 257278 598380
rect 257334 598324 257402 598380
rect 257458 598324 257526 598380
rect 257582 598324 257678 598380
rect 257058 598256 257678 598324
rect 257058 598200 257154 598256
rect 257210 598200 257278 598256
rect 257334 598200 257402 598256
rect 257458 598200 257526 598256
rect 257582 598200 257678 598256
rect 257058 598132 257678 598200
rect 257058 598076 257154 598132
rect 257210 598076 257278 598132
rect 257334 598076 257402 598132
rect 257458 598076 257526 598132
rect 257582 598076 257678 598132
rect 257058 598008 257678 598076
rect 257058 597952 257154 598008
rect 257210 597952 257278 598008
rect 257334 597952 257402 598008
rect 257458 597952 257526 598008
rect 257582 597952 257678 598008
rect 257058 596288 257678 597952
rect 260778 599340 261398 599436
rect 260778 599284 260874 599340
rect 260930 599284 260998 599340
rect 261054 599284 261122 599340
rect 261178 599284 261246 599340
rect 261302 599284 261398 599340
rect 260778 599216 261398 599284
rect 260778 599160 260874 599216
rect 260930 599160 260998 599216
rect 261054 599160 261122 599216
rect 261178 599160 261246 599216
rect 261302 599160 261398 599216
rect 260778 599092 261398 599160
rect 260778 599036 260874 599092
rect 260930 599036 260998 599092
rect 261054 599036 261122 599092
rect 261178 599036 261246 599092
rect 261302 599036 261398 599092
rect 260778 598968 261398 599036
rect 260778 598912 260874 598968
rect 260930 598912 260998 598968
rect 261054 598912 261122 598968
rect 261178 598912 261246 598968
rect 261302 598912 261398 598968
rect 260778 596288 261398 598912
rect 275058 598380 275678 599436
rect 275058 598324 275154 598380
rect 275210 598324 275278 598380
rect 275334 598324 275402 598380
rect 275458 598324 275526 598380
rect 275582 598324 275678 598380
rect 275058 598256 275678 598324
rect 275058 598200 275154 598256
rect 275210 598200 275278 598256
rect 275334 598200 275402 598256
rect 275458 598200 275526 598256
rect 275582 598200 275678 598256
rect 275058 598132 275678 598200
rect 275058 598076 275154 598132
rect 275210 598076 275278 598132
rect 275334 598076 275402 598132
rect 275458 598076 275526 598132
rect 275582 598076 275678 598132
rect 275058 598008 275678 598076
rect 275058 597952 275154 598008
rect 275210 597952 275278 598008
rect 275334 597952 275402 598008
rect 275458 597952 275526 598008
rect 275582 597952 275678 598008
rect 275058 596288 275678 597952
rect 278778 599340 279398 599436
rect 278778 599284 278874 599340
rect 278930 599284 278998 599340
rect 279054 599284 279122 599340
rect 279178 599284 279246 599340
rect 279302 599284 279398 599340
rect 278778 599216 279398 599284
rect 278778 599160 278874 599216
rect 278930 599160 278998 599216
rect 279054 599160 279122 599216
rect 279178 599160 279246 599216
rect 279302 599160 279398 599216
rect 278778 599092 279398 599160
rect 278778 599036 278874 599092
rect 278930 599036 278998 599092
rect 279054 599036 279122 599092
rect 279178 599036 279246 599092
rect 279302 599036 279398 599092
rect 278778 598968 279398 599036
rect 278778 598912 278874 598968
rect 278930 598912 278998 598968
rect 279054 598912 279122 598968
rect 279178 598912 279246 598968
rect 279302 598912 279398 598968
rect 278778 596288 279398 598912
rect 293058 598380 293678 599436
rect 293058 598324 293154 598380
rect 293210 598324 293278 598380
rect 293334 598324 293402 598380
rect 293458 598324 293526 598380
rect 293582 598324 293678 598380
rect 293058 598256 293678 598324
rect 293058 598200 293154 598256
rect 293210 598200 293278 598256
rect 293334 598200 293402 598256
rect 293458 598200 293526 598256
rect 293582 598200 293678 598256
rect 293058 598132 293678 598200
rect 293058 598076 293154 598132
rect 293210 598076 293278 598132
rect 293334 598076 293402 598132
rect 293458 598076 293526 598132
rect 293582 598076 293678 598132
rect 293058 598008 293678 598076
rect 293058 597952 293154 598008
rect 293210 597952 293278 598008
rect 293334 597952 293402 598008
rect 293458 597952 293526 598008
rect 293582 597952 293678 598008
rect 293058 596288 293678 597952
rect 296778 599340 297398 599436
rect 296778 599284 296874 599340
rect 296930 599284 296998 599340
rect 297054 599284 297122 599340
rect 297178 599284 297246 599340
rect 297302 599284 297398 599340
rect 296778 599216 297398 599284
rect 296778 599160 296874 599216
rect 296930 599160 296998 599216
rect 297054 599160 297122 599216
rect 297178 599160 297246 599216
rect 297302 599160 297398 599216
rect 296778 599092 297398 599160
rect 296778 599036 296874 599092
rect 296930 599036 296998 599092
rect 297054 599036 297122 599092
rect 297178 599036 297246 599092
rect 297302 599036 297398 599092
rect 296778 598968 297398 599036
rect 296778 598912 296874 598968
rect 296930 598912 296998 598968
rect 297054 598912 297122 598968
rect 297178 598912 297246 598968
rect 297302 598912 297398 598968
rect 296778 596288 297398 598912
rect 311058 598380 311678 599436
rect 311058 598324 311154 598380
rect 311210 598324 311278 598380
rect 311334 598324 311402 598380
rect 311458 598324 311526 598380
rect 311582 598324 311678 598380
rect 311058 598256 311678 598324
rect 311058 598200 311154 598256
rect 311210 598200 311278 598256
rect 311334 598200 311402 598256
rect 311458 598200 311526 598256
rect 311582 598200 311678 598256
rect 311058 598132 311678 598200
rect 311058 598076 311154 598132
rect 311210 598076 311278 598132
rect 311334 598076 311402 598132
rect 311458 598076 311526 598132
rect 311582 598076 311678 598132
rect 311058 598008 311678 598076
rect 311058 597952 311154 598008
rect 311210 597952 311278 598008
rect 311334 597952 311402 598008
rect 311458 597952 311526 598008
rect 311582 597952 311678 598008
rect 311058 596288 311678 597952
rect 314778 599340 315398 599436
rect 314778 599284 314874 599340
rect 314930 599284 314998 599340
rect 315054 599284 315122 599340
rect 315178 599284 315246 599340
rect 315302 599284 315398 599340
rect 314778 599216 315398 599284
rect 314778 599160 314874 599216
rect 314930 599160 314998 599216
rect 315054 599160 315122 599216
rect 315178 599160 315246 599216
rect 315302 599160 315398 599216
rect 314778 599092 315398 599160
rect 314778 599036 314874 599092
rect 314930 599036 314998 599092
rect 315054 599036 315122 599092
rect 315178 599036 315246 599092
rect 315302 599036 315398 599092
rect 314778 598968 315398 599036
rect 314778 598912 314874 598968
rect 314930 598912 314998 598968
rect 315054 598912 315122 598968
rect 315178 598912 315246 598968
rect 315302 598912 315398 598968
rect 314778 596288 315398 598912
rect 329058 598380 329678 599436
rect 329058 598324 329154 598380
rect 329210 598324 329278 598380
rect 329334 598324 329402 598380
rect 329458 598324 329526 598380
rect 329582 598324 329678 598380
rect 329058 598256 329678 598324
rect 329058 598200 329154 598256
rect 329210 598200 329278 598256
rect 329334 598200 329402 598256
rect 329458 598200 329526 598256
rect 329582 598200 329678 598256
rect 329058 598132 329678 598200
rect 329058 598076 329154 598132
rect 329210 598076 329278 598132
rect 329334 598076 329402 598132
rect 329458 598076 329526 598132
rect 329582 598076 329678 598132
rect 329058 598008 329678 598076
rect 329058 597952 329154 598008
rect 329210 597952 329278 598008
rect 329334 597952 329402 598008
rect 329458 597952 329526 598008
rect 329582 597952 329678 598008
rect 329058 596288 329678 597952
rect 332778 599340 333398 599436
rect 332778 599284 332874 599340
rect 332930 599284 332998 599340
rect 333054 599284 333122 599340
rect 333178 599284 333246 599340
rect 333302 599284 333398 599340
rect 332778 599216 333398 599284
rect 332778 599160 332874 599216
rect 332930 599160 332998 599216
rect 333054 599160 333122 599216
rect 333178 599160 333246 599216
rect 333302 599160 333398 599216
rect 332778 599092 333398 599160
rect 332778 599036 332874 599092
rect 332930 599036 332998 599092
rect 333054 599036 333122 599092
rect 333178 599036 333246 599092
rect 333302 599036 333398 599092
rect 332778 598968 333398 599036
rect 332778 598912 332874 598968
rect 332930 598912 332998 598968
rect 333054 598912 333122 598968
rect 333178 598912 333246 598968
rect 333302 598912 333398 598968
rect 332778 596288 333398 598912
rect 347058 598380 347678 599436
rect 347058 598324 347154 598380
rect 347210 598324 347278 598380
rect 347334 598324 347402 598380
rect 347458 598324 347526 598380
rect 347582 598324 347678 598380
rect 347058 598256 347678 598324
rect 347058 598200 347154 598256
rect 347210 598200 347278 598256
rect 347334 598200 347402 598256
rect 347458 598200 347526 598256
rect 347582 598200 347678 598256
rect 347058 598132 347678 598200
rect 347058 598076 347154 598132
rect 347210 598076 347278 598132
rect 347334 598076 347402 598132
rect 347458 598076 347526 598132
rect 347582 598076 347678 598132
rect 347058 598008 347678 598076
rect 347058 597952 347154 598008
rect 347210 597952 347278 598008
rect 347334 597952 347402 598008
rect 347458 597952 347526 598008
rect 347582 597952 347678 598008
rect 347058 596288 347678 597952
rect 350778 599340 351398 599436
rect 350778 599284 350874 599340
rect 350930 599284 350998 599340
rect 351054 599284 351122 599340
rect 351178 599284 351246 599340
rect 351302 599284 351398 599340
rect 350778 599216 351398 599284
rect 350778 599160 350874 599216
rect 350930 599160 350998 599216
rect 351054 599160 351122 599216
rect 351178 599160 351246 599216
rect 351302 599160 351398 599216
rect 350778 599092 351398 599160
rect 350778 599036 350874 599092
rect 350930 599036 350998 599092
rect 351054 599036 351122 599092
rect 351178 599036 351246 599092
rect 351302 599036 351398 599092
rect 350778 598968 351398 599036
rect 350778 598912 350874 598968
rect 350930 598912 350998 598968
rect 351054 598912 351122 598968
rect 351178 598912 351246 598968
rect 351302 598912 351398 598968
rect 350778 596288 351398 598912
rect 365058 598380 365678 599436
rect 365058 598324 365154 598380
rect 365210 598324 365278 598380
rect 365334 598324 365402 598380
rect 365458 598324 365526 598380
rect 365582 598324 365678 598380
rect 365058 598256 365678 598324
rect 365058 598200 365154 598256
rect 365210 598200 365278 598256
rect 365334 598200 365402 598256
rect 365458 598200 365526 598256
rect 365582 598200 365678 598256
rect 365058 598132 365678 598200
rect 365058 598076 365154 598132
rect 365210 598076 365278 598132
rect 365334 598076 365402 598132
rect 365458 598076 365526 598132
rect 365582 598076 365678 598132
rect 365058 598008 365678 598076
rect 365058 597952 365154 598008
rect 365210 597952 365278 598008
rect 365334 597952 365402 598008
rect 365458 597952 365526 598008
rect 365582 597952 365678 598008
rect 365058 596288 365678 597952
rect 368778 599340 369398 599436
rect 368778 599284 368874 599340
rect 368930 599284 368998 599340
rect 369054 599284 369122 599340
rect 369178 599284 369246 599340
rect 369302 599284 369398 599340
rect 368778 599216 369398 599284
rect 368778 599160 368874 599216
rect 368930 599160 368998 599216
rect 369054 599160 369122 599216
rect 369178 599160 369246 599216
rect 369302 599160 369398 599216
rect 368778 599092 369398 599160
rect 368778 599036 368874 599092
rect 368930 599036 368998 599092
rect 369054 599036 369122 599092
rect 369178 599036 369246 599092
rect 369302 599036 369398 599092
rect 368778 598968 369398 599036
rect 368778 598912 368874 598968
rect 368930 598912 368998 598968
rect 369054 598912 369122 598968
rect 369178 598912 369246 598968
rect 369302 598912 369398 598968
rect 368778 596288 369398 598912
rect 383058 598380 383678 599436
rect 383058 598324 383154 598380
rect 383210 598324 383278 598380
rect 383334 598324 383402 598380
rect 383458 598324 383526 598380
rect 383582 598324 383678 598380
rect 383058 598256 383678 598324
rect 383058 598200 383154 598256
rect 383210 598200 383278 598256
rect 383334 598200 383402 598256
rect 383458 598200 383526 598256
rect 383582 598200 383678 598256
rect 383058 598132 383678 598200
rect 383058 598076 383154 598132
rect 383210 598076 383278 598132
rect 383334 598076 383402 598132
rect 383458 598076 383526 598132
rect 383582 598076 383678 598132
rect 383058 598008 383678 598076
rect 383058 597952 383154 598008
rect 383210 597952 383278 598008
rect 383334 597952 383402 598008
rect 383458 597952 383526 598008
rect 383582 597952 383678 598008
rect 383058 596288 383678 597952
rect 386778 599340 387398 599436
rect 386778 599284 386874 599340
rect 386930 599284 386998 599340
rect 387054 599284 387122 599340
rect 387178 599284 387246 599340
rect 387302 599284 387398 599340
rect 386778 599216 387398 599284
rect 386778 599160 386874 599216
rect 386930 599160 386998 599216
rect 387054 599160 387122 599216
rect 387178 599160 387246 599216
rect 387302 599160 387398 599216
rect 386778 599092 387398 599160
rect 386778 599036 386874 599092
rect 386930 599036 386998 599092
rect 387054 599036 387122 599092
rect 387178 599036 387246 599092
rect 387302 599036 387398 599092
rect 386778 598968 387398 599036
rect 386778 598912 386874 598968
rect 386930 598912 386998 598968
rect 387054 598912 387122 598968
rect 387178 598912 387246 598968
rect 387302 598912 387398 598968
rect 386778 596288 387398 598912
rect 401058 598380 401678 599436
rect 401058 598324 401154 598380
rect 401210 598324 401278 598380
rect 401334 598324 401402 598380
rect 401458 598324 401526 598380
rect 401582 598324 401678 598380
rect 401058 598256 401678 598324
rect 401058 598200 401154 598256
rect 401210 598200 401278 598256
rect 401334 598200 401402 598256
rect 401458 598200 401526 598256
rect 401582 598200 401678 598256
rect 401058 598132 401678 598200
rect 401058 598076 401154 598132
rect 401210 598076 401278 598132
rect 401334 598076 401402 598132
rect 401458 598076 401526 598132
rect 401582 598076 401678 598132
rect 401058 598008 401678 598076
rect 401058 597952 401154 598008
rect 401210 597952 401278 598008
rect 401334 597952 401402 598008
rect 401458 597952 401526 598008
rect 401582 597952 401678 598008
rect 401058 596288 401678 597952
rect 404778 599340 405398 599436
rect 404778 599284 404874 599340
rect 404930 599284 404998 599340
rect 405054 599284 405122 599340
rect 405178 599284 405246 599340
rect 405302 599284 405398 599340
rect 404778 599216 405398 599284
rect 404778 599160 404874 599216
rect 404930 599160 404998 599216
rect 405054 599160 405122 599216
rect 405178 599160 405246 599216
rect 405302 599160 405398 599216
rect 404778 599092 405398 599160
rect 404778 599036 404874 599092
rect 404930 599036 404998 599092
rect 405054 599036 405122 599092
rect 405178 599036 405246 599092
rect 405302 599036 405398 599092
rect 404778 598968 405398 599036
rect 404778 598912 404874 598968
rect 404930 598912 404998 598968
rect 405054 598912 405122 598968
rect 405178 598912 405246 598968
rect 405302 598912 405398 598968
rect 404778 596288 405398 598912
rect 419058 598380 419678 599436
rect 419058 598324 419154 598380
rect 419210 598324 419278 598380
rect 419334 598324 419402 598380
rect 419458 598324 419526 598380
rect 419582 598324 419678 598380
rect 419058 598256 419678 598324
rect 419058 598200 419154 598256
rect 419210 598200 419278 598256
rect 419334 598200 419402 598256
rect 419458 598200 419526 598256
rect 419582 598200 419678 598256
rect 419058 598132 419678 598200
rect 419058 598076 419154 598132
rect 419210 598076 419278 598132
rect 419334 598076 419402 598132
rect 419458 598076 419526 598132
rect 419582 598076 419678 598132
rect 419058 598008 419678 598076
rect 419058 597952 419154 598008
rect 419210 597952 419278 598008
rect 419334 597952 419402 598008
rect 419458 597952 419526 598008
rect 419582 597952 419678 598008
rect 419058 596288 419678 597952
rect 422778 599340 423398 599436
rect 422778 599284 422874 599340
rect 422930 599284 422998 599340
rect 423054 599284 423122 599340
rect 423178 599284 423246 599340
rect 423302 599284 423398 599340
rect 422778 599216 423398 599284
rect 422778 599160 422874 599216
rect 422930 599160 422998 599216
rect 423054 599160 423122 599216
rect 423178 599160 423246 599216
rect 423302 599160 423398 599216
rect 422778 599092 423398 599160
rect 422778 599036 422874 599092
rect 422930 599036 422998 599092
rect 423054 599036 423122 599092
rect 423178 599036 423246 599092
rect 423302 599036 423398 599092
rect 422778 598968 423398 599036
rect 422778 598912 422874 598968
rect 422930 598912 422998 598968
rect 423054 598912 423122 598968
rect 423178 598912 423246 598968
rect 423302 598912 423398 598968
rect 422778 596288 423398 598912
rect 437058 598380 437678 599436
rect 437058 598324 437154 598380
rect 437210 598324 437278 598380
rect 437334 598324 437402 598380
rect 437458 598324 437526 598380
rect 437582 598324 437678 598380
rect 437058 598256 437678 598324
rect 437058 598200 437154 598256
rect 437210 598200 437278 598256
rect 437334 598200 437402 598256
rect 437458 598200 437526 598256
rect 437582 598200 437678 598256
rect 437058 598132 437678 598200
rect 437058 598076 437154 598132
rect 437210 598076 437278 598132
rect 437334 598076 437402 598132
rect 437458 598076 437526 598132
rect 437582 598076 437678 598132
rect 437058 598008 437678 598076
rect 437058 597952 437154 598008
rect 437210 597952 437278 598008
rect 437334 597952 437402 598008
rect 437458 597952 437526 598008
rect 437582 597952 437678 598008
rect 437058 596288 437678 597952
rect 440778 599340 441398 599436
rect 440778 599284 440874 599340
rect 440930 599284 440998 599340
rect 441054 599284 441122 599340
rect 441178 599284 441246 599340
rect 441302 599284 441398 599340
rect 440778 599216 441398 599284
rect 440778 599160 440874 599216
rect 440930 599160 440998 599216
rect 441054 599160 441122 599216
rect 441178 599160 441246 599216
rect 441302 599160 441398 599216
rect 440778 599092 441398 599160
rect 440778 599036 440874 599092
rect 440930 599036 440998 599092
rect 441054 599036 441122 599092
rect 441178 599036 441246 599092
rect 441302 599036 441398 599092
rect 440778 598968 441398 599036
rect 440778 598912 440874 598968
rect 440930 598912 440998 598968
rect 441054 598912 441122 598968
rect 441178 598912 441246 598968
rect 441302 598912 441398 598968
rect 440778 596288 441398 598912
rect 455058 598380 455678 599436
rect 455058 598324 455154 598380
rect 455210 598324 455278 598380
rect 455334 598324 455402 598380
rect 455458 598324 455526 598380
rect 455582 598324 455678 598380
rect 455058 598256 455678 598324
rect 455058 598200 455154 598256
rect 455210 598200 455278 598256
rect 455334 598200 455402 598256
rect 455458 598200 455526 598256
rect 455582 598200 455678 598256
rect 455058 598132 455678 598200
rect 455058 598076 455154 598132
rect 455210 598076 455278 598132
rect 455334 598076 455402 598132
rect 455458 598076 455526 598132
rect 455582 598076 455678 598132
rect 455058 598008 455678 598076
rect 455058 597952 455154 598008
rect 455210 597952 455278 598008
rect 455334 597952 455402 598008
rect 455458 597952 455526 598008
rect 455582 597952 455678 598008
rect 455058 596288 455678 597952
rect 458778 599340 459398 599436
rect 458778 599284 458874 599340
rect 458930 599284 458998 599340
rect 459054 599284 459122 599340
rect 459178 599284 459246 599340
rect 459302 599284 459398 599340
rect 458778 599216 459398 599284
rect 458778 599160 458874 599216
rect 458930 599160 458998 599216
rect 459054 599160 459122 599216
rect 459178 599160 459246 599216
rect 459302 599160 459398 599216
rect 458778 599092 459398 599160
rect 458778 599036 458874 599092
rect 458930 599036 458998 599092
rect 459054 599036 459122 599092
rect 459178 599036 459246 599092
rect 459302 599036 459398 599092
rect 458778 598968 459398 599036
rect 458778 598912 458874 598968
rect 458930 598912 458998 598968
rect 459054 598912 459122 598968
rect 459178 598912 459246 598968
rect 459302 598912 459398 598968
rect 458778 596288 459398 598912
rect 473058 598380 473678 599436
rect 473058 598324 473154 598380
rect 473210 598324 473278 598380
rect 473334 598324 473402 598380
rect 473458 598324 473526 598380
rect 473582 598324 473678 598380
rect 473058 598256 473678 598324
rect 473058 598200 473154 598256
rect 473210 598200 473278 598256
rect 473334 598200 473402 598256
rect 473458 598200 473526 598256
rect 473582 598200 473678 598256
rect 473058 598132 473678 598200
rect 473058 598076 473154 598132
rect 473210 598076 473278 598132
rect 473334 598076 473402 598132
rect 473458 598076 473526 598132
rect 473582 598076 473678 598132
rect 473058 598008 473678 598076
rect 473058 597952 473154 598008
rect 473210 597952 473278 598008
rect 473334 597952 473402 598008
rect 473458 597952 473526 598008
rect 473582 597952 473678 598008
rect 473058 596288 473678 597952
rect 476778 599340 477398 599436
rect 476778 599284 476874 599340
rect 476930 599284 476998 599340
rect 477054 599284 477122 599340
rect 477178 599284 477246 599340
rect 477302 599284 477398 599340
rect 476778 599216 477398 599284
rect 476778 599160 476874 599216
rect 476930 599160 476998 599216
rect 477054 599160 477122 599216
rect 477178 599160 477246 599216
rect 477302 599160 477398 599216
rect 476778 599092 477398 599160
rect 476778 599036 476874 599092
rect 476930 599036 476998 599092
rect 477054 599036 477122 599092
rect 477178 599036 477246 599092
rect 477302 599036 477398 599092
rect 476778 598968 477398 599036
rect 476778 598912 476874 598968
rect 476930 598912 476998 598968
rect 477054 598912 477122 598968
rect 477178 598912 477246 598968
rect 477302 598912 477398 598968
rect 476778 596288 477398 598912
rect 491058 598380 491678 599436
rect 491058 598324 491154 598380
rect 491210 598324 491278 598380
rect 491334 598324 491402 598380
rect 491458 598324 491526 598380
rect 491582 598324 491678 598380
rect 491058 598256 491678 598324
rect 491058 598200 491154 598256
rect 491210 598200 491278 598256
rect 491334 598200 491402 598256
rect 491458 598200 491526 598256
rect 491582 598200 491678 598256
rect 491058 598132 491678 598200
rect 491058 598076 491154 598132
rect 491210 598076 491278 598132
rect 491334 598076 491402 598132
rect 491458 598076 491526 598132
rect 491582 598076 491678 598132
rect 491058 598008 491678 598076
rect 491058 597952 491154 598008
rect 491210 597952 491278 598008
rect 491334 597952 491402 598008
rect 491458 597952 491526 598008
rect 491582 597952 491678 598008
rect 491058 596288 491678 597952
rect 494778 599340 495398 599436
rect 494778 599284 494874 599340
rect 494930 599284 494998 599340
rect 495054 599284 495122 599340
rect 495178 599284 495246 599340
rect 495302 599284 495398 599340
rect 494778 599216 495398 599284
rect 494778 599160 494874 599216
rect 494930 599160 494998 599216
rect 495054 599160 495122 599216
rect 495178 599160 495246 599216
rect 495302 599160 495398 599216
rect 494778 599092 495398 599160
rect 494778 599036 494874 599092
rect 494930 599036 494998 599092
rect 495054 599036 495122 599092
rect 495178 599036 495246 599092
rect 495302 599036 495398 599092
rect 494778 598968 495398 599036
rect 494778 598912 494874 598968
rect 494930 598912 494998 598968
rect 495054 598912 495122 598968
rect 495178 598912 495246 598968
rect 495302 598912 495398 598968
rect 494778 596288 495398 598912
rect 509058 598380 509678 599436
rect 509058 598324 509154 598380
rect 509210 598324 509278 598380
rect 509334 598324 509402 598380
rect 509458 598324 509526 598380
rect 509582 598324 509678 598380
rect 509058 598256 509678 598324
rect 509058 598200 509154 598256
rect 509210 598200 509278 598256
rect 509334 598200 509402 598256
rect 509458 598200 509526 598256
rect 509582 598200 509678 598256
rect 509058 598132 509678 598200
rect 509058 598076 509154 598132
rect 509210 598076 509278 598132
rect 509334 598076 509402 598132
rect 509458 598076 509526 598132
rect 509582 598076 509678 598132
rect 509058 598008 509678 598076
rect 509058 597952 509154 598008
rect 509210 597952 509278 598008
rect 509334 597952 509402 598008
rect 509458 597952 509526 598008
rect 509582 597952 509678 598008
rect 509058 596288 509678 597952
rect 512778 599340 513398 599436
rect 512778 599284 512874 599340
rect 512930 599284 512998 599340
rect 513054 599284 513122 599340
rect 513178 599284 513246 599340
rect 513302 599284 513398 599340
rect 512778 599216 513398 599284
rect 512778 599160 512874 599216
rect 512930 599160 512998 599216
rect 513054 599160 513122 599216
rect 513178 599160 513246 599216
rect 513302 599160 513398 599216
rect 512778 599092 513398 599160
rect 512778 599036 512874 599092
rect 512930 599036 512998 599092
rect 513054 599036 513122 599092
rect 513178 599036 513246 599092
rect 513302 599036 513398 599092
rect 512778 598968 513398 599036
rect 512778 598912 512874 598968
rect 512930 598912 512998 598968
rect 513054 598912 513122 598968
rect 513178 598912 513246 598968
rect 513302 598912 513398 598968
rect 512778 596288 513398 598912
rect 527058 598380 527678 599436
rect 527058 598324 527154 598380
rect 527210 598324 527278 598380
rect 527334 598324 527402 598380
rect 527458 598324 527526 598380
rect 527582 598324 527678 598380
rect 527058 598256 527678 598324
rect 527058 598200 527154 598256
rect 527210 598200 527278 598256
rect 527334 598200 527402 598256
rect 527458 598200 527526 598256
rect 527582 598200 527678 598256
rect 527058 598132 527678 598200
rect 527058 598076 527154 598132
rect 527210 598076 527278 598132
rect 527334 598076 527402 598132
rect 527458 598076 527526 598132
rect 527582 598076 527678 598132
rect 527058 598008 527678 598076
rect 527058 597952 527154 598008
rect 527210 597952 527278 598008
rect 527334 597952 527402 598008
rect 527458 597952 527526 598008
rect 527582 597952 527678 598008
rect 527058 596288 527678 597952
rect 530778 599340 531398 599436
rect 530778 599284 530874 599340
rect 530930 599284 530998 599340
rect 531054 599284 531122 599340
rect 531178 599284 531246 599340
rect 531302 599284 531398 599340
rect 530778 599216 531398 599284
rect 530778 599160 530874 599216
rect 530930 599160 530998 599216
rect 531054 599160 531122 599216
rect 531178 599160 531246 599216
rect 531302 599160 531398 599216
rect 530778 599092 531398 599160
rect 530778 599036 530874 599092
rect 530930 599036 530998 599092
rect 531054 599036 531122 599092
rect 531178 599036 531246 599092
rect 531302 599036 531398 599092
rect 530778 598968 531398 599036
rect 530778 598912 530874 598968
rect 530930 598912 530998 598968
rect 531054 598912 531122 598968
rect 531178 598912 531246 598968
rect 531302 598912 531398 598968
rect 530778 596288 531398 598912
rect 545058 598380 545678 599436
rect 545058 598324 545154 598380
rect 545210 598324 545278 598380
rect 545334 598324 545402 598380
rect 545458 598324 545526 598380
rect 545582 598324 545678 598380
rect 545058 598256 545678 598324
rect 545058 598200 545154 598256
rect 545210 598200 545278 598256
rect 545334 598200 545402 598256
rect 545458 598200 545526 598256
rect 545582 598200 545678 598256
rect 545058 598132 545678 598200
rect 545058 598076 545154 598132
rect 545210 598076 545278 598132
rect 545334 598076 545402 598132
rect 545458 598076 545526 598132
rect 545582 598076 545678 598132
rect 545058 598008 545678 598076
rect 545058 597952 545154 598008
rect 545210 597952 545278 598008
rect 545334 597952 545402 598008
rect 545458 597952 545526 598008
rect 545582 597952 545678 598008
rect 545058 596288 545678 597952
rect 548778 599340 549398 599436
rect 548778 599284 548874 599340
rect 548930 599284 548998 599340
rect 549054 599284 549122 599340
rect 549178 599284 549246 599340
rect 549302 599284 549398 599340
rect 548778 599216 549398 599284
rect 548778 599160 548874 599216
rect 548930 599160 548998 599216
rect 549054 599160 549122 599216
rect 549178 599160 549246 599216
rect 549302 599160 549398 599216
rect 548778 599092 549398 599160
rect 548778 599036 548874 599092
rect 548930 599036 548998 599092
rect 549054 599036 549122 599092
rect 549178 599036 549246 599092
rect 549302 599036 549398 599092
rect 548778 598968 549398 599036
rect 548778 598912 548874 598968
rect 548930 598912 548998 598968
rect 549054 598912 549122 598968
rect 549178 598912 549246 598968
rect 549302 598912 549398 598968
rect 548778 596288 549398 598912
rect 563058 598380 563678 599436
rect 563058 598324 563154 598380
rect 563210 598324 563278 598380
rect 563334 598324 563402 598380
rect 563458 598324 563526 598380
rect 563582 598324 563678 598380
rect 563058 598256 563678 598324
rect 563058 598200 563154 598256
rect 563210 598200 563278 598256
rect 563334 598200 563402 598256
rect 563458 598200 563526 598256
rect 563582 598200 563678 598256
rect 563058 598132 563678 598200
rect 563058 598076 563154 598132
rect 563210 598076 563278 598132
rect 563334 598076 563402 598132
rect 563458 598076 563526 598132
rect 563582 598076 563678 598132
rect 563058 598008 563678 598076
rect 563058 597952 563154 598008
rect 563210 597952 563278 598008
rect 563334 597952 563402 598008
rect 563458 597952 563526 598008
rect 563582 597952 563678 598008
rect 563058 596288 563678 597952
rect 566778 599340 567398 599436
rect 566778 599284 566874 599340
rect 566930 599284 566998 599340
rect 567054 599284 567122 599340
rect 567178 599284 567246 599340
rect 567302 599284 567398 599340
rect 566778 599216 567398 599284
rect 566778 599160 566874 599216
rect 566930 599160 566998 599216
rect 567054 599160 567122 599216
rect 567178 599160 567246 599216
rect 567302 599160 567398 599216
rect 566778 599092 567398 599160
rect 566778 599036 566874 599092
rect 566930 599036 566998 599092
rect 567054 599036 567122 599092
rect 567178 599036 567246 599092
rect 567302 599036 567398 599092
rect 566778 598968 567398 599036
rect 566778 598912 566874 598968
rect 566930 598912 566998 598968
rect 567054 598912 567122 598968
rect 567178 598912 567246 598968
rect 567302 598912 567398 598968
rect 566778 596288 567398 598912
rect 581058 598380 581678 599436
rect 581058 598324 581154 598380
rect 581210 598324 581278 598380
rect 581334 598324 581402 598380
rect 581458 598324 581526 598380
rect 581582 598324 581678 598380
rect 581058 598256 581678 598324
rect 581058 598200 581154 598256
rect 581210 598200 581278 598256
rect 581334 598200 581402 598256
rect 581458 598200 581526 598256
rect 581582 598200 581678 598256
rect 581058 598132 581678 598200
rect 581058 598076 581154 598132
rect 581210 598076 581278 598132
rect 581334 598076 581402 598132
rect 581458 598076 581526 598132
rect 581582 598076 581678 598132
rect 581058 598008 581678 598076
rect 581058 597952 581154 598008
rect 581210 597952 581278 598008
rect 581334 597952 581402 598008
rect 581458 597952 581526 598008
rect 581582 597952 581678 598008
rect 581058 596288 581678 597952
rect 584778 599340 585398 599436
rect 584778 599284 584874 599340
rect 584930 599284 584998 599340
rect 585054 599284 585122 599340
rect 585178 599284 585246 599340
rect 585302 599284 585398 599340
rect 584778 599216 585398 599284
rect 584778 599160 584874 599216
rect 584930 599160 584998 599216
rect 585054 599160 585122 599216
rect 585178 599160 585246 599216
rect 585302 599160 585398 599216
rect 584778 599092 585398 599160
rect 584778 599036 584874 599092
rect 584930 599036 584998 599092
rect 585054 599036 585122 599092
rect 585178 599036 585246 599092
rect 585302 599036 585398 599092
rect 584778 598968 585398 599036
rect 584778 598912 584874 598968
rect 584930 598912 584998 598968
rect 585054 598912 585122 598968
rect 585178 598912 585246 598968
rect 585302 598912 585398 598968
rect 584778 596288 585398 598912
rect 599376 599340 599996 599436
rect 599376 599284 599472 599340
rect 599528 599284 599596 599340
rect 599652 599284 599720 599340
rect 599776 599284 599844 599340
rect 599900 599284 599996 599340
rect 599376 599216 599996 599284
rect 599376 599160 599472 599216
rect 599528 599160 599596 599216
rect 599652 599160 599720 599216
rect 599776 599160 599844 599216
rect 599900 599160 599996 599216
rect 599376 599092 599996 599160
rect 599376 599036 599472 599092
rect 599528 599036 599596 599092
rect 599652 599036 599720 599092
rect 599776 599036 599844 599092
rect 599900 599036 599996 599092
rect 599376 598968 599996 599036
rect 599376 598912 599472 598968
rect 599528 598912 599596 598968
rect 599652 598912 599720 598968
rect 599776 598912 599844 598968
rect 599900 598912 599996 598968
rect 598416 598380 599036 598476
rect 598416 598324 598512 598380
rect 598568 598324 598636 598380
rect 598692 598324 598760 598380
rect 598816 598324 598884 598380
rect 598940 598324 599036 598380
rect 598416 598256 599036 598324
rect 598416 598200 598512 598256
rect 598568 598200 598636 598256
rect 598692 598200 598760 598256
rect 598816 598200 598884 598256
rect 598940 598200 599036 598256
rect 598416 598132 599036 598200
rect 598416 598076 598512 598132
rect 598568 598076 598636 598132
rect 598692 598076 598760 598132
rect 598816 598076 598884 598132
rect 598940 598076 599036 598132
rect 598416 598008 599036 598076
rect 598416 597952 598512 598008
rect 598568 597952 598636 598008
rect 598692 597952 598760 598008
rect 598816 597952 598884 598008
rect 598940 597952 599036 598008
rect 5058 581862 5154 581918
rect 5210 581862 5278 581918
rect 5334 581862 5402 581918
rect 5458 581862 5526 581918
rect 5582 581862 5678 581918
rect 5058 581794 5678 581862
rect 5058 581738 5154 581794
rect 5210 581738 5278 581794
rect 5334 581738 5402 581794
rect 5458 581738 5526 581794
rect 5582 581738 5678 581794
rect 5058 581670 5678 581738
rect 5058 581614 5154 581670
rect 5210 581614 5278 581670
rect 5334 581614 5402 581670
rect 5458 581614 5526 581670
rect 5582 581614 5678 581670
rect 5058 581546 5678 581614
rect 5058 581490 5154 581546
rect 5210 581490 5278 581546
rect 5334 581490 5402 581546
rect 5458 581490 5526 581546
rect 5582 581490 5678 581546
rect 5058 563918 5678 581490
rect 5058 563862 5154 563918
rect 5210 563862 5278 563918
rect 5334 563862 5402 563918
rect 5458 563862 5526 563918
rect 5582 563862 5678 563918
rect 5058 563794 5678 563862
rect 5058 563738 5154 563794
rect 5210 563738 5278 563794
rect 5334 563738 5402 563794
rect 5458 563738 5526 563794
rect 5582 563738 5678 563794
rect 5058 563670 5678 563738
rect 5058 563614 5154 563670
rect 5210 563614 5278 563670
rect 5334 563614 5402 563670
rect 5458 563614 5526 563670
rect 5582 563614 5678 563670
rect 5058 563546 5678 563614
rect 5058 563490 5154 563546
rect 5210 563490 5278 563546
rect 5334 563490 5402 563546
rect 5458 563490 5526 563546
rect 5582 563490 5678 563546
rect 5058 545918 5678 563490
rect 5058 545862 5154 545918
rect 5210 545862 5278 545918
rect 5334 545862 5402 545918
rect 5458 545862 5526 545918
rect 5582 545862 5678 545918
rect 5058 545794 5678 545862
rect 5058 545738 5154 545794
rect 5210 545738 5278 545794
rect 5334 545738 5402 545794
rect 5458 545738 5526 545794
rect 5582 545738 5678 545794
rect 5058 545670 5678 545738
rect 5058 545614 5154 545670
rect 5210 545614 5278 545670
rect 5334 545614 5402 545670
rect 5458 545614 5526 545670
rect 5582 545614 5678 545670
rect 5058 545546 5678 545614
rect 5058 545490 5154 545546
rect 5210 545490 5278 545546
rect 5334 545490 5402 545546
rect 5458 545490 5526 545546
rect 5582 545490 5678 545546
rect 5058 527918 5678 545490
rect 5058 527862 5154 527918
rect 5210 527862 5278 527918
rect 5334 527862 5402 527918
rect 5458 527862 5526 527918
rect 5582 527862 5678 527918
rect 5058 527794 5678 527862
rect 5058 527738 5154 527794
rect 5210 527738 5278 527794
rect 5334 527738 5402 527794
rect 5458 527738 5526 527794
rect 5582 527738 5678 527794
rect 5058 527670 5678 527738
rect 5058 527614 5154 527670
rect 5210 527614 5278 527670
rect 5334 527614 5402 527670
rect 5458 527614 5526 527670
rect 5582 527614 5678 527670
rect 5058 527546 5678 527614
rect 5058 527490 5154 527546
rect 5210 527490 5278 527546
rect 5334 527490 5402 527546
rect 5458 527490 5526 527546
rect 5582 527490 5678 527546
rect 5058 509918 5678 527490
rect 5058 509862 5154 509918
rect 5210 509862 5278 509918
rect 5334 509862 5402 509918
rect 5458 509862 5526 509918
rect 5582 509862 5678 509918
rect 5058 509794 5678 509862
rect 5058 509738 5154 509794
rect 5210 509738 5278 509794
rect 5334 509738 5402 509794
rect 5458 509738 5526 509794
rect 5582 509738 5678 509794
rect 5058 509670 5678 509738
rect 5058 509614 5154 509670
rect 5210 509614 5278 509670
rect 5334 509614 5402 509670
rect 5458 509614 5526 509670
rect 5582 509614 5678 509670
rect 5058 509546 5678 509614
rect 5058 509490 5154 509546
rect 5210 509490 5278 509546
rect 5334 509490 5402 509546
rect 5458 509490 5526 509546
rect 5582 509490 5678 509546
rect 5058 491918 5678 509490
rect 5058 491862 5154 491918
rect 5210 491862 5278 491918
rect 5334 491862 5402 491918
rect 5458 491862 5526 491918
rect 5582 491862 5678 491918
rect 5058 491794 5678 491862
rect 5058 491738 5154 491794
rect 5210 491738 5278 491794
rect 5334 491738 5402 491794
rect 5458 491738 5526 491794
rect 5582 491738 5678 491794
rect 5058 491670 5678 491738
rect 5058 491614 5154 491670
rect 5210 491614 5278 491670
rect 5334 491614 5402 491670
rect 5458 491614 5526 491670
rect 5582 491614 5678 491670
rect 5058 491546 5678 491614
rect 5058 491490 5154 491546
rect 5210 491490 5278 491546
rect 5334 491490 5402 491546
rect 5458 491490 5526 491546
rect 5582 491490 5678 491546
rect 5058 473918 5678 491490
rect 5058 473862 5154 473918
rect 5210 473862 5278 473918
rect 5334 473862 5402 473918
rect 5458 473862 5526 473918
rect 5582 473862 5678 473918
rect 5058 473794 5678 473862
rect 5058 473738 5154 473794
rect 5210 473738 5278 473794
rect 5334 473738 5402 473794
rect 5458 473738 5526 473794
rect 5582 473738 5678 473794
rect 5058 473670 5678 473738
rect 5058 473614 5154 473670
rect 5210 473614 5278 473670
rect 5334 473614 5402 473670
rect 5458 473614 5526 473670
rect 5582 473614 5678 473670
rect 5058 473546 5678 473614
rect 5058 473490 5154 473546
rect 5210 473490 5278 473546
rect 5334 473490 5402 473546
rect 5458 473490 5526 473546
rect 5582 473490 5678 473546
rect 5058 455918 5678 473490
rect 5058 455862 5154 455918
rect 5210 455862 5278 455918
rect 5334 455862 5402 455918
rect 5458 455862 5526 455918
rect 5582 455862 5678 455918
rect 5058 455794 5678 455862
rect 5058 455738 5154 455794
rect 5210 455738 5278 455794
rect 5334 455738 5402 455794
rect 5458 455738 5526 455794
rect 5582 455738 5678 455794
rect 5058 455670 5678 455738
rect 5058 455614 5154 455670
rect 5210 455614 5278 455670
rect 5334 455614 5402 455670
rect 5458 455614 5526 455670
rect 5582 455614 5678 455670
rect 5058 455546 5678 455614
rect 5058 455490 5154 455546
rect 5210 455490 5278 455546
rect 5334 455490 5402 455546
rect 5458 455490 5526 455546
rect 5582 455490 5678 455546
rect 5058 437918 5678 455490
rect 5058 437862 5154 437918
rect 5210 437862 5278 437918
rect 5334 437862 5402 437918
rect 5458 437862 5526 437918
rect 5582 437862 5678 437918
rect 5058 437794 5678 437862
rect 5058 437738 5154 437794
rect 5210 437738 5278 437794
rect 5334 437738 5402 437794
rect 5458 437738 5526 437794
rect 5582 437738 5678 437794
rect 5058 437670 5678 437738
rect 5058 437614 5154 437670
rect 5210 437614 5278 437670
rect 5334 437614 5402 437670
rect 5458 437614 5526 437670
rect 5582 437614 5678 437670
rect 5058 437546 5678 437614
rect 5058 437490 5154 437546
rect 5210 437490 5278 437546
rect 5334 437490 5402 437546
rect 5458 437490 5526 437546
rect 5582 437490 5678 437546
rect 5058 419918 5678 437490
rect 5058 419862 5154 419918
rect 5210 419862 5278 419918
rect 5334 419862 5402 419918
rect 5458 419862 5526 419918
rect 5582 419862 5678 419918
rect 5058 419794 5678 419862
rect 5058 419738 5154 419794
rect 5210 419738 5278 419794
rect 5334 419738 5402 419794
rect 5458 419738 5526 419794
rect 5582 419738 5678 419794
rect 5058 419670 5678 419738
rect 5058 419614 5154 419670
rect 5210 419614 5278 419670
rect 5334 419614 5402 419670
rect 5458 419614 5526 419670
rect 5582 419614 5678 419670
rect 5058 419546 5678 419614
rect 5058 419490 5154 419546
rect 5210 419490 5278 419546
rect 5334 419490 5402 419546
rect 5458 419490 5526 419546
rect 5582 419490 5678 419546
rect 5058 401918 5678 419490
rect 5058 401862 5154 401918
rect 5210 401862 5278 401918
rect 5334 401862 5402 401918
rect 5458 401862 5526 401918
rect 5582 401862 5678 401918
rect 5058 401794 5678 401862
rect 5058 401738 5154 401794
rect 5210 401738 5278 401794
rect 5334 401738 5402 401794
rect 5458 401738 5526 401794
rect 5582 401738 5678 401794
rect 5058 401670 5678 401738
rect 5058 401614 5154 401670
rect 5210 401614 5278 401670
rect 5334 401614 5402 401670
rect 5458 401614 5526 401670
rect 5582 401614 5678 401670
rect 5058 401546 5678 401614
rect 5058 401490 5154 401546
rect 5210 401490 5278 401546
rect 5334 401490 5402 401546
rect 5458 401490 5526 401546
rect 5582 401490 5678 401546
rect 5058 383918 5678 401490
rect 5058 383862 5154 383918
rect 5210 383862 5278 383918
rect 5334 383862 5402 383918
rect 5458 383862 5526 383918
rect 5582 383862 5678 383918
rect 5058 383794 5678 383862
rect 5058 383738 5154 383794
rect 5210 383738 5278 383794
rect 5334 383738 5402 383794
rect 5458 383738 5526 383794
rect 5582 383738 5678 383794
rect 5058 383670 5678 383738
rect 5058 383614 5154 383670
rect 5210 383614 5278 383670
rect 5334 383614 5402 383670
rect 5458 383614 5526 383670
rect 5582 383614 5678 383670
rect 5058 383546 5678 383614
rect 5058 383490 5154 383546
rect 5210 383490 5278 383546
rect 5334 383490 5402 383546
rect 5458 383490 5526 383546
rect 5582 383490 5678 383546
rect 5058 365918 5678 383490
rect 5058 365862 5154 365918
rect 5210 365862 5278 365918
rect 5334 365862 5402 365918
rect 5458 365862 5526 365918
rect 5582 365862 5678 365918
rect 5058 365794 5678 365862
rect 5058 365738 5154 365794
rect 5210 365738 5278 365794
rect 5334 365738 5402 365794
rect 5458 365738 5526 365794
rect 5582 365738 5678 365794
rect 5058 365670 5678 365738
rect 5058 365614 5154 365670
rect 5210 365614 5278 365670
rect 5334 365614 5402 365670
rect 5458 365614 5526 365670
rect 5582 365614 5678 365670
rect 5058 365546 5678 365614
rect 5058 365490 5154 365546
rect 5210 365490 5278 365546
rect 5334 365490 5402 365546
rect 5458 365490 5526 365546
rect 5582 365490 5678 365546
rect 5058 347918 5678 365490
rect 5058 347862 5154 347918
rect 5210 347862 5278 347918
rect 5334 347862 5402 347918
rect 5458 347862 5526 347918
rect 5582 347862 5678 347918
rect 5058 347794 5678 347862
rect 5058 347738 5154 347794
rect 5210 347738 5278 347794
rect 5334 347738 5402 347794
rect 5458 347738 5526 347794
rect 5582 347738 5678 347794
rect 5058 347670 5678 347738
rect 5058 347614 5154 347670
rect 5210 347614 5278 347670
rect 5334 347614 5402 347670
rect 5458 347614 5526 347670
rect 5582 347614 5678 347670
rect 5058 347546 5678 347614
rect 5058 347490 5154 347546
rect 5210 347490 5278 347546
rect 5334 347490 5402 347546
rect 5458 347490 5526 347546
rect 5582 347490 5678 347546
rect 5058 329918 5678 347490
rect 5058 329862 5154 329918
rect 5210 329862 5278 329918
rect 5334 329862 5402 329918
rect 5458 329862 5526 329918
rect 5582 329862 5678 329918
rect 5058 329794 5678 329862
rect 5058 329738 5154 329794
rect 5210 329738 5278 329794
rect 5334 329738 5402 329794
rect 5458 329738 5526 329794
rect 5582 329738 5678 329794
rect 5058 329670 5678 329738
rect 5058 329614 5154 329670
rect 5210 329614 5278 329670
rect 5334 329614 5402 329670
rect 5458 329614 5526 329670
rect 5582 329614 5678 329670
rect 5058 329546 5678 329614
rect 5058 329490 5154 329546
rect 5210 329490 5278 329546
rect 5334 329490 5402 329546
rect 5458 329490 5526 329546
rect 5582 329490 5678 329546
rect 5058 311918 5678 329490
rect 5058 311862 5154 311918
rect 5210 311862 5278 311918
rect 5334 311862 5402 311918
rect 5458 311862 5526 311918
rect 5582 311862 5678 311918
rect 5058 311794 5678 311862
rect 5058 311738 5154 311794
rect 5210 311738 5278 311794
rect 5334 311738 5402 311794
rect 5458 311738 5526 311794
rect 5582 311738 5678 311794
rect 5058 311670 5678 311738
rect 5058 311614 5154 311670
rect 5210 311614 5278 311670
rect 5334 311614 5402 311670
rect 5458 311614 5526 311670
rect 5582 311614 5678 311670
rect 5058 311546 5678 311614
rect 5058 311490 5154 311546
rect 5210 311490 5278 311546
rect 5334 311490 5402 311546
rect 5458 311490 5526 311546
rect 5582 311490 5678 311546
rect 5058 293918 5678 311490
rect 5058 293862 5154 293918
rect 5210 293862 5278 293918
rect 5334 293862 5402 293918
rect 5458 293862 5526 293918
rect 5582 293862 5678 293918
rect 5058 293794 5678 293862
rect 5058 293738 5154 293794
rect 5210 293738 5278 293794
rect 5334 293738 5402 293794
rect 5458 293738 5526 293794
rect 5582 293738 5678 293794
rect 5058 293670 5678 293738
rect 5058 293614 5154 293670
rect 5210 293614 5278 293670
rect 5334 293614 5402 293670
rect 5458 293614 5526 293670
rect 5582 293614 5678 293670
rect 5058 293546 5678 293614
rect 5058 293490 5154 293546
rect 5210 293490 5278 293546
rect 5334 293490 5402 293546
rect 5458 293490 5526 293546
rect 5582 293490 5678 293546
rect 5058 275918 5678 293490
rect 5058 275862 5154 275918
rect 5210 275862 5278 275918
rect 5334 275862 5402 275918
rect 5458 275862 5526 275918
rect 5582 275862 5678 275918
rect 5058 275794 5678 275862
rect 5058 275738 5154 275794
rect 5210 275738 5278 275794
rect 5334 275738 5402 275794
rect 5458 275738 5526 275794
rect 5582 275738 5678 275794
rect 5058 275670 5678 275738
rect 5058 275614 5154 275670
rect 5210 275614 5278 275670
rect 5334 275614 5402 275670
rect 5458 275614 5526 275670
rect 5582 275614 5678 275670
rect 5058 275546 5678 275614
rect 5058 275490 5154 275546
rect 5210 275490 5278 275546
rect 5334 275490 5402 275546
rect 5458 275490 5526 275546
rect 5582 275490 5678 275546
rect 5058 257918 5678 275490
rect 5058 257862 5154 257918
rect 5210 257862 5278 257918
rect 5334 257862 5402 257918
rect 5458 257862 5526 257918
rect 5582 257862 5678 257918
rect 5058 257794 5678 257862
rect 5058 257738 5154 257794
rect 5210 257738 5278 257794
rect 5334 257738 5402 257794
rect 5458 257738 5526 257794
rect 5582 257738 5678 257794
rect 5058 257670 5678 257738
rect 5058 257614 5154 257670
rect 5210 257614 5278 257670
rect 5334 257614 5402 257670
rect 5458 257614 5526 257670
rect 5582 257614 5678 257670
rect 5058 257546 5678 257614
rect 5058 257490 5154 257546
rect 5210 257490 5278 257546
rect 5334 257490 5402 257546
rect 5458 257490 5526 257546
rect 5582 257490 5678 257546
rect 5058 239918 5678 257490
rect 5058 239862 5154 239918
rect 5210 239862 5278 239918
rect 5334 239862 5402 239918
rect 5458 239862 5526 239918
rect 5582 239862 5678 239918
rect 5058 239794 5678 239862
rect 5058 239738 5154 239794
rect 5210 239738 5278 239794
rect 5334 239738 5402 239794
rect 5458 239738 5526 239794
rect 5582 239738 5678 239794
rect 5058 239670 5678 239738
rect 5058 239614 5154 239670
rect 5210 239614 5278 239670
rect 5334 239614 5402 239670
rect 5458 239614 5526 239670
rect 5582 239614 5678 239670
rect 5058 239546 5678 239614
rect 5058 239490 5154 239546
rect 5210 239490 5278 239546
rect 5334 239490 5402 239546
rect 5458 239490 5526 239546
rect 5582 239490 5678 239546
rect 5058 221918 5678 239490
rect 5058 221862 5154 221918
rect 5210 221862 5278 221918
rect 5334 221862 5402 221918
rect 5458 221862 5526 221918
rect 5582 221862 5678 221918
rect 5058 221794 5678 221862
rect 5058 221738 5154 221794
rect 5210 221738 5278 221794
rect 5334 221738 5402 221794
rect 5458 221738 5526 221794
rect 5582 221738 5678 221794
rect 5058 221670 5678 221738
rect 5058 221614 5154 221670
rect 5210 221614 5278 221670
rect 5334 221614 5402 221670
rect 5458 221614 5526 221670
rect 5582 221614 5678 221670
rect 5058 221546 5678 221614
rect 5058 221490 5154 221546
rect 5210 221490 5278 221546
rect 5334 221490 5402 221546
rect 5458 221490 5526 221546
rect 5582 221490 5678 221546
rect 5058 203918 5678 221490
rect 5058 203862 5154 203918
rect 5210 203862 5278 203918
rect 5334 203862 5402 203918
rect 5458 203862 5526 203918
rect 5582 203862 5678 203918
rect 5058 203794 5678 203862
rect 5058 203738 5154 203794
rect 5210 203738 5278 203794
rect 5334 203738 5402 203794
rect 5458 203738 5526 203794
rect 5582 203738 5678 203794
rect 5058 203670 5678 203738
rect 5058 203614 5154 203670
rect 5210 203614 5278 203670
rect 5334 203614 5402 203670
rect 5458 203614 5526 203670
rect 5582 203614 5678 203670
rect 5058 203546 5678 203614
rect 5058 203490 5154 203546
rect 5210 203490 5278 203546
rect 5334 203490 5402 203546
rect 5458 203490 5526 203546
rect 5582 203490 5678 203546
rect 5058 185918 5678 203490
rect 5058 185862 5154 185918
rect 5210 185862 5278 185918
rect 5334 185862 5402 185918
rect 5458 185862 5526 185918
rect 5582 185862 5678 185918
rect 5058 185794 5678 185862
rect 5058 185738 5154 185794
rect 5210 185738 5278 185794
rect 5334 185738 5402 185794
rect 5458 185738 5526 185794
rect 5582 185738 5678 185794
rect 5058 185670 5678 185738
rect 5058 185614 5154 185670
rect 5210 185614 5278 185670
rect 5334 185614 5402 185670
rect 5458 185614 5526 185670
rect 5582 185614 5678 185670
rect 5058 185546 5678 185614
rect 5058 185490 5154 185546
rect 5210 185490 5278 185546
rect 5334 185490 5402 185546
rect 5458 185490 5526 185546
rect 5582 185490 5678 185546
rect 5058 167918 5678 185490
rect 5058 167862 5154 167918
rect 5210 167862 5278 167918
rect 5334 167862 5402 167918
rect 5458 167862 5526 167918
rect 5582 167862 5678 167918
rect 5058 167794 5678 167862
rect 5058 167738 5154 167794
rect 5210 167738 5278 167794
rect 5334 167738 5402 167794
rect 5458 167738 5526 167794
rect 5582 167738 5678 167794
rect 5058 167670 5678 167738
rect 5058 167614 5154 167670
rect 5210 167614 5278 167670
rect 5334 167614 5402 167670
rect 5458 167614 5526 167670
rect 5582 167614 5678 167670
rect 5058 167546 5678 167614
rect 5058 167490 5154 167546
rect 5210 167490 5278 167546
rect 5334 167490 5402 167546
rect 5458 167490 5526 167546
rect 5582 167490 5678 167546
rect 5058 149918 5678 167490
rect 5058 149862 5154 149918
rect 5210 149862 5278 149918
rect 5334 149862 5402 149918
rect 5458 149862 5526 149918
rect 5582 149862 5678 149918
rect 5058 149794 5678 149862
rect 5058 149738 5154 149794
rect 5210 149738 5278 149794
rect 5334 149738 5402 149794
rect 5458 149738 5526 149794
rect 5582 149738 5678 149794
rect 5058 149670 5678 149738
rect 5058 149614 5154 149670
rect 5210 149614 5278 149670
rect 5334 149614 5402 149670
rect 5458 149614 5526 149670
rect 5582 149614 5678 149670
rect 5058 149546 5678 149614
rect 5058 149490 5154 149546
rect 5210 149490 5278 149546
rect 5334 149490 5402 149546
rect 5458 149490 5526 149546
rect 5582 149490 5678 149546
rect 5058 131918 5678 149490
rect 5058 131862 5154 131918
rect 5210 131862 5278 131918
rect 5334 131862 5402 131918
rect 5458 131862 5526 131918
rect 5582 131862 5678 131918
rect 5058 131794 5678 131862
rect 5058 131738 5154 131794
rect 5210 131738 5278 131794
rect 5334 131738 5402 131794
rect 5458 131738 5526 131794
rect 5582 131738 5678 131794
rect 5058 131670 5678 131738
rect 5058 131614 5154 131670
rect 5210 131614 5278 131670
rect 5334 131614 5402 131670
rect 5458 131614 5526 131670
rect 5582 131614 5678 131670
rect 5058 131546 5678 131614
rect 5058 131490 5154 131546
rect 5210 131490 5278 131546
rect 5334 131490 5402 131546
rect 5458 131490 5526 131546
rect 5582 131490 5678 131546
rect 5058 113918 5678 131490
rect 5058 113862 5154 113918
rect 5210 113862 5278 113918
rect 5334 113862 5402 113918
rect 5458 113862 5526 113918
rect 5582 113862 5678 113918
rect 5058 113794 5678 113862
rect 5058 113738 5154 113794
rect 5210 113738 5278 113794
rect 5334 113738 5402 113794
rect 5458 113738 5526 113794
rect 5582 113738 5678 113794
rect 5058 113670 5678 113738
rect 5058 113614 5154 113670
rect 5210 113614 5278 113670
rect 5334 113614 5402 113670
rect 5458 113614 5526 113670
rect 5582 113614 5678 113670
rect 5058 113546 5678 113614
rect 5058 113490 5154 113546
rect 5210 113490 5278 113546
rect 5334 113490 5402 113546
rect 5458 113490 5526 113546
rect 5582 113490 5678 113546
rect 5058 95918 5678 113490
rect 5058 95862 5154 95918
rect 5210 95862 5278 95918
rect 5334 95862 5402 95918
rect 5458 95862 5526 95918
rect 5582 95862 5678 95918
rect 5058 95794 5678 95862
rect 5058 95738 5154 95794
rect 5210 95738 5278 95794
rect 5334 95738 5402 95794
rect 5458 95738 5526 95794
rect 5582 95738 5678 95794
rect 5058 95670 5678 95738
rect 5058 95614 5154 95670
rect 5210 95614 5278 95670
rect 5334 95614 5402 95670
rect 5458 95614 5526 95670
rect 5582 95614 5678 95670
rect 5058 95546 5678 95614
rect 5058 95490 5154 95546
rect 5210 95490 5278 95546
rect 5334 95490 5402 95546
rect 5458 95490 5526 95546
rect 5582 95490 5678 95546
rect 5058 77918 5678 95490
rect 5058 77862 5154 77918
rect 5210 77862 5278 77918
rect 5334 77862 5402 77918
rect 5458 77862 5526 77918
rect 5582 77862 5678 77918
rect 5058 77794 5678 77862
rect 5058 77738 5154 77794
rect 5210 77738 5278 77794
rect 5334 77738 5402 77794
rect 5458 77738 5526 77794
rect 5582 77738 5678 77794
rect 5058 77670 5678 77738
rect 5058 77614 5154 77670
rect 5210 77614 5278 77670
rect 5334 77614 5402 77670
rect 5458 77614 5526 77670
rect 5582 77614 5678 77670
rect 5058 77546 5678 77614
rect 5058 77490 5154 77546
rect 5210 77490 5278 77546
rect 5334 77490 5402 77546
rect 5458 77490 5526 77546
rect 5582 77490 5678 77546
rect 5058 59918 5678 77490
rect 5058 59862 5154 59918
rect 5210 59862 5278 59918
rect 5334 59862 5402 59918
rect 5458 59862 5526 59918
rect 5582 59862 5678 59918
rect 5058 59794 5678 59862
rect 5058 59738 5154 59794
rect 5210 59738 5278 59794
rect 5334 59738 5402 59794
rect 5458 59738 5526 59794
rect 5582 59738 5678 59794
rect 5058 59670 5678 59738
rect 5058 59614 5154 59670
rect 5210 59614 5278 59670
rect 5334 59614 5402 59670
rect 5458 59614 5526 59670
rect 5582 59614 5678 59670
rect 5058 59546 5678 59614
rect 5058 59490 5154 59546
rect 5210 59490 5278 59546
rect 5334 59490 5402 59546
rect 5458 59490 5526 59546
rect 5582 59490 5678 59546
rect 5058 41918 5678 59490
rect 5058 41862 5154 41918
rect 5210 41862 5278 41918
rect 5334 41862 5402 41918
rect 5458 41862 5526 41918
rect 5582 41862 5678 41918
rect 5058 41794 5678 41862
rect 5058 41738 5154 41794
rect 5210 41738 5278 41794
rect 5334 41738 5402 41794
rect 5458 41738 5526 41794
rect 5582 41738 5678 41794
rect 5058 41670 5678 41738
rect 5058 41614 5154 41670
rect 5210 41614 5278 41670
rect 5334 41614 5402 41670
rect 5458 41614 5526 41670
rect 5582 41614 5678 41670
rect 5058 41546 5678 41614
rect 5058 41490 5154 41546
rect 5210 41490 5278 41546
rect 5334 41490 5402 41546
rect 5458 41490 5526 41546
rect 5582 41490 5678 41546
rect 5058 23918 5678 41490
rect 5058 23862 5154 23918
rect 5210 23862 5278 23918
rect 5334 23862 5402 23918
rect 5458 23862 5526 23918
rect 5582 23862 5678 23918
rect 5058 23794 5678 23862
rect 5058 23738 5154 23794
rect 5210 23738 5278 23794
rect 5334 23738 5402 23794
rect 5458 23738 5526 23794
rect 5582 23738 5678 23794
rect 5058 23670 5678 23738
rect 5058 23614 5154 23670
rect 5210 23614 5278 23670
rect 5334 23614 5402 23670
rect 5458 23614 5526 23670
rect 5582 23614 5678 23670
rect 5058 23546 5678 23614
rect 5058 23490 5154 23546
rect 5210 23490 5278 23546
rect 5334 23490 5402 23546
rect 5458 23490 5526 23546
rect 5582 23490 5678 23546
rect 5058 5918 5678 23490
rect 5058 5862 5154 5918
rect 5210 5862 5278 5918
rect 5334 5862 5402 5918
rect 5458 5862 5526 5918
rect 5582 5862 5678 5918
rect 5058 5794 5678 5862
rect 5058 5738 5154 5794
rect 5210 5738 5278 5794
rect 5334 5738 5402 5794
rect 5458 5738 5526 5794
rect 5582 5738 5678 5794
rect 5058 5670 5678 5738
rect 5058 5614 5154 5670
rect 5210 5614 5278 5670
rect 5334 5614 5402 5670
rect 5458 5614 5526 5670
rect 5582 5614 5678 5670
rect 5058 5546 5678 5614
rect 5058 5490 5154 5546
rect 5210 5490 5278 5546
rect 5334 5490 5402 5546
rect 5458 5490 5526 5546
rect 5582 5490 5678 5546
rect 5058 1808 5678 5490
rect 598416 581918 599036 597952
rect 598416 581862 598512 581918
rect 598568 581862 598636 581918
rect 598692 581862 598760 581918
rect 598816 581862 598884 581918
rect 598940 581862 599036 581918
rect 598416 581794 599036 581862
rect 598416 581738 598512 581794
rect 598568 581738 598636 581794
rect 598692 581738 598760 581794
rect 598816 581738 598884 581794
rect 598940 581738 599036 581794
rect 598416 581670 599036 581738
rect 598416 581614 598512 581670
rect 598568 581614 598636 581670
rect 598692 581614 598760 581670
rect 598816 581614 598884 581670
rect 598940 581614 599036 581670
rect 598416 581546 599036 581614
rect 598416 581490 598512 581546
rect 598568 581490 598636 581546
rect 598692 581490 598760 581546
rect 598816 581490 598884 581546
rect 598940 581490 599036 581546
rect 598416 563918 599036 581490
rect 598416 563862 598512 563918
rect 598568 563862 598636 563918
rect 598692 563862 598760 563918
rect 598816 563862 598884 563918
rect 598940 563862 599036 563918
rect 598416 563794 599036 563862
rect 598416 563738 598512 563794
rect 598568 563738 598636 563794
rect 598692 563738 598760 563794
rect 598816 563738 598884 563794
rect 598940 563738 599036 563794
rect 598416 563670 599036 563738
rect 598416 563614 598512 563670
rect 598568 563614 598636 563670
rect 598692 563614 598760 563670
rect 598816 563614 598884 563670
rect 598940 563614 599036 563670
rect 598416 563546 599036 563614
rect 598416 563490 598512 563546
rect 598568 563490 598636 563546
rect 598692 563490 598760 563546
rect 598816 563490 598884 563546
rect 598940 563490 599036 563546
rect 598416 545918 599036 563490
rect 598416 545862 598512 545918
rect 598568 545862 598636 545918
rect 598692 545862 598760 545918
rect 598816 545862 598884 545918
rect 598940 545862 599036 545918
rect 598416 545794 599036 545862
rect 598416 545738 598512 545794
rect 598568 545738 598636 545794
rect 598692 545738 598760 545794
rect 598816 545738 598884 545794
rect 598940 545738 599036 545794
rect 598416 545670 599036 545738
rect 598416 545614 598512 545670
rect 598568 545614 598636 545670
rect 598692 545614 598760 545670
rect 598816 545614 598884 545670
rect 598940 545614 599036 545670
rect 598416 545546 599036 545614
rect 598416 545490 598512 545546
rect 598568 545490 598636 545546
rect 598692 545490 598760 545546
rect 598816 545490 598884 545546
rect 598940 545490 599036 545546
rect 598416 527918 599036 545490
rect 598416 527862 598512 527918
rect 598568 527862 598636 527918
rect 598692 527862 598760 527918
rect 598816 527862 598884 527918
rect 598940 527862 599036 527918
rect 598416 527794 599036 527862
rect 598416 527738 598512 527794
rect 598568 527738 598636 527794
rect 598692 527738 598760 527794
rect 598816 527738 598884 527794
rect 598940 527738 599036 527794
rect 598416 527670 599036 527738
rect 598416 527614 598512 527670
rect 598568 527614 598636 527670
rect 598692 527614 598760 527670
rect 598816 527614 598884 527670
rect 598940 527614 599036 527670
rect 598416 527546 599036 527614
rect 598416 527490 598512 527546
rect 598568 527490 598636 527546
rect 598692 527490 598760 527546
rect 598816 527490 598884 527546
rect 598940 527490 599036 527546
rect 598416 509918 599036 527490
rect 598416 509862 598512 509918
rect 598568 509862 598636 509918
rect 598692 509862 598760 509918
rect 598816 509862 598884 509918
rect 598940 509862 599036 509918
rect 598416 509794 599036 509862
rect 598416 509738 598512 509794
rect 598568 509738 598636 509794
rect 598692 509738 598760 509794
rect 598816 509738 598884 509794
rect 598940 509738 599036 509794
rect 598416 509670 599036 509738
rect 598416 509614 598512 509670
rect 598568 509614 598636 509670
rect 598692 509614 598760 509670
rect 598816 509614 598884 509670
rect 598940 509614 599036 509670
rect 598416 509546 599036 509614
rect 598416 509490 598512 509546
rect 598568 509490 598636 509546
rect 598692 509490 598760 509546
rect 598816 509490 598884 509546
rect 598940 509490 599036 509546
rect 598416 491918 599036 509490
rect 598416 491862 598512 491918
rect 598568 491862 598636 491918
rect 598692 491862 598760 491918
rect 598816 491862 598884 491918
rect 598940 491862 599036 491918
rect 598416 491794 599036 491862
rect 598416 491738 598512 491794
rect 598568 491738 598636 491794
rect 598692 491738 598760 491794
rect 598816 491738 598884 491794
rect 598940 491738 599036 491794
rect 598416 491670 599036 491738
rect 598416 491614 598512 491670
rect 598568 491614 598636 491670
rect 598692 491614 598760 491670
rect 598816 491614 598884 491670
rect 598940 491614 599036 491670
rect 598416 491546 599036 491614
rect 598416 491490 598512 491546
rect 598568 491490 598636 491546
rect 598692 491490 598760 491546
rect 598816 491490 598884 491546
rect 598940 491490 599036 491546
rect 598416 473918 599036 491490
rect 598416 473862 598512 473918
rect 598568 473862 598636 473918
rect 598692 473862 598760 473918
rect 598816 473862 598884 473918
rect 598940 473862 599036 473918
rect 598416 473794 599036 473862
rect 598416 473738 598512 473794
rect 598568 473738 598636 473794
rect 598692 473738 598760 473794
rect 598816 473738 598884 473794
rect 598940 473738 599036 473794
rect 598416 473670 599036 473738
rect 598416 473614 598512 473670
rect 598568 473614 598636 473670
rect 598692 473614 598760 473670
rect 598816 473614 598884 473670
rect 598940 473614 599036 473670
rect 598416 473546 599036 473614
rect 598416 473490 598512 473546
rect 598568 473490 598636 473546
rect 598692 473490 598760 473546
rect 598816 473490 598884 473546
rect 598940 473490 599036 473546
rect 598416 455918 599036 473490
rect 598416 455862 598512 455918
rect 598568 455862 598636 455918
rect 598692 455862 598760 455918
rect 598816 455862 598884 455918
rect 598940 455862 599036 455918
rect 598416 455794 599036 455862
rect 598416 455738 598512 455794
rect 598568 455738 598636 455794
rect 598692 455738 598760 455794
rect 598816 455738 598884 455794
rect 598940 455738 599036 455794
rect 598416 455670 599036 455738
rect 598416 455614 598512 455670
rect 598568 455614 598636 455670
rect 598692 455614 598760 455670
rect 598816 455614 598884 455670
rect 598940 455614 599036 455670
rect 598416 455546 599036 455614
rect 598416 455490 598512 455546
rect 598568 455490 598636 455546
rect 598692 455490 598760 455546
rect 598816 455490 598884 455546
rect 598940 455490 599036 455546
rect 598416 437918 599036 455490
rect 598416 437862 598512 437918
rect 598568 437862 598636 437918
rect 598692 437862 598760 437918
rect 598816 437862 598884 437918
rect 598940 437862 599036 437918
rect 598416 437794 599036 437862
rect 598416 437738 598512 437794
rect 598568 437738 598636 437794
rect 598692 437738 598760 437794
rect 598816 437738 598884 437794
rect 598940 437738 599036 437794
rect 598416 437670 599036 437738
rect 598416 437614 598512 437670
rect 598568 437614 598636 437670
rect 598692 437614 598760 437670
rect 598816 437614 598884 437670
rect 598940 437614 599036 437670
rect 598416 437546 599036 437614
rect 598416 437490 598512 437546
rect 598568 437490 598636 437546
rect 598692 437490 598760 437546
rect 598816 437490 598884 437546
rect 598940 437490 599036 437546
rect 598416 419918 599036 437490
rect 598416 419862 598512 419918
rect 598568 419862 598636 419918
rect 598692 419862 598760 419918
rect 598816 419862 598884 419918
rect 598940 419862 599036 419918
rect 598416 419794 599036 419862
rect 598416 419738 598512 419794
rect 598568 419738 598636 419794
rect 598692 419738 598760 419794
rect 598816 419738 598884 419794
rect 598940 419738 599036 419794
rect 598416 419670 599036 419738
rect 598416 419614 598512 419670
rect 598568 419614 598636 419670
rect 598692 419614 598760 419670
rect 598816 419614 598884 419670
rect 598940 419614 599036 419670
rect 598416 419546 599036 419614
rect 598416 419490 598512 419546
rect 598568 419490 598636 419546
rect 598692 419490 598760 419546
rect 598816 419490 598884 419546
rect 598940 419490 599036 419546
rect 598416 401918 599036 419490
rect 598416 401862 598512 401918
rect 598568 401862 598636 401918
rect 598692 401862 598760 401918
rect 598816 401862 598884 401918
rect 598940 401862 599036 401918
rect 598416 401794 599036 401862
rect 598416 401738 598512 401794
rect 598568 401738 598636 401794
rect 598692 401738 598760 401794
rect 598816 401738 598884 401794
rect 598940 401738 599036 401794
rect 598416 401670 599036 401738
rect 598416 401614 598512 401670
rect 598568 401614 598636 401670
rect 598692 401614 598760 401670
rect 598816 401614 598884 401670
rect 598940 401614 599036 401670
rect 598416 401546 599036 401614
rect 598416 401490 598512 401546
rect 598568 401490 598636 401546
rect 598692 401490 598760 401546
rect 598816 401490 598884 401546
rect 598940 401490 599036 401546
rect 598416 383918 599036 401490
rect 598416 383862 598512 383918
rect 598568 383862 598636 383918
rect 598692 383862 598760 383918
rect 598816 383862 598884 383918
rect 598940 383862 599036 383918
rect 598416 383794 599036 383862
rect 598416 383738 598512 383794
rect 598568 383738 598636 383794
rect 598692 383738 598760 383794
rect 598816 383738 598884 383794
rect 598940 383738 599036 383794
rect 598416 383670 599036 383738
rect 598416 383614 598512 383670
rect 598568 383614 598636 383670
rect 598692 383614 598760 383670
rect 598816 383614 598884 383670
rect 598940 383614 599036 383670
rect 598416 383546 599036 383614
rect 598416 383490 598512 383546
rect 598568 383490 598636 383546
rect 598692 383490 598760 383546
rect 598816 383490 598884 383546
rect 598940 383490 599036 383546
rect 598416 365918 599036 383490
rect 598416 365862 598512 365918
rect 598568 365862 598636 365918
rect 598692 365862 598760 365918
rect 598816 365862 598884 365918
rect 598940 365862 599036 365918
rect 598416 365794 599036 365862
rect 598416 365738 598512 365794
rect 598568 365738 598636 365794
rect 598692 365738 598760 365794
rect 598816 365738 598884 365794
rect 598940 365738 599036 365794
rect 598416 365670 599036 365738
rect 598416 365614 598512 365670
rect 598568 365614 598636 365670
rect 598692 365614 598760 365670
rect 598816 365614 598884 365670
rect 598940 365614 599036 365670
rect 598416 365546 599036 365614
rect 598416 365490 598512 365546
rect 598568 365490 598636 365546
rect 598692 365490 598760 365546
rect 598816 365490 598884 365546
rect 598940 365490 599036 365546
rect 598416 347918 599036 365490
rect 598416 347862 598512 347918
rect 598568 347862 598636 347918
rect 598692 347862 598760 347918
rect 598816 347862 598884 347918
rect 598940 347862 599036 347918
rect 598416 347794 599036 347862
rect 598416 347738 598512 347794
rect 598568 347738 598636 347794
rect 598692 347738 598760 347794
rect 598816 347738 598884 347794
rect 598940 347738 599036 347794
rect 598416 347670 599036 347738
rect 598416 347614 598512 347670
rect 598568 347614 598636 347670
rect 598692 347614 598760 347670
rect 598816 347614 598884 347670
rect 598940 347614 599036 347670
rect 598416 347546 599036 347614
rect 598416 347490 598512 347546
rect 598568 347490 598636 347546
rect 598692 347490 598760 347546
rect 598816 347490 598884 347546
rect 598940 347490 599036 347546
rect 598416 329918 599036 347490
rect 598416 329862 598512 329918
rect 598568 329862 598636 329918
rect 598692 329862 598760 329918
rect 598816 329862 598884 329918
rect 598940 329862 599036 329918
rect 598416 329794 599036 329862
rect 598416 329738 598512 329794
rect 598568 329738 598636 329794
rect 598692 329738 598760 329794
rect 598816 329738 598884 329794
rect 598940 329738 599036 329794
rect 598416 329670 599036 329738
rect 598416 329614 598512 329670
rect 598568 329614 598636 329670
rect 598692 329614 598760 329670
rect 598816 329614 598884 329670
rect 598940 329614 599036 329670
rect 598416 329546 599036 329614
rect 598416 329490 598512 329546
rect 598568 329490 598636 329546
rect 598692 329490 598760 329546
rect 598816 329490 598884 329546
rect 598940 329490 599036 329546
rect 598416 311918 599036 329490
rect 598416 311862 598512 311918
rect 598568 311862 598636 311918
rect 598692 311862 598760 311918
rect 598816 311862 598884 311918
rect 598940 311862 599036 311918
rect 598416 311794 599036 311862
rect 598416 311738 598512 311794
rect 598568 311738 598636 311794
rect 598692 311738 598760 311794
rect 598816 311738 598884 311794
rect 598940 311738 599036 311794
rect 598416 311670 599036 311738
rect 598416 311614 598512 311670
rect 598568 311614 598636 311670
rect 598692 311614 598760 311670
rect 598816 311614 598884 311670
rect 598940 311614 599036 311670
rect 598416 311546 599036 311614
rect 598416 311490 598512 311546
rect 598568 311490 598636 311546
rect 598692 311490 598760 311546
rect 598816 311490 598884 311546
rect 598940 311490 599036 311546
rect 598416 293918 599036 311490
rect 598416 293862 598512 293918
rect 598568 293862 598636 293918
rect 598692 293862 598760 293918
rect 598816 293862 598884 293918
rect 598940 293862 599036 293918
rect 598416 293794 599036 293862
rect 598416 293738 598512 293794
rect 598568 293738 598636 293794
rect 598692 293738 598760 293794
rect 598816 293738 598884 293794
rect 598940 293738 599036 293794
rect 598416 293670 599036 293738
rect 598416 293614 598512 293670
rect 598568 293614 598636 293670
rect 598692 293614 598760 293670
rect 598816 293614 598884 293670
rect 598940 293614 599036 293670
rect 598416 293546 599036 293614
rect 598416 293490 598512 293546
rect 598568 293490 598636 293546
rect 598692 293490 598760 293546
rect 598816 293490 598884 293546
rect 598940 293490 599036 293546
rect 598416 275918 599036 293490
rect 598416 275862 598512 275918
rect 598568 275862 598636 275918
rect 598692 275862 598760 275918
rect 598816 275862 598884 275918
rect 598940 275862 599036 275918
rect 598416 275794 599036 275862
rect 598416 275738 598512 275794
rect 598568 275738 598636 275794
rect 598692 275738 598760 275794
rect 598816 275738 598884 275794
rect 598940 275738 599036 275794
rect 598416 275670 599036 275738
rect 598416 275614 598512 275670
rect 598568 275614 598636 275670
rect 598692 275614 598760 275670
rect 598816 275614 598884 275670
rect 598940 275614 599036 275670
rect 598416 275546 599036 275614
rect 598416 275490 598512 275546
rect 598568 275490 598636 275546
rect 598692 275490 598760 275546
rect 598816 275490 598884 275546
rect 598940 275490 599036 275546
rect 598416 257918 599036 275490
rect 598416 257862 598512 257918
rect 598568 257862 598636 257918
rect 598692 257862 598760 257918
rect 598816 257862 598884 257918
rect 598940 257862 599036 257918
rect 598416 257794 599036 257862
rect 598416 257738 598512 257794
rect 598568 257738 598636 257794
rect 598692 257738 598760 257794
rect 598816 257738 598884 257794
rect 598940 257738 599036 257794
rect 598416 257670 599036 257738
rect 598416 257614 598512 257670
rect 598568 257614 598636 257670
rect 598692 257614 598760 257670
rect 598816 257614 598884 257670
rect 598940 257614 599036 257670
rect 598416 257546 599036 257614
rect 598416 257490 598512 257546
rect 598568 257490 598636 257546
rect 598692 257490 598760 257546
rect 598816 257490 598884 257546
rect 598940 257490 599036 257546
rect 598416 239918 599036 257490
rect 598416 239862 598512 239918
rect 598568 239862 598636 239918
rect 598692 239862 598760 239918
rect 598816 239862 598884 239918
rect 598940 239862 599036 239918
rect 598416 239794 599036 239862
rect 598416 239738 598512 239794
rect 598568 239738 598636 239794
rect 598692 239738 598760 239794
rect 598816 239738 598884 239794
rect 598940 239738 599036 239794
rect 598416 239670 599036 239738
rect 598416 239614 598512 239670
rect 598568 239614 598636 239670
rect 598692 239614 598760 239670
rect 598816 239614 598884 239670
rect 598940 239614 599036 239670
rect 598416 239546 599036 239614
rect 598416 239490 598512 239546
rect 598568 239490 598636 239546
rect 598692 239490 598760 239546
rect 598816 239490 598884 239546
rect 598940 239490 599036 239546
rect 598416 221918 599036 239490
rect 598416 221862 598512 221918
rect 598568 221862 598636 221918
rect 598692 221862 598760 221918
rect 598816 221862 598884 221918
rect 598940 221862 599036 221918
rect 598416 221794 599036 221862
rect 598416 221738 598512 221794
rect 598568 221738 598636 221794
rect 598692 221738 598760 221794
rect 598816 221738 598884 221794
rect 598940 221738 599036 221794
rect 598416 221670 599036 221738
rect 598416 221614 598512 221670
rect 598568 221614 598636 221670
rect 598692 221614 598760 221670
rect 598816 221614 598884 221670
rect 598940 221614 599036 221670
rect 598416 221546 599036 221614
rect 598416 221490 598512 221546
rect 598568 221490 598636 221546
rect 598692 221490 598760 221546
rect 598816 221490 598884 221546
rect 598940 221490 599036 221546
rect 598416 203918 599036 221490
rect 598416 203862 598512 203918
rect 598568 203862 598636 203918
rect 598692 203862 598760 203918
rect 598816 203862 598884 203918
rect 598940 203862 599036 203918
rect 598416 203794 599036 203862
rect 598416 203738 598512 203794
rect 598568 203738 598636 203794
rect 598692 203738 598760 203794
rect 598816 203738 598884 203794
rect 598940 203738 599036 203794
rect 598416 203670 599036 203738
rect 598416 203614 598512 203670
rect 598568 203614 598636 203670
rect 598692 203614 598760 203670
rect 598816 203614 598884 203670
rect 598940 203614 599036 203670
rect 598416 203546 599036 203614
rect 598416 203490 598512 203546
rect 598568 203490 598636 203546
rect 598692 203490 598760 203546
rect 598816 203490 598884 203546
rect 598940 203490 599036 203546
rect 598416 185918 599036 203490
rect 598416 185862 598512 185918
rect 598568 185862 598636 185918
rect 598692 185862 598760 185918
rect 598816 185862 598884 185918
rect 598940 185862 599036 185918
rect 598416 185794 599036 185862
rect 598416 185738 598512 185794
rect 598568 185738 598636 185794
rect 598692 185738 598760 185794
rect 598816 185738 598884 185794
rect 598940 185738 599036 185794
rect 598416 185670 599036 185738
rect 598416 185614 598512 185670
rect 598568 185614 598636 185670
rect 598692 185614 598760 185670
rect 598816 185614 598884 185670
rect 598940 185614 599036 185670
rect 598416 185546 599036 185614
rect 598416 185490 598512 185546
rect 598568 185490 598636 185546
rect 598692 185490 598760 185546
rect 598816 185490 598884 185546
rect 598940 185490 599036 185546
rect 598416 167918 599036 185490
rect 598416 167862 598512 167918
rect 598568 167862 598636 167918
rect 598692 167862 598760 167918
rect 598816 167862 598884 167918
rect 598940 167862 599036 167918
rect 598416 167794 599036 167862
rect 598416 167738 598512 167794
rect 598568 167738 598636 167794
rect 598692 167738 598760 167794
rect 598816 167738 598884 167794
rect 598940 167738 599036 167794
rect 598416 167670 599036 167738
rect 598416 167614 598512 167670
rect 598568 167614 598636 167670
rect 598692 167614 598760 167670
rect 598816 167614 598884 167670
rect 598940 167614 599036 167670
rect 598416 167546 599036 167614
rect 598416 167490 598512 167546
rect 598568 167490 598636 167546
rect 598692 167490 598760 167546
rect 598816 167490 598884 167546
rect 598940 167490 599036 167546
rect 598416 149918 599036 167490
rect 598416 149862 598512 149918
rect 598568 149862 598636 149918
rect 598692 149862 598760 149918
rect 598816 149862 598884 149918
rect 598940 149862 599036 149918
rect 598416 149794 599036 149862
rect 598416 149738 598512 149794
rect 598568 149738 598636 149794
rect 598692 149738 598760 149794
rect 598816 149738 598884 149794
rect 598940 149738 599036 149794
rect 598416 149670 599036 149738
rect 598416 149614 598512 149670
rect 598568 149614 598636 149670
rect 598692 149614 598760 149670
rect 598816 149614 598884 149670
rect 598940 149614 599036 149670
rect 598416 149546 599036 149614
rect 598416 149490 598512 149546
rect 598568 149490 598636 149546
rect 598692 149490 598760 149546
rect 598816 149490 598884 149546
rect 598940 149490 599036 149546
rect 598416 131918 599036 149490
rect 598416 131862 598512 131918
rect 598568 131862 598636 131918
rect 598692 131862 598760 131918
rect 598816 131862 598884 131918
rect 598940 131862 599036 131918
rect 598416 131794 599036 131862
rect 598416 131738 598512 131794
rect 598568 131738 598636 131794
rect 598692 131738 598760 131794
rect 598816 131738 598884 131794
rect 598940 131738 599036 131794
rect 598416 131670 599036 131738
rect 598416 131614 598512 131670
rect 598568 131614 598636 131670
rect 598692 131614 598760 131670
rect 598816 131614 598884 131670
rect 598940 131614 599036 131670
rect 598416 131546 599036 131614
rect 598416 131490 598512 131546
rect 598568 131490 598636 131546
rect 598692 131490 598760 131546
rect 598816 131490 598884 131546
rect 598940 131490 599036 131546
rect 598416 113918 599036 131490
rect 598416 113862 598512 113918
rect 598568 113862 598636 113918
rect 598692 113862 598760 113918
rect 598816 113862 598884 113918
rect 598940 113862 599036 113918
rect 598416 113794 599036 113862
rect 598416 113738 598512 113794
rect 598568 113738 598636 113794
rect 598692 113738 598760 113794
rect 598816 113738 598884 113794
rect 598940 113738 599036 113794
rect 598416 113670 599036 113738
rect 598416 113614 598512 113670
rect 598568 113614 598636 113670
rect 598692 113614 598760 113670
rect 598816 113614 598884 113670
rect 598940 113614 599036 113670
rect 598416 113546 599036 113614
rect 598416 113490 598512 113546
rect 598568 113490 598636 113546
rect 598692 113490 598760 113546
rect 598816 113490 598884 113546
rect 598940 113490 599036 113546
rect 598416 95918 599036 113490
rect 598416 95862 598512 95918
rect 598568 95862 598636 95918
rect 598692 95862 598760 95918
rect 598816 95862 598884 95918
rect 598940 95862 599036 95918
rect 598416 95794 599036 95862
rect 598416 95738 598512 95794
rect 598568 95738 598636 95794
rect 598692 95738 598760 95794
rect 598816 95738 598884 95794
rect 598940 95738 599036 95794
rect 598416 95670 599036 95738
rect 598416 95614 598512 95670
rect 598568 95614 598636 95670
rect 598692 95614 598760 95670
rect 598816 95614 598884 95670
rect 598940 95614 599036 95670
rect 598416 95546 599036 95614
rect 598416 95490 598512 95546
rect 598568 95490 598636 95546
rect 598692 95490 598760 95546
rect 598816 95490 598884 95546
rect 598940 95490 599036 95546
rect 598416 77918 599036 95490
rect 598416 77862 598512 77918
rect 598568 77862 598636 77918
rect 598692 77862 598760 77918
rect 598816 77862 598884 77918
rect 598940 77862 599036 77918
rect 598416 77794 599036 77862
rect 598416 77738 598512 77794
rect 598568 77738 598636 77794
rect 598692 77738 598760 77794
rect 598816 77738 598884 77794
rect 598940 77738 599036 77794
rect 598416 77670 599036 77738
rect 598416 77614 598512 77670
rect 598568 77614 598636 77670
rect 598692 77614 598760 77670
rect 598816 77614 598884 77670
rect 598940 77614 599036 77670
rect 598416 77546 599036 77614
rect 598416 77490 598512 77546
rect 598568 77490 598636 77546
rect 598692 77490 598760 77546
rect 598816 77490 598884 77546
rect 598940 77490 599036 77546
rect 598416 59918 599036 77490
rect 598416 59862 598512 59918
rect 598568 59862 598636 59918
rect 598692 59862 598760 59918
rect 598816 59862 598884 59918
rect 598940 59862 599036 59918
rect 598416 59794 599036 59862
rect 598416 59738 598512 59794
rect 598568 59738 598636 59794
rect 598692 59738 598760 59794
rect 598816 59738 598884 59794
rect 598940 59738 599036 59794
rect 598416 59670 599036 59738
rect 598416 59614 598512 59670
rect 598568 59614 598636 59670
rect 598692 59614 598760 59670
rect 598816 59614 598884 59670
rect 598940 59614 599036 59670
rect 598416 59546 599036 59614
rect 598416 59490 598512 59546
rect 598568 59490 598636 59546
rect 598692 59490 598760 59546
rect 598816 59490 598884 59546
rect 598940 59490 599036 59546
rect 598416 41918 599036 59490
rect 598416 41862 598512 41918
rect 598568 41862 598636 41918
rect 598692 41862 598760 41918
rect 598816 41862 598884 41918
rect 598940 41862 599036 41918
rect 598416 41794 599036 41862
rect 598416 41738 598512 41794
rect 598568 41738 598636 41794
rect 598692 41738 598760 41794
rect 598816 41738 598884 41794
rect 598940 41738 599036 41794
rect 598416 41670 599036 41738
rect 598416 41614 598512 41670
rect 598568 41614 598636 41670
rect 598692 41614 598760 41670
rect 598816 41614 598884 41670
rect 598940 41614 599036 41670
rect 598416 41546 599036 41614
rect 598416 41490 598512 41546
rect 598568 41490 598636 41546
rect 598692 41490 598760 41546
rect 598816 41490 598884 41546
rect 598940 41490 599036 41546
rect 598416 23918 599036 41490
rect 598416 23862 598512 23918
rect 598568 23862 598636 23918
rect 598692 23862 598760 23918
rect 598816 23862 598884 23918
rect 598940 23862 599036 23918
rect 598416 23794 599036 23862
rect 598416 23738 598512 23794
rect 598568 23738 598636 23794
rect 598692 23738 598760 23794
rect 598816 23738 598884 23794
rect 598940 23738 599036 23794
rect 598416 23670 599036 23738
rect 598416 23614 598512 23670
rect 598568 23614 598636 23670
rect 598692 23614 598760 23670
rect 598816 23614 598884 23670
rect 598940 23614 599036 23670
rect 598416 23546 599036 23614
rect 598416 23490 598512 23546
rect 598568 23490 598636 23546
rect 598692 23490 598760 23546
rect 598816 23490 598884 23546
rect 598940 23490 599036 23546
rect 598416 5918 599036 23490
rect 598416 5862 598512 5918
rect 598568 5862 598636 5918
rect 598692 5862 598760 5918
rect 598816 5862 598884 5918
rect 598940 5862 599036 5918
rect 598416 5794 599036 5862
rect 598416 5738 598512 5794
rect 598568 5738 598636 5794
rect 598692 5738 598760 5794
rect 598816 5738 598884 5794
rect 598940 5738 599036 5794
rect 598416 5670 599036 5738
rect 598416 5614 598512 5670
rect 598568 5614 598636 5670
rect 598692 5614 598760 5670
rect 598816 5614 598884 5670
rect 598940 5614 599036 5670
rect 598416 5546 599036 5614
rect 598416 5490 598512 5546
rect 598568 5490 598636 5546
rect 598692 5490 598760 5546
rect 598816 5490 598884 5546
rect 598940 5490 599036 5546
rect 5058 1752 5154 1808
rect 5210 1752 5278 1808
rect 5334 1752 5402 1808
rect 5458 1752 5526 1808
rect 5582 1752 5678 1808
rect 5058 1684 5678 1752
rect 5058 1628 5154 1684
rect 5210 1628 5278 1684
rect 5334 1628 5402 1684
rect 5458 1628 5526 1684
rect 5582 1628 5678 1684
rect 5058 1560 5678 1628
rect 5058 1504 5154 1560
rect 5210 1504 5278 1560
rect 5334 1504 5402 1560
rect 5458 1504 5526 1560
rect 5582 1504 5678 1560
rect 5058 1436 5678 1504
rect 5058 1380 5154 1436
rect 5210 1380 5278 1436
rect 5334 1380 5402 1436
rect 5458 1380 5526 1436
rect 5582 1380 5678 1436
rect -12 792 84 848
rect 140 792 208 848
rect 264 792 332 848
rect 388 792 456 848
rect 512 792 608 848
rect -12 724 608 792
rect -12 668 84 724
rect 140 668 208 724
rect 264 668 332 724
rect 388 668 456 724
rect 512 668 608 724
rect -12 600 608 668
rect -12 544 84 600
rect 140 544 208 600
rect 264 544 332 600
rect 388 544 456 600
rect 512 544 608 600
rect -12 476 608 544
rect -12 420 84 476
rect 140 420 208 476
rect 264 420 332 476
rect 388 420 456 476
rect 512 420 608 476
rect -12 324 608 420
rect 5058 324 5678 1380
rect 8778 848 9398 2326
rect 8778 792 8874 848
rect 8930 792 8998 848
rect 9054 792 9122 848
rect 9178 792 9246 848
rect 9302 792 9398 848
rect 8778 724 9398 792
rect 8778 668 8874 724
rect 8930 668 8998 724
rect 9054 668 9122 724
rect 9178 668 9246 724
rect 9302 668 9398 724
rect 8778 600 9398 668
rect 8778 544 8874 600
rect 8930 544 8998 600
rect 9054 544 9122 600
rect 9178 544 9246 600
rect 9302 544 9398 600
rect 8778 476 9398 544
rect 8778 420 8874 476
rect 8930 420 8998 476
rect 9054 420 9122 476
rect 9178 420 9246 476
rect 9302 420 9398 476
rect 8778 324 9398 420
rect 23058 1808 23678 2326
rect 23058 1752 23154 1808
rect 23210 1752 23278 1808
rect 23334 1752 23402 1808
rect 23458 1752 23526 1808
rect 23582 1752 23678 1808
rect 23058 1684 23678 1752
rect 23058 1628 23154 1684
rect 23210 1628 23278 1684
rect 23334 1628 23402 1684
rect 23458 1628 23526 1684
rect 23582 1628 23678 1684
rect 23058 1560 23678 1628
rect 23058 1504 23154 1560
rect 23210 1504 23278 1560
rect 23334 1504 23402 1560
rect 23458 1504 23526 1560
rect 23582 1504 23678 1560
rect 23058 1436 23678 1504
rect 23058 1380 23154 1436
rect 23210 1380 23278 1436
rect 23334 1380 23402 1436
rect 23458 1380 23526 1436
rect 23582 1380 23678 1436
rect 23058 324 23678 1380
rect 26778 848 27398 2326
rect 26778 792 26874 848
rect 26930 792 26998 848
rect 27054 792 27122 848
rect 27178 792 27246 848
rect 27302 792 27398 848
rect 26778 724 27398 792
rect 26778 668 26874 724
rect 26930 668 26998 724
rect 27054 668 27122 724
rect 27178 668 27246 724
rect 27302 668 27398 724
rect 26778 600 27398 668
rect 26778 544 26874 600
rect 26930 544 26998 600
rect 27054 544 27122 600
rect 27178 544 27246 600
rect 27302 544 27398 600
rect 26778 476 27398 544
rect 26778 420 26874 476
rect 26930 420 26998 476
rect 27054 420 27122 476
rect 27178 420 27246 476
rect 27302 420 27398 476
rect 26778 324 27398 420
rect 41058 1808 41678 2326
rect 41058 1752 41154 1808
rect 41210 1752 41278 1808
rect 41334 1752 41402 1808
rect 41458 1752 41526 1808
rect 41582 1752 41678 1808
rect 41058 1684 41678 1752
rect 41058 1628 41154 1684
rect 41210 1628 41278 1684
rect 41334 1628 41402 1684
rect 41458 1628 41526 1684
rect 41582 1628 41678 1684
rect 41058 1560 41678 1628
rect 41058 1504 41154 1560
rect 41210 1504 41278 1560
rect 41334 1504 41402 1560
rect 41458 1504 41526 1560
rect 41582 1504 41678 1560
rect 41058 1436 41678 1504
rect 41058 1380 41154 1436
rect 41210 1380 41278 1436
rect 41334 1380 41402 1436
rect 41458 1380 41526 1436
rect 41582 1380 41678 1436
rect 41058 324 41678 1380
rect 44778 848 45398 2326
rect 44778 792 44874 848
rect 44930 792 44998 848
rect 45054 792 45122 848
rect 45178 792 45246 848
rect 45302 792 45398 848
rect 44778 724 45398 792
rect 44778 668 44874 724
rect 44930 668 44998 724
rect 45054 668 45122 724
rect 45178 668 45246 724
rect 45302 668 45398 724
rect 44778 600 45398 668
rect 44778 544 44874 600
rect 44930 544 44998 600
rect 45054 544 45122 600
rect 45178 544 45246 600
rect 45302 544 45398 600
rect 44778 476 45398 544
rect 44778 420 44874 476
rect 44930 420 44998 476
rect 45054 420 45122 476
rect 45178 420 45246 476
rect 45302 420 45398 476
rect 44778 324 45398 420
rect 59058 1808 59678 2326
rect 59058 1752 59154 1808
rect 59210 1752 59278 1808
rect 59334 1752 59402 1808
rect 59458 1752 59526 1808
rect 59582 1752 59678 1808
rect 59058 1684 59678 1752
rect 59058 1628 59154 1684
rect 59210 1628 59278 1684
rect 59334 1628 59402 1684
rect 59458 1628 59526 1684
rect 59582 1628 59678 1684
rect 59058 1560 59678 1628
rect 59058 1504 59154 1560
rect 59210 1504 59278 1560
rect 59334 1504 59402 1560
rect 59458 1504 59526 1560
rect 59582 1504 59678 1560
rect 59058 1436 59678 1504
rect 59058 1380 59154 1436
rect 59210 1380 59278 1436
rect 59334 1380 59402 1436
rect 59458 1380 59526 1436
rect 59582 1380 59678 1436
rect 59058 324 59678 1380
rect 62778 848 63398 2326
rect 62778 792 62874 848
rect 62930 792 62998 848
rect 63054 792 63122 848
rect 63178 792 63246 848
rect 63302 792 63398 848
rect 62778 724 63398 792
rect 62778 668 62874 724
rect 62930 668 62998 724
rect 63054 668 63122 724
rect 63178 668 63246 724
rect 63302 668 63398 724
rect 62778 600 63398 668
rect 62778 544 62874 600
rect 62930 544 62998 600
rect 63054 544 63122 600
rect 63178 544 63246 600
rect 63302 544 63398 600
rect 62778 476 63398 544
rect 62778 420 62874 476
rect 62930 420 62998 476
rect 63054 420 63122 476
rect 63178 420 63246 476
rect 63302 420 63398 476
rect 62778 324 63398 420
rect 77058 1808 77678 2326
rect 77058 1752 77154 1808
rect 77210 1752 77278 1808
rect 77334 1752 77402 1808
rect 77458 1752 77526 1808
rect 77582 1752 77678 1808
rect 77058 1684 77678 1752
rect 77058 1628 77154 1684
rect 77210 1628 77278 1684
rect 77334 1628 77402 1684
rect 77458 1628 77526 1684
rect 77582 1628 77678 1684
rect 77058 1560 77678 1628
rect 77058 1504 77154 1560
rect 77210 1504 77278 1560
rect 77334 1504 77402 1560
rect 77458 1504 77526 1560
rect 77582 1504 77678 1560
rect 77058 1436 77678 1504
rect 77058 1380 77154 1436
rect 77210 1380 77278 1436
rect 77334 1380 77402 1436
rect 77458 1380 77526 1436
rect 77582 1380 77678 1436
rect 77058 324 77678 1380
rect 80778 848 81398 2326
rect 80778 792 80874 848
rect 80930 792 80998 848
rect 81054 792 81122 848
rect 81178 792 81246 848
rect 81302 792 81398 848
rect 80778 724 81398 792
rect 80778 668 80874 724
rect 80930 668 80998 724
rect 81054 668 81122 724
rect 81178 668 81246 724
rect 81302 668 81398 724
rect 80778 600 81398 668
rect 80778 544 80874 600
rect 80930 544 80998 600
rect 81054 544 81122 600
rect 81178 544 81246 600
rect 81302 544 81398 600
rect 80778 476 81398 544
rect 80778 420 80874 476
rect 80930 420 80998 476
rect 81054 420 81122 476
rect 81178 420 81246 476
rect 81302 420 81398 476
rect 80778 324 81398 420
rect 95058 1808 95678 2326
rect 95058 1752 95154 1808
rect 95210 1752 95278 1808
rect 95334 1752 95402 1808
rect 95458 1752 95526 1808
rect 95582 1752 95678 1808
rect 95058 1684 95678 1752
rect 95058 1628 95154 1684
rect 95210 1628 95278 1684
rect 95334 1628 95402 1684
rect 95458 1628 95526 1684
rect 95582 1628 95678 1684
rect 95058 1560 95678 1628
rect 95058 1504 95154 1560
rect 95210 1504 95278 1560
rect 95334 1504 95402 1560
rect 95458 1504 95526 1560
rect 95582 1504 95678 1560
rect 95058 1436 95678 1504
rect 95058 1380 95154 1436
rect 95210 1380 95278 1436
rect 95334 1380 95402 1436
rect 95458 1380 95526 1436
rect 95582 1380 95678 1436
rect 95058 324 95678 1380
rect 98778 848 99398 2326
rect 98778 792 98874 848
rect 98930 792 98998 848
rect 99054 792 99122 848
rect 99178 792 99246 848
rect 99302 792 99398 848
rect 98778 724 99398 792
rect 98778 668 98874 724
rect 98930 668 98998 724
rect 99054 668 99122 724
rect 99178 668 99246 724
rect 99302 668 99398 724
rect 98778 600 99398 668
rect 98778 544 98874 600
rect 98930 544 98998 600
rect 99054 544 99122 600
rect 99178 544 99246 600
rect 99302 544 99398 600
rect 98778 476 99398 544
rect 98778 420 98874 476
rect 98930 420 98998 476
rect 99054 420 99122 476
rect 99178 420 99246 476
rect 99302 420 99398 476
rect 98778 324 99398 420
rect 113058 1808 113678 2326
rect 113058 1752 113154 1808
rect 113210 1752 113278 1808
rect 113334 1752 113402 1808
rect 113458 1752 113526 1808
rect 113582 1752 113678 1808
rect 113058 1684 113678 1752
rect 113058 1628 113154 1684
rect 113210 1628 113278 1684
rect 113334 1628 113402 1684
rect 113458 1628 113526 1684
rect 113582 1628 113678 1684
rect 113058 1560 113678 1628
rect 113058 1504 113154 1560
rect 113210 1504 113278 1560
rect 113334 1504 113402 1560
rect 113458 1504 113526 1560
rect 113582 1504 113678 1560
rect 113058 1436 113678 1504
rect 113058 1380 113154 1436
rect 113210 1380 113278 1436
rect 113334 1380 113402 1436
rect 113458 1380 113526 1436
rect 113582 1380 113678 1436
rect 113058 324 113678 1380
rect 116778 848 117398 2326
rect 116778 792 116874 848
rect 116930 792 116998 848
rect 117054 792 117122 848
rect 117178 792 117246 848
rect 117302 792 117398 848
rect 116778 724 117398 792
rect 116778 668 116874 724
rect 116930 668 116998 724
rect 117054 668 117122 724
rect 117178 668 117246 724
rect 117302 668 117398 724
rect 116778 600 117398 668
rect 116778 544 116874 600
rect 116930 544 116998 600
rect 117054 544 117122 600
rect 117178 544 117246 600
rect 117302 544 117398 600
rect 116778 476 117398 544
rect 116778 420 116874 476
rect 116930 420 116998 476
rect 117054 420 117122 476
rect 117178 420 117246 476
rect 117302 420 117398 476
rect 116778 324 117398 420
rect 131058 1808 131678 2326
rect 131058 1752 131154 1808
rect 131210 1752 131278 1808
rect 131334 1752 131402 1808
rect 131458 1752 131526 1808
rect 131582 1752 131678 1808
rect 131058 1684 131678 1752
rect 131058 1628 131154 1684
rect 131210 1628 131278 1684
rect 131334 1628 131402 1684
rect 131458 1628 131526 1684
rect 131582 1628 131678 1684
rect 131058 1560 131678 1628
rect 131058 1504 131154 1560
rect 131210 1504 131278 1560
rect 131334 1504 131402 1560
rect 131458 1504 131526 1560
rect 131582 1504 131678 1560
rect 131058 1436 131678 1504
rect 131058 1380 131154 1436
rect 131210 1380 131278 1436
rect 131334 1380 131402 1436
rect 131458 1380 131526 1436
rect 131582 1380 131678 1436
rect 131058 324 131678 1380
rect 134778 848 135398 2326
rect 134778 792 134874 848
rect 134930 792 134998 848
rect 135054 792 135122 848
rect 135178 792 135246 848
rect 135302 792 135398 848
rect 134778 724 135398 792
rect 134778 668 134874 724
rect 134930 668 134998 724
rect 135054 668 135122 724
rect 135178 668 135246 724
rect 135302 668 135398 724
rect 134778 600 135398 668
rect 134778 544 134874 600
rect 134930 544 134998 600
rect 135054 544 135122 600
rect 135178 544 135246 600
rect 135302 544 135398 600
rect 134778 476 135398 544
rect 134778 420 134874 476
rect 134930 420 134998 476
rect 135054 420 135122 476
rect 135178 420 135246 476
rect 135302 420 135398 476
rect 134778 324 135398 420
rect 149058 1808 149678 2326
rect 149058 1752 149154 1808
rect 149210 1752 149278 1808
rect 149334 1752 149402 1808
rect 149458 1752 149526 1808
rect 149582 1752 149678 1808
rect 149058 1684 149678 1752
rect 149058 1628 149154 1684
rect 149210 1628 149278 1684
rect 149334 1628 149402 1684
rect 149458 1628 149526 1684
rect 149582 1628 149678 1684
rect 149058 1560 149678 1628
rect 149058 1504 149154 1560
rect 149210 1504 149278 1560
rect 149334 1504 149402 1560
rect 149458 1504 149526 1560
rect 149582 1504 149678 1560
rect 149058 1436 149678 1504
rect 149058 1380 149154 1436
rect 149210 1380 149278 1436
rect 149334 1380 149402 1436
rect 149458 1380 149526 1436
rect 149582 1380 149678 1436
rect 149058 324 149678 1380
rect 152778 848 153398 2326
rect 152778 792 152874 848
rect 152930 792 152998 848
rect 153054 792 153122 848
rect 153178 792 153246 848
rect 153302 792 153398 848
rect 152778 724 153398 792
rect 152778 668 152874 724
rect 152930 668 152998 724
rect 153054 668 153122 724
rect 153178 668 153246 724
rect 153302 668 153398 724
rect 152778 600 153398 668
rect 152778 544 152874 600
rect 152930 544 152998 600
rect 153054 544 153122 600
rect 153178 544 153246 600
rect 153302 544 153398 600
rect 152778 476 153398 544
rect 152778 420 152874 476
rect 152930 420 152998 476
rect 153054 420 153122 476
rect 153178 420 153246 476
rect 153302 420 153398 476
rect 152778 324 153398 420
rect 167058 1808 167678 2326
rect 167058 1752 167154 1808
rect 167210 1752 167278 1808
rect 167334 1752 167402 1808
rect 167458 1752 167526 1808
rect 167582 1752 167678 1808
rect 167058 1684 167678 1752
rect 167058 1628 167154 1684
rect 167210 1628 167278 1684
rect 167334 1628 167402 1684
rect 167458 1628 167526 1684
rect 167582 1628 167678 1684
rect 167058 1560 167678 1628
rect 167058 1504 167154 1560
rect 167210 1504 167278 1560
rect 167334 1504 167402 1560
rect 167458 1504 167526 1560
rect 167582 1504 167678 1560
rect 167058 1436 167678 1504
rect 167058 1380 167154 1436
rect 167210 1380 167278 1436
rect 167334 1380 167402 1436
rect 167458 1380 167526 1436
rect 167582 1380 167678 1436
rect 167058 324 167678 1380
rect 170778 848 171398 2326
rect 170778 792 170874 848
rect 170930 792 170998 848
rect 171054 792 171122 848
rect 171178 792 171246 848
rect 171302 792 171398 848
rect 170778 724 171398 792
rect 170778 668 170874 724
rect 170930 668 170998 724
rect 171054 668 171122 724
rect 171178 668 171246 724
rect 171302 668 171398 724
rect 170778 600 171398 668
rect 170778 544 170874 600
rect 170930 544 170998 600
rect 171054 544 171122 600
rect 171178 544 171246 600
rect 171302 544 171398 600
rect 170778 476 171398 544
rect 170778 420 170874 476
rect 170930 420 170998 476
rect 171054 420 171122 476
rect 171178 420 171246 476
rect 171302 420 171398 476
rect 170778 324 171398 420
rect 185058 1808 185678 2326
rect 185058 1752 185154 1808
rect 185210 1752 185278 1808
rect 185334 1752 185402 1808
rect 185458 1752 185526 1808
rect 185582 1752 185678 1808
rect 185058 1684 185678 1752
rect 185058 1628 185154 1684
rect 185210 1628 185278 1684
rect 185334 1628 185402 1684
rect 185458 1628 185526 1684
rect 185582 1628 185678 1684
rect 185058 1560 185678 1628
rect 185058 1504 185154 1560
rect 185210 1504 185278 1560
rect 185334 1504 185402 1560
rect 185458 1504 185526 1560
rect 185582 1504 185678 1560
rect 185058 1436 185678 1504
rect 185058 1380 185154 1436
rect 185210 1380 185278 1436
rect 185334 1380 185402 1436
rect 185458 1380 185526 1436
rect 185582 1380 185678 1436
rect 185058 324 185678 1380
rect 188778 848 189398 2326
rect 188778 792 188874 848
rect 188930 792 188998 848
rect 189054 792 189122 848
rect 189178 792 189246 848
rect 189302 792 189398 848
rect 188778 724 189398 792
rect 188778 668 188874 724
rect 188930 668 188998 724
rect 189054 668 189122 724
rect 189178 668 189246 724
rect 189302 668 189398 724
rect 188778 600 189398 668
rect 188778 544 188874 600
rect 188930 544 188998 600
rect 189054 544 189122 600
rect 189178 544 189246 600
rect 189302 544 189398 600
rect 188778 476 189398 544
rect 188778 420 188874 476
rect 188930 420 188998 476
rect 189054 420 189122 476
rect 189178 420 189246 476
rect 189302 420 189398 476
rect 188778 324 189398 420
rect 203058 1808 203678 2326
rect 203058 1752 203154 1808
rect 203210 1752 203278 1808
rect 203334 1752 203402 1808
rect 203458 1752 203526 1808
rect 203582 1752 203678 1808
rect 203058 1684 203678 1752
rect 203058 1628 203154 1684
rect 203210 1628 203278 1684
rect 203334 1628 203402 1684
rect 203458 1628 203526 1684
rect 203582 1628 203678 1684
rect 203058 1560 203678 1628
rect 203058 1504 203154 1560
rect 203210 1504 203278 1560
rect 203334 1504 203402 1560
rect 203458 1504 203526 1560
rect 203582 1504 203678 1560
rect 203058 1436 203678 1504
rect 203058 1380 203154 1436
rect 203210 1380 203278 1436
rect 203334 1380 203402 1436
rect 203458 1380 203526 1436
rect 203582 1380 203678 1436
rect 203058 324 203678 1380
rect 206778 848 207398 2326
rect 206778 792 206874 848
rect 206930 792 206998 848
rect 207054 792 207122 848
rect 207178 792 207246 848
rect 207302 792 207398 848
rect 206778 724 207398 792
rect 206778 668 206874 724
rect 206930 668 206998 724
rect 207054 668 207122 724
rect 207178 668 207246 724
rect 207302 668 207398 724
rect 206778 600 207398 668
rect 206778 544 206874 600
rect 206930 544 206998 600
rect 207054 544 207122 600
rect 207178 544 207246 600
rect 207302 544 207398 600
rect 206778 476 207398 544
rect 206778 420 206874 476
rect 206930 420 206998 476
rect 207054 420 207122 476
rect 207178 420 207246 476
rect 207302 420 207398 476
rect 206778 324 207398 420
rect 221058 1808 221678 2326
rect 221058 1752 221154 1808
rect 221210 1752 221278 1808
rect 221334 1752 221402 1808
rect 221458 1752 221526 1808
rect 221582 1752 221678 1808
rect 221058 1684 221678 1752
rect 221058 1628 221154 1684
rect 221210 1628 221278 1684
rect 221334 1628 221402 1684
rect 221458 1628 221526 1684
rect 221582 1628 221678 1684
rect 221058 1560 221678 1628
rect 221058 1504 221154 1560
rect 221210 1504 221278 1560
rect 221334 1504 221402 1560
rect 221458 1504 221526 1560
rect 221582 1504 221678 1560
rect 221058 1436 221678 1504
rect 221058 1380 221154 1436
rect 221210 1380 221278 1436
rect 221334 1380 221402 1436
rect 221458 1380 221526 1436
rect 221582 1380 221678 1436
rect 221058 324 221678 1380
rect 224778 848 225398 2326
rect 224778 792 224874 848
rect 224930 792 224998 848
rect 225054 792 225122 848
rect 225178 792 225246 848
rect 225302 792 225398 848
rect 224778 724 225398 792
rect 224778 668 224874 724
rect 224930 668 224998 724
rect 225054 668 225122 724
rect 225178 668 225246 724
rect 225302 668 225398 724
rect 224778 600 225398 668
rect 224778 544 224874 600
rect 224930 544 224998 600
rect 225054 544 225122 600
rect 225178 544 225246 600
rect 225302 544 225398 600
rect 224778 476 225398 544
rect 224778 420 224874 476
rect 224930 420 224998 476
rect 225054 420 225122 476
rect 225178 420 225246 476
rect 225302 420 225398 476
rect 224778 324 225398 420
rect 239058 1808 239678 2326
rect 239058 1752 239154 1808
rect 239210 1752 239278 1808
rect 239334 1752 239402 1808
rect 239458 1752 239526 1808
rect 239582 1752 239678 1808
rect 239058 1684 239678 1752
rect 239058 1628 239154 1684
rect 239210 1628 239278 1684
rect 239334 1628 239402 1684
rect 239458 1628 239526 1684
rect 239582 1628 239678 1684
rect 239058 1560 239678 1628
rect 239058 1504 239154 1560
rect 239210 1504 239278 1560
rect 239334 1504 239402 1560
rect 239458 1504 239526 1560
rect 239582 1504 239678 1560
rect 239058 1436 239678 1504
rect 239058 1380 239154 1436
rect 239210 1380 239278 1436
rect 239334 1380 239402 1436
rect 239458 1380 239526 1436
rect 239582 1380 239678 1436
rect 239058 324 239678 1380
rect 242778 848 243398 2326
rect 242778 792 242874 848
rect 242930 792 242998 848
rect 243054 792 243122 848
rect 243178 792 243246 848
rect 243302 792 243398 848
rect 242778 724 243398 792
rect 242778 668 242874 724
rect 242930 668 242998 724
rect 243054 668 243122 724
rect 243178 668 243246 724
rect 243302 668 243398 724
rect 242778 600 243398 668
rect 242778 544 242874 600
rect 242930 544 242998 600
rect 243054 544 243122 600
rect 243178 544 243246 600
rect 243302 544 243398 600
rect 242778 476 243398 544
rect 242778 420 242874 476
rect 242930 420 242998 476
rect 243054 420 243122 476
rect 243178 420 243246 476
rect 243302 420 243398 476
rect 242778 324 243398 420
rect 257058 1808 257678 2326
rect 257058 1752 257154 1808
rect 257210 1752 257278 1808
rect 257334 1752 257402 1808
rect 257458 1752 257526 1808
rect 257582 1752 257678 1808
rect 257058 1684 257678 1752
rect 257058 1628 257154 1684
rect 257210 1628 257278 1684
rect 257334 1628 257402 1684
rect 257458 1628 257526 1684
rect 257582 1628 257678 1684
rect 257058 1560 257678 1628
rect 257058 1504 257154 1560
rect 257210 1504 257278 1560
rect 257334 1504 257402 1560
rect 257458 1504 257526 1560
rect 257582 1504 257678 1560
rect 257058 1436 257678 1504
rect 257058 1380 257154 1436
rect 257210 1380 257278 1436
rect 257334 1380 257402 1436
rect 257458 1380 257526 1436
rect 257582 1380 257678 1436
rect 257058 324 257678 1380
rect 260778 848 261398 2326
rect 260778 792 260874 848
rect 260930 792 260998 848
rect 261054 792 261122 848
rect 261178 792 261246 848
rect 261302 792 261398 848
rect 260778 724 261398 792
rect 260778 668 260874 724
rect 260930 668 260998 724
rect 261054 668 261122 724
rect 261178 668 261246 724
rect 261302 668 261398 724
rect 260778 600 261398 668
rect 260778 544 260874 600
rect 260930 544 260998 600
rect 261054 544 261122 600
rect 261178 544 261246 600
rect 261302 544 261398 600
rect 260778 476 261398 544
rect 260778 420 260874 476
rect 260930 420 260998 476
rect 261054 420 261122 476
rect 261178 420 261246 476
rect 261302 420 261398 476
rect 260778 324 261398 420
rect 275058 1808 275678 2326
rect 275058 1752 275154 1808
rect 275210 1752 275278 1808
rect 275334 1752 275402 1808
rect 275458 1752 275526 1808
rect 275582 1752 275678 1808
rect 275058 1684 275678 1752
rect 275058 1628 275154 1684
rect 275210 1628 275278 1684
rect 275334 1628 275402 1684
rect 275458 1628 275526 1684
rect 275582 1628 275678 1684
rect 275058 1560 275678 1628
rect 275058 1504 275154 1560
rect 275210 1504 275278 1560
rect 275334 1504 275402 1560
rect 275458 1504 275526 1560
rect 275582 1504 275678 1560
rect 275058 1436 275678 1504
rect 275058 1380 275154 1436
rect 275210 1380 275278 1436
rect 275334 1380 275402 1436
rect 275458 1380 275526 1436
rect 275582 1380 275678 1436
rect 275058 324 275678 1380
rect 278778 848 279398 2326
rect 278778 792 278874 848
rect 278930 792 278998 848
rect 279054 792 279122 848
rect 279178 792 279246 848
rect 279302 792 279398 848
rect 278778 724 279398 792
rect 278778 668 278874 724
rect 278930 668 278998 724
rect 279054 668 279122 724
rect 279178 668 279246 724
rect 279302 668 279398 724
rect 278778 600 279398 668
rect 278778 544 278874 600
rect 278930 544 278998 600
rect 279054 544 279122 600
rect 279178 544 279246 600
rect 279302 544 279398 600
rect 278778 476 279398 544
rect 278778 420 278874 476
rect 278930 420 278998 476
rect 279054 420 279122 476
rect 279178 420 279246 476
rect 279302 420 279398 476
rect 278778 324 279398 420
rect 293058 1808 293678 2326
rect 293058 1752 293154 1808
rect 293210 1752 293278 1808
rect 293334 1752 293402 1808
rect 293458 1752 293526 1808
rect 293582 1752 293678 1808
rect 293058 1684 293678 1752
rect 293058 1628 293154 1684
rect 293210 1628 293278 1684
rect 293334 1628 293402 1684
rect 293458 1628 293526 1684
rect 293582 1628 293678 1684
rect 293058 1560 293678 1628
rect 293058 1504 293154 1560
rect 293210 1504 293278 1560
rect 293334 1504 293402 1560
rect 293458 1504 293526 1560
rect 293582 1504 293678 1560
rect 293058 1436 293678 1504
rect 293058 1380 293154 1436
rect 293210 1380 293278 1436
rect 293334 1380 293402 1436
rect 293458 1380 293526 1436
rect 293582 1380 293678 1436
rect 293058 324 293678 1380
rect 296778 848 297398 2326
rect 296778 792 296874 848
rect 296930 792 296998 848
rect 297054 792 297122 848
rect 297178 792 297246 848
rect 297302 792 297398 848
rect 296778 724 297398 792
rect 296778 668 296874 724
rect 296930 668 296998 724
rect 297054 668 297122 724
rect 297178 668 297246 724
rect 297302 668 297398 724
rect 296778 600 297398 668
rect 296778 544 296874 600
rect 296930 544 296998 600
rect 297054 544 297122 600
rect 297178 544 297246 600
rect 297302 544 297398 600
rect 296778 476 297398 544
rect 296778 420 296874 476
rect 296930 420 296998 476
rect 297054 420 297122 476
rect 297178 420 297246 476
rect 297302 420 297398 476
rect 296778 324 297398 420
rect 311058 1808 311678 2326
rect 311058 1752 311154 1808
rect 311210 1752 311278 1808
rect 311334 1752 311402 1808
rect 311458 1752 311526 1808
rect 311582 1752 311678 1808
rect 311058 1684 311678 1752
rect 311058 1628 311154 1684
rect 311210 1628 311278 1684
rect 311334 1628 311402 1684
rect 311458 1628 311526 1684
rect 311582 1628 311678 1684
rect 311058 1560 311678 1628
rect 311058 1504 311154 1560
rect 311210 1504 311278 1560
rect 311334 1504 311402 1560
rect 311458 1504 311526 1560
rect 311582 1504 311678 1560
rect 311058 1436 311678 1504
rect 311058 1380 311154 1436
rect 311210 1380 311278 1436
rect 311334 1380 311402 1436
rect 311458 1380 311526 1436
rect 311582 1380 311678 1436
rect 311058 324 311678 1380
rect 314778 848 315398 2326
rect 314778 792 314874 848
rect 314930 792 314998 848
rect 315054 792 315122 848
rect 315178 792 315246 848
rect 315302 792 315398 848
rect 314778 724 315398 792
rect 314778 668 314874 724
rect 314930 668 314998 724
rect 315054 668 315122 724
rect 315178 668 315246 724
rect 315302 668 315398 724
rect 314778 600 315398 668
rect 314778 544 314874 600
rect 314930 544 314998 600
rect 315054 544 315122 600
rect 315178 544 315246 600
rect 315302 544 315398 600
rect 314778 476 315398 544
rect 314778 420 314874 476
rect 314930 420 314998 476
rect 315054 420 315122 476
rect 315178 420 315246 476
rect 315302 420 315398 476
rect 314778 324 315398 420
rect 329058 1808 329678 2326
rect 329058 1752 329154 1808
rect 329210 1752 329278 1808
rect 329334 1752 329402 1808
rect 329458 1752 329526 1808
rect 329582 1752 329678 1808
rect 329058 1684 329678 1752
rect 329058 1628 329154 1684
rect 329210 1628 329278 1684
rect 329334 1628 329402 1684
rect 329458 1628 329526 1684
rect 329582 1628 329678 1684
rect 329058 1560 329678 1628
rect 329058 1504 329154 1560
rect 329210 1504 329278 1560
rect 329334 1504 329402 1560
rect 329458 1504 329526 1560
rect 329582 1504 329678 1560
rect 329058 1436 329678 1504
rect 329058 1380 329154 1436
rect 329210 1380 329278 1436
rect 329334 1380 329402 1436
rect 329458 1380 329526 1436
rect 329582 1380 329678 1436
rect 329058 324 329678 1380
rect 332778 848 333398 2326
rect 332778 792 332874 848
rect 332930 792 332998 848
rect 333054 792 333122 848
rect 333178 792 333246 848
rect 333302 792 333398 848
rect 332778 724 333398 792
rect 332778 668 332874 724
rect 332930 668 332998 724
rect 333054 668 333122 724
rect 333178 668 333246 724
rect 333302 668 333398 724
rect 332778 600 333398 668
rect 332778 544 332874 600
rect 332930 544 332998 600
rect 333054 544 333122 600
rect 333178 544 333246 600
rect 333302 544 333398 600
rect 332778 476 333398 544
rect 332778 420 332874 476
rect 332930 420 332998 476
rect 333054 420 333122 476
rect 333178 420 333246 476
rect 333302 420 333398 476
rect 332778 324 333398 420
rect 347058 1808 347678 2326
rect 347058 1752 347154 1808
rect 347210 1752 347278 1808
rect 347334 1752 347402 1808
rect 347458 1752 347526 1808
rect 347582 1752 347678 1808
rect 347058 1684 347678 1752
rect 347058 1628 347154 1684
rect 347210 1628 347278 1684
rect 347334 1628 347402 1684
rect 347458 1628 347526 1684
rect 347582 1628 347678 1684
rect 347058 1560 347678 1628
rect 347058 1504 347154 1560
rect 347210 1504 347278 1560
rect 347334 1504 347402 1560
rect 347458 1504 347526 1560
rect 347582 1504 347678 1560
rect 347058 1436 347678 1504
rect 347058 1380 347154 1436
rect 347210 1380 347278 1436
rect 347334 1380 347402 1436
rect 347458 1380 347526 1436
rect 347582 1380 347678 1436
rect 347058 324 347678 1380
rect 350778 848 351398 2326
rect 350778 792 350874 848
rect 350930 792 350998 848
rect 351054 792 351122 848
rect 351178 792 351246 848
rect 351302 792 351398 848
rect 350778 724 351398 792
rect 350778 668 350874 724
rect 350930 668 350998 724
rect 351054 668 351122 724
rect 351178 668 351246 724
rect 351302 668 351398 724
rect 350778 600 351398 668
rect 350778 544 350874 600
rect 350930 544 350998 600
rect 351054 544 351122 600
rect 351178 544 351246 600
rect 351302 544 351398 600
rect 350778 476 351398 544
rect 350778 420 350874 476
rect 350930 420 350998 476
rect 351054 420 351122 476
rect 351178 420 351246 476
rect 351302 420 351398 476
rect 350778 324 351398 420
rect 365058 1808 365678 2326
rect 365058 1752 365154 1808
rect 365210 1752 365278 1808
rect 365334 1752 365402 1808
rect 365458 1752 365526 1808
rect 365582 1752 365678 1808
rect 365058 1684 365678 1752
rect 365058 1628 365154 1684
rect 365210 1628 365278 1684
rect 365334 1628 365402 1684
rect 365458 1628 365526 1684
rect 365582 1628 365678 1684
rect 365058 1560 365678 1628
rect 365058 1504 365154 1560
rect 365210 1504 365278 1560
rect 365334 1504 365402 1560
rect 365458 1504 365526 1560
rect 365582 1504 365678 1560
rect 365058 1436 365678 1504
rect 365058 1380 365154 1436
rect 365210 1380 365278 1436
rect 365334 1380 365402 1436
rect 365458 1380 365526 1436
rect 365582 1380 365678 1436
rect 365058 324 365678 1380
rect 368778 848 369398 2326
rect 368778 792 368874 848
rect 368930 792 368998 848
rect 369054 792 369122 848
rect 369178 792 369246 848
rect 369302 792 369398 848
rect 368778 724 369398 792
rect 368778 668 368874 724
rect 368930 668 368998 724
rect 369054 668 369122 724
rect 369178 668 369246 724
rect 369302 668 369398 724
rect 368778 600 369398 668
rect 368778 544 368874 600
rect 368930 544 368998 600
rect 369054 544 369122 600
rect 369178 544 369246 600
rect 369302 544 369398 600
rect 368778 476 369398 544
rect 368778 420 368874 476
rect 368930 420 368998 476
rect 369054 420 369122 476
rect 369178 420 369246 476
rect 369302 420 369398 476
rect 368778 324 369398 420
rect 383058 1808 383678 2326
rect 383058 1752 383154 1808
rect 383210 1752 383278 1808
rect 383334 1752 383402 1808
rect 383458 1752 383526 1808
rect 383582 1752 383678 1808
rect 383058 1684 383678 1752
rect 383058 1628 383154 1684
rect 383210 1628 383278 1684
rect 383334 1628 383402 1684
rect 383458 1628 383526 1684
rect 383582 1628 383678 1684
rect 383058 1560 383678 1628
rect 383058 1504 383154 1560
rect 383210 1504 383278 1560
rect 383334 1504 383402 1560
rect 383458 1504 383526 1560
rect 383582 1504 383678 1560
rect 383058 1436 383678 1504
rect 383058 1380 383154 1436
rect 383210 1380 383278 1436
rect 383334 1380 383402 1436
rect 383458 1380 383526 1436
rect 383582 1380 383678 1436
rect 383058 324 383678 1380
rect 386778 848 387398 2326
rect 386778 792 386874 848
rect 386930 792 386998 848
rect 387054 792 387122 848
rect 387178 792 387246 848
rect 387302 792 387398 848
rect 386778 724 387398 792
rect 386778 668 386874 724
rect 386930 668 386998 724
rect 387054 668 387122 724
rect 387178 668 387246 724
rect 387302 668 387398 724
rect 386778 600 387398 668
rect 386778 544 386874 600
rect 386930 544 386998 600
rect 387054 544 387122 600
rect 387178 544 387246 600
rect 387302 544 387398 600
rect 386778 476 387398 544
rect 386778 420 386874 476
rect 386930 420 386998 476
rect 387054 420 387122 476
rect 387178 420 387246 476
rect 387302 420 387398 476
rect 386778 324 387398 420
rect 401058 1808 401678 2326
rect 401058 1752 401154 1808
rect 401210 1752 401278 1808
rect 401334 1752 401402 1808
rect 401458 1752 401526 1808
rect 401582 1752 401678 1808
rect 401058 1684 401678 1752
rect 401058 1628 401154 1684
rect 401210 1628 401278 1684
rect 401334 1628 401402 1684
rect 401458 1628 401526 1684
rect 401582 1628 401678 1684
rect 401058 1560 401678 1628
rect 401058 1504 401154 1560
rect 401210 1504 401278 1560
rect 401334 1504 401402 1560
rect 401458 1504 401526 1560
rect 401582 1504 401678 1560
rect 401058 1436 401678 1504
rect 401058 1380 401154 1436
rect 401210 1380 401278 1436
rect 401334 1380 401402 1436
rect 401458 1380 401526 1436
rect 401582 1380 401678 1436
rect 401058 324 401678 1380
rect 404778 848 405398 2326
rect 404778 792 404874 848
rect 404930 792 404998 848
rect 405054 792 405122 848
rect 405178 792 405246 848
rect 405302 792 405398 848
rect 404778 724 405398 792
rect 404778 668 404874 724
rect 404930 668 404998 724
rect 405054 668 405122 724
rect 405178 668 405246 724
rect 405302 668 405398 724
rect 404778 600 405398 668
rect 404778 544 404874 600
rect 404930 544 404998 600
rect 405054 544 405122 600
rect 405178 544 405246 600
rect 405302 544 405398 600
rect 404778 476 405398 544
rect 404778 420 404874 476
rect 404930 420 404998 476
rect 405054 420 405122 476
rect 405178 420 405246 476
rect 405302 420 405398 476
rect 404778 324 405398 420
rect 419058 1808 419678 2326
rect 419058 1752 419154 1808
rect 419210 1752 419278 1808
rect 419334 1752 419402 1808
rect 419458 1752 419526 1808
rect 419582 1752 419678 1808
rect 419058 1684 419678 1752
rect 419058 1628 419154 1684
rect 419210 1628 419278 1684
rect 419334 1628 419402 1684
rect 419458 1628 419526 1684
rect 419582 1628 419678 1684
rect 419058 1560 419678 1628
rect 419058 1504 419154 1560
rect 419210 1504 419278 1560
rect 419334 1504 419402 1560
rect 419458 1504 419526 1560
rect 419582 1504 419678 1560
rect 419058 1436 419678 1504
rect 419058 1380 419154 1436
rect 419210 1380 419278 1436
rect 419334 1380 419402 1436
rect 419458 1380 419526 1436
rect 419582 1380 419678 1436
rect 419058 324 419678 1380
rect 422778 848 423398 2326
rect 422778 792 422874 848
rect 422930 792 422998 848
rect 423054 792 423122 848
rect 423178 792 423246 848
rect 423302 792 423398 848
rect 422778 724 423398 792
rect 422778 668 422874 724
rect 422930 668 422998 724
rect 423054 668 423122 724
rect 423178 668 423246 724
rect 423302 668 423398 724
rect 422778 600 423398 668
rect 422778 544 422874 600
rect 422930 544 422998 600
rect 423054 544 423122 600
rect 423178 544 423246 600
rect 423302 544 423398 600
rect 422778 476 423398 544
rect 422778 420 422874 476
rect 422930 420 422998 476
rect 423054 420 423122 476
rect 423178 420 423246 476
rect 423302 420 423398 476
rect 422778 324 423398 420
rect 437058 1808 437678 2326
rect 437058 1752 437154 1808
rect 437210 1752 437278 1808
rect 437334 1752 437402 1808
rect 437458 1752 437526 1808
rect 437582 1752 437678 1808
rect 437058 1684 437678 1752
rect 437058 1628 437154 1684
rect 437210 1628 437278 1684
rect 437334 1628 437402 1684
rect 437458 1628 437526 1684
rect 437582 1628 437678 1684
rect 437058 1560 437678 1628
rect 437058 1504 437154 1560
rect 437210 1504 437278 1560
rect 437334 1504 437402 1560
rect 437458 1504 437526 1560
rect 437582 1504 437678 1560
rect 437058 1436 437678 1504
rect 437058 1380 437154 1436
rect 437210 1380 437278 1436
rect 437334 1380 437402 1436
rect 437458 1380 437526 1436
rect 437582 1380 437678 1436
rect 437058 324 437678 1380
rect 440778 848 441398 2326
rect 440778 792 440874 848
rect 440930 792 440998 848
rect 441054 792 441122 848
rect 441178 792 441246 848
rect 441302 792 441398 848
rect 440778 724 441398 792
rect 440778 668 440874 724
rect 440930 668 440998 724
rect 441054 668 441122 724
rect 441178 668 441246 724
rect 441302 668 441398 724
rect 440778 600 441398 668
rect 440778 544 440874 600
rect 440930 544 440998 600
rect 441054 544 441122 600
rect 441178 544 441246 600
rect 441302 544 441398 600
rect 440778 476 441398 544
rect 440778 420 440874 476
rect 440930 420 440998 476
rect 441054 420 441122 476
rect 441178 420 441246 476
rect 441302 420 441398 476
rect 440778 324 441398 420
rect 455058 1808 455678 2326
rect 455058 1752 455154 1808
rect 455210 1752 455278 1808
rect 455334 1752 455402 1808
rect 455458 1752 455526 1808
rect 455582 1752 455678 1808
rect 455058 1684 455678 1752
rect 455058 1628 455154 1684
rect 455210 1628 455278 1684
rect 455334 1628 455402 1684
rect 455458 1628 455526 1684
rect 455582 1628 455678 1684
rect 455058 1560 455678 1628
rect 455058 1504 455154 1560
rect 455210 1504 455278 1560
rect 455334 1504 455402 1560
rect 455458 1504 455526 1560
rect 455582 1504 455678 1560
rect 455058 1436 455678 1504
rect 455058 1380 455154 1436
rect 455210 1380 455278 1436
rect 455334 1380 455402 1436
rect 455458 1380 455526 1436
rect 455582 1380 455678 1436
rect 455058 324 455678 1380
rect 458778 848 459398 2326
rect 458778 792 458874 848
rect 458930 792 458998 848
rect 459054 792 459122 848
rect 459178 792 459246 848
rect 459302 792 459398 848
rect 458778 724 459398 792
rect 458778 668 458874 724
rect 458930 668 458998 724
rect 459054 668 459122 724
rect 459178 668 459246 724
rect 459302 668 459398 724
rect 458778 600 459398 668
rect 458778 544 458874 600
rect 458930 544 458998 600
rect 459054 544 459122 600
rect 459178 544 459246 600
rect 459302 544 459398 600
rect 458778 476 459398 544
rect 458778 420 458874 476
rect 458930 420 458998 476
rect 459054 420 459122 476
rect 459178 420 459246 476
rect 459302 420 459398 476
rect 458778 324 459398 420
rect 473058 1808 473678 2326
rect 473058 1752 473154 1808
rect 473210 1752 473278 1808
rect 473334 1752 473402 1808
rect 473458 1752 473526 1808
rect 473582 1752 473678 1808
rect 473058 1684 473678 1752
rect 473058 1628 473154 1684
rect 473210 1628 473278 1684
rect 473334 1628 473402 1684
rect 473458 1628 473526 1684
rect 473582 1628 473678 1684
rect 473058 1560 473678 1628
rect 473058 1504 473154 1560
rect 473210 1504 473278 1560
rect 473334 1504 473402 1560
rect 473458 1504 473526 1560
rect 473582 1504 473678 1560
rect 473058 1436 473678 1504
rect 473058 1380 473154 1436
rect 473210 1380 473278 1436
rect 473334 1380 473402 1436
rect 473458 1380 473526 1436
rect 473582 1380 473678 1436
rect 473058 324 473678 1380
rect 476778 848 477398 2326
rect 476778 792 476874 848
rect 476930 792 476998 848
rect 477054 792 477122 848
rect 477178 792 477246 848
rect 477302 792 477398 848
rect 476778 724 477398 792
rect 476778 668 476874 724
rect 476930 668 476998 724
rect 477054 668 477122 724
rect 477178 668 477246 724
rect 477302 668 477398 724
rect 476778 600 477398 668
rect 476778 544 476874 600
rect 476930 544 476998 600
rect 477054 544 477122 600
rect 477178 544 477246 600
rect 477302 544 477398 600
rect 476778 476 477398 544
rect 476778 420 476874 476
rect 476930 420 476998 476
rect 477054 420 477122 476
rect 477178 420 477246 476
rect 477302 420 477398 476
rect 476778 324 477398 420
rect 491058 1808 491678 2326
rect 491058 1752 491154 1808
rect 491210 1752 491278 1808
rect 491334 1752 491402 1808
rect 491458 1752 491526 1808
rect 491582 1752 491678 1808
rect 491058 1684 491678 1752
rect 491058 1628 491154 1684
rect 491210 1628 491278 1684
rect 491334 1628 491402 1684
rect 491458 1628 491526 1684
rect 491582 1628 491678 1684
rect 491058 1560 491678 1628
rect 491058 1504 491154 1560
rect 491210 1504 491278 1560
rect 491334 1504 491402 1560
rect 491458 1504 491526 1560
rect 491582 1504 491678 1560
rect 491058 1436 491678 1504
rect 491058 1380 491154 1436
rect 491210 1380 491278 1436
rect 491334 1380 491402 1436
rect 491458 1380 491526 1436
rect 491582 1380 491678 1436
rect 491058 324 491678 1380
rect 494778 848 495398 2326
rect 494778 792 494874 848
rect 494930 792 494998 848
rect 495054 792 495122 848
rect 495178 792 495246 848
rect 495302 792 495398 848
rect 494778 724 495398 792
rect 494778 668 494874 724
rect 494930 668 494998 724
rect 495054 668 495122 724
rect 495178 668 495246 724
rect 495302 668 495398 724
rect 494778 600 495398 668
rect 494778 544 494874 600
rect 494930 544 494998 600
rect 495054 544 495122 600
rect 495178 544 495246 600
rect 495302 544 495398 600
rect 494778 476 495398 544
rect 494778 420 494874 476
rect 494930 420 494998 476
rect 495054 420 495122 476
rect 495178 420 495246 476
rect 495302 420 495398 476
rect 494778 324 495398 420
rect 509058 1808 509678 2326
rect 509058 1752 509154 1808
rect 509210 1752 509278 1808
rect 509334 1752 509402 1808
rect 509458 1752 509526 1808
rect 509582 1752 509678 1808
rect 509058 1684 509678 1752
rect 509058 1628 509154 1684
rect 509210 1628 509278 1684
rect 509334 1628 509402 1684
rect 509458 1628 509526 1684
rect 509582 1628 509678 1684
rect 509058 1560 509678 1628
rect 509058 1504 509154 1560
rect 509210 1504 509278 1560
rect 509334 1504 509402 1560
rect 509458 1504 509526 1560
rect 509582 1504 509678 1560
rect 509058 1436 509678 1504
rect 509058 1380 509154 1436
rect 509210 1380 509278 1436
rect 509334 1380 509402 1436
rect 509458 1380 509526 1436
rect 509582 1380 509678 1436
rect 509058 324 509678 1380
rect 512778 848 513398 2326
rect 512778 792 512874 848
rect 512930 792 512998 848
rect 513054 792 513122 848
rect 513178 792 513246 848
rect 513302 792 513398 848
rect 512778 724 513398 792
rect 512778 668 512874 724
rect 512930 668 512998 724
rect 513054 668 513122 724
rect 513178 668 513246 724
rect 513302 668 513398 724
rect 512778 600 513398 668
rect 512778 544 512874 600
rect 512930 544 512998 600
rect 513054 544 513122 600
rect 513178 544 513246 600
rect 513302 544 513398 600
rect 512778 476 513398 544
rect 512778 420 512874 476
rect 512930 420 512998 476
rect 513054 420 513122 476
rect 513178 420 513246 476
rect 513302 420 513398 476
rect 512778 324 513398 420
rect 527058 1808 527678 2326
rect 527058 1752 527154 1808
rect 527210 1752 527278 1808
rect 527334 1752 527402 1808
rect 527458 1752 527526 1808
rect 527582 1752 527678 1808
rect 527058 1684 527678 1752
rect 527058 1628 527154 1684
rect 527210 1628 527278 1684
rect 527334 1628 527402 1684
rect 527458 1628 527526 1684
rect 527582 1628 527678 1684
rect 527058 1560 527678 1628
rect 527058 1504 527154 1560
rect 527210 1504 527278 1560
rect 527334 1504 527402 1560
rect 527458 1504 527526 1560
rect 527582 1504 527678 1560
rect 527058 1436 527678 1504
rect 527058 1380 527154 1436
rect 527210 1380 527278 1436
rect 527334 1380 527402 1436
rect 527458 1380 527526 1436
rect 527582 1380 527678 1436
rect 527058 324 527678 1380
rect 530778 848 531398 2326
rect 530778 792 530874 848
rect 530930 792 530998 848
rect 531054 792 531122 848
rect 531178 792 531246 848
rect 531302 792 531398 848
rect 530778 724 531398 792
rect 530778 668 530874 724
rect 530930 668 530998 724
rect 531054 668 531122 724
rect 531178 668 531246 724
rect 531302 668 531398 724
rect 530778 600 531398 668
rect 530778 544 530874 600
rect 530930 544 530998 600
rect 531054 544 531122 600
rect 531178 544 531246 600
rect 531302 544 531398 600
rect 530778 476 531398 544
rect 530778 420 530874 476
rect 530930 420 530998 476
rect 531054 420 531122 476
rect 531178 420 531246 476
rect 531302 420 531398 476
rect 530778 324 531398 420
rect 545058 1808 545678 2326
rect 545058 1752 545154 1808
rect 545210 1752 545278 1808
rect 545334 1752 545402 1808
rect 545458 1752 545526 1808
rect 545582 1752 545678 1808
rect 545058 1684 545678 1752
rect 545058 1628 545154 1684
rect 545210 1628 545278 1684
rect 545334 1628 545402 1684
rect 545458 1628 545526 1684
rect 545582 1628 545678 1684
rect 545058 1560 545678 1628
rect 545058 1504 545154 1560
rect 545210 1504 545278 1560
rect 545334 1504 545402 1560
rect 545458 1504 545526 1560
rect 545582 1504 545678 1560
rect 545058 1436 545678 1504
rect 545058 1380 545154 1436
rect 545210 1380 545278 1436
rect 545334 1380 545402 1436
rect 545458 1380 545526 1436
rect 545582 1380 545678 1436
rect 545058 324 545678 1380
rect 548778 848 549398 2326
rect 548778 792 548874 848
rect 548930 792 548998 848
rect 549054 792 549122 848
rect 549178 792 549246 848
rect 549302 792 549398 848
rect 548778 724 549398 792
rect 548778 668 548874 724
rect 548930 668 548998 724
rect 549054 668 549122 724
rect 549178 668 549246 724
rect 549302 668 549398 724
rect 548778 600 549398 668
rect 548778 544 548874 600
rect 548930 544 548998 600
rect 549054 544 549122 600
rect 549178 544 549246 600
rect 549302 544 549398 600
rect 548778 476 549398 544
rect 548778 420 548874 476
rect 548930 420 548998 476
rect 549054 420 549122 476
rect 549178 420 549246 476
rect 549302 420 549398 476
rect 548778 324 549398 420
rect 563058 1808 563678 2326
rect 563058 1752 563154 1808
rect 563210 1752 563278 1808
rect 563334 1752 563402 1808
rect 563458 1752 563526 1808
rect 563582 1752 563678 1808
rect 563058 1684 563678 1752
rect 563058 1628 563154 1684
rect 563210 1628 563278 1684
rect 563334 1628 563402 1684
rect 563458 1628 563526 1684
rect 563582 1628 563678 1684
rect 563058 1560 563678 1628
rect 563058 1504 563154 1560
rect 563210 1504 563278 1560
rect 563334 1504 563402 1560
rect 563458 1504 563526 1560
rect 563582 1504 563678 1560
rect 563058 1436 563678 1504
rect 563058 1380 563154 1436
rect 563210 1380 563278 1436
rect 563334 1380 563402 1436
rect 563458 1380 563526 1436
rect 563582 1380 563678 1436
rect 563058 324 563678 1380
rect 566778 848 567398 2326
rect 566778 792 566874 848
rect 566930 792 566998 848
rect 567054 792 567122 848
rect 567178 792 567246 848
rect 567302 792 567398 848
rect 566778 724 567398 792
rect 566778 668 566874 724
rect 566930 668 566998 724
rect 567054 668 567122 724
rect 567178 668 567246 724
rect 567302 668 567398 724
rect 566778 600 567398 668
rect 566778 544 566874 600
rect 566930 544 566998 600
rect 567054 544 567122 600
rect 567178 544 567246 600
rect 567302 544 567398 600
rect 566778 476 567398 544
rect 566778 420 566874 476
rect 566930 420 566998 476
rect 567054 420 567122 476
rect 567178 420 567246 476
rect 567302 420 567398 476
rect 566778 324 567398 420
rect 581058 1808 581678 2326
rect 581058 1752 581154 1808
rect 581210 1752 581278 1808
rect 581334 1752 581402 1808
rect 581458 1752 581526 1808
rect 581582 1752 581678 1808
rect 581058 1684 581678 1752
rect 581058 1628 581154 1684
rect 581210 1628 581278 1684
rect 581334 1628 581402 1684
rect 581458 1628 581526 1684
rect 581582 1628 581678 1684
rect 581058 1560 581678 1628
rect 581058 1504 581154 1560
rect 581210 1504 581278 1560
rect 581334 1504 581402 1560
rect 581458 1504 581526 1560
rect 581582 1504 581678 1560
rect 581058 1436 581678 1504
rect 581058 1380 581154 1436
rect 581210 1380 581278 1436
rect 581334 1380 581402 1436
rect 581458 1380 581526 1436
rect 581582 1380 581678 1436
rect 581058 324 581678 1380
rect 584778 848 585398 2326
rect 598416 1808 599036 5490
rect 598416 1752 598512 1808
rect 598568 1752 598636 1808
rect 598692 1752 598760 1808
rect 598816 1752 598884 1808
rect 598940 1752 599036 1808
rect 598416 1684 599036 1752
rect 598416 1628 598512 1684
rect 598568 1628 598636 1684
rect 598692 1628 598760 1684
rect 598816 1628 598884 1684
rect 598940 1628 599036 1684
rect 598416 1560 599036 1628
rect 598416 1504 598512 1560
rect 598568 1504 598636 1560
rect 598692 1504 598760 1560
rect 598816 1504 598884 1560
rect 598940 1504 599036 1560
rect 598416 1436 599036 1504
rect 598416 1380 598512 1436
rect 598568 1380 598636 1436
rect 598692 1380 598760 1436
rect 598816 1380 598884 1436
rect 598940 1380 599036 1436
rect 598416 1284 599036 1380
rect 599376 587918 599996 598912
rect 599376 587862 599472 587918
rect 599528 587862 599596 587918
rect 599652 587862 599720 587918
rect 599776 587862 599844 587918
rect 599900 587862 599996 587918
rect 599376 587794 599996 587862
rect 599376 587738 599472 587794
rect 599528 587738 599596 587794
rect 599652 587738 599720 587794
rect 599776 587738 599844 587794
rect 599900 587738 599996 587794
rect 599376 587670 599996 587738
rect 599376 587614 599472 587670
rect 599528 587614 599596 587670
rect 599652 587614 599720 587670
rect 599776 587614 599844 587670
rect 599900 587614 599996 587670
rect 599376 587546 599996 587614
rect 599376 587490 599472 587546
rect 599528 587490 599596 587546
rect 599652 587490 599720 587546
rect 599776 587490 599844 587546
rect 599900 587490 599996 587546
rect 599376 569918 599996 587490
rect 599376 569862 599472 569918
rect 599528 569862 599596 569918
rect 599652 569862 599720 569918
rect 599776 569862 599844 569918
rect 599900 569862 599996 569918
rect 599376 569794 599996 569862
rect 599376 569738 599472 569794
rect 599528 569738 599596 569794
rect 599652 569738 599720 569794
rect 599776 569738 599844 569794
rect 599900 569738 599996 569794
rect 599376 569670 599996 569738
rect 599376 569614 599472 569670
rect 599528 569614 599596 569670
rect 599652 569614 599720 569670
rect 599776 569614 599844 569670
rect 599900 569614 599996 569670
rect 599376 569546 599996 569614
rect 599376 569490 599472 569546
rect 599528 569490 599596 569546
rect 599652 569490 599720 569546
rect 599776 569490 599844 569546
rect 599900 569490 599996 569546
rect 599376 551918 599996 569490
rect 599376 551862 599472 551918
rect 599528 551862 599596 551918
rect 599652 551862 599720 551918
rect 599776 551862 599844 551918
rect 599900 551862 599996 551918
rect 599376 551794 599996 551862
rect 599376 551738 599472 551794
rect 599528 551738 599596 551794
rect 599652 551738 599720 551794
rect 599776 551738 599844 551794
rect 599900 551738 599996 551794
rect 599376 551670 599996 551738
rect 599376 551614 599472 551670
rect 599528 551614 599596 551670
rect 599652 551614 599720 551670
rect 599776 551614 599844 551670
rect 599900 551614 599996 551670
rect 599376 551546 599996 551614
rect 599376 551490 599472 551546
rect 599528 551490 599596 551546
rect 599652 551490 599720 551546
rect 599776 551490 599844 551546
rect 599900 551490 599996 551546
rect 599376 533918 599996 551490
rect 599376 533862 599472 533918
rect 599528 533862 599596 533918
rect 599652 533862 599720 533918
rect 599776 533862 599844 533918
rect 599900 533862 599996 533918
rect 599376 533794 599996 533862
rect 599376 533738 599472 533794
rect 599528 533738 599596 533794
rect 599652 533738 599720 533794
rect 599776 533738 599844 533794
rect 599900 533738 599996 533794
rect 599376 533670 599996 533738
rect 599376 533614 599472 533670
rect 599528 533614 599596 533670
rect 599652 533614 599720 533670
rect 599776 533614 599844 533670
rect 599900 533614 599996 533670
rect 599376 533546 599996 533614
rect 599376 533490 599472 533546
rect 599528 533490 599596 533546
rect 599652 533490 599720 533546
rect 599776 533490 599844 533546
rect 599900 533490 599996 533546
rect 599376 515918 599996 533490
rect 599376 515862 599472 515918
rect 599528 515862 599596 515918
rect 599652 515862 599720 515918
rect 599776 515862 599844 515918
rect 599900 515862 599996 515918
rect 599376 515794 599996 515862
rect 599376 515738 599472 515794
rect 599528 515738 599596 515794
rect 599652 515738 599720 515794
rect 599776 515738 599844 515794
rect 599900 515738 599996 515794
rect 599376 515670 599996 515738
rect 599376 515614 599472 515670
rect 599528 515614 599596 515670
rect 599652 515614 599720 515670
rect 599776 515614 599844 515670
rect 599900 515614 599996 515670
rect 599376 515546 599996 515614
rect 599376 515490 599472 515546
rect 599528 515490 599596 515546
rect 599652 515490 599720 515546
rect 599776 515490 599844 515546
rect 599900 515490 599996 515546
rect 599376 497918 599996 515490
rect 599376 497862 599472 497918
rect 599528 497862 599596 497918
rect 599652 497862 599720 497918
rect 599776 497862 599844 497918
rect 599900 497862 599996 497918
rect 599376 497794 599996 497862
rect 599376 497738 599472 497794
rect 599528 497738 599596 497794
rect 599652 497738 599720 497794
rect 599776 497738 599844 497794
rect 599900 497738 599996 497794
rect 599376 497670 599996 497738
rect 599376 497614 599472 497670
rect 599528 497614 599596 497670
rect 599652 497614 599720 497670
rect 599776 497614 599844 497670
rect 599900 497614 599996 497670
rect 599376 497546 599996 497614
rect 599376 497490 599472 497546
rect 599528 497490 599596 497546
rect 599652 497490 599720 497546
rect 599776 497490 599844 497546
rect 599900 497490 599996 497546
rect 599376 479918 599996 497490
rect 599376 479862 599472 479918
rect 599528 479862 599596 479918
rect 599652 479862 599720 479918
rect 599776 479862 599844 479918
rect 599900 479862 599996 479918
rect 599376 479794 599996 479862
rect 599376 479738 599472 479794
rect 599528 479738 599596 479794
rect 599652 479738 599720 479794
rect 599776 479738 599844 479794
rect 599900 479738 599996 479794
rect 599376 479670 599996 479738
rect 599376 479614 599472 479670
rect 599528 479614 599596 479670
rect 599652 479614 599720 479670
rect 599776 479614 599844 479670
rect 599900 479614 599996 479670
rect 599376 479546 599996 479614
rect 599376 479490 599472 479546
rect 599528 479490 599596 479546
rect 599652 479490 599720 479546
rect 599776 479490 599844 479546
rect 599900 479490 599996 479546
rect 599376 461918 599996 479490
rect 599376 461862 599472 461918
rect 599528 461862 599596 461918
rect 599652 461862 599720 461918
rect 599776 461862 599844 461918
rect 599900 461862 599996 461918
rect 599376 461794 599996 461862
rect 599376 461738 599472 461794
rect 599528 461738 599596 461794
rect 599652 461738 599720 461794
rect 599776 461738 599844 461794
rect 599900 461738 599996 461794
rect 599376 461670 599996 461738
rect 599376 461614 599472 461670
rect 599528 461614 599596 461670
rect 599652 461614 599720 461670
rect 599776 461614 599844 461670
rect 599900 461614 599996 461670
rect 599376 461546 599996 461614
rect 599376 461490 599472 461546
rect 599528 461490 599596 461546
rect 599652 461490 599720 461546
rect 599776 461490 599844 461546
rect 599900 461490 599996 461546
rect 599376 443918 599996 461490
rect 599376 443862 599472 443918
rect 599528 443862 599596 443918
rect 599652 443862 599720 443918
rect 599776 443862 599844 443918
rect 599900 443862 599996 443918
rect 599376 443794 599996 443862
rect 599376 443738 599472 443794
rect 599528 443738 599596 443794
rect 599652 443738 599720 443794
rect 599776 443738 599844 443794
rect 599900 443738 599996 443794
rect 599376 443670 599996 443738
rect 599376 443614 599472 443670
rect 599528 443614 599596 443670
rect 599652 443614 599720 443670
rect 599776 443614 599844 443670
rect 599900 443614 599996 443670
rect 599376 443546 599996 443614
rect 599376 443490 599472 443546
rect 599528 443490 599596 443546
rect 599652 443490 599720 443546
rect 599776 443490 599844 443546
rect 599900 443490 599996 443546
rect 599376 425918 599996 443490
rect 599376 425862 599472 425918
rect 599528 425862 599596 425918
rect 599652 425862 599720 425918
rect 599776 425862 599844 425918
rect 599900 425862 599996 425918
rect 599376 425794 599996 425862
rect 599376 425738 599472 425794
rect 599528 425738 599596 425794
rect 599652 425738 599720 425794
rect 599776 425738 599844 425794
rect 599900 425738 599996 425794
rect 599376 425670 599996 425738
rect 599376 425614 599472 425670
rect 599528 425614 599596 425670
rect 599652 425614 599720 425670
rect 599776 425614 599844 425670
rect 599900 425614 599996 425670
rect 599376 425546 599996 425614
rect 599376 425490 599472 425546
rect 599528 425490 599596 425546
rect 599652 425490 599720 425546
rect 599776 425490 599844 425546
rect 599900 425490 599996 425546
rect 599376 407918 599996 425490
rect 599376 407862 599472 407918
rect 599528 407862 599596 407918
rect 599652 407862 599720 407918
rect 599776 407862 599844 407918
rect 599900 407862 599996 407918
rect 599376 407794 599996 407862
rect 599376 407738 599472 407794
rect 599528 407738 599596 407794
rect 599652 407738 599720 407794
rect 599776 407738 599844 407794
rect 599900 407738 599996 407794
rect 599376 407670 599996 407738
rect 599376 407614 599472 407670
rect 599528 407614 599596 407670
rect 599652 407614 599720 407670
rect 599776 407614 599844 407670
rect 599900 407614 599996 407670
rect 599376 407546 599996 407614
rect 599376 407490 599472 407546
rect 599528 407490 599596 407546
rect 599652 407490 599720 407546
rect 599776 407490 599844 407546
rect 599900 407490 599996 407546
rect 599376 389918 599996 407490
rect 599376 389862 599472 389918
rect 599528 389862 599596 389918
rect 599652 389862 599720 389918
rect 599776 389862 599844 389918
rect 599900 389862 599996 389918
rect 599376 389794 599996 389862
rect 599376 389738 599472 389794
rect 599528 389738 599596 389794
rect 599652 389738 599720 389794
rect 599776 389738 599844 389794
rect 599900 389738 599996 389794
rect 599376 389670 599996 389738
rect 599376 389614 599472 389670
rect 599528 389614 599596 389670
rect 599652 389614 599720 389670
rect 599776 389614 599844 389670
rect 599900 389614 599996 389670
rect 599376 389546 599996 389614
rect 599376 389490 599472 389546
rect 599528 389490 599596 389546
rect 599652 389490 599720 389546
rect 599776 389490 599844 389546
rect 599900 389490 599996 389546
rect 599376 371918 599996 389490
rect 599376 371862 599472 371918
rect 599528 371862 599596 371918
rect 599652 371862 599720 371918
rect 599776 371862 599844 371918
rect 599900 371862 599996 371918
rect 599376 371794 599996 371862
rect 599376 371738 599472 371794
rect 599528 371738 599596 371794
rect 599652 371738 599720 371794
rect 599776 371738 599844 371794
rect 599900 371738 599996 371794
rect 599376 371670 599996 371738
rect 599376 371614 599472 371670
rect 599528 371614 599596 371670
rect 599652 371614 599720 371670
rect 599776 371614 599844 371670
rect 599900 371614 599996 371670
rect 599376 371546 599996 371614
rect 599376 371490 599472 371546
rect 599528 371490 599596 371546
rect 599652 371490 599720 371546
rect 599776 371490 599844 371546
rect 599900 371490 599996 371546
rect 599376 353918 599996 371490
rect 599376 353862 599472 353918
rect 599528 353862 599596 353918
rect 599652 353862 599720 353918
rect 599776 353862 599844 353918
rect 599900 353862 599996 353918
rect 599376 353794 599996 353862
rect 599376 353738 599472 353794
rect 599528 353738 599596 353794
rect 599652 353738 599720 353794
rect 599776 353738 599844 353794
rect 599900 353738 599996 353794
rect 599376 353670 599996 353738
rect 599376 353614 599472 353670
rect 599528 353614 599596 353670
rect 599652 353614 599720 353670
rect 599776 353614 599844 353670
rect 599900 353614 599996 353670
rect 599376 353546 599996 353614
rect 599376 353490 599472 353546
rect 599528 353490 599596 353546
rect 599652 353490 599720 353546
rect 599776 353490 599844 353546
rect 599900 353490 599996 353546
rect 599376 335918 599996 353490
rect 599376 335862 599472 335918
rect 599528 335862 599596 335918
rect 599652 335862 599720 335918
rect 599776 335862 599844 335918
rect 599900 335862 599996 335918
rect 599376 335794 599996 335862
rect 599376 335738 599472 335794
rect 599528 335738 599596 335794
rect 599652 335738 599720 335794
rect 599776 335738 599844 335794
rect 599900 335738 599996 335794
rect 599376 335670 599996 335738
rect 599376 335614 599472 335670
rect 599528 335614 599596 335670
rect 599652 335614 599720 335670
rect 599776 335614 599844 335670
rect 599900 335614 599996 335670
rect 599376 335546 599996 335614
rect 599376 335490 599472 335546
rect 599528 335490 599596 335546
rect 599652 335490 599720 335546
rect 599776 335490 599844 335546
rect 599900 335490 599996 335546
rect 599376 317918 599996 335490
rect 599376 317862 599472 317918
rect 599528 317862 599596 317918
rect 599652 317862 599720 317918
rect 599776 317862 599844 317918
rect 599900 317862 599996 317918
rect 599376 317794 599996 317862
rect 599376 317738 599472 317794
rect 599528 317738 599596 317794
rect 599652 317738 599720 317794
rect 599776 317738 599844 317794
rect 599900 317738 599996 317794
rect 599376 317670 599996 317738
rect 599376 317614 599472 317670
rect 599528 317614 599596 317670
rect 599652 317614 599720 317670
rect 599776 317614 599844 317670
rect 599900 317614 599996 317670
rect 599376 317546 599996 317614
rect 599376 317490 599472 317546
rect 599528 317490 599596 317546
rect 599652 317490 599720 317546
rect 599776 317490 599844 317546
rect 599900 317490 599996 317546
rect 599376 299918 599996 317490
rect 599376 299862 599472 299918
rect 599528 299862 599596 299918
rect 599652 299862 599720 299918
rect 599776 299862 599844 299918
rect 599900 299862 599996 299918
rect 599376 299794 599996 299862
rect 599376 299738 599472 299794
rect 599528 299738 599596 299794
rect 599652 299738 599720 299794
rect 599776 299738 599844 299794
rect 599900 299738 599996 299794
rect 599376 299670 599996 299738
rect 599376 299614 599472 299670
rect 599528 299614 599596 299670
rect 599652 299614 599720 299670
rect 599776 299614 599844 299670
rect 599900 299614 599996 299670
rect 599376 299546 599996 299614
rect 599376 299490 599472 299546
rect 599528 299490 599596 299546
rect 599652 299490 599720 299546
rect 599776 299490 599844 299546
rect 599900 299490 599996 299546
rect 599376 281918 599996 299490
rect 599376 281862 599472 281918
rect 599528 281862 599596 281918
rect 599652 281862 599720 281918
rect 599776 281862 599844 281918
rect 599900 281862 599996 281918
rect 599376 281794 599996 281862
rect 599376 281738 599472 281794
rect 599528 281738 599596 281794
rect 599652 281738 599720 281794
rect 599776 281738 599844 281794
rect 599900 281738 599996 281794
rect 599376 281670 599996 281738
rect 599376 281614 599472 281670
rect 599528 281614 599596 281670
rect 599652 281614 599720 281670
rect 599776 281614 599844 281670
rect 599900 281614 599996 281670
rect 599376 281546 599996 281614
rect 599376 281490 599472 281546
rect 599528 281490 599596 281546
rect 599652 281490 599720 281546
rect 599776 281490 599844 281546
rect 599900 281490 599996 281546
rect 599376 263918 599996 281490
rect 599376 263862 599472 263918
rect 599528 263862 599596 263918
rect 599652 263862 599720 263918
rect 599776 263862 599844 263918
rect 599900 263862 599996 263918
rect 599376 263794 599996 263862
rect 599376 263738 599472 263794
rect 599528 263738 599596 263794
rect 599652 263738 599720 263794
rect 599776 263738 599844 263794
rect 599900 263738 599996 263794
rect 599376 263670 599996 263738
rect 599376 263614 599472 263670
rect 599528 263614 599596 263670
rect 599652 263614 599720 263670
rect 599776 263614 599844 263670
rect 599900 263614 599996 263670
rect 599376 263546 599996 263614
rect 599376 263490 599472 263546
rect 599528 263490 599596 263546
rect 599652 263490 599720 263546
rect 599776 263490 599844 263546
rect 599900 263490 599996 263546
rect 599376 245918 599996 263490
rect 599376 245862 599472 245918
rect 599528 245862 599596 245918
rect 599652 245862 599720 245918
rect 599776 245862 599844 245918
rect 599900 245862 599996 245918
rect 599376 245794 599996 245862
rect 599376 245738 599472 245794
rect 599528 245738 599596 245794
rect 599652 245738 599720 245794
rect 599776 245738 599844 245794
rect 599900 245738 599996 245794
rect 599376 245670 599996 245738
rect 599376 245614 599472 245670
rect 599528 245614 599596 245670
rect 599652 245614 599720 245670
rect 599776 245614 599844 245670
rect 599900 245614 599996 245670
rect 599376 245546 599996 245614
rect 599376 245490 599472 245546
rect 599528 245490 599596 245546
rect 599652 245490 599720 245546
rect 599776 245490 599844 245546
rect 599900 245490 599996 245546
rect 599376 227918 599996 245490
rect 599376 227862 599472 227918
rect 599528 227862 599596 227918
rect 599652 227862 599720 227918
rect 599776 227862 599844 227918
rect 599900 227862 599996 227918
rect 599376 227794 599996 227862
rect 599376 227738 599472 227794
rect 599528 227738 599596 227794
rect 599652 227738 599720 227794
rect 599776 227738 599844 227794
rect 599900 227738 599996 227794
rect 599376 227670 599996 227738
rect 599376 227614 599472 227670
rect 599528 227614 599596 227670
rect 599652 227614 599720 227670
rect 599776 227614 599844 227670
rect 599900 227614 599996 227670
rect 599376 227546 599996 227614
rect 599376 227490 599472 227546
rect 599528 227490 599596 227546
rect 599652 227490 599720 227546
rect 599776 227490 599844 227546
rect 599900 227490 599996 227546
rect 599376 209918 599996 227490
rect 599376 209862 599472 209918
rect 599528 209862 599596 209918
rect 599652 209862 599720 209918
rect 599776 209862 599844 209918
rect 599900 209862 599996 209918
rect 599376 209794 599996 209862
rect 599376 209738 599472 209794
rect 599528 209738 599596 209794
rect 599652 209738 599720 209794
rect 599776 209738 599844 209794
rect 599900 209738 599996 209794
rect 599376 209670 599996 209738
rect 599376 209614 599472 209670
rect 599528 209614 599596 209670
rect 599652 209614 599720 209670
rect 599776 209614 599844 209670
rect 599900 209614 599996 209670
rect 599376 209546 599996 209614
rect 599376 209490 599472 209546
rect 599528 209490 599596 209546
rect 599652 209490 599720 209546
rect 599776 209490 599844 209546
rect 599900 209490 599996 209546
rect 599376 191918 599996 209490
rect 599376 191862 599472 191918
rect 599528 191862 599596 191918
rect 599652 191862 599720 191918
rect 599776 191862 599844 191918
rect 599900 191862 599996 191918
rect 599376 191794 599996 191862
rect 599376 191738 599472 191794
rect 599528 191738 599596 191794
rect 599652 191738 599720 191794
rect 599776 191738 599844 191794
rect 599900 191738 599996 191794
rect 599376 191670 599996 191738
rect 599376 191614 599472 191670
rect 599528 191614 599596 191670
rect 599652 191614 599720 191670
rect 599776 191614 599844 191670
rect 599900 191614 599996 191670
rect 599376 191546 599996 191614
rect 599376 191490 599472 191546
rect 599528 191490 599596 191546
rect 599652 191490 599720 191546
rect 599776 191490 599844 191546
rect 599900 191490 599996 191546
rect 599376 173918 599996 191490
rect 599376 173862 599472 173918
rect 599528 173862 599596 173918
rect 599652 173862 599720 173918
rect 599776 173862 599844 173918
rect 599900 173862 599996 173918
rect 599376 173794 599996 173862
rect 599376 173738 599472 173794
rect 599528 173738 599596 173794
rect 599652 173738 599720 173794
rect 599776 173738 599844 173794
rect 599900 173738 599996 173794
rect 599376 173670 599996 173738
rect 599376 173614 599472 173670
rect 599528 173614 599596 173670
rect 599652 173614 599720 173670
rect 599776 173614 599844 173670
rect 599900 173614 599996 173670
rect 599376 173546 599996 173614
rect 599376 173490 599472 173546
rect 599528 173490 599596 173546
rect 599652 173490 599720 173546
rect 599776 173490 599844 173546
rect 599900 173490 599996 173546
rect 599376 155918 599996 173490
rect 599376 155862 599472 155918
rect 599528 155862 599596 155918
rect 599652 155862 599720 155918
rect 599776 155862 599844 155918
rect 599900 155862 599996 155918
rect 599376 155794 599996 155862
rect 599376 155738 599472 155794
rect 599528 155738 599596 155794
rect 599652 155738 599720 155794
rect 599776 155738 599844 155794
rect 599900 155738 599996 155794
rect 599376 155670 599996 155738
rect 599376 155614 599472 155670
rect 599528 155614 599596 155670
rect 599652 155614 599720 155670
rect 599776 155614 599844 155670
rect 599900 155614 599996 155670
rect 599376 155546 599996 155614
rect 599376 155490 599472 155546
rect 599528 155490 599596 155546
rect 599652 155490 599720 155546
rect 599776 155490 599844 155546
rect 599900 155490 599996 155546
rect 599376 137918 599996 155490
rect 599376 137862 599472 137918
rect 599528 137862 599596 137918
rect 599652 137862 599720 137918
rect 599776 137862 599844 137918
rect 599900 137862 599996 137918
rect 599376 137794 599996 137862
rect 599376 137738 599472 137794
rect 599528 137738 599596 137794
rect 599652 137738 599720 137794
rect 599776 137738 599844 137794
rect 599900 137738 599996 137794
rect 599376 137670 599996 137738
rect 599376 137614 599472 137670
rect 599528 137614 599596 137670
rect 599652 137614 599720 137670
rect 599776 137614 599844 137670
rect 599900 137614 599996 137670
rect 599376 137546 599996 137614
rect 599376 137490 599472 137546
rect 599528 137490 599596 137546
rect 599652 137490 599720 137546
rect 599776 137490 599844 137546
rect 599900 137490 599996 137546
rect 599376 119918 599996 137490
rect 599376 119862 599472 119918
rect 599528 119862 599596 119918
rect 599652 119862 599720 119918
rect 599776 119862 599844 119918
rect 599900 119862 599996 119918
rect 599376 119794 599996 119862
rect 599376 119738 599472 119794
rect 599528 119738 599596 119794
rect 599652 119738 599720 119794
rect 599776 119738 599844 119794
rect 599900 119738 599996 119794
rect 599376 119670 599996 119738
rect 599376 119614 599472 119670
rect 599528 119614 599596 119670
rect 599652 119614 599720 119670
rect 599776 119614 599844 119670
rect 599900 119614 599996 119670
rect 599376 119546 599996 119614
rect 599376 119490 599472 119546
rect 599528 119490 599596 119546
rect 599652 119490 599720 119546
rect 599776 119490 599844 119546
rect 599900 119490 599996 119546
rect 599376 101918 599996 119490
rect 599376 101862 599472 101918
rect 599528 101862 599596 101918
rect 599652 101862 599720 101918
rect 599776 101862 599844 101918
rect 599900 101862 599996 101918
rect 599376 101794 599996 101862
rect 599376 101738 599472 101794
rect 599528 101738 599596 101794
rect 599652 101738 599720 101794
rect 599776 101738 599844 101794
rect 599900 101738 599996 101794
rect 599376 101670 599996 101738
rect 599376 101614 599472 101670
rect 599528 101614 599596 101670
rect 599652 101614 599720 101670
rect 599776 101614 599844 101670
rect 599900 101614 599996 101670
rect 599376 101546 599996 101614
rect 599376 101490 599472 101546
rect 599528 101490 599596 101546
rect 599652 101490 599720 101546
rect 599776 101490 599844 101546
rect 599900 101490 599996 101546
rect 599376 83918 599996 101490
rect 599376 83862 599472 83918
rect 599528 83862 599596 83918
rect 599652 83862 599720 83918
rect 599776 83862 599844 83918
rect 599900 83862 599996 83918
rect 599376 83794 599996 83862
rect 599376 83738 599472 83794
rect 599528 83738 599596 83794
rect 599652 83738 599720 83794
rect 599776 83738 599844 83794
rect 599900 83738 599996 83794
rect 599376 83670 599996 83738
rect 599376 83614 599472 83670
rect 599528 83614 599596 83670
rect 599652 83614 599720 83670
rect 599776 83614 599844 83670
rect 599900 83614 599996 83670
rect 599376 83546 599996 83614
rect 599376 83490 599472 83546
rect 599528 83490 599596 83546
rect 599652 83490 599720 83546
rect 599776 83490 599844 83546
rect 599900 83490 599996 83546
rect 599376 65918 599996 83490
rect 599376 65862 599472 65918
rect 599528 65862 599596 65918
rect 599652 65862 599720 65918
rect 599776 65862 599844 65918
rect 599900 65862 599996 65918
rect 599376 65794 599996 65862
rect 599376 65738 599472 65794
rect 599528 65738 599596 65794
rect 599652 65738 599720 65794
rect 599776 65738 599844 65794
rect 599900 65738 599996 65794
rect 599376 65670 599996 65738
rect 599376 65614 599472 65670
rect 599528 65614 599596 65670
rect 599652 65614 599720 65670
rect 599776 65614 599844 65670
rect 599900 65614 599996 65670
rect 599376 65546 599996 65614
rect 599376 65490 599472 65546
rect 599528 65490 599596 65546
rect 599652 65490 599720 65546
rect 599776 65490 599844 65546
rect 599900 65490 599996 65546
rect 599376 47918 599996 65490
rect 599376 47862 599472 47918
rect 599528 47862 599596 47918
rect 599652 47862 599720 47918
rect 599776 47862 599844 47918
rect 599900 47862 599996 47918
rect 599376 47794 599996 47862
rect 599376 47738 599472 47794
rect 599528 47738 599596 47794
rect 599652 47738 599720 47794
rect 599776 47738 599844 47794
rect 599900 47738 599996 47794
rect 599376 47670 599996 47738
rect 599376 47614 599472 47670
rect 599528 47614 599596 47670
rect 599652 47614 599720 47670
rect 599776 47614 599844 47670
rect 599900 47614 599996 47670
rect 599376 47546 599996 47614
rect 599376 47490 599472 47546
rect 599528 47490 599596 47546
rect 599652 47490 599720 47546
rect 599776 47490 599844 47546
rect 599900 47490 599996 47546
rect 599376 29918 599996 47490
rect 599376 29862 599472 29918
rect 599528 29862 599596 29918
rect 599652 29862 599720 29918
rect 599776 29862 599844 29918
rect 599900 29862 599996 29918
rect 599376 29794 599996 29862
rect 599376 29738 599472 29794
rect 599528 29738 599596 29794
rect 599652 29738 599720 29794
rect 599776 29738 599844 29794
rect 599900 29738 599996 29794
rect 599376 29670 599996 29738
rect 599376 29614 599472 29670
rect 599528 29614 599596 29670
rect 599652 29614 599720 29670
rect 599776 29614 599844 29670
rect 599900 29614 599996 29670
rect 599376 29546 599996 29614
rect 599376 29490 599472 29546
rect 599528 29490 599596 29546
rect 599652 29490 599720 29546
rect 599776 29490 599844 29546
rect 599900 29490 599996 29546
rect 599376 11918 599996 29490
rect 599376 11862 599472 11918
rect 599528 11862 599596 11918
rect 599652 11862 599720 11918
rect 599776 11862 599844 11918
rect 599900 11862 599996 11918
rect 599376 11794 599996 11862
rect 599376 11738 599472 11794
rect 599528 11738 599596 11794
rect 599652 11738 599720 11794
rect 599776 11738 599844 11794
rect 599900 11738 599996 11794
rect 599376 11670 599996 11738
rect 599376 11614 599472 11670
rect 599528 11614 599596 11670
rect 599652 11614 599720 11670
rect 599776 11614 599844 11670
rect 599900 11614 599996 11670
rect 599376 11546 599996 11614
rect 599376 11490 599472 11546
rect 599528 11490 599596 11546
rect 599652 11490 599720 11546
rect 599776 11490 599844 11546
rect 599900 11490 599996 11546
rect 584778 792 584874 848
rect 584930 792 584998 848
rect 585054 792 585122 848
rect 585178 792 585246 848
rect 585302 792 585398 848
rect 584778 724 585398 792
rect 584778 668 584874 724
rect 584930 668 584998 724
rect 585054 668 585122 724
rect 585178 668 585246 724
rect 585302 668 585398 724
rect 584778 600 585398 668
rect 584778 544 584874 600
rect 584930 544 584998 600
rect 585054 544 585122 600
rect 585178 544 585246 600
rect 585302 544 585398 600
rect 584778 476 585398 544
rect 584778 420 584874 476
rect 584930 420 584998 476
rect 585054 420 585122 476
rect 585178 420 585246 476
rect 585302 420 585398 476
rect 584778 324 585398 420
rect 599376 848 599996 11490
rect 599376 792 599472 848
rect 599528 792 599596 848
rect 599652 792 599720 848
rect 599776 792 599844 848
rect 599900 792 599996 848
rect 599376 724 599996 792
rect 599376 668 599472 724
rect 599528 668 599596 724
rect 599652 668 599720 724
rect 599776 668 599844 724
rect 599900 668 599996 724
rect 599376 600 599996 668
rect 599376 544 599472 600
rect 599528 544 599596 600
rect 599652 544 599720 600
rect 599776 544 599844 600
rect 599900 544 599996 600
rect 599376 476 599996 544
rect 599376 420 599472 476
rect 599528 420 599596 476
rect 599652 420 599720 476
rect 599776 420 599844 476
rect 599900 420 599996 476
rect 599376 324 599996 420
<< via4 >>
rect 84 599284 140 599340
rect 208 599284 264 599340
rect 332 599284 388 599340
rect 456 599284 512 599340
rect 84 599160 140 599216
rect 208 599160 264 599216
rect 332 599160 388 599216
rect 456 599160 512 599216
rect 84 599036 140 599092
rect 208 599036 264 599092
rect 332 599036 388 599092
rect 456 599036 512 599092
rect 84 598912 140 598968
rect 208 598912 264 598968
rect 332 598912 388 598968
rect 456 598912 512 598968
rect 84 587862 140 587918
rect 208 587862 264 587918
rect 332 587862 388 587918
rect 456 587862 512 587918
rect 84 587738 140 587794
rect 208 587738 264 587794
rect 332 587738 388 587794
rect 456 587738 512 587794
rect 84 587614 140 587670
rect 208 587614 264 587670
rect 332 587614 388 587670
rect 456 587614 512 587670
rect 84 587490 140 587546
rect 208 587490 264 587546
rect 332 587490 388 587546
rect 456 587490 512 587546
rect 84 569862 140 569918
rect 208 569862 264 569918
rect 332 569862 388 569918
rect 456 569862 512 569918
rect 84 569738 140 569794
rect 208 569738 264 569794
rect 332 569738 388 569794
rect 456 569738 512 569794
rect 84 569614 140 569670
rect 208 569614 264 569670
rect 332 569614 388 569670
rect 456 569614 512 569670
rect 84 569490 140 569546
rect 208 569490 264 569546
rect 332 569490 388 569546
rect 456 569490 512 569546
rect 84 551862 140 551918
rect 208 551862 264 551918
rect 332 551862 388 551918
rect 456 551862 512 551918
rect 84 551738 140 551794
rect 208 551738 264 551794
rect 332 551738 388 551794
rect 456 551738 512 551794
rect 84 551614 140 551670
rect 208 551614 264 551670
rect 332 551614 388 551670
rect 456 551614 512 551670
rect 84 551490 140 551546
rect 208 551490 264 551546
rect 332 551490 388 551546
rect 456 551490 512 551546
rect 84 533862 140 533918
rect 208 533862 264 533918
rect 332 533862 388 533918
rect 456 533862 512 533918
rect 84 533738 140 533794
rect 208 533738 264 533794
rect 332 533738 388 533794
rect 456 533738 512 533794
rect 84 533614 140 533670
rect 208 533614 264 533670
rect 332 533614 388 533670
rect 456 533614 512 533670
rect 84 533490 140 533546
rect 208 533490 264 533546
rect 332 533490 388 533546
rect 456 533490 512 533546
rect 84 515862 140 515918
rect 208 515862 264 515918
rect 332 515862 388 515918
rect 456 515862 512 515918
rect 84 515738 140 515794
rect 208 515738 264 515794
rect 332 515738 388 515794
rect 456 515738 512 515794
rect 84 515614 140 515670
rect 208 515614 264 515670
rect 332 515614 388 515670
rect 456 515614 512 515670
rect 84 515490 140 515546
rect 208 515490 264 515546
rect 332 515490 388 515546
rect 456 515490 512 515546
rect 84 497862 140 497918
rect 208 497862 264 497918
rect 332 497862 388 497918
rect 456 497862 512 497918
rect 84 497738 140 497794
rect 208 497738 264 497794
rect 332 497738 388 497794
rect 456 497738 512 497794
rect 84 497614 140 497670
rect 208 497614 264 497670
rect 332 497614 388 497670
rect 456 497614 512 497670
rect 84 497490 140 497546
rect 208 497490 264 497546
rect 332 497490 388 497546
rect 456 497490 512 497546
rect 84 479862 140 479918
rect 208 479862 264 479918
rect 332 479862 388 479918
rect 456 479862 512 479918
rect 84 479738 140 479794
rect 208 479738 264 479794
rect 332 479738 388 479794
rect 456 479738 512 479794
rect 84 479614 140 479670
rect 208 479614 264 479670
rect 332 479614 388 479670
rect 456 479614 512 479670
rect 84 479490 140 479546
rect 208 479490 264 479546
rect 332 479490 388 479546
rect 456 479490 512 479546
rect 84 461862 140 461918
rect 208 461862 264 461918
rect 332 461862 388 461918
rect 456 461862 512 461918
rect 84 461738 140 461794
rect 208 461738 264 461794
rect 332 461738 388 461794
rect 456 461738 512 461794
rect 84 461614 140 461670
rect 208 461614 264 461670
rect 332 461614 388 461670
rect 456 461614 512 461670
rect 84 461490 140 461546
rect 208 461490 264 461546
rect 332 461490 388 461546
rect 456 461490 512 461546
rect 84 443862 140 443918
rect 208 443862 264 443918
rect 332 443862 388 443918
rect 456 443862 512 443918
rect 84 443738 140 443794
rect 208 443738 264 443794
rect 332 443738 388 443794
rect 456 443738 512 443794
rect 84 443614 140 443670
rect 208 443614 264 443670
rect 332 443614 388 443670
rect 456 443614 512 443670
rect 84 443490 140 443546
rect 208 443490 264 443546
rect 332 443490 388 443546
rect 456 443490 512 443546
rect 84 425862 140 425918
rect 208 425862 264 425918
rect 332 425862 388 425918
rect 456 425862 512 425918
rect 84 425738 140 425794
rect 208 425738 264 425794
rect 332 425738 388 425794
rect 456 425738 512 425794
rect 84 425614 140 425670
rect 208 425614 264 425670
rect 332 425614 388 425670
rect 456 425614 512 425670
rect 84 425490 140 425546
rect 208 425490 264 425546
rect 332 425490 388 425546
rect 456 425490 512 425546
rect 84 407862 140 407918
rect 208 407862 264 407918
rect 332 407862 388 407918
rect 456 407862 512 407918
rect 84 407738 140 407794
rect 208 407738 264 407794
rect 332 407738 388 407794
rect 456 407738 512 407794
rect 84 407614 140 407670
rect 208 407614 264 407670
rect 332 407614 388 407670
rect 456 407614 512 407670
rect 84 407490 140 407546
rect 208 407490 264 407546
rect 332 407490 388 407546
rect 456 407490 512 407546
rect 84 389862 140 389918
rect 208 389862 264 389918
rect 332 389862 388 389918
rect 456 389862 512 389918
rect 84 389738 140 389794
rect 208 389738 264 389794
rect 332 389738 388 389794
rect 456 389738 512 389794
rect 84 389614 140 389670
rect 208 389614 264 389670
rect 332 389614 388 389670
rect 456 389614 512 389670
rect 84 389490 140 389546
rect 208 389490 264 389546
rect 332 389490 388 389546
rect 456 389490 512 389546
rect 84 371862 140 371918
rect 208 371862 264 371918
rect 332 371862 388 371918
rect 456 371862 512 371918
rect 84 371738 140 371794
rect 208 371738 264 371794
rect 332 371738 388 371794
rect 456 371738 512 371794
rect 84 371614 140 371670
rect 208 371614 264 371670
rect 332 371614 388 371670
rect 456 371614 512 371670
rect 84 371490 140 371546
rect 208 371490 264 371546
rect 332 371490 388 371546
rect 456 371490 512 371546
rect 84 353862 140 353918
rect 208 353862 264 353918
rect 332 353862 388 353918
rect 456 353862 512 353918
rect 84 353738 140 353794
rect 208 353738 264 353794
rect 332 353738 388 353794
rect 456 353738 512 353794
rect 84 353614 140 353670
rect 208 353614 264 353670
rect 332 353614 388 353670
rect 456 353614 512 353670
rect 84 353490 140 353546
rect 208 353490 264 353546
rect 332 353490 388 353546
rect 456 353490 512 353546
rect 84 335862 140 335918
rect 208 335862 264 335918
rect 332 335862 388 335918
rect 456 335862 512 335918
rect 84 335738 140 335794
rect 208 335738 264 335794
rect 332 335738 388 335794
rect 456 335738 512 335794
rect 84 335614 140 335670
rect 208 335614 264 335670
rect 332 335614 388 335670
rect 456 335614 512 335670
rect 84 335490 140 335546
rect 208 335490 264 335546
rect 332 335490 388 335546
rect 456 335490 512 335546
rect 84 317862 140 317918
rect 208 317862 264 317918
rect 332 317862 388 317918
rect 456 317862 512 317918
rect 84 317738 140 317794
rect 208 317738 264 317794
rect 332 317738 388 317794
rect 456 317738 512 317794
rect 84 317614 140 317670
rect 208 317614 264 317670
rect 332 317614 388 317670
rect 456 317614 512 317670
rect 84 317490 140 317546
rect 208 317490 264 317546
rect 332 317490 388 317546
rect 456 317490 512 317546
rect 84 299862 140 299918
rect 208 299862 264 299918
rect 332 299862 388 299918
rect 456 299862 512 299918
rect 84 299738 140 299794
rect 208 299738 264 299794
rect 332 299738 388 299794
rect 456 299738 512 299794
rect 84 299614 140 299670
rect 208 299614 264 299670
rect 332 299614 388 299670
rect 456 299614 512 299670
rect 84 299490 140 299546
rect 208 299490 264 299546
rect 332 299490 388 299546
rect 456 299490 512 299546
rect 84 281862 140 281918
rect 208 281862 264 281918
rect 332 281862 388 281918
rect 456 281862 512 281918
rect 84 281738 140 281794
rect 208 281738 264 281794
rect 332 281738 388 281794
rect 456 281738 512 281794
rect 84 281614 140 281670
rect 208 281614 264 281670
rect 332 281614 388 281670
rect 456 281614 512 281670
rect 84 281490 140 281546
rect 208 281490 264 281546
rect 332 281490 388 281546
rect 456 281490 512 281546
rect 84 263862 140 263918
rect 208 263862 264 263918
rect 332 263862 388 263918
rect 456 263862 512 263918
rect 84 263738 140 263794
rect 208 263738 264 263794
rect 332 263738 388 263794
rect 456 263738 512 263794
rect 84 263614 140 263670
rect 208 263614 264 263670
rect 332 263614 388 263670
rect 456 263614 512 263670
rect 84 263490 140 263546
rect 208 263490 264 263546
rect 332 263490 388 263546
rect 456 263490 512 263546
rect 84 245862 140 245918
rect 208 245862 264 245918
rect 332 245862 388 245918
rect 456 245862 512 245918
rect 84 245738 140 245794
rect 208 245738 264 245794
rect 332 245738 388 245794
rect 456 245738 512 245794
rect 84 245614 140 245670
rect 208 245614 264 245670
rect 332 245614 388 245670
rect 456 245614 512 245670
rect 84 245490 140 245546
rect 208 245490 264 245546
rect 332 245490 388 245546
rect 456 245490 512 245546
rect 84 227862 140 227918
rect 208 227862 264 227918
rect 332 227862 388 227918
rect 456 227862 512 227918
rect 84 227738 140 227794
rect 208 227738 264 227794
rect 332 227738 388 227794
rect 456 227738 512 227794
rect 84 227614 140 227670
rect 208 227614 264 227670
rect 332 227614 388 227670
rect 456 227614 512 227670
rect 84 227490 140 227546
rect 208 227490 264 227546
rect 332 227490 388 227546
rect 456 227490 512 227546
rect 84 209862 140 209918
rect 208 209862 264 209918
rect 332 209862 388 209918
rect 456 209862 512 209918
rect 84 209738 140 209794
rect 208 209738 264 209794
rect 332 209738 388 209794
rect 456 209738 512 209794
rect 84 209614 140 209670
rect 208 209614 264 209670
rect 332 209614 388 209670
rect 456 209614 512 209670
rect 84 209490 140 209546
rect 208 209490 264 209546
rect 332 209490 388 209546
rect 456 209490 512 209546
rect 84 191862 140 191918
rect 208 191862 264 191918
rect 332 191862 388 191918
rect 456 191862 512 191918
rect 84 191738 140 191794
rect 208 191738 264 191794
rect 332 191738 388 191794
rect 456 191738 512 191794
rect 84 191614 140 191670
rect 208 191614 264 191670
rect 332 191614 388 191670
rect 456 191614 512 191670
rect 84 191490 140 191546
rect 208 191490 264 191546
rect 332 191490 388 191546
rect 456 191490 512 191546
rect 84 173862 140 173918
rect 208 173862 264 173918
rect 332 173862 388 173918
rect 456 173862 512 173918
rect 84 173738 140 173794
rect 208 173738 264 173794
rect 332 173738 388 173794
rect 456 173738 512 173794
rect 84 173614 140 173670
rect 208 173614 264 173670
rect 332 173614 388 173670
rect 456 173614 512 173670
rect 84 173490 140 173546
rect 208 173490 264 173546
rect 332 173490 388 173546
rect 456 173490 512 173546
rect 84 155862 140 155918
rect 208 155862 264 155918
rect 332 155862 388 155918
rect 456 155862 512 155918
rect 84 155738 140 155794
rect 208 155738 264 155794
rect 332 155738 388 155794
rect 456 155738 512 155794
rect 84 155614 140 155670
rect 208 155614 264 155670
rect 332 155614 388 155670
rect 456 155614 512 155670
rect 84 155490 140 155546
rect 208 155490 264 155546
rect 332 155490 388 155546
rect 456 155490 512 155546
rect 84 137862 140 137918
rect 208 137862 264 137918
rect 332 137862 388 137918
rect 456 137862 512 137918
rect 84 137738 140 137794
rect 208 137738 264 137794
rect 332 137738 388 137794
rect 456 137738 512 137794
rect 84 137614 140 137670
rect 208 137614 264 137670
rect 332 137614 388 137670
rect 456 137614 512 137670
rect 84 137490 140 137546
rect 208 137490 264 137546
rect 332 137490 388 137546
rect 456 137490 512 137546
rect 84 119862 140 119918
rect 208 119862 264 119918
rect 332 119862 388 119918
rect 456 119862 512 119918
rect 84 119738 140 119794
rect 208 119738 264 119794
rect 332 119738 388 119794
rect 456 119738 512 119794
rect 84 119614 140 119670
rect 208 119614 264 119670
rect 332 119614 388 119670
rect 456 119614 512 119670
rect 84 119490 140 119546
rect 208 119490 264 119546
rect 332 119490 388 119546
rect 456 119490 512 119546
rect 84 101862 140 101918
rect 208 101862 264 101918
rect 332 101862 388 101918
rect 456 101862 512 101918
rect 84 101738 140 101794
rect 208 101738 264 101794
rect 332 101738 388 101794
rect 456 101738 512 101794
rect 84 101614 140 101670
rect 208 101614 264 101670
rect 332 101614 388 101670
rect 456 101614 512 101670
rect 84 101490 140 101546
rect 208 101490 264 101546
rect 332 101490 388 101546
rect 456 101490 512 101546
rect 84 83862 140 83918
rect 208 83862 264 83918
rect 332 83862 388 83918
rect 456 83862 512 83918
rect 84 83738 140 83794
rect 208 83738 264 83794
rect 332 83738 388 83794
rect 456 83738 512 83794
rect 84 83614 140 83670
rect 208 83614 264 83670
rect 332 83614 388 83670
rect 456 83614 512 83670
rect 84 83490 140 83546
rect 208 83490 264 83546
rect 332 83490 388 83546
rect 456 83490 512 83546
rect 84 65862 140 65918
rect 208 65862 264 65918
rect 332 65862 388 65918
rect 456 65862 512 65918
rect 84 65738 140 65794
rect 208 65738 264 65794
rect 332 65738 388 65794
rect 456 65738 512 65794
rect 84 65614 140 65670
rect 208 65614 264 65670
rect 332 65614 388 65670
rect 456 65614 512 65670
rect 84 65490 140 65546
rect 208 65490 264 65546
rect 332 65490 388 65546
rect 456 65490 512 65546
rect 84 47862 140 47918
rect 208 47862 264 47918
rect 332 47862 388 47918
rect 456 47862 512 47918
rect 84 47738 140 47794
rect 208 47738 264 47794
rect 332 47738 388 47794
rect 456 47738 512 47794
rect 84 47614 140 47670
rect 208 47614 264 47670
rect 332 47614 388 47670
rect 456 47614 512 47670
rect 84 47490 140 47546
rect 208 47490 264 47546
rect 332 47490 388 47546
rect 456 47490 512 47546
rect 84 29862 140 29918
rect 208 29862 264 29918
rect 332 29862 388 29918
rect 456 29862 512 29918
rect 84 29738 140 29794
rect 208 29738 264 29794
rect 332 29738 388 29794
rect 456 29738 512 29794
rect 84 29614 140 29670
rect 208 29614 264 29670
rect 332 29614 388 29670
rect 456 29614 512 29670
rect 84 29490 140 29546
rect 208 29490 264 29546
rect 332 29490 388 29546
rect 456 29490 512 29546
rect 84 11862 140 11918
rect 208 11862 264 11918
rect 332 11862 388 11918
rect 456 11862 512 11918
rect 84 11738 140 11794
rect 208 11738 264 11794
rect 332 11738 388 11794
rect 456 11738 512 11794
rect 84 11614 140 11670
rect 208 11614 264 11670
rect 332 11614 388 11670
rect 456 11614 512 11670
rect 84 11490 140 11546
rect 208 11490 264 11546
rect 332 11490 388 11546
rect 456 11490 512 11546
rect 1044 598324 1100 598380
rect 1168 598324 1224 598380
rect 1292 598324 1348 598380
rect 1416 598324 1472 598380
rect 1044 598200 1100 598256
rect 1168 598200 1224 598256
rect 1292 598200 1348 598256
rect 1416 598200 1472 598256
rect 1044 598076 1100 598132
rect 1168 598076 1224 598132
rect 1292 598076 1348 598132
rect 1416 598076 1472 598132
rect 1044 597952 1100 598008
rect 1168 597952 1224 598008
rect 1292 597952 1348 598008
rect 1416 597952 1472 598008
rect 1044 581862 1100 581918
rect 1168 581862 1224 581918
rect 1292 581862 1348 581918
rect 1416 581862 1472 581918
rect 1044 581738 1100 581794
rect 1168 581738 1224 581794
rect 1292 581738 1348 581794
rect 1416 581738 1472 581794
rect 1044 581614 1100 581670
rect 1168 581614 1224 581670
rect 1292 581614 1348 581670
rect 1416 581614 1472 581670
rect 1044 581490 1100 581546
rect 1168 581490 1224 581546
rect 1292 581490 1348 581546
rect 1416 581490 1472 581546
rect 1044 563862 1100 563918
rect 1168 563862 1224 563918
rect 1292 563862 1348 563918
rect 1416 563862 1472 563918
rect 1044 563738 1100 563794
rect 1168 563738 1224 563794
rect 1292 563738 1348 563794
rect 1416 563738 1472 563794
rect 1044 563614 1100 563670
rect 1168 563614 1224 563670
rect 1292 563614 1348 563670
rect 1416 563614 1472 563670
rect 1044 563490 1100 563546
rect 1168 563490 1224 563546
rect 1292 563490 1348 563546
rect 1416 563490 1472 563546
rect 1044 545862 1100 545918
rect 1168 545862 1224 545918
rect 1292 545862 1348 545918
rect 1416 545862 1472 545918
rect 1044 545738 1100 545794
rect 1168 545738 1224 545794
rect 1292 545738 1348 545794
rect 1416 545738 1472 545794
rect 1044 545614 1100 545670
rect 1168 545614 1224 545670
rect 1292 545614 1348 545670
rect 1416 545614 1472 545670
rect 1044 545490 1100 545546
rect 1168 545490 1224 545546
rect 1292 545490 1348 545546
rect 1416 545490 1472 545546
rect 1044 527862 1100 527918
rect 1168 527862 1224 527918
rect 1292 527862 1348 527918
rect 1416 527862 1472 527918
rect 1044 527738 1100 527794
rect 1168 527738 1224 527794
rect 1292 527738 1348 527794
rect 1416 527738 1472 527794
rect 1044 527614 1100 527670
rect 1168 527614 1224 527670
rect 1292 527614 1348 527670
rect 1416 527614 1472 527670
rect 1044 527490 1100 527546
rect 1168 527490 1224 527546
rect 1292 527490 1348 527546
rect 1416 527490 1472 527546
rect 1044 509862 1100 509918
rect 1168 509862 1224 509918
rect 1292 509862 1348 509918
rect 1416 509862 1472 509918
rect 1044 509738 1100 509794
rect 1168 509738 1224 509794
rect 1292 509738 1348 509794
rect 1416 509738 1472 509794
rect 1044 509614 1100 509670
rect 1168 509614 1224 509670
rect 1292 509614 1348 509670
rect 1416 509614 1472 509670
rect 1044 509490 1100 509546
rect 1168 509490 1224 509546
rect 1292 509490 1348 509546
rect 1416 509490 1472 509546
rect 1044 491862 1100 491918
rect 1168 491862 1224 491918
rect 1292 491862 1348 491918
rect 1416 491862 1472 491918
rect 1044 491738 1100 491794
rect 1168 491738 1224 491794
rect 1292 491738 1348 491794
rect 1416 491738 1472 491794
rect 1044 491614 1100 491670
rect 1168 491614 1224 491670
rect 1292 491614 1348 491670
rect 1416 491614 1472 491670
rect 1044 491490 1100 491546
rect 1168 491490 1224 491546
rect 1292 491490 1348 491546
rect 1416 491490 1472 491546
rect 1044 473862 1100 473918
rect 1168 473862 1224 473918
rect 1292 473862 1348 473918
rect 1416 473862 1472 473918
rect 1044 473738 1100 473794
rect 1168 473738 1224 473794
rect 1292 473738 1348 473794
rect 1416 473738 1472 473794
rect 1044 473614 1100 473670
rect 1168 473614 1224 473670
rect 1292 473614 1348 473670
rect 1416 473614 1472 473670
rect 1044 473490 1100 473546
rect 1168 473490 1224 473546
rect 1292 473490 1348 473546
rect 1416 473490 1472 473546
rect 1044 455862 1100 455918
rect 1168 455862 1224 455918
rect 1292 455862 1348 455918
rect 1416 455862 1472 455918
rect 1044 455738 1100 455794
rect 1168 455738 1224 455794
rect 1292 455738 1348 455794
rect 1416 455738 1472 455794
rect 1044 455614 1100 455670
rect 1168 455614 1224 455670
rect 1292 455614 1348 455670
rect 1416 455614 1472 455670
rect 1044 455490 1100 455546
rect 1168 455490 1224 455546
rect 1292 455490 1348 455546
rect 1416 455490 1472 455546
rect 1044 437862 1100 437918
rect 1168 437862 1224 437918
rect 1292 437862 1348 437918
rect 1416 437862 1472 437918
rect 1044 437738 1100 437794
rect 1168 437738 1224 437794
rect 1292 437738 1348 437794
rect 1416 437738 1472 437794
rect 1044 437614 1100 437670
rect 1168 437614 1224 437670
rect 1292 437614 1348 437670
rect 1416 437614 1472 437670
rect 1044 437490 1100 437546
rect 1168 437490 1224 437546
rect 1292 437490 1348 437546
rect 1416 437490 1472 437546
rect 1044 419862 1100 419918
rect 1168 419862 1224 419918
rect 1292 419862 1348 419918
rect 1416 419862 1472 419918
rect 1044 419738 1100 419794
rect 1168 419738 1224 419794
rect 1292 419738 1348 419794
rect 1416 419738 1472 419794
rect 1044 419614 1100 419670
rect 1168 419614 1224 419670
rect 1292 419614 1348 419670
rect 1416 419614 1472 419670
rect 1044 419490 1100 419546
rect 1168 419490 1224 419546
rect 1292 419490 1348 419546
rect 1416 419490 1472 419546
rect 1044 401862 1100 401918
rect 1168 401862 1224 401918
rect 1292 401862 1348 401918
rect 1416 401862 1472 401918
rect 1044 401738 1100 401794
rect 1168 401738 1224 401794
rect 1292 401738 1348 401794
rect 1416 401738 1472 401794
rect 1044 401614 1100 401670
rect 1168 401614 1224 401670
rect 1292 401614 1348 401670
rect 1416 401614 1472 401670
rect 1044 401490 1100 401546
rect 1168 401490 1224 401546
rect 1292 401490 1348 401546
rect 1416 401490 1472 401546
rect 1044 383862 1100 383918
rect 1168 383862 1224 383918
rect 1292 383862 1348 383918
rect 1416 383862 1472 383918
rect 1044 383738 1100 383794
rect 1168 383738 1224 383794
rect 1292 383738 1348 383794
rect 1416 383738 1472 383794
rect 1044 383614 1100 383670
rect 1168 383614 1224 383670
rect 1292 383614 1348 383670
rect 1416 383614 1472 383670
rect 1044 383490 1100 383546
rect 1168 383490 1224 383546
rect 1292 383490 1348 383546
rect 1416 383490 1472 383546
rect 1044 365862 1100 365918
rect 1168 365862 1224 365918
rect 1292 365862 1348 365918
rect 1416 365862 1472 365918
rect 1044 365738 1100 365794
rect 1168 365738 1224 365794
rect 1292 365738 1348 365794
rect 1416 365738 1472 365794
rect 1044 365614 1100 365670
rect 1168 365614 1224 365670
rect 1292 365614 1348 365670
rect 1416 365614 1472 365670
rect 1044 365490 1100 365546
rect 1168 365490 1224 365546
rect 1292 365490 1348 365546
rect 1416 365490 1472 365546
rect 1044 347862 1100 347918
rect 1168 347862 1224 347918
rect 1292 347862 1348 347918
rect 1416 347862 1472 347918
rect 1044 347738 1100 347794
rect 1168 347738 1224 347794
rect 1292 347738 1348 347794
rect 1416 347738 1472 347794
rect 1044 347614 1100 347670
rect 1168 347614 1224 347670
rect 1292 347614 1348 347670
rect 1416 347614 1472 347670
rect 1044 347490 1100 347546
rect 1168 347490 1224 347546
rect 1292 347490 1348 347546
rect 1416 347490 1472 347546
rect 1044 329862 1100 329918
rect 1168 329862 1224 329918
rect 1292 329862 1348 329918
rect 1416 329862 1472 329918
rect 1044 329738 1100 329794
rect 1168 329738 1224 329794
rect 1292 329738 1348 329794
rect 1416 329738 1472 329794
rect 1044 329614 1100 329670
rect 1168 329614 1224 329670
rect 1292 329614 1348 329670
rect 1416 329614 1472 329670
rect 1044 329490 1100 329546
rect 1168 329490 1224 329546
rect 1292 329490 1348 329546
rect 1416 329490 1472 329546
rect 1044 311862 1100 311918
rect 1168 311862 1224 311918
rect 1292 311862 1348 311918
rect 1416 311862 1472 311918
rect 1044 311738 1100 311794
rect 1168 311738 1224 311794
rect 1292 311738 1348 311794
rect 1416 311738 1472 311794
rect 1044 311614 1100 311670
rect 1168 311614 1224 311670
rect 1292 311614 1348 311670
rect 1416 311614 1472 311670
rect 1044 311490 1100 311546
rect 1168 311490 1224 311546
rect 1292 311490 1348 311546
rect 1416 311490 1472 311546
rect 1044 293862 1100 293918
rect 1168 293862 1224 293918
rect 1292 293862 1348 293918
rect 1416 293862 1472 293918
rect 1044 293738 1100 293794
rect 1168 293738 1224 293794
rect 1292 293738 1348 293794
rect 1416 293738 1472 293794
rect 1044 293614 1100 293670
rect 1168 293614 1224 293670
rect 1292 293614 1348 293670
rect 1416 293614 1472 293670
rect 1044 293490 1100 293546
rect 1168 293490 1224 293546
rect 1292 293490 1348 293546
rect 1416 293490 1472 293546
rect 1044 275862 1100 275918
rect 1168 275862 1224 275918
rect 1292 275862 1348 275918
rect 1416 275862 1472 275918
rect 1044 275738 1100 275794
rect 1168 275738 1224 275794
rect 1292 275738 1348 275794
rect 1416 275738 1472 275794
rect 1044 275614 1100 275670
rect 1168 275614 1224 275670
rect 1292 275614 1348 275670
rect 1416 275614 1472 275670
rect 1044 275490 1100 275546
rect 1168 275490 1224 275546
rect 1292 275490 1348 275546
rect 1416 275490 1472 275546
rect 1044 257862 1100 257918
rect 1168 257862 1224 257918
rect 1292 257862 1348 257918
rect 1416 257862 1472 257918
rect 1044 257738 1100 257794
rect 1168 257738 1224 257794
rect 1292 257738 1348 257794
rect 1416 257738 1472 257794
rect 1044 257614 1100 257670
rect 1168 257614 1224 257670
rect 1292 257614 1348 257670
rect 1416 257614 1472 257670
rect 1044 257490 1100 257546
rect 1168 257490 1224 257546
rect 1292 257490 1348 257546
rect 1416 257490 1472 257546
rect 1044 239862 1100 239918
rect 1168 239862 1224 239918
rect 1292 239862 1348 239918
rect 1416 239862 1472 239918
rect 1044 239738 1100 239794
rect 1168 239738 1224 239794
rect 1292 239738 1348 239794
rect 1416 239738 1472 239794
rect 1044 239614 1100 239670
rect 1168 239614 1224 239670
rect 1292 239614 1348 239670
rect 1416 239614 1472 239670
rect 1044 239490 1100 239546
rect 1168 239490 1224 239546
rect 1292 239490 1348 239546
rect 1416 239490 1472 239546
rect 1044 221862 1100 221918
rect 1168 221862 1224 221918
rect 1292 221862 1348 221918
rect 1416 221862 1472 221918
rect 1044 221738 1100 221794
rect 1168 221738 1224 221794
rect 1292 221738 1348 221794
rect 1416 221738 1472 221794
rect 1044 221614 1100 221670
rect 1168 221614 1224 221670
rect 1292 221614 1348 221670
rect 1416 221614 1472 221670
rect 1044 221490 1100 221546
rect 1168 221490 1224 221546
rect 1292 221490 1348 221546
rect 1416 221490 1472 221546
rect 1044 203862 1100 203918
rect 1168 203862 1224 203918
rect 1292 203862 1348 203918
rect 1416 203862 1472 203918
rect 1044 203738 1100 203794
rect 1168 203738 1224 203794
rect 1292 203738 1348 203794
rect 1416 203738 1472 203794
rect 1044 203614 1100 203670
rect 1168 203614 1224 203670
rect 1292 203614 1348 203670
rect 1416 203614 1472 203670
rect 1044 203490 1100 203546
rect 1168 203490 1224 203546
rect 1292 203490 1348 203546
rect 1416 203490 1472 203546
rect 1044 185862 1100 185918
rect 1168 185862 1224 185918
rect 1292 185862 1348 185918
rect 1416 185862 1472 185918
rect 1044 185738 1100 185794
rect 1168 185738 1224 185794
rect 1292 185738 1348 185794
rect 1416 185738 1472 185794
rect 1044 185614 1100 185670
rect 1168 185614 1224 185670
rect 1292 185614 1348 185670
rect 1416 185614 1472 185670
rect 1044 185490 1100 185546
rect 1168 185490 1224 185546
rect 1292 185490 1348 185546
rect 1416 185490 1472 185546
rect 1044 167862 1100 167918
rect 1168 167862 1224 167918
rect 1292 167862 1348 167918
rect 1416 167862 1472 167918
rect 1044 167738 1100 167794
rect 1168 167738 1224 167794
rect 1292 167738 1348 167794
rect 1416 167738 1472 167794
rect 1044 167614 1100 167670
rect 1168 167614 1224 167670
rect 1292 167614 1348 167670
rect 1416 167614 1472 167670
rect 1044 167490 1100 167546
rect 1168 167490 1224 167546
rect 1292 167490 1348 167546
rect 1416 167490 1472 167546
rect 1044 149862 1100 149918
rect 1168 149862 1224 149918
rect 1292 149862 1348 149918
rect 1416 149862 1472 149918
rect 1044 149738 1100 149794
rect 1168 149738 1224 149794
rect 1292 149738 1348 149794
rect 1416 149738 1472 149794
rect 1044 149614 1100 149670
rect 1168 149614 1224 149670
rect 1292 149614 1348 149670
rect 1416 149614 1472 149670
rect 1044 149490 1100 149546
rect 1168 149490 1224 149546
rect 1292 149490 1348 149546
rect 1416 149490 1472 149546
rect 1044 131862 1100 131918
rect 1168 131862 1224 131918
rect 1292 131862 1348 131918
rect 1416 131862 1472 131918
rect 1044 131738 1100 131794
rect 1168 131738 1224 131794
rect 1292 131738 1348 131794
rect 1416 131738 1472 131794
rect 1044 131614 1100 131670
rect 1168 131614 1224 131670
rect 1292 131614 1348 131670
rect 1416 131614 1472 131670
rect 1044 131490 1100 131546
rect 1168 131490 1224 131546
rect 1292 131490 1348 131546
rect 1416 131490 1472 131546
rect 1044 113862 1100 113918
rect 1168 113862 1224 113918
rect 1292 113862 1348 113918
rect 1416 113862 1472 113918
rect 1044 113738 1100 113794
rect 1168 113738 1224 113794
rect 1292 113738 1348 113794
rect 1416 113738 1472 113794
rect 1044 113614 1100 113670
rect 1168 113614 1224 113670
rect 1292 113614 1348 113670
rect 1416 113614 1472 113670
rect 1044 113490 1100 113546
rect 1168 113490 1224 113546
rect 1292 113490 1348 113546
rect 1416 113490 1472 113546
rect 1044 95862 1100 95918
rect 1168 95862 1224 95918
rect 1292 95862 1348 95918
rect 1416 95862 1472 95918
rect 1044 95738 1100 95794
rect 1168 95738 1224 95794
rect 1292 95738 1348 95794
rect 1416 95738 1472 95794
rect 1044 95614 1100 95670
rect 1168 95614 1224 95670
rect 1292 95614 1348 95670
rect 1416 95614 1472 95670
rect 1044 95490 1100 95546
rect 1168 95490 1224 95546
rect 1292 95490 1348 95546
rect 1416 95490 1472 95546
rect 1044 77862 1100 77918
rect 1168 77862 1224 77918
rect 1292 77862 1348 77918
rect 1416 77862 1472 77918
rect 1044 77738 1100 77794
rect 1168 77738 1224 77794
rect 1292 77738 1348 77794
rect 1416 77738 1472 77794
rect 1044 77614 1100 77670
rect 1168 77614 1224 77670
rect 1292 77614 1348 77670
rect 1416 77614 1472 77670
rect 1044 77490 1100 77546
rect 1168 77490 1224 77546
rect 1292 77490 1348 77546
rect 1416 77490 1472 77546
rect 1044 59862 1100 59918
rect 1168 59862 1224 59918
rect 1292 59862 1348 59918
rect 1416 59862 1472 59918
rect 1044 59738 1100 59794
rect 1168 59738 1224 59794
rect 1292 59738 1348 59794
rect 1416 59738 1472 59794
rect 1044 59614 1100 59670
rect 1168 59614 1224 59670
rect 1292 59614 1348 59670
rect 1416 59614 1472 59670
rect 1044 59490 1100 59546
rect 1168 59490 1224 59546
rect 1292 59490 1348 59546
rect 1416 59490 1472 59546
rect 1044 41862 1100 41918
rect 1168 41862 1224 41918
rect 1292 41862 1348 41918
rect 1416 41862 1472 41918
rect 1044 41738 1100 41794
rect 1168 41738 1224 41794
rect 1292 41738 1348 41794
rect 1416 41738 1472 41794
rect 1044 41614 1100 41670
rect 1168 41614 1224 41670
rect 1292 41614 1348 41670
rect 1416 41614 1472 41670
rect 1044 41490 1100 41546
rect 1168 41490 1224 41546
rect 1292 41490 1348 41546
rect 1416 41490 1472 41546
rect 1044 23862 1100 23918
rect 1168 23862 1224 23918
rect 1292 23862 1348 23918
rect 1416 23862 1472 23918
rect 1044 23738 1100 23794
rect 1168 23738 1224 23794
rect 1292 23738 1348 23794
rect 1416 23738 1472 23794
rect 1044 23614 1100 23670
rect 1168 23614 1224 23670
rect 1292 23614 1348 23670
rect 1416 23614 1472 23670
rect 1044 23490 1100 23546
rect 1168 23490 1224 23546
rect 1292 23490 1348 23546
rect 1416 23490 1472 23546
rect 1044 5862 1100 5918
rect 1168 5862 1224 5918
rect 1292 5862 1348 5918
rect 1416 5862 1472 5918
rect 1044 5738 1100 5794
rect 1168 5738 1224 5794
rect 1292 5738 1348 5794
rect 1416 5738 1472 5794
rect 1044 5614 1100 5670
rect 1168 5614 1224 5670
rect 1292 5614 1348 5670
rect 1416 5614 1472 5670
rect 1044 5490 1100 5546
rect 1168 5490 1224 5546
rect 1292 5490 1348 5546
rect 1416 5490 1472 5546
rect 1044 1752 1100 1808
rect 1168 1752 1224 1808
rect 1292 1752 1348 1808
rect 1416 1752 1472 1808
rect 1044 1628 1100 1684
rect 1168 1628 1224 1684
rect 1292 1628 1348 1684
rect 1416 1628 1472 1684
rect 1044 1504 1100 1560
rect 1168 1504 1224 1560
rect 1292 1504 1348 1560
rect 1416 1504 1472 1560
rect 1044 1380 1100 1436
rect 1168 1380 1224 1436
rect 1292 1380 1348 1436
rect 1416 1380 1472 1436
rect 5154 598324 5210 598380
rect 5278 598324 5334 598380
rect 5402 598324 5458 598380
rect 5526 598324 5582 598380
rect 5154 598200 5210 598256
rect 5278 598200 5334 598256
rect 5402 598200 5458 598256
rect 5526 598200 5582 598256
rect 5154 598076 5210 598132
rect 5278 598076 5334 598132
rect 5402 598076 5458 598132
rect 5526 598076 5582 598132
rect 5154 597952 5210 598008
rect 5278 597952 5334 598008
rect 5402 597952 5458 598008
rect 5526 597952 5582 598008
rect 8874 599284 8930 599340
rect 8998 599284 9054 599340
rect 9122 599284 9178 599340
rect 9246 599284 9302 599340
rect 8874 599160 8930 599216
rect 8998 599160 9054 599216
rect 9122 599160 9178 599216
rect 9246 599160 9302 599216
rect 8874 599036 8930 599092
rect 8998 599036 9054 599092
rect 9122 599036 9178 599092
rect 9246 599036 9302 599092
rect 8874 598912 8930 598968
rect 8998 598912 9054 598968
rect 9122 598912 9178 598968
rect 9246 598912 9302 598968
rect 23154 598324 23210 598380
rect 23278 598324 23334 598380
rect 23402 598324 23458 598380
rect 23526 598324 23582 598380
rect 23154 598200 23210 598256
rect 23278 598200 23334 598256
rect 23402 598200 23458 598256
rect 23526 598200 23582 598256
rect 23154 598076 23210 598132
rect 23278 598076 23334 598132
rect 23402 598076 23458 598132
rect 23526 598076 23582 598132
rect 23154 597952 23210 598008
rect 23278 597952 23334 598008
rect 23402 597952 23458 598008
rect 23526 597952 23582 598008
rect 26874 599284 26930 599340
rect 26998 599284 27054 599340
rect 27122 599284 27178 599340
rect 27246 599284 27302 599340
rect 26874 599160 26930 599216
rect 26998 599160 27054 599216
rect 27122 599160 27178 599216
rect 27246 599160 27302 599216
rect 26874 599036 26930 599092
rect 26998 599036 27054 599092
rect 27122 599036 27178 599092
rect 27246 599036 27302 599092
rect 26874 598912 26930 598968
rect 26998 598912 27054 598968
rect 27122 598912 27178 598968
rect 27246 598912 27302 598968
rect 41154 598324 41210 598380
rect 41278 598324 41334 598380
rect 41402 598324 41458 598380
rect 41526 598324 41582 598380
rect 41154 598200 41210 598256
rect 41278 598200 41334 598256
rect 41402 598200 41458 598256
rect 41526 598200 41582 598256
rect 41154 598076 41210 598132
rect 41278 598076 41334 598132
rect 41402 598076 41458 598132
rect 41526 598076 41582 598132
rect 41154 597952 41210 598008
rect 41278 597952 41334 598008
rect 41402 597952 41458 598008
rect 41526 597952 41582 598008
rect 44874 599284 44930 599340
rect 44998 599284 45054 599340
rect 45122 599284 45178 599340
rect 45246 599284 45302 599340
rect 44874 599160 44930 599216
rect 44998 599160 45054 599216
rect 45122 599160 45178 599216
rect 45246 599160 45302 599216
rect 44874 599036 44930 599092
rect 44998 599036 45054 599092
rect 45122 599036 45178 599092
rect 45246 599036 45302 599092
rect 44874 598912 44930 598968
rect 44998 598912 45054 598968
rect 45122 598912 45178 598968
rect 45246 598912 45302 598968
rect 59154 598324 59210 598380
rect 59278 598324 59334 598380
rect 59402 598324 59458 598380
rect 59526 598324 59582 598380
rect 59154 598200 59210 598256
rect 59278 598200 59334 598256
rect 59402 598200 59458 598256
rect 59526 598200 59582 598256
rect 59154 598076 59210 598132
rect 59278 598076 59334 598132
rect 59402 598076 59458 598132
rect 59526 598076 59582 598132
rect 59154 597952 59210 598008
rect 59278 597952 59334 598008
rect 59402 597952 59458 598008
rect 59526 597952 59582 598008
rect 62874 599284 62930 599340
rect 62998 599284 63054 599340
rect 63122 599284 63178 599340
rect 63246 599284 63302 599340
rect 62874 599160 62930 599216
rect 62998 599160 63054 599216
rect 63122 599160 63178 599216
rect 63246 599160 63302 599216
rect 62874 599036 62930 599092
rect 62998 599036 63054 599092
rect 63122 599036 63178 599092
rect 63246 599036 63302 599092
rect 62874 598912 62930 598968
rect 62998 598912 63054 598968
rect 63122 598912 63178 598968
rect 63246 598912 63302 598968
rect 77154 598324 77210 598380
rect 77278 598324 77334 598380
rect 77402 598324 77458 598380
rect 77526 598324 77582 598380
rect 77154 598200 77210 598256
rect 77278 598200 77334 598256
rect 77402 598200 77458 598256
rect 77526 598200 77582 598256
rect 77154 598076 77210 598132
rect 77278 598076 77334 598132
rect 77402 598076 77458 598132
rect 77526 598076 77582 598132
rect 77154 597952 77210 598008
rect 77278 597952 77334 598008
rect 77402 597952 77458 598008
rect 77526 597952 77582 598008
rect 80874 599284 80930 599340
rect 80998 599284 81054 599340
rect 81122 599284 81178 599340
rect 81246 599284 81302 599340
rect 80874 599160 80930 599216
rect 80998 599160 81054 599216
rect 81122 599160 81178 599216
rect 81246 599160 81302 599216
rect 80874 599036 80930 599092
rect 80998 599036 81054 599092
rect 81122 599036 81178 599092
rect 81246 599036 81302 599092
rect 80874 598912 80930 598968
rect 80998 598912 81054 598968
rect 81122 598912 81178 598968
rect 81246 598912 81302 598968
rect 95154 598324 95210 598380
rect 95278 598324 95334 598380
rect 95402 598324 95458 598380
rect 95526 598324 95582 598380
rect 95154 598200 95210 598256
rect 95278 598200 95334 598256
rect 95402 598200 95458 598256
rect 95526 598200 95582 598256
rect 95154 598076 95210 598132
rect 95278 598076 95334 598132
rect 95402 598076 95458 598132
rect 95526 598076 95582 598132
rect 95154 597952 95210 598008
rect 95278 597952 95334 598008
rect 95402 597952 95458 598008
rect 95526 597952 95582 598008
rect 98874 599284 98930 599340
rect 98998 599284 99054 599340
rect 99122 599284 99178 599340
rect 99246 599284 99302 599340
rect 98874 599160 98930 599216
rect 98998 599160 99054 599216
rect 99122 599160 99178 599216
rect 99246 599160 99302 599216
rect 98874 599036 98930 599092
rect 98998 599036 99054 599092
rect 99122 599036 99178 599092
rect 99246 599036 99302 599092
rect 98874 598912 98930 598968
rect 98998 598912 99054 598968
rect 99122 598912 99178 598968
rect 99246 598912 99302 598968
rect 113154 598324 113210 598380
rect 113278 598324 113334 598380
rect 113402 598324 113458 598380
rect 113526 598324 113582 598380
rect 113154 598200 113210 598256
rect 113278 598200 113334 598256
rect 113402 598200 113458 598256
rect 113526 598200 113582 598256
rect 113154 598076 113210 598132
rect 113278 598076 113334 598132
rect 113402 598076 113458 598132
rect 113526 598076 113582 598132
rect 113154 597952 113210 598008
rect 113278 597952 113334 598008
rect 113402 597952 113458 598008
rect 113526 597952 113582 598008
rect 116874 599284 116930 599340
rect 116998 599284 117054 599340
rect 117122 599284 117178 599340
rect 117246 599284 117302 599340
rect 116874 599160 116930 599216
rect 116998 599160 117054 599216
rect 117122 599160 117178 599216
rect 117246 599160 117302 599216
rect 116874 599036 116930 599092
rect 116998 599036 117054 599092
rect 117122 599036 117178 599092
rect 117246 599036 117302 599092
rect 116874 598912 116930 598968
rect 116998 598912 117054 598968
rect 117122 598912 117178 598968
rect 117246 598912 117302 598968
rect 131154 598324 131210 598380
rect 131278 598324 131334 598380
rect 131402 598324 131458 598380
rect 131526 598324 131582 598380
rect 131154 598200 131210 598256
rect 131278 598200 131334 598256
rect 131402 598200 131458 598256
rect 131526 598200 131582 598256
rect 131154 598076 131210 598132
rect 131278 598076 131334 598132
rect 131402 598076 131458 598132
rect 131526 598076 131582 598132
rect 131154 597952 131210 598008
rect 131278 597952 131334 598008
rect 131402 597952 131458 598008
rect 131526 597952 131582 598008
rect 134874 599284 134930 599340
rect 134998 599284 135054 599340
rect 135122 599284 135178 599340
rect 135246 599284 135302 599340
rect 134874 599160 134930 599216
rect 134998 599160 135054 599216
rect 135122 599160 135178 599216
rect 135246 599160 135302 599216
rect 134874 599036 134930 599092
rect 134998 599036 135054 599092
rect 135122 599036 135178 599092
rect 135246 599036 135302 599092
rect 134874 598912 134930 598968
rect 134998 598912 135054 598968
rect 135122 598912 135178 598968
rect 135246 598912 135302 598968
rect 149154 598324 149210 598380
rect 149278 598324 149334 598380
rect 149402 598324 149458 598380
rect 149526 598324 149582 598380
rect 149154 598200 149210 598256
rect 149278 598200 149334 598256
rect 149402 598200 149458 598256
rect 149526 598200 149582 598256
rect 149154 598076 149210 598132
rect 149278 598076 149334 598132
rect 149402 598076 149458 598132
rect 149526 598076 149582 598132
rect 149154 597952 149210 598008
rect 149278 597952 149334 598008
rect 149402 597952 149458 598008
rect 149526 597952 149582 598008
rect 152874 599284 152930 599340
rect 152998 599284 153054 599340
rect 153122 599284 153178 599340
rect 153246 599284 153302 599340
rect 152874 599160 152930 599216
rect 152998 599160 153054 599216
rect 153122 599160 153178 599216
rect 153246 599160 153302 599216
rect 152874 599036 152930 599092
rect 152998 599036 153054 599092
rect 153122 599036 153178 599092
rect 153246 599036 153302 599092
rect 152874 598912 152930 598968
rect 152998 598912 153054 598968
rect 153122 598912 153178 598968
rect 153246 598912 153302 598968
rect 167154 598324 167210 598380
rect 167278 598324 167334 598380
rect 167402 598324 167458 598380
rect 167526 598324 167582 598380
rect 167154 598200 167210 598256
rect 167278 598200 167334 598256
rect 167402 598200 167458 598256
rect 167526 598200 167582 598256
rect 167154 598076 167210 598132
rect 167278 598076 167334 598132
rect 167402 598076 167458 598132
rect 167526 598076 167582 598132
rect 167154 597952 167210 598008
rect 167278 597952 167334 598008
rect 167402 597952 167458 598008
rect 167526 597952 167582 598008
rect 170874 599284 170930 599340
rect 170998 599284 171054 599340
rect 171122 599284 171178 599340
rect 171246 599284 171302 599340
rect 170874 599160 170930 599216
rect 170998 599160 171054 599216
rect 171122 599160 171178 599216
rect 171246 599160 171302 599216
rect 170874 599036 170930 599092
rect 170998 599036 171054 599092
rect 171122 599036 171178 599092
rect 171246 599036 171302 599092
rect 170874 598912 170930 598968
rect 170998 598912 171054 598968
rect 171122 598912 171178 598968
rect 171246 598912 171302 598968
rect 185154 598324 185210 598380
rect 185278 598324 185334 598380
rect 185402 598324 185458 598380
rect 185526 598324 185582 598380
rect 185154 598200 185210 598256
rect 185278 598200 185334 598256
rect 185402 598200 185458 598256
rect 185526 598200 185582 598256
rect 185154 598076 185210 598132
rect 185278 598076 185334 598132
rect 185402 598076 185458 598132
rect 185526 598076 185582 598132
rect 185154 597952 185210 598008
rect 185278 597952 185334 598008
rect 185402 597952 185458 598008
rect 185526 597952 185582 598008
rect 188874 599284 188930 599340
rect 188998 599284 189054 599340
rect 189122 599284 189178 599340
rect 189246 599284 189302 599340
rect 188874 599160 188930 599216
rect 188998 599160 189054 599216
rect 189122 599160 189178 599216
rect 189246 599160 189302 599216
rect 188874 599036 188930 599092
rect 188998 599036 189054 599092
rect 189122 599036 189178 599092
rect 189246 599036 189302 599092
rect 188874 598912 188930 598968
rect 188998 598912 189054 598968
rect 189122 598912 189178 598968
rect 189246 598912 189302 598968
rect 203154 598324 203210 598380
rect 203278 598324 203334 598380
rect 203402 598324 203458 598380
rect 203526 598324 203582 598380
rect 203154 598200 203210 598256
rect 203278 598200 203334 598256
rect 203402 598200 203458 598256
rect 203526 598200 203582 598256
rect 203154 598076 203210 598132
rect 203278 598076 203334 598132
rect 203402 598076 203458 598132
rect 203526 598076 203582 598132
rect 203154 597952 203210 598008
rect 203278 597952 203334 598008
rect 203402 597952 203458 598008
rect 203526 597952 203582 598008
rect 206874 599284 206930 599340
rect 206998 599284 207054 599340
rect 207122 599284 207178 599340
rect 207246 599284 207302 599340
rect 206874 599160 206930 599216
rect 206998 599160 207054 599216
rect 207122 599160 207178 599216
rect 207246 599160 207302 599216
rect 206874 599036 206930 599092
rect 206998 599036 207054 599092
rect 207122 599036 207178 599092
rect 207246 599036 207302 599092
rect 206874 598912 206930 598968
rect 206998 598912 207054 598968
rect 207122 598912 207178 598968
rect 207246 598912 207302 598968
rect 221154 598324 221210 598380
rect 221278 598324 221334 598380
rect 221402 598324 221458 598380
rect 221526 598324 221582 598380
rect 221154 598200 221210 598256
rect 221278 598200 221334 598256
rect 221402 598200 221458 598256
rect 221526 598200 221582 598256
rect 221154 598076 221210 598132
rect 221278 598076 221334 598132
rect 221402 598076 221458 598132
rect 221526 598076 221582 598132
rect 221154 597952 221210 598008
rect 221278 597952 221334 598008
rect 221402 597952 221458 598008
rect 221526 597952 221582 598008
rect 224874 599284 224930 599340
rect 224998 599284 225054 599340
rect 225122 599284 225178 599340
rect 225246 599284 225302 599340
rect 224874 599160 224930 599216
rect 224998 599160 225054 599216
rect 225122 599160 225178 599216
rect 225246 599160 225302 599216
rect 224874 599036 224930 599092
rect 224998 599036 225054 599092
rect 225122 599036 225178 599092
rect 225246 599036 225302 599092
rect 224874 598912 224930 598968
rect 224998 598912 225054 598968
rect 225122 598912 225178 598968
rect 225246 598912 225302 598968
rect 239154 598324 239210 598380
rect 239278 598324 239334 598380
rect 239402 598324 239458 598380
rect 239526 598324 239582 598380
rect 239154 598200 239210 598256
rect 239278 598200 239334 598256
rect 239402 598200 239458 598256
rect 239526 598200 239582 598256
rect 239154 598076 239210 598132
rect 239278 598076 239334 598132
rect 239402 598076 239458 598132
rect 239526 598076 239582 598132
rect 239154 597952 239210 598008
rect 239278 597952 239334 598008
rect 239402 597952 239458 598008
rect 239526 597952 239582 598008
rect 242874 599284 242930 599340
rect 242998 599284 243054 599340
rect 243122 599284 243178 599340
rect 243246 599284 243302 599340
rect 242874 599160 242930 599216
rect 242998 599160 243054 599216
rect 243122 599160 243178 599216
rect 243246 599160 243302 599216
rect 242874 599036 242930 599092
rect 242998 599036 243054 599092
rect 243122 599036 243178 599092
rect 243246 599036 243302 599092
rect 242874 598912 242930 598968
rect 242998 598912 243054 598968
rect 243122 598912 243178 598968
rect 243246 598912 243302 598968
rect 257154 598324 257210 598380
rect 257278 598324 257334 598380
rect 257402 598324 257458 598380
rect 257526 598324 257582 598380
rect 257154 598200 257210 598256
rect 257278 598200 257334 598256
rect 257402 598200 257458 598256
rect 257526 598200 257582 598256
rect 257154 598076 257210 598132
rect 257278 598076 257334 598132
rect 257402 598076 257458 598132
rect 257526 598076 257582 598132
rect 257154 597952 257210 598008
rect 257278 597952 257334 598008
rect 257402 597952 257458 598008
rect 257526 597952 257582 598008
rect 260874 599284 260930 599340
rect 260998 599284 261054 599340
rect 261122 599284 261178 599340
rect 261246 599284 261302 599340
rect 260874 599160 260930 599216
rect 260998 599160 261054 599216
rect 261122 599160 261178 599216
rect 261246 599160 261302 599216
rect 260874 599036 260930 599092
rect 260998 599036 261054 599092
rect 261122 599036 261178 599092
rect 261246 599036 261302 599092
rect 260874 598912 260930 598968
rect 260998 598912 261054 598968
rect 261122 598912 261178 598968
rect 261246 598912 261302 598968
rect 275154 598324 275210 598380
rect 275278 598324 275334 598380
rect 275402 598324 275458 598380
rect 275526 598324 275582 598380
rect 275154 598200 275210 598256
rect 275278 598200 275334 598256
rect 275402 598200 275458 598256
rect 275526 598200 275582 598256
rect 275154 598076 275210 598132
rect 275278 598076 275334 598132
rect 275402 598076 275458 598132
rect 275526 598076 275582 598132
rect 275154 597952 275210 598008
rect 275278 597952 275334 598008
rect 275402 597952 275458 598008
rect 275526 597952 275582 598008
rect 278874 599284 278930 599340
rect 278998 599284 279054 599340
rect 279122 599284 279178 599340
rect 279246 599284 279302 599340
rect 278874 599160 278930 599216
rect 278998 599160 279054 599216
rect 279122 599160 279178 599216
rect 279246 599160 279302 599216
rect 278874 599036 278930 599092
rect 278998 599036 279054 599092
rect 279122 599036 279178 599092
rect 279246 599036 279302 599092
rect 278874 598912 278930 598968
rect 278998 598912 279054 598968
rect 279122 598912 279178 598968
rect 279246 598912 279302 598968
rect 293154 598324 293210 598380
rect 293278 598324 293334 598380
rect 293402 598324 293458 598380
rect 293526 598324 293582 598380
rect 293154 598200 293210 598256
rect 293278 598200 293334 598256
rect 293402 598200 293458 598256
rect 293526 598200 293582 598256
rect 293154 598076 293210 598132
rect 293278 598076 293334 598132
rect 293402 598076 293458 598132
rect 293526 598076 293582 598132
rect 293154 597952 293210 598008
rect 293278 597952 293334 598008
rect 293402 597952 293458 598008
rect 293526 597952 293582 598008
rect 296874 599284 296930 599340
rect 296998 599284 297054 599340
rect 297122 599284 297178 599340
rect 297246 599284 297302 599340
rect 296874 599160 296930 599216
rect 296998 599160 297054 599216
rect 297122 599160 297178 599216
rect 297246 599160 297302 599216
rect 296874 599036 296930 599092
rect 296998 599036 297054 599092
rect 297122 599036 297178 599092
rect 297246 599036 297302 599092
rect 296874 598912 296930 598968
rect 296998 598912 297054 598968
rect 297122 598912 297178 598968
rect 297246 598912 297302 598968
rect 311154 598324 311210 598380
rect 311278 598324 311334 598380
rect 311402 598324 311458 598380
rect 311526 598324 311582 598380
rect 311154 598200 311210 598256
rect 311278 598200 311334 598256
rect 311402 598200 311458 598256
rect 311526 598200 311582 598256
rect 311154 598076 311210 598132
rect 311278 598076 311334 598132
rect 311402 598076 311458 598132
rect 311526 598076 311582 598132
rect 311154 597952 311210 598008
rect 311278 597952 311334 598008
rect 311402 597952 311458 598008
rect 311526 597952 311582 598008
rect 314874 599284 314930 599340
rect 314998 599284 315054 599340
rect 315122 599284 315178 599340
rect 315246 599284 315302 599340
rect 314874 599160 314930 599216
rect 314998 599160 315054 599216
rect 315122 599160 315178 599216
rect 315246 599160 315302 599216
rect 314874 599036 314930 599092
rect 314998 599036 315054 599092
rect 315122 599036 315178 599092
rect 315246 599036 315302 599092
rect 314874 598912 314930 598968
rect 314998 598912 315054 598968
rect 315122 598912 315178 598968
rect 315246 598912 315302 598968
rect 329154 598324 329210 598380
rect 329278 598324 329334 598380
rect 329402 598324 329458 598380
rect 329526 598324 329582 598380
rect 329154 598200 329210 598256
rect 329278 598200 329334 598256
rect 329402 598200 329458 598256
rect 329526 598200 329582 598256
rect 329154 598076 329210 598132
rect 329278 598076 329334 598132
rect 329402 598076 329458 598132
rect 329526 598076 329582 598132
rect 329154 597952 329210 598008
rect 329278 597952 329334 598008
rect 329402 597952 329458 598008
rect 329526 597952 329582 598008
rect 332874 599284 332930 599340
rect 332998 599284 333054 599340
rect 333122 599284 333178 599340
rect 333246 599284 333302 599340
rect 332874 599160 332930 599216
rect 332998 599160 333054 599216
rect 333122 599160 333178 599216
rect 333246 599160 333302 599216
rect 332874 599036 332930 599092
rect 332998 599036 333054 599092
rect 333122 599036 333178 599092
rect 333246 599036 333302 599092
rect 332874 598912 332930 598968
rect 332998 598912 333054 598968
rect 333122 598912 333178 598968
rect 333246 598912 333302 598968
rect 347154 598324 347210 598380
rect 347278 598324 347334 598380
rect 347402 598324 347458 598380
rect 347526 598324 347582 598380
rect 347154 598200 347210 598256
rect 347278 598200 347334 598256
rect 347402 598200 347458 598256
rect 347526 598200 347582 598256
rect 347154 598076 347210 598132
rect 347278 598076 347334 598132
rect 347402 598076 347458 598132
rect 347526 598076 347582 598132
rect 347154 597952 347210 598008
rect 347278 597952 347334 598008
rect 347402 597952 347458 598008
rect 347526 597952 347582 598008
rect 350874 599284 350930 599340
rect 350998 599284 351054 599340
rect 351122 599284 351178 599340
rect 351246 599284 351302 599340
rect 350874 599160 350930 599216
rect 350998 599160 351054 599216
rect 351122 599160 351178 599216
rect 351246 599160 351302 599216
rect 350874 599036 350930 599092
rect 350998 599036 351054 599092
rect 351122 599036 351178 599092
rect 351246 599036 351302 599092
rect 350874 598912 350930 598968
rect 350998 598912 351054 598968
rect 351122 598912 351178 598968
rect 351246 598912 351302 598968
rect 365154 598324 365210 598380
rect 365278 598324 365334 598380
rect 365402 598324 365458 598380
rect 365526 598324 365582 598380
rect 365154 598200 365210 598256
rect 365278 598200 365334 598256
rect 365402 598200 365458 598256
rect 365526 598200 365582 598256
rect 365154 598076 365210 598132
rect 365278 598076 365334 598132
rect 365402 598076 365458 598132
rect 365526 598076 365582 598132
rect 365154 597952 365210 598008
rect 365278 597952 365334 598008
rect 365402 597952 365458 598008
rect 365526 597952 365582 598008
rect 368874 599284 368930 599340
rect 368998 599284 369054 599340
rect 369122 599284 369178 599340
rect 369246 599284 369302 599340
rect 368874 599160 368930 599216
rect 368998 599160 369054 599216
rect 369122 599160 369178 599216
rect 369246 599160 369302 599216
rect 368874 599036 368930 599092
rect 368998 599036 369054 599092
rect 369122 599036 369178 599092
rect 369246 599036 369302 599092
rect 368874 598912 368930 598968
rect 368998 598912 369054 598968
rect 369122 598912 369178 598968
rect 369246 598912 369302 598968
rect 383154 598324 383210 598380
rect 383278 598324 383334 598380
rect 383402 598324 383458 598380
rect 383526 598324 383582 598380
rect 383154 598200 383210 598256
rect 383278 598200 383334 598256
rect 383402 598200 383458 598256
rect 383526 598200 383582 598256
rect 383154 598076 383210 598132
rect 383278 598076 383334 598132
rect 383402 598076 383458 598132
rect 383526 598076 383582 598132
rect 383154 597952 383210 598008
rect 383278 597952 383334 598008
rect 383402 597952 383458 598008
rect 383526 597952 383582 598008
rect 386874 599284 386930 599340
rect 386998 599284 387054 599340
rect 387122 599284 387178 599340
rect 387246 599284 387302 599340
rect 386874 599160 386930 599216
rect 386998 599160 387054 599216
rect 387122 599160 387178 599216
rect 387246 599160 387302 599216
rect 386874 599036 386930 599092
rect 386998 599036 387054 599092
rect 387122 599036 387178 599092
rect 387246 599036 387302 599092
rect 386874 598912 386930 598968
rect 386998 598912 387054 598968
rect 387122 598912 387178 598968
rect 387246 598912 387302 598968
rect 401154 598324 401210 598380
rect 401278 598324 401334 598380
rect 401402 598324 401458 598380
rect 401526 598324 401582 598380
rect 401154 598200 401210 598256
rect 401278 598200 401334 598256
rect 401402 598200 401458 598256
rect 401526 598200 401582 598256
rect 401154 598076 401210 598132
rect 401278 598076 401334 598132
rect 401402 598076 401458 598132
rect 401526 598076 401582 598132
rect 401154 597952 401210 598008
rect 401278 597952 401334 598008
rect 401402 597952 401458 598008
rect 401526 597952 401582 598008
rect 404874 599284 404930 599340
rect 404998 599284 405054 599340
rect 405122 599284 405178 599340
rect 405246 599284 405302 599340
rect 404874 599160 404930 599216
rect 404998 599160 405054 599216
rect 405122 599160 405178 599216
rect 405246 599160 405302 599216
rect 404874 599036 404930 599092
rect 404998 599036 405054 599092
rect 405122 599036 405178 599092
rect 405246 599036 405302 599092
rect 404874 598912 404930 598968
rect 404998 598912 405054 598968
rect 405122 598912 405178 598968
rect 405246 598912 405302 598968
rect 419154 598324 419210 598380
rect 419278 598324 419334 598380
rect 419402 598324 419458 598380
rect 419526 598324 419582 598380
rect 419154 598200 419210 598256
rect 419278 598200 419334 598256
rect 419402 598200 419458 598256
rect 419526 598200 419582 598256
rect 419154 598076 419210 598132
rect 419278 598076 419334 598132
rect 419402 598076 419458 598132
rect 419526 598076 419582 598132
rect 419154 597952 419210 598008
rect 419278 597952 419334 598008
rect 419402 597952 419458 598008
rect 419526 597952 419582 598008
rect 422874 599284 422930 599340
rect 422998 599284 423054 599340
rect 423122 599284 423178 599340
rect 423246 599284 423302 599340
rect 422874 599160 422930 599216
rect 422998 599160 423054 599216
rect 423122 599160 423178 599216
rect 423246 599160 423302 599216
rect 422874 599036 422930 599092
rect 422998 599036 423054 599092
rect 423122 599036 423178 599092
rect 423246 599036 423302 599092
rect 422874 598912 422930 598968
rect 422998 598912 423054 598968
rect 423122 598912 423178 598968
rect 423246 598912 423302 598968
rect 437154 598324 437210 598380
rect 437278 598324 437334 598380
rect 437402 598324 437458 598380
rect 437526 598324 437582 598380
rect 437154 598200 437210 598256
rect 437278 598200 437334 598256
rect 437402 598200 437458 598256
rect 437526 598200 437582 598256
rect 437154 598076 437210 598132
rect 437278 598076 437334 598132
rect 437402 598076 437458 598132
rect 437526 598076 437582 598132
rect 437154 597952 437210 598008
rect 437278 597952 437334 598008
rect 437402 597952 437458 598008
rect 437526 597952 437582 598008
rect 440874 599284 440930 599340
rect 440998 599284 441054 599340
rect 441122 599284 441178 599340
rect 441246 599284 441302 599340
rect 440874 599160 440930 599216
rect 440998 599160 441054 599216
rect 441122 599160 441178 599216
rect 441246 599160 441302 599216
rect 440874 599036 440930 599092
rect 440998 599036 441054 599092
rect 441122 599036 441178 599092
rect 441246 599036 441302 599092
rect 440874 598912 440930 598968
rect 440998 598912 441054 598968
rect 441122 598912 441178 598968
rect 441246 598912 441302 598968
rect 455154 598324 455210 598380
rect 455278 598324 455334 598380
rect 455402 598324 455458 598380
rect 455526 598324 455582 598380
rect 455154 598200 455210 598256
rect 455278 598200 455334 598256
rect 455402 598200 455458 598256
rect 455526 598200 455582 598256
rect 455154 598076 455210 598132
rect 455278 598076 455334 598132
rect 455402 598076 455458 598132
rect 455526 598076 455582 598132
rect 455154 597952 455210 598008
rect 455278 597952 455334 598008
rect 455402 597952 455458 598008
rect 455526 597952 455582 598008
rect 458874 599284 458930 599340
rect 458998 599284 459054 599340
rect 459122 599284 459178 599340
rect 459246 599284 459302 599340
rect 458874 599160 458930 599216
rect 458998 599160 459054 599216
rect 459122 599160 459178 599216
rect 459246 599160 459302 599216
rect 458874 599036 458930 599092
rect 458998 599036 459054 599092
rect 459122 599036 459178 599092
rect 459246 599036 459302 599092
rect 458874 598912 458930 598968
rect 458998 598912 459054 598968
rect 459122 598912 459178 598968
rect 459246 598912 459302 598968
rect 473154 598324 473210 598380
rect 473278 598324 473334 598380
rect 473402 598324 473458 598380
rect 473526 598324 473582 598380
rect 473154 598200 473210 598256
rect 473278 598200 473334 598256
rect 473402 598200 473458 598256
rect 473526 598200 473582 598256
rect 473154 598076 473210 598132
rect 473278 598076 473334 598132
rect 473402 598076 473458 598132
rect 473526 598076 473582 598132
rect 473154 597952 473210 598008
rect 473278 597952 473334 598008
rect 473402 597952 473458 598008
rect 473526 597952 473582 598008
rect 476874 599284 476930 599340
rect 476998 599284 477054 599340
rect 477122 599284 477178 599340
rect 477246 599284 477302 599340
rect 476874 599160 476930 599216
rect 476998 599160 477054 599216
rect 477122 599160 477178 599216
rect 477246 599160 477302 599216
rect 476874 599036 476930 599092
rect 476998 599036 477054 599092
rect 477122 599036 477178 599092
rect 477246 599036 477302 599092
rect 476874 598912 476930 598968
rect 476998 598912 477054 598968
rect 477122 598912 477178 598968
rect 477246 598912 477302 598968
rect 491154 598324 491210 598380
rect 491278 598324 491334 598380
rect 491402 598324 491458 598380
rect 491526 598324 491582 598380
rect 491154 598200 491210 598256
rect 491278 598200 491334 598256
rect 491402 598200 491458 598256
rect 491526 598200 491582 598256
rect 491154 598076 491210 598132
rect 491278 598076 491334 598132
rect 491402 598076 491458 598132
rect 491526 598076 491582 598132
rect 491154 597952 491210 598008
rect 491278 597952 491334 598008
rect 491402 597952 491458 598008
rect 491526 597952 491582 598008
rect 494874 599284 494930 599340
rect 494998 599284 495054 599340
rect 495122 599284 495178 599340
rect 495246 599284 495302 599340
rect 494874 599160 494930 599216
rect 494998 599160 495054 599216
rect 495122 599160 495178 599216
rect 495246 599160 495302 599216
rect 494874 599036 494930 599092
rect 494998 599036 495054 599092
rect 495122 599036 495178 599092
rect 495246 599036 495302 599092
rect 494874 598912 494930 598968
rect 494998 598912 495054 598968
rect 495122 598912 495178 598968
rect 495246 598912 495302 598968
rect 509154 598324 509210 598380
rect 509278 598324 509334 598380
rect 509402 598324 509458 598380
rect 509526 598324 509582 598380
rect 509154 598200 509210 598256
rect 509278 598200 509334 598256
rect 509402 598200 509458 598256
rect 509526 598200 509582 598256
rect 509154 598076 509210 598132
rect 509278 598076 509334 598132
rect 509402 598076 509458 598132
rect 509526 598076 509582 598132
rect 509154 597952 509210 598008
rect 509278 597952 509334 598008
rect 509402 597952 509458 598008
rect 509526 597952 509582 598008
rect 512874 599284 512930 599340
rect 512998 599284 513054 599340
rect 513122 599284 513178 599340
rect 513246 599284 513302 599340
rect 512874 599160 512930 599216
rect 512998 599160 513054 599216
rect 513122 599160 513178 599216
rect 513246 599160 513302 599216
rect 512874 599036 512930 599092
rect 512998 599036 513054 599092
rect 513122 599036 513178 599092
rect 513246 599036 513302 599092
rect 512874 598912 512930 598968
rect 512998 598912 513054 598968
rect 513122 598912 513178 598968
rect 513246 598912 513302 598968
rect 527154 598324 527210 598380
rect 527278 598324 527334 598380
rect 527402 598324 527458 598380
rect 527526 598324 527582 598380
rect 527154 598200 527210 598256
rect 527278 598200 527334 598256
rect 527402 598200 527458 598256
rect 527526 598200 527582 598256
rect 527154 598076 527210 598132
rect 527278 598076 527334 598132
rect 527402 598076 527458 598132
rect 527526 598076 527582 598132
rect 527154 597952 527210 598008
rect 527278 597952 527334 598008
rect 527402 597952 527458 598008
rect 527526 597952 527582 598008
rect 530874 599284 530930 599340
rect 530998 599284 531054 599340
rect 531122 599284 531178 599340
rect 531246 599284 531302 599340
rect 530874 599160 530930 599216
rect 530998 599160 531054 599216
rect 531122 599160 531178 599216
rect 531246 599160 531302 599216
rect 530874 599036 530930 599092
rect 530998 599036 531054 599092
rect 531122 599036 531178 599092
rect 531246 599036 531302 599092
rect 530874 598912 530930 598968
rect 530998 598912 531054 598968
rect 531122 598912 531178 598968
rect 531246 598912 531302 598968
rect 545154 598324 545210 598380
rect 545278 598324 545334 598380
rect 545402 598324 545458 598380
rect 545526 598324 545582 598380
rect 545154 598200 545210 598256
rect 545278 598200 545334 598256
rect 545402 598200 545458 598256
rect 545526 598200 545582 598256
rect 545154 598076 545210 598132
rect 545278 598076 545334 598132
rect 545402 598076 545458 598132
rect 545526 598076 545582 598132
rect 545154 597952 545210 598008
rect 545278 597952 545334 598008
rect 545402 597952 545458 598008
rect 545526 597952 545582 598008
rect 548874 599284 548930 599340
rect 548998 599284 549054 599340
rect 549122 599284 549178 599340
rect 549246 599284 549302 599340
rect 548874 599160 548930 599216
rect 548998 599160 549054 599216
rect 549122 599160 549178 599216
rect 549246 599160 549302 599216
rect 548874 599036 548930 599092
rect 548998 599036 549054 599092
rect 549122 599036 549178 599092
rect 549246 599036 549302 599092
rect 548874 598912 548930 598968
rect 548998 598912 549054 598968
rect 549122 598912 549178 598968
rect 549246 598912 549302 598968
rect 563154 598324 563210 598380
rect 563278 598324 563334 598380
rect 563402 598324 563458 598380
rect 563526 598324 563582 598380
rect 563154 598200 563210 598256
rect 563278 598200 563334 598256
rect 563402 598200 563458 598256
rect 563526 598200 563582 598256
rect 563154 598076 563210 598132
rect 563278 598076 563334 598132
rect 563402 598076 563458 598132
rect 563526 598076 563582 598132
rect 563154 597952 563210 598008
rect 563278 597952 563334 598008
rect 563402 597952 563458 598008
rect 563526 597952 563582 598008
rect 566874 599284 566930 599340
rect 566998 599284 567054 599340
rect 567122 599284 567178 599340
rect 567246 599284 567302 599340
rect 566874 599160 566930 599216
rect 566998 599160 567054 599216
rect 567122 599160 567178 599216
rect 567246 599160 567302 599216
rect 566874 599036 566930 599092
rect 566998 599036 567054 599092
rect 567122 599036 567178 599092
rect 567246 599036 567302 599092
rect 566874 598912 566930 598968
rect 566998 598912 567054 598968
rect 567122 598912 567178 598968
rect 567246 598912 567302 598968
rect 581154 598324 581210 598380
rect 581278 598324 581334 598380
rect 581402 598324 581458 598380
rect 581526 598324 581582 598380
rect 581154 598200 581210 598256
rect 581278 598200 581334 598256
rect 581402 598200 581458 598256
rect 581526 598200 581582 598256
rect 581154 598076 581210 598132
rect 581278 598076 581334 598132
rect 581402 598076 581458 598132
rect 581526 598076 581582 598132
rect 581154 597952 581210 598008
rect 581278 597952 581334 598008
rect 581402 597952 581458 598008
rect 581526 597952 581582 598008
rect 584874 599284 584930 599340
rect 584998 599284 585054 599340
rect 585122 599284 585178 599340
rect 585246 599284 585302 599340
rect 584874 599160 584930 599216
rect 584998 599160 585054 599216
rect 585122 599160 585178 599216
rect 585246 599160 585302 599216
rect 584874 599036 584930 599092
rect 584998 599036 585054 599092
rect 585122 599036 585178 599092
rect 585246 599036 585302 599092
rect 584874 598912 584930 598968
rect 584998 598912 585054 598968
rect 585122 598912 585178 598968
rect 585246 598912 585302 598968
rect 599472 599284 599528 599340
rect 599596 599284 599652 599340
rect 599720 599284 599776 599340
rect 599844 599284 599900 599340
rect 599472 599160 599528 599216
rect 599596 599160 599652 599216
rect 599720 599160 599776 599216
rect 599844 599160 599900 599216
rect 599472 599036 599528 599092
rect 599596 599036 599652 599092
rect 599720 599036 599776 599092
rect 599844 599036 599900 599092
rect 599472 598912 599528 598968
rect 599596 598912 599652 598968
rect 599720 598912 599776 598968
rect 599844 598912 599900 598968
rect 598512 598324 598568 598380
rect 598636 598324 598692 598380
rect 598760 598324 598816 598380
rect 598884 598324 598940 598380
rect 598512 598200 598568 598256
rect 598636 598200 598692 598256
rect 598760 598200 598816 598256
rect 598884 598200 598940 598256
rect 598512 598076 598568 598132
rect 598636 598076 598692 598132
rect 598760 598076 598816 598132
rect 598884 598076 598940 598132
rect 598512 597952 598568 598008
rect 598636 597952 598692 598008
rect 598760 597952 598816 598008
rect 598884 597952 598940 598008
rect 5154 581862 5210 581918
rect 5278 581862 5334 581918
rect 5402 581862 5458 581918
rect 5526 581862 5582 581918
rect 5154 581738 5210 581794
rect 5278 581738 5334 581794
rect 5402 581738 5458 581794
rect 5526 581738 5582 581794
rect 5154 581614 5210 581670
rect 5278 581614 5334 581670
rect 5402 581614 5458 581670
rect 5526 581614 5582 581670
rect 5154 581490 5210 581546
rect 5278 581490 5334 581546
rect 5402 581490 5458 581546
rect 5526 581490 5582 581546
rect 5154 563862 5210 563918
rect 5278 563862 5334 563918
rect 5402 563862 5458 563918
rect 5526 563862 5582 563918
rect 5154 563738 5210 563794
rect 5278 563738 5334 563794
rect 5402 563738 5458 563794
rect 5526 563738 5582 563794
rect 5154 563614 5210 563670
rect 5278 563614 5334 563670
rect 5402 563614 5458 563670
rect 5526 563614 5582 563670
rect 5154 563490 5210 563546
rect 5278 563490 5334 563546
rect 5402 563490 5458 563546
rect 5526 563490 5582 563546
rect 5154 545862 5210 545918
rect 5278 545862 5334 545918
rect 5402 545862 5458 545918
rect 5526 545862 5582 545918
rect 5154 545738 5210 545794
rect 5278 545738 5334 545794
rect 5402 545738 5458 545794
rect 5526 545738 5582 545794
rect 5154 545614 5210 545670
rect 5278 545614 5334 545670
rect 5402 545614 5458 545670
rect 5526 545614 5582 545670
rect 5154 545490 5210 545546
rect 5278 545490 5334 545546
rect 5402 545490 5458 545546
rect 5526 545490 5582 545546
rect 5154 527862 5210 527918
rect 5278 527862 5334 527918
rect 5402 527862 5458 527918
rect 5526 527862 5582 527918
rect 5154 527738 5210 527794
rect 5278 527738 5334 527794
rect 5402 527738 5458 527794
rect 5526 527738 5582 527794
rect 5154 527614 5210 527670
rect 5278 527614 5334 527670
rect 5402 527614 5458 527670
rect 5526 527614 5582 527670
rect 5154 527490 5210 527546
rect 5278 527490 5334 527546
rect 5402 527490 5458 527546
rect 5526 527490 5582 527546
rect 5154 509862 5210 509918
rect 5278 509862 5334 509918
rect 5402 509862 5458 509918
rect 5526 509862 5582 509918
rect 5154 509738 5210 509794
rect 5278 509738 5334 509794
rect 5402 509738 5458 509794
rect 5526 509738 5582 509794
rect 5154 509614 5210 509670
rect 5278 509614 5334 509670
rect 5402 509614 5458 509670
rect 5526 509614 5582 509670
rect 5154 509490 5210 509546
rect 5278 509490 5334 509546
rect 5402 509490 5458 509546
rect 5526 509490 5582 509546
rect 5154 491862 5210 491918
rect 5278 491862 5334 491918
rect 5402 491862 5458 491918
rect 5526 491862 5582 491918
rect 5154 491738 5210 491794
rect 5278 491738 5334 491794
rect 5402 491738 5458 491794
rect 5526 491738 5582 491794
rect 5154 491614 5210 491670
rect 5278 491614 5334 491670
rect 5402 491614 5458 491670
rect 5526 491614 5582 491670
rect 5154 491490 5210 491546
rect 5278 491490 5334 491546
rect 5402 491490 5458 491546
rect 5526 491490 5582 491546
rect 5154 473862 5210 473918
rect 5278 473862 5334 473918
rect 5402 473862 5458 473918
rect 5526 473862 5582 473918
rect 5154 473738 5210 473794
rect 5278 473738 5334 473794
rect 5402 473738 5458 473794
rect 5526 473738 5582 473794
rect 5154 473614 5210 473670
rect 5278 473614 5334 473670
rect 5402 473614 5458 473670
rect 5526 473614 5582 473670
rect 5154 473490 5210 473546
rect 5278 473490 5334 473546
rect 5402 473490 5458 473546
rect 5526 473490 5582 473546
rect 5154 455862 5210 455918
rect 5278 455862 5334 455918
rect 5402 455862 5458 455918
rect 5526 455862 5582 455918
rect 5154 455738 5210 455794
rect 5278 455738 5334 455794
rect 5402 455738 5458 455794
rect 5526 455738 5582 455794
rect 5154 455614 5210 455670
rect 5278 455614 5334 455670
rect 5402 455614 5458 455670
rect 5526 455614 5582 455670
rect 5154 455490 5210 455546
rect 5278 455490 5334 455546
rect 5402 455490 5458 455546
rect 5526 455490 5582 455546
rect 5154 437862 5210 437918
rect 5278 437862 5334 437918
rect 5402 437862 5458 437918
rect 5526 437862 5582 437918
rect 5154 437738 5210 437794
rect 5278 437738 5334 437794
rect 5402 437738 5458 437794
rect 5526 437738 5582 437794
rect 5154 437614 5210 437670
rect 5278 437614 5334 437670
rect 5402 437614 5458 437670
rect 5526 437614 5582 437670
rect 5154 437490 5210 437546
rect 5278 437490 5334 437546
rect 5402 437490 5458 437546
rect 5526 437490 5582 437546
rect 5154 419862 5210 419918
rect 5278 419862 5334 419918
rect 5402 419862 5458 419918
rect 5526 419862 5582 419918
rect 5154 419738 5210 419794
rect 5278 419738 5334 419794
rect 5402 419738 5458 419794
rect 5526 419738 5582 419794
rect 5154 419614 5210 419670
rect 5278 419614 5334 419670
rect 5402 419614 5458 419670
rect 5526 419614 5582 419670
rect 5154 419490 5210 419546
rect 5278 419490 5334 419546
rect 5402 419490 5458 419546
rect 5526 419490 5582 419546
rect 5154 401862 5210 401918
rect 5278 401862 5334 401918
rect 5402 401862 5458 401918
rect 5526 401862 5582 401918
rect 5154 401738 5210 401794
rect 5278 401738 5334 401794
rect 5402 401738 5458 401794
rect 5526 401738 5582 401794
rect 5154 401614 5210 401670
rect 5278 401614 5334 401670
rect 5402 401614 5458 401670
rect 5526 401614 5582 401670
rect 5154 401490 5210 401546
rect 5278 401490 5334 401546
rect 5402 401490 5458 401546
rect 5526 401490 5582 401546
rect 5154 383862 5210 383918
rect 5278 383862 5334 383918
rect 5402 383862 5458 383918
rect 5526 383862 5582 383918
rect 5154 383738 5210 383794
rect 5278 383738 5334 383794
rect 5402 383738 5458 383794
rect 5526 383738 5582 383794
rect 5154 383614 5210 383670
rect 5278 383614 5334 383670
rect 5402 383614 5458 383670
rect 5526 383614 5582 383670
rect 5154 383490 5210 383546
rect 5278 383490 5334 383546
rect 5402 383490 5458 383546
rect 5526 383490 5582 383546
rect 5154 365862 5210 365918
rect 5278 365862 5334 365918
rect 5402 365862 5458 365918
rect 5526 365862 5582 365918
rect 5154 365738 5210 365794
rect 5278 365738 5334 365794
rect 5402 365738 5458 365794
rect 5526 365738 5582 365794
rect 5154 365614 5210 365670
rect 5278 365614 5334 365670
rect 5402 365614 5458 365670
rect 5526 365614 5582 365670
rect 5154 365490 5210 365546
rect 5278 365490 5334 365546
rect 5402 365490 5458 365546
rect 5526 365490 5582 365546
rect 5154 347862 5210 347918
rect 5278 347862 5334 347918
rect 5402 347862 5458 347918
rect 5526 347862 5582 347918
rect 5154 347738 5210 347794
rect 5278 347738 5334 347794
rect 5402 347738 5458 347794
rect 5526 347738 5582 347794
rect 5154 347614 5210 347670
rect 5278 347614 5334 347670
rect 5402 347614 5458 347670
rect 5526 347614 5582 347670
rect 5154 347490 5210 347546
rect 5278 347490 5334 347546
rect 5402 347490 5458 347546
rect 5526 347490 5582 347546
rect 5154 329862 5210 329918
rect 5278 329862 5334 329918
rect 5402 329862 5458 329918
rect 5526 329862 5582 329918
rect 5154 329738 5210 329794
rect 5278 329738 5334 329794
rect 5402 329738 5458 329794
rect 5526 329738 5582 329794
rect 5154 329614 5210 329670
rect 5278 329614 5334 329670
rect 5402 329614 5458 329670
rect 5526 329614 5582 329670
rect 5154 329490 5210 329546
rect 5278 329490 5334 329546
rect 5402 329490 5458 329546
rect 5526 329490 5582 329546
rect 5154 311862 5210 311918
rect 5278 311862 5334 311918
rect 5402 311862 5458 311918
rect 5526 311862 5582 311918
rect 5154 311738 5210 311794
rect 5278 311738 5334 311794
rect 5402 311738 5458 311794
rect 5526 311738 5582 311794
rect 5154 311614 5210 311670
rect 5278 311614 5334 311670
rect 5402 311614 5458 311670
rect 5526 311614 5582 311670
rect 5154 311490 5210 311546
rect 5278 311490 5334 311546
rect 5402 311490 5458 311546
rect 5526 311490 5582 311546
rect 5154 293862 5210 293918
rect 5278 293862 5334 293918
rect 5402 293862 5458 293918
rect 5526 293862 5582 293918
rect 5154 293738 5210 293794
rect 5278 293738 5334 293794
rect 5402 293738 5458 293794
rect 5526 293738 5582 293794
rect 5154 293614 5210 293670
rect 5278 293614 5334 293670
rect 5402 293614 5458 293670
rect 5526 293614 5582 293670
rect 5154 293490 5210 293546
rect 5278 293490 5334 293546
rect 5402 293490 5458 293546
rect 5526 293490 5582 293546
rect 5154 275862 5210 275918
rect 5278 275862 5334 275918
rect 5402 275862 5458 275918
rect 5526 275862 5582 275918
rect 5154 275738 5210 275794
rect 5278 275738 5334 275794
rect 5402 275738 5458 275794
rect 5526 275738 5582 275794
rect 5154 275614 5210 275670
rect 5278 275614 5334 275670
rect 5402 275614 5458 275670
rect 5526 275614 5582 275670
rect 5154 275490 5210 275546
rect 5278 275490 5334 275546
rect 5402 275490 5458 275546
rect 5526 275490 5582 275546
rect 5154 257862 5210 257918
rect 5278 257862 5334 257918
rect 5402 257862 5458 257918
rect 5526 257862 5582 257918
rect 5154 257738 5210 257794
rect 5278 257738 5334 257794
rect 5402 257738 5458 257794
rect 5526 257738 5582 257794
rect 5154 257614 5210 257670
rect 5278 257614 5334 257670
rect 5402 257614 5458 257670
rect 5526 257614 5582 257670
rect 5154 257490 5210 257546
rect 5278 257490 5334 257546
rect 5402 257490 5458 257546
rect 5526 257490 5582 257546
rect 5154 239862 5210 239918
rect 5278 239862 5334 239918
rect 5402 239862 5458 239918
rect 5526 239862 5582 239918
rect 5154 239738 5210 239794
rect 5278 239738 5334 239794
rect 5402 239738 5458 239794
rect 5526 239738 5582 239794
rect 5154 239614 5210 239670
rect 5278 239614 5334 239670
rect 5402 239614 5458 239670
rect 5526 239614 5582 239670
rect 5154 239490 5210 239546
rect 5278 239490 5334 239546
rect 5402 239490 5458 239546
rect 5526 239490 5582 239546
rect 5154 221862 5210 221918
rect 5278 221862 5334 221918
rect 5402 221862 5458 221918
rect 5526 221862 5582 221918
rect 5154 221738 5210 221794
rect 5278 221738 5334 221794
rect 5402 221738 5458 221794
rect 5526 221738 5582 221794
rect 5154 221614 5210 221670
rect 5278 221614 5334 221670
rect 5402 221614 5458 221670
rect 5526 221614 5582 221670
rect 5154 221490 5210 221546
rect 5278 221490 5334 221546
rect 5402 221490 5458 221546
rect 5526 221490 5582 221546
rect 5154 203862 5210 203918
rect 5278 203862 5334 203918
rect 5402 203862 5458 203918
rect 5526 203862 5582 203918
rect 5154 203738 5210 203794
rect 5278 203738 5334 203794
rect 5402 203738 5458 203794
rect 5526 203738 5582 203794
rect 5154 203614 5210 203670
rect 5278 203614 5334 203670
rect 5402 203614 5458 203670
rect 5526 203614 5582 203670
rect 5154 203490 5210 203546
rect 5278 203490 5334 203546
rect 5402 203490 5458 203546
rect 5526 203490 5582 203546
rect 5154 185862 5210 185918
rect 5278 185862 5334 185918
rect 5402 185862 5458 185918
rect 5526 185862 5582 185918
rect 5154 185738 5210 185794
rect 5278 185738 5334 185794
rect 5402 185738 5458 185794
rect 5526 185738 5582 185794
rect 5154 185614 5210 185670
rect 5278 185614 5334 185670
rect 5402 185614 5458 185670
rect 5526 185614 5582 185670
rect 5154 185490 5210 185546
rect 5278 185490 5334 185546
rect 5402 185490 5458 185546
rect 5526 185490 5582 185546
rect 5154 167862 5210 167918
rect 5278 167862 5334 167918
rect 5402 167862 5458 167918
rect 5526 167862 5582 167918
rect 5154 167738 5210 167794
rect 5278 167738 5334 167794
rect 5402 167738 5458 167794
rect 5526 167738 5582 167794
rect 5154 167614 5210 167670
rect 5278 167614 5334 167670
rect 5402 167614 5458 167670
rect 5526 167614 5582 167670
rect 5154 167490 5210 167546
rect 5278 167490 5334 167546
rect 5402 167490 5458 167546
rect 5526 167490 5582 167546
rect 5154 149862 5210 149918
rect 5278 149862 5334 149918
rect 5402 149862 5458 149918
rect 5526 149862 5582 149918
rect 5154 149738 5210 149794
rect 5278 149738 5334 149794
rect 5402 149738 5458 149794
rect 5526 149738 5582 149794
rect 5154 149614 5210 149670
rect 5278 149614 5334 149670
rect 5402 149614 5458 149670
rect 5526 149614 5582 149670
rect 5154 149490 5210 149546
rect 5278 149490 5334 149546
rect 5402 149490 5458 149546
rect 5526 149490 5582 149546
rect 5154 131862 5210 131918
rect 5278 131862 5334 131918
rect 5402 131862 5458 131918
rect 5526 131862 5582 131918
rect 5154 131738 5210 131794
rect 5278 131738 5334 131794
rect 5402 131738 5458 131794
rect 5526 131738 5582 131794
rect 5154 131614 5210 131670
rect 5278 131614 5334 131670
rect 5402 131614 5458 131670
rect 5526 131614 5582 131670
rect 5154 131490 5210 131546
rect 5278 131490 5334 131546
rect 5402 131490 5458 131546
rect 5526 131490 5582 131546
rect 5154 113862 5210 113918
rect 5278 113862 5334 113918
rect 5402 113862 5458 113918
rect 5526 113862 5582 113918
rect 5154 113738 5210 113794
rect 5278 113738 5334 113794
rect 5402 113738 5458 113794
rect 5526 113738 5582 113794
rect 5154 113614 5210 113670
rect 5278 113614 5334 113670
rect 5402 113614 5458 113670
rect 5526 113614 5582 113670
rect 5154 113490 5210 113546
rect 5278 113490 5334 113546
rect 5402 113490 5458 113546
rect 5526 113490 5582 113546
rect 5154 95862 5210 95918
rect 5278 95862 5334 95918
rect 5402 95862 5458 95918
rect 5526 95862 5582 95918
rect 5154 95738 5210 95794
rect 5278 95738 5334 95794
rect 5402 95738 5458 95794
rect 5526 95738 5582 95794
rect 5154 95614 5210 95670
rect 5278 95614 5334 95670
rect 5402 95614 5458 95670
rect 5526 95614 5582 95670
rect 5154 95490 5210 95546
rect 5278 95490 5334 95546
rect 5402 95490 5458 95546
rect 5526 95490 5582 95546
rect 5154 77862 5210 77918
rect 5278 77862 5334 77918
rect 5402 77862 5458 77918
rect 5526 77862 5582 77918
rect 5154 77738 5210 77794
rect 5278 77738 5334 77794
rect 5402 77738 5458 77794
rect 5526 77738 5582 77794
rect 5154 77614 5210 77670
rect 5278 77614 5334 77670
rect 5402 77614 5458 77670
rect 5526 77614 5582 77670
rect 5154 77490 5210 77546
rect 5278 77490 5334 77546
rect 5402 77490 5458 77546
rect 5526 77490 5582 77546
rect 5154 59862 5210 59918
rect 5278 59862 5334 59918
rect 5402 59862 5458 59918
rect 5526 59862 5582 59918
rect 5154 59738 5210 59794
rect 5278 59738 5334 59794
rect 5402 59738 5458 59794
rect 5526 59738 5582 59794
rect 5154 59614 5210 59670
rect 5278 59614 5334 59670
rect 5402 59614 5458 59670
rect 5526 59614 5582 59670
rect 5154 59490 5210 59546
rect 5278 59490 5334 59546
rect 5402 59490 5458 59546
rect 5526 59490 5582 59546
rect 5154 41862 5210 41918
rect 5278 41862 5334 41918
rect 5402 41862 5458 41918
rect 5526 41862 5582 41918
rect 5154 41738 5210 41794
rect 5278 41738 5334 41794
rect 5402 41738 5458 41794
rect 5526 41738 5582 41794
rect 5154 41614 5210 41670
rect 5278 41614 5334 41670
rect 5402 41614 5458 41670
rect 5526 41614 5582 41670
rect 5154 41490 5210 41546
rect 5278 41490 5334 41546
rect 5402 41490 5458 41546
rect 5526 41490 5582 41546
rect 5154 23862 5210 23918
rect 5278 23862 5334 23918
rect 5402 23862 5458 23918
rect 5526 23862 5582 23918
rect 5154 23738 5210 23794
rect 5278 23738 5334 23794
rect 5402 23738 5458 23794
rect 5526 23738 5582 23794
rect 5154 23614 5210 23670
rect 5278 23614 5334 23670
rect 5402 23614 5458 23670
rect 5526 23614 5582 23670
rect 5154 23490 5210 23546
rect 5278 23490 5334 23546
rect 5402 23490 5458 23546
rect 5526 23490 5582 23546
rect 5154 5862 5210 5918
rect 5278 5862 5334 5918
rect 5402 5862 5458 5918
rect 5526 5862 5582 5918
rect 5154 5738 5210 5794
rect 5278 5738 5334 5794
rect 5402 5738 5458 5794
rect 5526 5738 5582 5794
rect 5154 5614 5210 5670
rect 5278 5614 5334 5670
rect 5402 5614 5458 5670
rect 5526 5614 5582 5670
rect 5154 5490 5210 5546
rect 5278 5490 5334 5546
rect 5402 5490 5458 5546
rect 5526 5490 5582 5546
rect 598512 581862 598568 581918
rect 598636 581862 598692 581918
rect 598760 581862 598816 581918
rect 598884 581862 598940 581918
rect 598512 581738 598568 581794
rect 598636 581738 598692 581794
rect 598760 581738 598816 581794
rect 598884 581738 598940 581794
rect 598512 581614 598568 581670
rect 598636 581614 598692 581670
rect 598760 581614 598816 581670
rect 598884 581614 598940 581670
rect 598512 581490 598568 581546
rect 598636 581490 598692 581546
rect 598760 581490 598816 581546
rect 598884 581490 598940 581546
rect 598512 563862 598568 563918
rect 598636 563862 598692 563918
rect 598760 563862 598816 563918
rect 598884 563862 598940 563918
rect 598512 563738 598568 563794
rect 598636 563738 598692 563794
rect 598760 563738 598816 563794
rect 598884 563738 598940 563794
rect 598512 563614 598568 563670
rect 598636 563614 598692 563670
rect 598760 563614 598816 563670
rect 598884 563614 598940 563670
rect 598512 563490 598568 563546
rect 598636 563490 598692 563546
rect 598760 563490 598816 563546
rect 598884 563490 598940 563546
rect 598512 545862 598568 545918
rect 598636 545862 598692 545918
rect 598760 545862 598816 545918
rect 598884 545862 598940 545918
rect 598512 545738 598568 545794
rect 598636 545738 598692 545794
rect 598760 545738 598816 545794
rect 598884 545738 598940 545794
rect 598512 545614 598568 545670
rect 598636 545614 598692 545670
rect 598760 545614 598816 545670
rect 598884 545614 598940 545670
rect 598512 545490 598568 545546
rect 598636 545490 598692 545546
rect 598760 545490 598816 545546
rect 598884 545490 598940 545546
rect 598512 527862 598568 527918
rect 598636 527862 598692 527918
rect 598760 527862 598816 527918
rect 598884 527862 598940 527918
rect 598512 527738 598568 527794
rect 598636 527738 598692 527794
rect 598760 527738 598816 527794
rect 598884 527738 598940 527794
rect 598512 527614 598568 527670
rect 598636 527614 598692 527670
rect 598760 527614 598816 527670
rect 598884 527614 598940 527670
rect 598512 527490 598568 527546
rect 598636 527490 598692 527546
rect 598760 527490 598816 527546
rect 598884 527490 598940 527546
rect 598512 509862 598568 509918
rect 598636 509862 598692 509918
rect 598760 509862 598816 509918
rect 598884 509862 598940 509918
rect 598512 509738 598568 509794
rect 598636 509738 598692 509794
rect 598760 509738 598816 509794
rect 598884 509738 598940 509794
rect 598512 509614 598568 509670
rect 598636 509614 598692 509670
rect 598760 509614 598816 509670
rect 598884 509614 598940 509670
rect 598512 509490 598568 509546
rect 598636 509490 598692 509546
rect 598760 509490 598816 509546
rect 598884 509490 598940 509546
rect 598512 491862 598568 491918
rect 598636 491862 598692 491918
rect 598760 491862 598816 491918
rect 598884 491862 598940 491918
rect 598512 491738 598568 491794
rect 598636 491738 598692 491794
rect 598760 491738 598816 491794
rect 598884 491738 598940 491794
rect 598512 491614 598568 491670
rect 598636 491614 598692 491670
rect 598760 491614 598816 491670
rect 598884 491614 598940 491670
rect 598512 491490 598568 491546
rect 598636 491490 598692 491546
rect 598760 491490 598816 491546
rect 598884 491490 598940 491546
rect 598512 473862 598568 473918
rect 598636 473862 598692 473918
rect 598760 473862 598816 473918
rect 598884 473862 598940 473918
rect 598512 473738 598568 473794
rect 598636 473738 598692 473794
rect 598760 473738 598816 473794
rect 598884 473738 598940 473794
rect 598512 473614 598568 473670
rect 598636 473614 598692 473670
rect 598760 473614 598816 473670
rect 598884 473614 598940 473670
rect 598512 473490 598568 473546
rect 598636 473490 598692 473546
rect 598760 473490 598816 473546
rect 598884 473490 598940 473546
rect 598512 455862 598568 455918
rect 598636 455862 598692 455918
rect 598760 455862 598816 455918
rect 598884 455862 598940 455918
rect 598512 455738 598568 455794
rect 598636 455738 598692 455794
rect 598760 455738 598816 455794
rect 598884 455738 598940 455794
rect 598512 455614 598568 455670
rect 598636 455614 598692 455670
rect 598760 455614 598816 455670
rect 598884 455614 598940 455670
rect 598512 455490 598568 455546
rect 598636 455490 598692 455546
rect 598760 455490 598816 455546
rect 598884 455490 598940 455546
rect 598512 437862 598568 437918
rect 598636 437862 598692 437918
rect 598760 437862 598816 437918
rect 598884 437862 598940 437918
rect 598512 437738 598568 437794
rect 598636 437738 598692 437794
rect 598760 437738 598816 437794
rect 598884 437738 598940 437794
rect 598512 437614 598568 437670
rect 598636 437614 598692 437670
rect 598760 437614 598816 437670
rect 598884 437614 598940 437670
rect 598512 437490 598568 437546
rect 598636 437490 598692 437546
rect 598760 437490 598816 437546
rect 598884 437490 598940 437546
rect 598512 419862 598568 419918
rect 598636 419862 598692 419918
rect 598760 419862 598816 419918
rect 598884 419862 598940 419918
rect 598512 419738 598568 419794
rect 598636 419738 598692 419794
rect 598760 419738 598816 419794
rect 598884 419738 598940 419794
rect 598512 419614 598568 419670
rect 598636 419614 598692 419670
rect 598760 419614 598816 419670
rect 598884 419614 598940 419670
rect 598512 419490 598568 419546
rect 598636 419490 598692 419546
rect 598760 419490 598816 419546
rect 598884 419490 598940 419546
rect 598512 401862 598568 401918
rect 598636 401862 598692 401918
rect 598760 401862 598816 401918
rect 598884 401862 598940 401918
rect 598512 401738 598568 401794
rect 598636 401738 598692 401794
rect 598760 401738 598816 401794
rect 598884 401738 598940 401794
rect 598512 401614 598568 401670
rect 598636 401614 598692 401670
rect 598760 401614 598816 401670
rect 598884 401614 598940 401670
rect 598512 401490 598568 401546
rect 598636 401490 598692 401546
rect 598760 401490 598816 401546
rect 598884 401490 598940 401546
rect 598512 383862 598568 383918
rect 598636 383862 598692 383918
rect 598760 383862 598816 383918
rect 598884 383862 598940 383918
rect 598512 383738 598568 383794
rect 598636 383738 598692 383794
rect 598760 383738 598816 383794
rect 598884 383738 598940 383794
rect 598512 383614 598568 383670
rect 598636 383614 598692 383670
rect 598760 383614 598816 383670
rect 598884 383614 598940 383670
rect 598512 383490 598568 383546
rect 598636 383490 598692 383546
rect 598760 383490 598816 383546
rect 598884 383490 598940 383546
rect 598512 365862 598568 365918
rect 598636 365862 598692 365918
rect 598760 365862 598816 365918
rect 598884 365862 598940 365918
rect 598512 365738 598568 365794
rect 598636 365738 598692 365794
rect 598760 365738 598816 365794
rect 598884 365738 598940 365794
rect 598512 365614 598568 365670
rect 598636 365614 598692 365670
rect 598760 365614 598816 365670
rect 598884 365614 598940 365670
rect 598512 365490 598568 365546
rect 598636 365490 598692 365546
rect 598760 365490 598816 365546
rect 598884 365490 598940 365546
rect 598512 347862 598568 347918
rect 598636 347862 598692 347918
rect 598760 347862 598816 347918
rect 598884 347862 598940 347918
rect 598512 347738 598568 347794
rect 598636 347738 598692 347794
rect 598760 347738 598816 347794
rect 598884 347738 598940 347794
rect 598512 347614 598568 347670
rect 598636 347614 598692 347670
rect 598760 347614 598816 347670
rect 598884 347614 598940 347670
rect 598512 347490 598568 347546
rect 598636 347490 598692 347546
rect 598760 347490 598816 347546
rect 598884 347490 598940 347546
rect 598512 329862 598568 329918
rect 598636 329862 598692 329918
rect 598760 329862 598816 329918
rect 598884 329862 598940 329918
rect 598512 329738 598568 329794
rect 598636 329738 598692 329794
rect 598760 329738 598816 329794
rect 598884 329738 598940 329794
rect 598512 329614 598568 329670
rect 598636 329614 598692 329670
rect 598760 329614 598816 329670
rect 598884 329614 598940 329670
rect 598512 329490 598568 329546
rect 598636 329490 598692 329546
rect 598760 329490 598816 329546
rect 598884 329490 598940 329546
rect 598512 311862 598568 311918
rect 598636 311862 598692 311918
rect 598760 311862 598816 311918
rect 598884 311862 598940 311918
rect 598512 311738 598568 311794
rect 598636 311738 598692 311794
rect 598760 311738 598816 311794
rect 598884 311738 598940 311794
rect 598512 311614 598568 311670
rect 598636 311614 598692 311670
rect 598760 311614 598816 311670
rect 598884 311614 598940 311670
rect 598512 311490 598568 311546
rect 598636 311490 598692 311546
rect 598760 311490 598816 311546
rect 598884 311490 598940 311546
rect 598512 293862 598568 293918
rect 598636 293862 598692 293918
rect 598760 293862 598816 293918
rect 598884 293862 598940 293918
rect 598512 293738 598568 293794
rect 598636 293738 598692 293794
rect 598760 293738 598816 293794
rect 598884 293738 598940 293794
rect 598512 293614 598568 293670
rect 598636 293614 598692 293670
rect 598760 293614 598816 293670
rect 598884 293614 598940 293670
rect 598512 293490 598568 293546
rect 598636 293490 598692 293546
rect 598760 293490 598816 293546
rect 598884 293490 598940 293546
rect 598512 275862 598568 275918
rect 598636 275862 598692 275918
rect 598760 275862 598816 275918
rect 598884 275862 598940 275918
rect 598512 275738 598568 275794
rect 598636 275738 598692 275794
rect 598760 275738 598816 275794
rect 598884 275738 598940 275794
rect 598512 275614 598568 275670
rect 598636 275614 598692 275670
rect 598760 275614 598816 275670
rect 598884 275614 598940 275670
rect 598512 275490 598568 275546
rect 598636 275490 598692 275546
rect 598760 275490 598816 275546
rect 598884 275490 598940 275546
rect 598512 257862 598568 257918
rect 598636 257862 598692 257918
rect 598760 257862 598816 257918
rect 598884 257862 598940 257918
rect 598512 257738 598568 257794
rect 598636 257738 598692 257794
rect 598760 257738 598816 257794
rect 598884 257738 598940 257794
rect 598512 257614 598568 257670
rect 598636 257614 598692 257670
rect 598760 257614 598816 257670
rect 598884 257614 598940 257670
rect 598512 257490 598568 257546
rect 598636 257490 598692 257546
rect 598760 257490 598816 257546
rect 598884 257490 598940 257546
rect 598512 239862 598568 239918
rect 598636 239862 598692 239918
rect 598760 239862 598816 239918
rect 598884 239862 598940 239918
rect 598512 239738 598568 239794
rect 598636 239738 598692 239794
rect 598760 239738 598816 239794
rect 598884 239738 598940 239794
rect 598512 239614 598568 239670
rect 598636 239614 598692 239670
rect 598760 239614 598816 239670
rect 598884 239614 598940 239670
rect 598512 239490 598568 239546
rect 598636 239490 598692 239546
rect 598760 239490 598816 239546
rect 598884 239490 598940 239546
rect 598512 221862 598568 221918
rect 598636 221862 598692 221918
rect 598760 221862 598816 221918
rect 598884 221862 598940 221918
rect 598512 221738 598568 221794
rect 598636 221738 598692 221794
rect 598760 221738 598816 221794
rect 598884 221738 598940 221794
rect 598512 221614 598568 221670
rect 598636 221614 598692 221670
rect 598760 221614 598816 221670
rect 598884 221614 598940 221670
rect 598512 221490 598568 221546
rect 598636 221490 598692 221546
rect 598760 221490 598816 221546
rect 598884 221490 598940 221546
rect 598512 203862 598568 203918
rect 598636 203862 598692 203918
rect 598760 203862 598816 203918
rect 598884 203862 598940 203918
rect 598512 203738 598568 203794
rect 598636 203738 598692 203794
rect 598760 203738 598816 203794
rect 598884 203738 598940 203794
rect 598512 203614 598568 203670
rect 598636 203614 598692 203670
rect 598760 203614 598816 203670
rect 598884 203614 598940 203670
rect 598512 203490 598568 203546
rect 598636 203490 598692 203546
rect 598760 203490 598816 203546
rect 598884 203490 598940 203546
rect 598512 185862 598568 185918
rect 598636 185862 598692 185918
rect 598760 185862 598816 185918
rect 598884 185862 598940 185918
rect 598512 185738 598568 185794
rect 598636 185738 598692 185794
rect 598760 185738 598816 185794
rect 598884 185738 598940 185794
rect 598512 185614 598568 185670
rect 598636 185614 598692 185670
rect 598760 185614 598816 185670
rect 598884 185614 598940 185670
rect 598512 185490 598568 185546
rect 598636 185490 598692 185546
rect 598760 185490 598816 185546
rect 598884 185490 598940 185546
rect 598512 167862 598568 167918
rect 598636 167862 598692 167918
rect 598760 167862 598816 167918
rect 598884 167862 598940 167918
rect 598512 167738 598568 167794
rect 598636 167738 598692 167794
rect 598760 167738 598816 167794
rect 598884 167738 598940 167794
rect 598512 167614 598568 167670
rect 598636 167614 598692 167670
rect 598760 167614 598816 167670
rect 598884 167614 598940 167670
rect 598512 167490 598568 167546
rect 598636 167490 598692 167546
rect 598760 167490 598816 167546
rect 598884 167490 598940 167546
rect 598512 149862 598568 149918
rect 598636 149862 598692 149918
rect 598760 149862 598816 149918
rect 598884 149862 598940 149918
rect 598512 149738 598568 149794
rect 598636 149738 598692 149794
rect 598760 149738 598816 149794
rect 598884 149738 598940 149794
rect 598512 149614 598568 149670
rect 598636 149614 598692 149670
rect 598760 149614 598816 149670
rect 598884 149614 598940 149670
rect 598512 149490 598568 149546
rect 598636 149490 598692 149546
rect 598760 149490 598816 149546
rect 598884 149490 598940 149546
rect 598512 131862 598568 131918
rect 598636 131862 598692 131918
rect 598760 131862 598816 131918
rect 598884 131862 598940 131918
rect 598512 131738 598568 131794
rect 598636 131738 598692 131794
rect 598760 131738 598816 131794
rect 598884 131738 598940 131794
rect 598512 131614 598568 131670
rect 598636 131614 598692 131670
rect 598760 131614 598816 131670
rect 598884 131614 598940 131670
rect 598512 131490 598568 131546
rect 598636 131490 598692 131546
rect 598760 131490 598816 131546
rect 598884 131490 598940 131546
rect 598512 113862 598568 113918
rect 598636 113862 598692 113918
rect 598760 113862 598816 113918
rect 598884 113862 598940 113918
rect 598512 113738 598568 113794
rect 598636 113738 598692 113794
rect 598760 113738 598816 113794
rect 598884 113738 598940 113794
rect 598512 113614 598568 113670
rect 598636 113614 598692 113670
rect 598760 113614 598816 113670
rect 598884 113614 598940 113670
rect 598512 113490 598568 113546
rect 598636 113490 598692 113546
rect 598760 113490 598816 113546
rect 598884 113490 598940 113546
rect 598512 95862 598568 95918
rect 598636 95862 598692 95918
rect 598760 95862 598816 95918
rect 598884 95862 598940 95918
rect 598512 95738 598568 95794
rect 598636 95738 598692 95794
rect 598760 95738 598816 95794
rect 598884 95738 598940 95794
rect 598512 95614 598568 95670
rect 598636 95614 598692 95670
rect 598760 95614 598816 95670
rect 598884 95614 598940 95670
rect 598512 95490 598568 95546
rect 598636 95490 598692 95546
rect 598760 95490 598816 95546
rect 598884 95490 598940 95546
rect 598512 77862 598568 77918
rect 598636 77862 598692 77918
rect 598760 77862 598816 77918
rect 598884 77862 598940 77918
rect 598512 77738 598568 77794
rect 598636 77738 598692 77794
rect 598760 77738 598816 77794
rect 598884 77738 598940 77794
rect 598512 77614 598568 77670
rect 598636 77614 598692 77670
rect 598760 77614 598816 77670
rect 598884 77614 598940 77670
rect 598512 77490 598568 77546
rect 598636 77490 598692 77546
rect 598760 77490 598816 77546
rect 598884 77490 598940 77546
rect 598512 59862 598568 59918
rect 598636 59862 598692 59918
rect 598760 59862 598816 59918
rect 598884 59862 598940 59918
rect 598512 59738 598568 59794
rect 598636 59738 598692 59794
rect 598760 59738 598816 59794
rect 598884 59738 598940 59794
rect 598512 59614 598568 59670
rect 598636 59614 598692 59670
rect 598760 59614 598816 59670
rect 598884 59614 598940 59670
rect 598512 59490 598568 59546
rect 598636 59490 598692 59546
rect 598760 59490 598816 59546
rect 598884 59490 598940 59546
rect 598512 41862 598568 41918
rect 598636 41862 598692 41918
rect 598760 41862 598816 41918
rect 598884 41862 598940 41918
rect 598512 41738 598568 41794
rect 598636 41738 598692 41794
rect 598760 41738 598816 41794
rect 598884 41738 598940 41794
rect 598512 41614 598568 41670
rect 598636 41614 598692 41670
rect 598760 41614 598816 41670
rect 598884 41614 598940 41670
rect 598512 41490 598568 41546
rect 598636 41490 598692 41546
rect 598760 41490 598816 41546
rect 598884 41490 598940 41546
rect 598512 23862 598568 23918
rect 598636 23862 598692 23918
rect 598760 23862 598816 23918
rect 598884 23862 598940 23918
rect 598512 23738 598568 23794
rect 598636 23738 598692 23794
rect 598760 23738 598816 23794
rect 598884 23738 598940 23794
rect 598512 23614 598568 23670
rect 598636 23614 598692 23670
rect 598760 23614 598816 23670
rect 598884 23614 598940 23670
rect 598512 23490 598568 23546
rect 598636 23490 598692 23546
rect 598760 23490 598816 23546
rect 598884 23490 598940 23546
rect 598512 5862 598568 5918
rect 598636 5862 598692 5918
rect 598760 5862 598816 5918
rect 598884 5862 598940 5918
rect 598512 5738 598568 5794
rect 598636 5738 598692 5794
rect 598760 5738 598816 5794
rect 598884 5738 598940 5794
rect 598512 5614 598568 5670
rect 598636 5614 598692 5670
rect 598760 5614 598816 5670
rect 598884 5614 598940 5670
rect 598512 5490 598568 5546
rect 598636 5490 598692 5546
rect 598760 5490 598816 5546
rect 598884 5490 598940 5546
rect 5154 1752 5210 1808
rect 5278 1752 5334 1808
rect 5402 1752 5458 1808
rect 5526 1752 5582 1808
rect 5154 1628 5210 1684
rect 5278 1628 5334 1684
rect 5402 1628 5458 1684
rect 5526 1628 5582 1684
rect 5154 1504 5210 1560
rect 5278 1504 5334 1560
rect 5402 1504 5458 1560
rect 5526 1504 5582 1560
rect 5154 1380 5210 1436
rect 5278 1380 5334 1436
rect 5402 1380 5458 1436
rect 5526 1380 5582 1436
rect 84 792 140 848
rect 208 792 264 848
rect 332 792 388 848
rect 456 792 512 848
rect 84 668 140 724
rect 208 668 264 724
rect 332 668 388 724
rect 456 668 512 724
rect 84 544 140 600
rect 208 544 264 600
rect 332 544 388 600
rect 456 544 512 600
rect 84 420 140 476
rect 208 420 264 476
rect 332 420 388 476
rect 456 420 512 476
rect 8874 792 8930 848
rect 8998 792 9054 848
rect 9122 792 9178 848
rect 9246 792 9302 848
rect 8874 668 8930 724
rect 8998 668 9054 724
rect 9122 668 9178 724
rect 9246 668 9302 724
rect 8874 544 8930 600
rect 8998 544 9054 600
rect 9122 544 9178 600
rect 9246 544 9302 600
rect 8874 420 8930 476
rect 8998 420 9054 476
rect 9122 420 9178 476
rect 9246 420 9302 476
rect 23154 1752 23210 1808
rect 23278 1752 23334 1808
rect 23402 1752 23458 1808
rect 23526 1752 23582 1808
rect 23154 1628 23210 1684
rect 23278 1628 23334 1684
rect 23402 1628 23458 1684
rect 23526 1628 23582 1684
rect 23154 1504 23210 1560
rect 23278 1504 23334 1560
rect 23402 1504 23458 1560
rect 23526 1504 23582 1560
rect 23154 1380 23210 1436
rect 23278 1380 23334 1436
rect 23402 1380 23458 1436
rect 23526 1380 23582 1436
rect 26874 792 26930 848
rect 26998 792 27054 848
rect 27122 792 27178 848
rect 27246 792 27302 848
rect 26874 668 26930 724
rect 26998 668 27054 724
rect 27122 668 27178 724
rect 27246 668 27302 724
rect 26874 544 26930 600
rect 26998 544 27054 600
rect 27122 544 27178 600
rect 27246 544 27302 600
rect 26874 420 26930 476
rect 26998 420 27054 476
rect 27122 420 27178 476
rect 27246 420 27302 476
rect 41154 1752 41210 1808
rect 41278 1752 41334 1808
rect 41402 1752 41458 1808
rect 41526 1752 41582 1808
rect 41154 1628 41210 1684
rect 41278 1628 41334 1684
rect 41402 1628 41458 1684
rect 41526 1628 41582 1684
rect 41154 1504 41210 1560
rect 41278 1504 41334 1560
rect 41402 1504 41458 1560
rect 41526 1504 41582 1560
rect 41154 1380 41210 1436
rect 41278 1380 41334 1436
rect 41402 1380 41458 1436
rect 41526 1380 41582 1436
rect 44874 792 44930 848
rect 44998 792 45054 848
rect 45122 792 45178 848
rect 45246 792 45302 848
rect 44874 668 44930 724
rect 44998 668 45054 724
rect 45122 668 45178 724
rect 45246 668 45302 724
rect 44874 544 44930 600
rect 44998 544 45054 600
rect 45122 544 45178 600
rect 45246 544 45302 600
rect 44874 420 44930 476
rect 44998 420 45054 476
rect 45122 420 45178 476
rect 45246 420 45302 476
rect 59154 1752 59210 1808
rect 59278 1752 59334 1808
rect 59402 1752 59458 1808
rect 59526 1752 59582 1808
rect 59154 1628 59210 1684
rect 59278 1628 59334 1684
rect 59402 1628 59458 1684
rect 59526 1628 59582 1684
rect 59154 1504 59210 1560
rect 59278 1504 59334 1560
rect 59402 1504 59458 1560
rect 59526 1504 59582 1560
rect 59154 1380 59210 1436
rect 59278 1380 59334 1436
rect 59402 1380 59458 1436
rect 59526 1380 59582 1436
rect 62874 792 62930 848
rect 62998 792 63054 848
rect 63122 792 63178 848
rect 63246 792 63302 848
rect 62874 668 62930 724
rect 62998 668 63054 724
rect 63122 668 63178 724
rect 63246 668 63302 724
rect 62874 544 62930 600
rect 62998 544 63054 600
rect 63122 544 63178 600
rect 63246 544 63302 600
rect 62874 420 62930 476
rect 62998 420 63054 476
rect 63122 420 63178 476
rect 63246 420 63302 476
rect 77154 1752 77210 1808
rect 77278 1752 77334 1808
rect 77402 1752 77458 1808
rect 77526 1752 77582 1808
rect 77154 1628 77210 1684
rect 77278 1628 77334 1684
rect 77402 1628 77458 1684
rect 77526 1628 77582 1684
rect 77154 1504 77210 1560
rect 77278 1504 77334 1560
rect 77402 1504 77458 1560
rect 77526 1504 77582 1560
rect 77154 1380 77210 1436
rect 77278 1380 77334 1436
rect 77402 1380 77458 1436
rect 77526 1380 77582 1436
rect 80874 792 80930 848
rect 80998 792 81054 848
rect 81122 792 81178 848
rect 81246 792 81302 848
rect 80874 668 80930 724
rect 80998 668 81054 724
rect 81122 668 81178 724
rect 81246 668 81302 724
rect 80874 544 80930 600
rect 80998 544 81054 600
rect 81122 544 81178 600
rect 81246 544 81302 600
rect 80874 420 80930 476
rect 80998 420 81054 476
rect 81122 420 81178 476
rect 81246 420 81302 476
rect 95154 1752 95210 1808
rect 95278 1752 95334 1808
rect 95402 1752 95458 1808
rect 95526 1752 95582 1808
rect 95154 1628 95210 1684
rect 95278 1628 95334 1684
rect 95402 1628 95458 1684
rect 95526 1628 95582 1684
rect 95154 1504 95210 1560
rect 95278 1504 95334 1560
rect 95402 1504 95458 1560
rect 95526 1504 95582 1560
rect 95154 1380 95210 1436
rect 95278 1380 95334 1436
rect 95402 1380 95458 1436
rect 95526 1380 95582 1436
rect 98874 792 98930 848
rect 98998 792 99054 848
rect 99122 792 99178 848
rect 99246 792 99302 848
rect 98874 668 98930 724
rect 98998 668 99054 724
rect 99122 668 99178 724
rect 99246 668 99302 724
rect 98874 544 98930 600
rect 98998 544 99054 600
rect 99122 544 99178 600
rect 99246 544 99302 600
rect 98874 420 98930 476
rect 98998 420 99054 476
rect 99122 420 99178 476
rect 99246 420 99302 476
rect 113154 1752 113210 1808
rect 113278 1752 113334 1808
rect 113402 1752 113458 1808
rect 113526 1752 113582 1808
rect 113154 1628 113210 1684
rect 113278 1628 113334 1684
rect 113402 1628 113458 1684
rect 113526 1628 113582 1684
rect 113154 1504 113210 1560
rect 113278 1504 113334 1560
rect 113402 1504 113458 1560
rect 113526 1504 113582 1560
rect 113154 1380 113210 1436
rect 113278 1380 113334 1436
rect 113402 1380 113458 1436
rect 113526 1380 113582 1436
rect 116874 792 116930 848
rect 116998 792 117054 848
rect 117122 792 117178 848
rect 117246 792 117302 848
rect 116874 668 116930 724
rect 116998 668 117054 724
rect 117122 668 117178 724
rect 117246 668 117302 724
rect 116874 544 116930 600
rect 116998 544 117054 600
rect 117122 544 117178 600
rect 117246 544 117302 600
rect 116874 420 116930 476
rect 116998 420 117054 476
rect 117122 420 117178 476
rect 117246 420 117302 476
rect 131154 1752 131210 1808
rect 131278 1752 131334 1808
rect 131402 1752 131458 1808
rect 131526 1752 131582 1808
rect 131154 1628 131210 1684
rect 131278 1628 131334 1684
rect 131402 1628 131458 1684
rect 131526 1628 131582 1684
rect 131154 1504 131210 1560
rect 131278 1504 131334 1560
rect 131402 1504 131458 1560
rect 131526 1504 131582 1560
rect 131154 1380 131210 1436
rect 131278 1380 131334 1436
rect 131402 1380 131458 1436
rect 131526 1380 131582 1436
rect 134874 792 134930 848
rect 134998 792 135054 848
rect 135122 792 135178 848
rect 135246 792 135302 848
rect 134874 668 134930 724
rect 134998 668 135054 724
rect 135122 668 135178 724
rect 135246 668 135302 724
rect 134874 544 134930 600
rect 134998 544 135054 600
rect 135122 544 135178 600
rect 135246 544 135302 600
rect 134874 420 134930 476
rect 134998 420 135054 476
rect 135122 420 135178 476
rect 135246 420 135302 476
rect 149154 1752 149210 1808
rect 149278 1752 149334 1808
rect 149402 1752 149458 1808
rect 149526 1752 149582 1808
rect 149154 1628 149210 1684
rect 149278 1628 149334 1684
rect 149402 1628 149458 1684
rect 149526 1628 149582 1684
rect 149154 1504 149210 1560
rect 149278 1504 149334 1560
rect 149402 1504 149458 1560
rect 149526 1504 149582 1560
rect 149154 1380 149210 1436
rect 149278 1380 149334 1436
rect 149402 1380 149458 1436
rect 149526 1380 149582 1436
rect 152874 792 152930 848
rect 152998 792 153054 848
rect 153122 792 153178 848
rect 153246 792 153302 848
rect 152874 668 152930 724
rect 152998 668 153054 724
rect 153122 668 153178 724
rect 153246 668 153302 724
rect 152874 544 152930 600
rect 152998 544 153054 600
rect 153122 544 153178 600
rect 153246 544 153302 600
rect 152874 420 152930 476
rect 152998 420 153054 476
rect 153122 420 153178 476
rect 153246 420 153302 476
rect 167154 1752 167210 1808
rect 167278 1752 167334 1808
rect 167402 1752 167458 1808
rect 167526 1752 167582 1808
rect 167154 1628 167210 1684
rect 167278 1628 167334 1684
rect 167402 1628 167458 1684
rect 167526 1628 167582 1684
rect 167154 1504 167210 1560
rect 167278 1504 167334 1560
rect 167402 1504 167458 1560
rect 167526 1504 167582 1560
rect 167154 1380 167210 1436
rect 167278 1380 167334 1436
rect 167402 1380 167458 1436
rect 167526 1380 167582 1436
rect 170874 792 170930 848
rect 170998 792 171054 848
rect 171122 792 171178 848
rect 171246 792 171302 848
rect 170874 668 170930 724
rect 170998 668 171054 724
rect 171122 668 171178 724
rect 171246 668 171302 724
rect 170874 544 170930 600
rect 170998 544 171054 600
rect 171122 544 171178 600
rect 171246 544 171302 600
rect 170874 420 170930 476
rect 170998 420 171054 476
rect 171122 420 171178 476
rect 171246 420 171302 476
rect 185154 1752 185210 1808
rect 185278 1752 185334 1808
rect 185402 1752 185458 1808
rect 185526 1752 185582 1808
rect 185154 1628 185210 1684
rect 185278 1628 185334 1684
rect 185402 1628 185458 1684
rect 185526 1628 185582 1684
rect 185154 1504 185210 1560
rect 185278 1504 185334 1560
rect 185402 1504 185458 1560
rect 185526 1504 185582 1560
rect 185154 1380 185210 1436
rect 185278 1380 185334 1436
rect 185402 1380 185458 1436
rect 185526 1380 185582 1436
rect 188874 792 188930 848
rect 188998 792 189054 848
rect 189122 792 189178 848
rect 189246 792 189302 848
rect 188874 668 188930 724
rect 188998 668 189054 724
rect 189122 668 189178 724
rect 189246 668 189302 724
rect 188874 544 188930 600
rect 188998 544 189054 600
rect 189122 544 189178 600
rect 189246 544 189302 600
rect 188874 420 188930 476
rect 188998 420 189054 476
rect 189122 420 189178 476
rect 189246 420 189302 476
rect 203154 1752 203210 1808
rect 203278 1752 203334 1808
rect 203402 1752 203458 1808
rect 203526 1752 203582 1808
rect 203154 1628 203210 1684
rect 203278 1628 203334 1684
rect 203402 1628 203458 1684
rect 203526 1628 203582 1684
rect 203154 1504 203210 1560
rect 203278 1504 203334 1560
rect 203402 1504 203458 1560
rect 203526 1504 203582 1560
rect 203154 1380 203210 1436
rect 203278 1380 203334 1436
rect 203402 1380 203458 1436
rect 203526 1380 203582 1436
rect 206874 792 206930 848
rect 206998 792 207054 848
rect 207122 792 207178 848
rect 207246 792 207302 848
rect 206874 668 206930 724
rect 206998 668 207054 724
rect 207122 668 207178 724
rect 207246 668 207302 724
rect 206874 544 206930 600
rect 206998 544 207054 600
rect 207122 544 207178 600
rect 207246 544 207302 600
rect 206874 420 206930 476
rect 206998 420 207054 476
rect 207122 420 207178 476
rect 207246 420 207302 476
rect 221154 1752 221210 1808
rect 221278 1752 221334 1808
rect 221402 1752 221458 1808
rect 221526 1752 221582 1808
rect 221154 1628 221210 1684
rect 221278 1628 221334 1684
rect 221402 1628 221458 1684
rect 221526 1628 221582 1684
rect 221154 1504 221210 1560
rect 221278 1504 221334 1560
rect 221402 1504 221458 1560
rect 221526 1504 221582 1560
rect 221154 1380 221210 1436
rect 221278 1380 221334 1436
rect 221402 1380 221458 1436
rect 221526 1380 221582 1436
rect 224874 792 224930 848
rect 224998 792 225054 848
rect 225122 792 225178 848
rect 225246 792 225302 848
rect 224874 668 224930 724
rect 224998 668 225054 724
rect 225122 668 225178 724
rect 225246 668 225302 724
rect 224874 544 224930 600
rect 224998 544 225054 600
rect 225122 544 225178 600
rect 225246 544 225302 600
rect 224874 420 224930 476
rect 224998 420 225054 476
rect 225122 420 225178 476
rect 225246 420 225302 476
rect 239154 1752 239210 1808
rect 239278 1752 239334 1808
rect 239402 1752 239458 1808
rect 239526 1752 239582 1808
rect 239154 1628 239210 1684
rect 239278 1628 239334 1684
rect 239402 1628 239458 1684
rect 239526 1628 239582 1684
rect 239154 1504 239210 1560
rect 239278 1504 239334 1560
rect 239402 1504 239458 1560
rect 239526 1504 239582 1560
rect 239154 1380 239210 1436
rect 239278 1380 239334 1436
rect 239402 1380 239458 1436
rect 239526 1380 239582 1436
rect 242874 792 242930 848
rect 242998 792 243054 848
rect 243122 792 243178 848
rect 243246 792 243302 848
rect 242874 668 242930 724
rect 242998 668 243054 724
rect 243122 668 243178 724
rect 243246 668 243302 724
rect 242874 544 242930 600
rect 242998 544 243054 600
rect 243122 544 243178 600
rect 243246 544 243302 600
rect 242874 420 242930 476
rect 242998 420 243054 476
rect 243122 420 243178 476
rect 243246 420 243302 476
rect 257154 1752 257210 1808
rect 257278 1752 257334 1808
rect 257402 1752 257458 1808
rect 257526 1752 257582 1808
rect 257154 1628 257210 1684
rect 257278 1628 257334 1684
rect 257402 1628 257458 1684
rect 257526 1628 257582 1684
rect 257154 1504 257210 1560
rect 257278 1504 257334 1560
rect 257402 1504 257458 1560
rect 257526 1504 257582 1560
rect 257154 1380 257210 1436
rect 257278 1380 257334 1436
rect 257402 1380 257458 1436
rect 257526 1380 257582 1436
rect 260874 792 260930 848
rect 260998 792 261054 848
rect 261122 792 261178 848
rect 261246 792 261302 848
rect 260874 668 260930 724
rect 260998 668 261054 724
rect 261122 668 261178 724
rect 261246 668 261302 724
rect 260874 544 260930 600
rect 260998 544 261054 600
rect 261122 544 261178 600
rect 261246 544 261302 600
rect 260874 420 260930 476
rect 260998 420 261054 476
rect 261122 420 261178 476
rect 261246 420 261302 476
rect 275154 1752 275210 1808
rect 275278 1752 275334 1808
rect 275402 1752 275458 1808
rect 275526 1752 275582 1808
rect 275154 1628 275210 1684
rect 275278 1628 275334 1684
rect 275402 1628 275458 1684
rect 275526 1628 275582 1684
rect 275154 1504 275210 1560
rect 275278 1504 275334 1560
rect 275402 1504 275458 1560
rect 275526 1504 275582 1560
rect 275154 1380 275210 1436
rect 275278 1380 275334 1436
rect 275402 1380 275458 1436
rect 275526 1380 275582 1436
rect 278874 792 278930 848
rect 278998 792 279054 848
rect 279122 792 279178 848
rect 279246 792 279302 848
rect 278874 668 278930 724
rect 278998 668 279054 724
rect 279122 668 279178 724
rect 279246 668 279302 724
rect 278874 544 278930 600
rect 278998 544 279054 600
rect 279122 544 279178 600
rect 279246 544 279302 600
rect 278874 420 278930 476
rect 278998 420 279054 476
rect 279122 420 279178 476
rect 279246 420 279302 476
rect 293154 1752 293210 1808
rect 293278 1752 293334 1808
rect 293402 1752 293458 1808
rect 293526 1752 293582 1808
rect 293154 1628 293210 1684
rect 293278 1628 293334 1684
rect 293402 1628 293458 1684
rect 293526 1628 293582 1684
rect 293154 1504 293210 1560
rect 293278 1504 293334 1560
rect 293402 1504 293458 1560
rect 293526 1504 293582 1560
rect 293154 1380 293210 1436
rect 293278 1380 293334 1436
rect 293402 1380 293458 1436
rect 293526 1380 293582 1436
rect 296874 792 296930 848
rect 296998 792 297054 848
rect 297122 792 297178 848
rect 297246 792 297302 848
rect 296874 668 296930 724
rect 296998 668 297054 724
rect 297122 668 297178 724
rect 297246 668 297302 724
rect 296874 544 296930 600
rect 296998 544 297054 600
rect 297122 544 297178 600
rect 297246 544 297302 600
rect 296874 420 296930 476
rect 296998 420 297054 476
rect 297122 420 297178 476
rect 297246 420 297302 476
rect 311154 1752 311210 1808
rect 311278 1752 311334 1808
rect 311402 1752 311458 1808
rect 311526 1752 311582 1808
rect 311154 1628 311210 1684
rect 311278 1628 311334 1684
rect 311402 1628 311458 1684
rect 311526 1628 311582 1684
rect 311154 1504 311210 1560
rect 311278 1504 311334 1560
rect 311402 1504 311458 1560
rect 311526 1504 311582 1560
rect 311154 1380 311210 1436
rect 311278 1380 311334 1436
rect 311402 1380 311458 1436
rect 311526 1380 311582 1436
rect 314874 792 314930 848
rect 314998 792 315054 848
rect 315122 792 315178 848
rect 315246 792 315302 848
rect 314874 668 314930 724
rect 314998 668 315054 724
rect 315122 668 315178 724
rect 315246 668 315302 724
rect 314874 544 314930 600
rect 314998 544 315054 600
rect 315122 544 315178 600
rect 315246 544 315302 600
rect 314874 420 314930 476
rect 314998 420 315054 476
rect 315122 420 315178 476
rect 315246 420 315302 476
rect 329154 1752 329210 1808
rect 329278 1752 329334 1808
rect 329402 1752 329458 1808
rect 329526 1752 329582 1808
rect 329154 1628 329210 1684
rect 329278 1628 329334 1684
rect 329402 1628 329458 1684
rect 329526 1628 329582 1684
rect 329154 1504 329210 1560
rect 329278 1504 329334 1560
rect 329402 1504 329458 1560
rect 329526 1504 329582 1560
rect 329154 1380 329210 1436
rect 329278 1380 329334 1436
rect 329402 1380 329458 1436
rect 329526 1380 329582 1436
rect 332874 792 332930 848
rect 332998 792 333054 848
rect 333122 792 333178 848
rect 333246 792 333302 848
rect 332874 668 332930 724
rect 332998 668 333054 724
rect 333122 668 333178 724
rect 333246 668 333302 724
rect 332874 544 332930 600
rect 332998 544 333054 600
rect 333122 544 333178 600
rect 333246 544 333302 600
rect 332874 420 332930 476
rect 332998 420 333054 476
rect 333122 420 333178 476
rect 333246 420 333302 476
rect 347154 1752 347210 1808
rect 347278 1752 347334 1808
rect 347402 1752 347458 1808
rect 347526 1752 347582 1808
rect 347154 1628 347210 1684
rect 347278 1628 347334 1684
rect 347402 1628 347458 1684
rect 347526 1628 347582 1684
rect 347154 1504 347210 1560
rect 347278 1504 347334 1560
rect 347402 1504 347458 1560
rect 347526 1504 347582 1560
rect 347154 1380 347210 1436
rect 347278 1380 347334 1436
rect 347402 1380 347458 1436
rect 347526 1380 347582 1436
rect 350874 792 350930 848
rect 350998 792 351054 848
rect 351122 792 351178 848
rect 351246 792 351302 848
rect 350874 668 350930 724
rect 350998 668 351054 724
rect 351122 668 351178 724
rect 351246 668 351302 724
rect 350874 544 350930 600
rect 350998 544 351054 600
rect 351122 544 351178 600
rect 351246 544 351302 600
rect 350874 420 350930 476
rect 350998 420 351054 476
rect 351122 420 351178 476
rect 351246 420 351302 476
rect 365154 1752 365210 1808
rect 365278 1752 365334 1808
rect 365402 1752 365458 1808
rect 365526 1752 365582 1808
rect 365154 1628 365210 1684
rect 365278 1628 365334 1684
rect 365402 1628 365458 1684
rect 365526 1628 365582 1684
rect 365154 1504 365210 1560
rect 365278 1504 365334 1560
rect 365402 1504 365458 1560
rect 365526 1504 365582 1560
rect 365154 1380 365210 1436
rect 365278 1380 365334 1436
rect 365402 1380 365458 1436
rect 365526 1380 365582 1436
rect 368874 792 368930 848
rect 368998 792 369054 848
rect 369122 792 369178 848
rect 369246 792 369302 848
rect 368874 668 368930 724
rect 368998 668 369054 724
rect 369122 668 369178 724
rect 369246 668 369302 724
rect 368874 544 368930 600
rect 368998 544 369054 600
rect 369122 544 369178 600
rect 369246 544 369302 600
rect 368874 420 368930 476
rect 368998 420 369054 476
rect 369122 420 369178 476
rect 369246 420 369302 476
rect 383154 1752 383210 1808
rect 383278 1752 383334 1808
rect 383402 1752 383458 1808
rect 383526 1752 383582 1808
rect 383154 1628 383210 1684
rect 383278 1628 383334 1684
rect 383402 1628 383458 1684
rect 383526 1628 383582 1684
rect 383154 1504 383210 1560
rect 383278 1504 383334 1560
rect 383402 1504 383458 1560
rect 383526 1504 383582 1560
rect 383154 1380 383210 1436
rect 383278 1380 383334 1436
rect 383402 1380 383458 1436
rect 383526 1380 383582 1436
rect 386874 792 386930 848
rect 386998 792 387054 848
rect 387122 792 387178 848
rect 387246 792 387302 848
rect 386874 668 386930 724
rect 386998 668 387054 724
rect 387122 668 387178 724
rect 387246 668 387302 724
rect 386874 544 386930 600
rect 386998 544 387054 600
rect 387122 544 387178 600
rect 387246 544 387302 600
rect 386874 420 386930 476
rect 386998 420 387054 476
rect 387122 420 387178 476
rect 387246 420 387302 476
rect 401154 1752 401210 1808
rect 401278 1752 401334 1808
rect 401402 1752 401458 1808
rect 401526 1752 401582 1808
rect 401154 1628 401210 1684
rect 401278 1628 401334 1684
rect 401402 1628 401458 1684
rect 401526 1628 401582 1684
rect 401154 1504 401210 1560
rect 401278 1504 401334 1560
rect 401402 1504 401458 1560
rect 401526 1504 401582 1560
rect 401154 1380 401210 1436
rect 401278 1380 401334 1436
rect 401402 1380 401458 1436
rect 401526 1380 401582 1436
rect 404874 792 404930 848
rect 404998 792 405054 848
rect 405122 792 405178 848
rect 405246 792 405302 848
rect 404874 668 404930 724
rect 404998 668 405054 724
rect 405122 668 405178 724
rect 405246 668 405302 724
rect 404874 544 404930 600
rect 404998 544 405054 600
rect 405122 544 405178 600
rect 405246 544 405302 600
rect 404874 420 404930 476
rect 404998 420 405054 476
rect 405122 420 405178 476
rect 405246 420 405302 476
rect 419154 1752 419210 1808
rect 419278 1752 419334 1808
rect 419402 1752 419458 1808
rect 419526 1752 419582 1808
rect 419154 1628 419210 1684
rect 419278 1628 419334 1684
rect 419402 1628 419458 1684
rect 419526 1628 419582 1684
rect 419154 1504 419210 1560
rect 419278 1504 419334 1560
rect 419402 1504 419458 1560
rect 419526 1504 419582 1560
rect 419154 1380 419210 1436
rect 419278 1380 419334 1436
rect 419402 1380 419458 1436
rect 419526 1380 419582 1436
rect 422874 792 422930 848
rect 422998 792 423054 848
rect 423122 792 423178 848
rect 423246 792 423302 848
rect 422874 668 422930 724
rect 422998 668 423054 724
rect 423122 668 423178 724
rect 423246 668 423302 724
rect 422874 544 422930 600
rect 422998 544 423054 600
rect 423122 544 423178 600
rect 423246 544 423302 600
rect 422874 420 422930 476
rect 422998 420 423054 476
rect 423122 420 423178 476
rect 423246 420 423302 476
rect 437154 1752 437210 1808
rect 437278 1752 437334 1808
rect 437402 1752 437458 1808
rect 437526 1752 437582 1808
rect 437154 1628 437210 1684
rect 437278 1628 437334 1684
rect 437402 1628 437458 1684
rect 437526 1628 437582 1684
rect 437154 1504 437210 1560
rect 437278 1504 437334 1560
rect 437402 1504 437458 1560
rect 437526 1504 437582 1560
rect 437154 1380 437210 1436
rect 437278 1380 437334 1436
rect 437402 1380 437458 1436
rect 437526 1380 437582 1436
rect 440874 792 440930 848
rect 440998 792 441054 848
rect 441122 792 441178 848
rect 441246 792 441302 848
rect 440874 668 440930 724
rect 440998 668 441054 724
rect 441122 668 441178 724
rect 441246 668 441302 724
rect 440874 544 440930 600
rect 440998 544 441054 600
rect 441122 544 441178 600
rect 441246 544 441302 600
rect 440874 420 440930 476
rect 440998 420 441054 476
rect 441122 420 441178 476
rect 441246 420 441302 476
rect 455154 1752 455210 1808
rect 455278 1752 455334 1808
rect 455402 1752 455458 1808
rect 455526 1752 455582 1808
rect 455154 1628 455210 1684
rect 455278 1628 455334 1684
rect 455402 1628 455458 1684
rect 455526 1628 455582 1684
rect 455154 1504 455210 1560
rect 455278 1504 455334 1560
rect 455402 1504 455458 1560
rect 455526 1504 455582 1560
rect 455154 1380 455210 1436
rect 455278 1380 455334 1436
rect 455402 1380 455458 1436
rect 455526 1380 455582 1436
rect 458874 792 458930 848
rect 458998 792 459054 848
rect 459122 792 459178 848
rect 459246 792 459302 848
rect 458874 668 458930 724
rect 458998 668 459054 724
rect 459122 668 459178 724
rect 459246 668 459302 724
rect 458874 544 458930 600
rect 458998 544 459054 600
rect 459122 544 459178 600
rect 459246 544 459302 600
rect 458874 420 458930 476
rect 458998 420 459054 476
rect 459122 420 459178 476
rect 459246 420 459302 476
rect 473154 1752 473210 1808
rect 473278 1752 473334 1808
rect 473402 1752 473458 1808
rect 473526 1752 473582 1808
rect 473154 1628 473210 1684
rect 473278 1628 473334 1684
rect 473402 1628 473458 1684
rect 473526 1628 473582 1684
rect 473154 1504 473210 1560
rect 473278 1504 473334 1560
rect 473402 1504 473458 1560
rect 473526 1504 473582 1560
rect 473154 1380 473210 1436
rect 473278 1380 473334 1436
rect 473402 1380 473458 1436
rect 473526 1380 473582 1436
rect 476874 792 476930 848
rect 476998 792 477054 848
rect 477122 792 477178 848
rect 477246 792 477302 848
rect 476874 668 476930 724
rect 476998 668 477054 724
rect 477122 668 477178 724
rect 477246 668 477302 724
rect 476874 544 476930 600
rect 476998 544 477054 600
rect 477122 544 477178 600
rect 477246 544 477302 600
rect 476874 420 476930 476
rect 476998 420 477054 476
rect 477122 420 477178 476
rect 477246 420 477302 476
rect 491154 1752 491210 1808
rect 491278 1752 491334 1808
rect 491402 1752 491458 1808
rect 491526 1752 491582 1808
rect 491154 1628 491210 1684
rect 491278 1628 491334 1684
rect 491402 1628 491458 1684
rect 491526 1628 491582 1684
rect 491154 1504 491210 1560
rect 491278 1504 491334 1560
rect 491402 1504 491458 1560
rect 491526 1504 491582 1560
rect 491154 1380 491210 1436
rect 491278 1380 491334 1436
rect 491402 1380 491458 1436
rect 491526 1380 491582 1436
rect 494874 792 494930 848
rect 494998 792 495054 848
rect 495122 792 495178 848
rect 495246 792 495302 848
rect 494874 668 494930 724
rect 494998 668 495054 724
rect 495122 668 495178 724
rect 495246 668 495302 724
rect 494874 544 494930 600
rect 494998 544 495054 600
rect 495122 544 495178 600
rect 495246 544 495302 600
rect 494874 420 494930 476
rect 494998 420 495054 476
rect 495122 420 495178 476
rect 495246 420 495302 476
rect 509154 1752 509210 1808
rect 509278 1752 509334 1808
rect 509402 1752 509458 1808
rect 509526 1752 509582 1808
rect 509154 1628 509210 1684
rect 509278 1628 509334 1684
rect 509402 1628 509458 1684
rect 509526 1628 509582 1684
rect 509154 1504 509210 1560
rect 509278 1504 509334 1560
rect 509402 1504 509458 1560
rect 509526 1504 509582 1560
rect 509154 1380 509210 1436
rect 509278 1380 509334 1436
rect 509402 1380 509458 1436
rect 509526 1380 509582 1436
rect 512874 792 512930 848
rect 512998 792 513054 848
rect 513122 792 513178 848
rect 513246 792 513302 848
rect 512874 668 512930 724
rect 512998 668 513054 724
rect 513122 668 513178 724
rect 513246 668 513302 724
rect 512874 544 512930 600
rect 512998 544 513054 600
rect 513122 544 513178 600
rect 513246 544 513302 600
rect 512874 420 512930 476
rect 512998 420 513054 476
rect 513122 420 513178 476
rect 513246 420 513302 476
rect 527154 1752 527210 1808
rect 527278 1752 527334 1808
rect 527402 1752 527458 1808
rect 527526 1752 527582 1808
rect 527154 1628 527210 1684
rect 527278 1628 527334 1684
rect 527402 1628 527458 1684
rect 527526 1628 527582 1684
rect 527154 1504 527210 1560
rect 527278 1504 527334 1560
rect 527402 1504 527458 1560
rect 527526 1504 527582 1560
rect 527154 1380 527210 1436
rect 527278 1380 527334 1436
rect 527402 1380 527458 1436
rect 527526 1380 527582 1436
rect 530874 792 530930 848
rect 530998 792 531054 848
rect 531122 792 531178 848
rect 531246 792 531302 848
rect 530874 668 530930 724
rect 530998 668 531054 724
rect 531122 668 531178 724
rect 531246 668 531302 724
rect 530874 544 530930 600
rect 530998 544 531054 600
rect 531122 544 531178 600
rect 531246 544 531302 600
rect 530874 420 530930 476
rect 530998 420 531054 476
rect 531122 420 531178 476
rect 531246 420 531302 476
rect 545154 1752 545210 1808
rect 545278 1752 545334 1808
rect 545402 1752 545458 1808
rect 545526 1752 545582 1808
rect 545154 1628 545210 1684
rect 545278 1628 545334 1684
rect 545402 1628 545458 1684
rect 545526 1628 545582 1684
rect 545154 1504 545210 1560
rect 545278 1504 545334 1560
rect 545402 1504 545458 1560
rect 545526 1504 545582 1560
rect 545154 1380 545210 1436
rect 545278 1380 545334 1436
rect 545402 1380 545458 1436
rect 545526 1380 545582 1436
rect 548874 792 548930 848
rect 548998 792 549054 848
rect 549122 792 549178 848
rect 549246 792 549302 848
rect 548874 668 548930 724
rect 548998 668 549054 724
rect 549122 668 549178 724
rect 549246 668 549302 724
rect 548874 544 548930 600
rect 548998 544 549054 600
rect 549122 544 549178 600
rect 549246 544 549302 600
rect 548874 420 548930 476
rect 548998 420 549054 476
rect 549122 420 549178 476
rect 549246 420 549302 476
rect 563154 1752 563210 1808
rect 563278 1752 563334 1808
rect 563402 1752 563458 1808
rect 563526 1752 563582 1808
rect 563154 1628 563210 1684
rect 563278 1628 563334 1684
rect 563402 1628 563458 1684
rect 563526 1628 563582 1684
rect 563154 1504 563210 1560
rect 563278 1504 563334 1560
rect 563402 1504 563458 1560
rect 563526 1504 563582 1560
rect 563154 1380 563210 1436
rect 563278 1380 563334 1436
rect 563402 1380 563458 1436
rect 563526 1380 563582 1436
rect 566874 792 566930 848
rect 566998 792 567054 848
rect 567122 792 567178 848
rect 567246 792 567302 848
rect 566874 668 566930 724
rect 566998 668 567054 724
rect 567122 668 567178 724
rect 567246 668 567302 724
rect 566874 544 566930 600
rect 566998 544 567054 600
rect 567122 544 567178 600
rect 567246 544 567302 600
rect 566874 420 566930 476
rect 566998 420 567054 476
rect 567122 420 567178 476
rect 567246 420 567302 476
rect 581154 1752 581210 1808
rect 581278 1752 581334 1808
rect 581402 1752 581458 1808
rect 581526 1752 581582 1808
rect 581154 1628 581210 1684
rect 581278 1628 581334 1684
rect 581402 1628 581458 1684
rect 581526 1628 581582 1684
rect 581154 1504 581210 1560
rect 581278 1504 581334 1560
rect 581402 1504 581458 1560
rect 581526 1504 581582 1560
rect 581154 1380 581210 1436
rect 581278 1380 581334 1436
rect 581402 1380 581458 1436
rect 581526 1380 581582 1436
rect 598512 1752 598568 1808
rect 598636 1752 598692 1808
rect 598760 1752 598816 1808
rect 598884 1752 598940 1808
rect 598512 1628 598568 1684
rect 598636 1628 598692 1684
rect 598760 1628 598816 1684
rect 598884 1628 598940 1684
rect 598512 1504 598568 1560
rect 598636 1504 598692 1560
rect 598760 1504 598816 1560
rect 598884 1504 598940 1560
rect 598512 1380 598568 1436
rect 598636 1380 598692 1436
rect 598760 1380 598816 1436
rect 598884 1380 598940 1436
rect 599472 587862 599528 587918
rect 599596 587862 599652 587918
rect 599720 587862 599776 587918
rect 599844 587862 599900 587918
rect 599472 587738 599528 587794
rect 599596 587738 599652 587794
rect 599720 587738 599776 587794
rect 599844 587738 599900 587794
rect 599472 587614 599528 587670
rect 599596 587614 599652 587670
rect 599720 587614 599776 587670
rect 599844 587614 599900 587670
rect 599472 587490 599528 587546
rect 599596 587490 599652 587546
rect 599720 587490 599776 587546
rect 599844 587490 599900 587546
rect 599472 569862 599528 569918
rect 599596 569862 599652 569918
rect 599720 569862 599776 569918
rect 599844 569862 599900 569918
rect 599472 569738 599528 569794
rect 599596 569738 599652 569794
rect 599720 569738 599776 569794
rect 599844 569738 599900 569794
rect 599472 569614 599528 569670
rect 599596 569614 599652 569670
rect 599720 569614 599776 569670
rect 599844 569614 599900 569670
rect 599472 569490 599528 569546
rect 599596 569490 599652 569546
rect 599720 569490 599776 569546
rect 599844 569490 599900 569546
rect 599472 551862 599528 551918
rect 599596 551862 599652 551918
rect 599720 551862 599776 551918
rect 599844 551862 599900 551918
rect 599472 551738 599528 551794
rect 599596 551738 599652 551794
rect 599720 551738 599776 551794
rect 599844 551738 599900 551794
rect 599472 551614 599528 551670
rect 599596 551614 599652 551670
rect 599720 551614 599776 551670
rect 599844 551614 599900 551670
rect 599472 551490 599528 551546
rect 599596 551490 599652 551546
rect 599720 551490 599776 551546
rect 599844 551490 599900 551546
rect 599472 533862 599528 533918
rect 599596 533862 599652 533918
rect 599720 533862 599776 533918
rect 599844 533862 599900 533918
rect 599472 533738 599528 533794
rect 599596 533738 599652 533794
rect 599720 533738 599776 533794
rect 599844 533738 599900 533794
rect 599472 533614 599528 533670
rect 599596 533614 599652 533670
rect 599720 533614 599776 533670
rect 599844 533614 599900 533670
rect 599472 533490 599528 533546
rect 599596 533490 599652 533546
rect 599720 533490 599776 533546
rect 599844 533490 599900 533546
rect 599472 515862 599528 515918
rect 599596 515862 599652 515918
rect 599720 515862 599776 515918
rect 599844 515862 599900 515918
rect 599472 515738 599528 515794
rect 599596 515738 599652 515794
rect 599720 515738 599776 515794
rect 599844 515738 599900 515794
rect 599472 515614 599528 515670
rect 599596 515614 599652 515670
rect 599720 515614 599776 515670
rect 599844 515614 599900 515670
rect 599472 515490 599528 515546
rect 599596 515490 599652 515546
rect 599720 515490 599776 515546
rect 599844 515490 599900 515546
rect 599472 497862 599528 497918
rect 599596 497862 599652 497918
rect 599720 497862 599776 497918
rect 599844 497862 599900 497918
rect 599472 497738 599528 497794
rect 599596 497738 599652 497794
rect 599720 497738 599776 497794
rect 599844 497738 599900 497794
rect 599472 497614 599528 497670
rect 599596 497614 599652 497670
rect 599720 497614 599776 497670
rect 599844 497614 599900 497670
rect 599472 497490 599528 497546
rect 599596 497490 599652 497546
rect 599720 497490 599776 497546
rect 599844 497490 599900 497546
rect 599472 479862 599528 479918
rect 599596 479862 599652 479918
rect 599720 479862 599776 479918
rect 599844 479862 599900 479918
rect 599472 479738 599528 479794
rect 599596 479738 599652 479794
rect 599720 479738 599776 479794
rect 599844 479738 599900 479794
rect 599472 479614 599528 479670
rect 599596 479614 599652 479670
rect 599720 479614 599776 479670
rect 599844 479614 599900 479670
rect 599472 479490 599528 479546
rect 599596 479490 599652 479546
rect 599720 479490 599776 479546
rect 599844 479490 599900 479546
rect 599472 461862 599528 461918
rect 599596 461862 599652 461918
rect 599720 461862 599776 461918
rect 599844 461862 599900 461918
rect 599472 461738 599528 461794
rect 599596 461738 599652 461794
rect 599720 461738 599776 461794
rect 599844 461738 599900 461794
rect 599472 461614 599528 461670
rect 599596 461614 599652 461670
rect 599720 461614 599776 461670
rect 599844 461614 599900 461670
rect 599472 461490 599528 461546
rect 599596 461490 599652 461546
rect 599720 461490 599776 461546
rect 599844 461490 599900 461546
rect 599472 443862 599528 443918
rect 599596 443862 599652 443918
rect 599720 443862 599776 443918
rect 599844 443862 599900 443918
rect 599472 443738 599528 443794
rect 599596 443738 599652 443794
rect 599720 443738 599776 443794
rect 599844 443738 599900 443794
rect 599472 443614 599528 443670
rect 599596 443614 599652 443670
rect 599720 443614 599776 443670
rect 599844 443614 599900 443670
rect 599472 443490 599528 443546
rect 599596 443490 599652 443546
rect 599720 443490 599776 443546
rect 599844 443490 599900 443546
rect 599472 425862 599528 425918
rect 599596 425862 599652 425918
rect 599720 425862 599776 425918
rect 599844 425862 599900 425918
rect 599472 425738 599528 425794
rect 599596 425738 599652 425794
rect 599720 425738 599776 425794
rect 599844 425738 599900 425794
rect 599472 425614 599528 425670
rect 599596 425614 599652 425670
rect 599720 425614 599776 425670
rect 599844 425614 599900 425670
rect 599472 425490 599528 425546
rect 599596 425490 599652 425546
rect 599720 425490 599776 425546
rect 599844 425490 599900 425546
rect 599472 407862 599528 407918
rect 599596 407862 599652 407918
rect 599720 407862 599776 407918
rect 599844 407862 599900 407918
rect 599472 407738 599528 407794
rect 599596 407738 599652 407794
rect 599720 407738 599776 407794
rect 599844 407738 599900 407794
rect 599472 407614 599528 407670
rect 599596 407614 599652 407670
rect 599720 407614 599776 407670
rect 599844 407614 599900 407670
rect 599472 407490 599528 407546
rect 599596 407490 599652 407546
rect 599720 407490 599776 407546
rect 599844 407490 599900 407546
rect 599472 389862 599528 389918
rect 599596 389862 599652 389918
rect 599720 389862 599776 389918
rect 599844 389862 599900 389918
rect 599472 389738 599528 389794
rect 599596 389738 599652 389794
rect 599720 389738 599776 389794
rect 599844 389738 599900 389794
rect 599472 389614 599528 389670
rect 599596 389614 599652 389670
rect 599720 389614 599776 389670
rect 599844 389614 599900 389670
rect 599472 389490 599528 389546
rect 599596 389490 599652 389546
rect 599720 389490 599776 389546
rect 599844 389490 599900 389546
rect 599472 371862 599528 371918
rect 599596 371862 599652 371918
rect 599720 371862 599776 371918
rect 599844 371862 599900 371918
rect 599472 371738 599528 371794
rect 599596 371738 599652 371794
rect 599720 371738 599776 371794
rect 599844 371738 599900 371794
rect 599472 371614 599528 371670
rect 599596 371614 599652 371670
rect 599720 371614 599776 371670
rect 599844 371614 599900 371670
rect 599472 371490 599528 371546
rect 599596 371490 599652 371546
rect 599720 371490 599776 371546
rect 599844 371490 599900 371546
rect 599472 353862 599528 353918
rect 599596 353862 599652 353918
rect 599720 353862 599776 353918
rect 599844 353862 599900 353918
rect 599472 353738 599528 353794
rect 599596 353738 599652 353794
rect 599720 353738 599776 353794
rect 599844 353738 599900 353794
rect 599472 353614 599528 353670
rect 599596 353614 599652 353670
rect 599720 353614 599776 353670
rect 599844 353614 599900 353670
rect 599472 353490 599528 353546
rect 599596 353490 599652 353546
rect 599720 353490 599776 353546
rect 599844 353490 599900 353546
rect 599472 335862 599528 335918
rect 599596 335862 599652 335918
rect 599720 335862 599776 335918
rect 599844 335862 599900 335918
rect 599472 335738 599528 335794
rect 599596 335738 599652 335794
rect 599720 335738 599776 335794
rect 599844 335738 599900 335794
rect 599472 335614 599528 335670
rect 599596 335614 599652 335670
rect 599720 335614 599776 335670
rect 599844 335614 599900 335670
rect 599472 335490 599528 335546
rect 599596 335490 599652 335546
rect 599720 335490 599776 335546
rect 599844 335490 599900 335546
rect 599472 317862 599528 317918
rect 599596 317862 599652 317918
rect 599720 317862 599776 317918
rect 599844 317862 599900 317918
rect 599472 317738 599528 317794
rect 599596 317738 599652 317794
rect 599720 317738 599776 317794
rect 599844 317738 599900 317794
rect 599472 317614 599528 317670
rect 599596 317614 599652 317670
rect 599720 317614 599776 317670
rect 599844 317614 599900 317670
rect 599472 317490 599528 317546
rect 599596 317490 599652 317546
rect 599720 317490 599776 317546
rect 599844 317490 599900 317546
rect 599472 299862 599528 299918
rect 599596 299862 599652 299918
rect 599720 299862 599776 299918
rect 599844 299862 599900 299918
rect 599472 299738 599528 299794
rect 599596 299738 599652 299794
rect 599720 299738 599776 299794
rect 599844 299738 599900 299794
rect 599472 299614 599528 299670
rect 599596 299614 599652 299670
rect 599720 299614 599776 299670
rect 599844 299614 599900 299670
rect 599472 299490 599528 299546
rect 599596 299490 599652 299546
rect 599720 299490 599776 299546
rect 599844 299490 599900 299546
rect 599472 281862 599528 281918
rect 599596 281862 599652 281918
rect 599720 281862 599776 281918
rect 599844 281862 599900 281918
rect 599472 281738 599528 281794
rect 599596 281738 599652 281794
rect 599720 281738 599776 281794
rect 599844 281738 599900 281794
rect 599472 281614 599528 281670
rect 599596 281614 599652 281670
rect 599720 281614 599776 281670
rect 599844 281614 599900 281670
rect 599472 281490 599528 281546
rect 599596 281490 599652 281546
rect 599720 281490 599776 281546
rect 599844 281490 599900 281546
rect 599472 263862 599528 263918
rect 599596 263862 599652 263918
rect 599720 263862 599776 263918
rect 599844 263862 599900 263918
rect 599472 263738 599528 263794
rect 599596 263738 599652 263794
rect 599720 263738 599776 263794
rect 599844 263738 599900 263794
rect 599472 263614 599528 263670
rect 599596 263614 599652 263670
rect 599720 263614 599776 263670
rect 599844 263614 599900 263670
rect 599472 263490 599528 263546
rect 599596 263490 599652 263546
rect 599720 263490 599776 263546
rect 599844 263490 599900 263546
rect 599472 245862 599528 245918
rect 599596 245862 599652 245918
rect 599720 245862 599776 245918
rect 599844 245862 599900 245918
rect 599472 245738 599528 245794
rect 599596 245738 599652 245794
rect 599720 245738 599776 245794
rect 599844 245738 599900 245794
rect 599472 245614 599528 245670
rect 599596 245614 599652 245670
rect 599720 245614 599776 245670
rect 599844 245614 599900 245670
rect 599472 245490 599528 245546
rect 599596 245490 599652 245546
rect 599720 245490 599776 245546
rect 599844 245490 599900 245546
rect 599472 227862 599528 227918
rect 599596 227862 599652 227918
rect 599720 227862 599776 227918
rect 599844 227862 599900 227918
rect 599472 227738 599528 227794
rect 599596 227738 599652 227794
rect 599720 227738 599776 227794
rect 599844 227738 599900 227794
rect 599472 227614 599528 227670
rect 599596 227614 599652 227670
rect 599720 227614 599776 227670
rect 599844 227614 599900 227670
rect 599472 227490 599528 227546
rect 599596 227490 599652 227546
rect 599720 227490 599776 227546
rect 599844 227490 599900 227546
rect 599472 209862 599528 209918
rect 599596 209862 599652 209918
rect 599720 209862 599776 209918
rect 599844 209862 599900 209918
rect 599472 209738 599528 209794
rect 599596 209738 599652 209794
rect 599720 209738 599776 209794
rect 599844 209738 599900 209794
rect 599472 209614 599528 209670
rect 599596 209614 599652 209670
rect 599720 209614 599776 209670
rect 599844 209614 599900 209670
rect 599472 209490 599528 209546
rect 599596 209490 599652 209546
rect 599720 209490 599776 209546
rect 599844 209490 599900 209546
rect 599472 191862 599528 191918
rect 599596 191862 599652 191918
rect 599720 191862 599776 191918
rect 599844 191862 599900 191918
rect 599472 191738 599528 191794
rect 599596 191738 599652 191794
rect 599720 191738 599776 191794
rect 599844 191738 599900 191794
rect 599472 191614 599528 191670
rect 599596 191614 599652 191670
rect 599720 191614 599776 191670
rect 599844 191614 599900 191670
rect 599472 191490 599528 191546
rect 599596 191490 599652 191546
rect 599720 191490 599776 191546
rect 599844 191490 599900 191546
rect 599472 173862 599528 173918
rect 599596 173862 599652 173918
rect 599720 173862 599776 173918
rect 599844 173862 599900 173918
rect 599472 173738 599528 173794
rect 599596 173738 599652 173794
rect 599720 173738 599776 173794
rect 599844 173738 599900 173794
rect 599472 173614 599528 173670
rect 599596 173614 599652 173670
rect 599720 173614 599776 173670
rect 599844 173614 599900 173670
rect 599472 173490 599528 173546
rect 599596 173490 599652 173546
rect 599720 173490 599776 173546
rect 599844 173490 599900 173546
rect 599472 155862 599528 155918
rect 599596 155862 599652 155918
rect 599720 155862 599776 155918
rect 599844 155862 599900 155918
rect 599472 155738 599528 155794
rect 599596 155738 599652 155794
rect 599720 155738 599776 155794
rect 599844 155738 599900 155794
rect 599472 155614 599528 155670
rect 599596 155614 599652 155670
rect 599720 155614 599776 155670
rect 599844 155614 599900 155670
rect 599472 155490 599528 155546
rect 599596 155490 599652 155546
rect 599720 155490 599776 155546
rect 599844 155490 599900 155546
rect 599472 137862 599528 137918
rect 599596 137862 599652 137918
rect 599720 137862 599776 137918
rect 599844 137862 599900 137918
rect 599472 137738 599528 137794
rect 599596 137738 599652 137794
rect 599720 137738 599776 137794
rect 599844 137738 599900 137794
rect 599472 137614 599528 137670
rect 599596 137614 599652 137670
rect 599720 137614 599776 137670
rect 599844 137614 599900 137670
rect 599472 137490 599528 137546
rect 599596 137490 599652 137546
rect 599720 137490 599776 137546
rect 599844 137490 599900 137546
rect 599472 119862 599528 119918
rect 599596 119862 599652 119918
rect 599720 119862 599776 119918
rect 599844 119862 599900 119918
rect 599472 119738 599528 119794
rect 599596 119738 599652 119794
rect 599720 119738 599776 119794
rect 599844 119738 599900 119794
rect 599472 119614 599528 119670
rect 599596 119614 599652 119670
rect 599720 119614 599776 119670
rect 599844 119614 599900 119670
rect 599472 119490 599528 119546
rect 599596 119490 599652 119546
rect 599720 119490 599776 119546
rect 599844 119490 599900 119546
rect 599472 101862 599528 101918
rect 599596 101862 599652 101918
rect 599720 101862 599776 101918
rect 599844 101862 599900 101918
rect 599472 101738 599528 101794
rect 599596 101738 599652 101794
rect 599720 101738 599776 101794
rect 599844 101738 599900 101794
rect 599472 101614 599528 101670
rect 599596 101614 599652 101670
rect 599720 101614 599776 101670
rect 599844 101614 599900 101670
rect 599472 101490 599528 101546
rect 599596 101490 599652 101546
rect 599720 101490 599776 101546
rect 599844 101490 599900 101546
rect 599472 83862 599528 83918
rect 599596 83862 599652 83918
rect 599720 83862 599776 83918
rect 599844 83862 599900 83918
rect 599472 83738 599528 83794
rect 599596 83738 599652 83794
rect 599720 83738 599776 83794
rect 599844 83738 599900 83794
rect 599472 83614 599528 83670
rect 599596 83614 599652 83670
rect 599720 83614 599776 83670
rect 599844 83614 599900 83670
rect 599472 83490 599528 83546
rect 599596 83490 599652 83546
rect 599720 83490 599776 83546
rect 599844 83490 599900 83546
rect 599472 65862 599528 65918
rect 599596 65862 599652 65918
rect 599720 65862 599776 65918
rect 599844 65862 599900 65918
rect 599472 65738 599528 65794
rect 599596 65738 599652 65794
rect 599720 65738 599776 65794
rect 599844 65738 599900 65794
rect 599472 65614 599528 65670
rect 599596 65614 599652 65670
rect 599720 65614 599776 65670
rect 599844 65614 599900 65670
rect 599472 65490 599528 65546
rect 599596 65490 599652 65546
rect 599720 65490 599776 65546
rect 599844 65490 599900 65546
rect 599472 47862 599528 47918
rect 599596 47862 599652 47918
rect 599720 47862 599776 47918
rect 599844 47862 599900 47918
rect 599472 47738 599528 47794
rect 599596 47738 599652 47794
rect 599720 47738 599776 47794
rect 599844 47738 599900 47794
rect 599472 47614 599528 47670
rect 599596 47614 599652 47670
rect 599720 47614 599776 47670
rect 599844 47614 599900 47670
rect 599472 47490 599528 47546
rect 599596 47490 599652 47546
rect 599720 47490 599776 47546
rect 599844 47490 599900 47546
rect 599472 29862 599528 29918
rect 599596 29862 599652 29918
rect 599720 29862 599776 29918
rect 599844 29862 599900 29918
rect 599472 29738 599528 29794
rect 599596 29738 599652 29794
rect 599720 29738 599776 29794
rect 599844 29738 599900 29794
rect 599472 29614 599528 29670
rect 599596 29614 599652 29670
rect 599720 29614 599776 29670
rect 599844 29614 599900 29670
rect 599472 29490 599528 29546
rect 599596 29490 599652 29546
rect 599720 29490 599776 29546
rect 599844 29490 599900 29546
rect 599472 11862 599528 11918
rect 599596 11862 599652 11918
rect 599720 11862 599776 11918
rect 599844 11862 599900 11918
rect 599472 11738 599528 11794
rect 599596 11738 599652 11794
rect 599720 11738 599776 11794
rect 599844 11738 599900 11794
rect 599472 11614 599528 11670
rect 599596 11614 599652 11670
rect 599720 11614 599776 11670
rect 599844 11614 599900 11670
rect 599472 11490 599528 11546
rect 599596 11490 599652 11546
rect 599720 11490 599776 11546
rect 599844 11490 599900 11546
rect 584874 792 584930 848
rect 584998 792 585054 848
rect 585122 792 585178 848
rect 585246 792 585302 848
rect 584874 668 584930 724
rect 584998 668 585054 724
rect 585122 668 585178 724
rect 585246 668 585302 724
rect 584874 544 584930 600
rect 584998 544 585054 600
rect 585122 544 585178 600
rect 585246 544 585302 600
rect 584874 420 584930 476
rect 584998 420 585054 476
rect 585122 420 585178 476
rect 585246 420 585302 476
rect 599472 792 599528 848
rect 599596 792 599652 848
rect 599720 792 599776 848
rect 599844 792 599900 848
rect 599472 668 599528 724
rect 599596 668 599652 724
rect 599720 668 599776 724
rect 599844 668 599900 724
rect 599472 544 599528 600
rect 599596 544 599652 600
rect 599720 544 599776 600
rect 599844 544 599900 600
rect 599472 420 599528 476
rect 599596 420 599652 476
rect 599720 420 599776 476
rect 599844 420 599900 476
<< metal5 >>
rect -12 599340 599996 599436
rect -12 599284 84 599340
rect 140 599284 208 599340
rect 264 599284 332 599340
rect 388 599284 456 599340
rect 512 599284 8874 599340
rect 8930 599284 8998 599340
rect 9054 599284 9122 599340
rect 9178 599284 9246 599340
rect 9302 599284 26874 599340
rect 26930 599284 26998 599340
rect 27054 599284 27122 599340
rect 27178 599284 27246 599340
rect 27302 599284 44874 599340
rect 44930 599284 44998 599340
rect 45054 599284 45122 599340
rect 45178 599284 45246 599340
rect 45302 599284 62874 599340
rect 62930 599284 62998 599340
rect 63054 599284 63122 599340
rect 63178 599284 63246 599340
rect 63302 599284 80874 599340
rect 80930 599284 80998 599340
rect 81054 599284 81122 599340
rect 81178 599284 81246 599340
rect 81302 599284 98874 599340
rect 98930 599284 98998 599340
rect 99054 599284 99122 599340
rect 99178 599284 99246 599340
rect 99302 599284 116874 599340
rect 116930 599284 116998 599340
rect 117054 599284 117122 599340
rect 117178 599284 117246 599340
rect 117302 599284 134874 599340
rect 134930 599284 134998 599340
rect 135054 599284 135122 599340
rect 135178 599284 135246 599340
rect 135302 599284 152874 599340
rect 152930 599284 152998 599340
rect 153054 599284 153122 599340
rect 153178 599284 153246 599340
rect 153302 599284 170874 599340
rect 170930 599284 170998 599340
rect 171054 599284 171122 599340
rect 171178 599284 171246 599340
rect 171302 599284 188874 599340
rect 188930 599284 188998 599340
rect 189054 599284 189122 599340
rect 189178 599284 189246 599340
rect 189302 599284 206874 599340
rect 206930 599284 206998 599340
rect 207054 599284 207122 599340
rect 207178 599284 207246 599340
rect 207302 599284 224874 599340
rect 224930 599284 224998 599340
rect 225054 599284 225122 599340
rect 225178 599284 225246 599340
rect 225302 599284 242874 599340
rect 242930 599284 242998 599340
rect 243054 599284 243122 599340
rect 243178 599284 243246 599340
rect 243302 599284 260874 599340
rect 260930 599284 260998 599340
rect 261054 599284 261122 599340
rect 261178 599284 261246 599340
rect 261302 599284 278874 599340
rect 278930 599284 278998 599340
rect 279054 599284 279122 599340
rect 279178 599284 279246 599340
rect 279302 599284 296874 599340
rect 296930 599284 296998 599340
rect 297054 599284 297122 599340
rect 297178 599284 297246 599340
rect 297302 599284 314874 599340
rect 314930 599284 314998 599340
rect 315054 599284 315122 599340
rect 315178 599284 315246 599340
rect 315302 599284 332874 599340
rect 332930 599284 332998 599340
rect 333054 599284 333122 599340
rect 333178 599284 333246 599340
rect 333302 599284 350874 599340
rect 350930 599284 350998 599340
rect 351054 599284 351122 599340
rect 351178 599284 351246 599340
rect 351302 599284 368874 599340
rect 368930 599284 368998 599340
rect 369054 599284 369122 599340
rect 369178 599284 369246 599340
rect 369302 599284 386874 599340
rect 386930 599284 386998 599340
rect 387054 599284 387122 599340
rect 387178 599284 387246 599340
rect 387302 599284 404874 599340
rect 404930 599284 404998 599340
rect 405054 599284 405122 599340
rect 405178 599284 405246 599340
rect 405302 599284 422874 599340
rect 422930 599284 422998 599340
rect 423054 599284 423122 599340
rect 423178 599284 423246 599340
rect 423302 599284 440874 599340
rect 440930 599284 440998 599340
rect 441054 599284 441122 599340
rect 441178 599284 441246 599340
rect 441302 599284 458874 599340
rect 458930 599284 458998 599340
rect 459054 599284 459122 599340
rect 459178 599284 459246 599340
rect 459302 599284 476874 599340
rect 476930 599284 476998 599340
rect 477054 599284 477122 599340
rect 477178 599284 477246 599340
rect 477302 599284 494874 599340
rect 494930 599284 494998 599340
rect 495054 599284 495122 599340
rect 495178 599284 495246 599340
rect 495302 599284 512874 599340
rect 512930 599284 512998 599340
rect 513054 599284 513122 599340
rect 513178 599284 513246 599340
rect 513302 599284 530874 599340
rect 530930 599284 530998 599340
rect 531054 599284 531122 599340
rect 531178 599284 531246 599340
rect 531302 599284 548874 599340
rect 548930 599284 548998 599340
rect 549054 599284 549122 599340
rect 549178 599284 549246 599340
rect 549302 599284 566874 599340
rect 566930 599284 566998 599340
rect 567054 599284 567122 599340
rect 567178 599284 567246 599340
rect 567302 599284 584874 599340
rect 584930 599284 584998 599340
rect 585054 599284 585122 599340
rect 585178 599284 585246 599340
rect 585302 599284 599472 599340
rect 599528 599284 599596 599340
rect 599652 599284 599720 599340
rect 599776 599284 599844 599340
rect 599900 599284 599996 599340
rect -12 599216 599996 599284
rect -12 599160 84 599216
rect 140 599160 208 599216
rect 264 599160 332 599216
rect 388 599160 456 599216
rect 512 599160 8874 599216
rect 8930 599160 8998 599216
rect 9054 599160 9122 599216
rect 9178 599160 9246 599216
rect 9302 599160 26874 599216
rect 26930 599160 26998 599216
rect 27054 599160 27122 599216
rect 27178 599160 27246 599216
rect 27302 599160 44874 599216
rect 44930 599160 44998 599216
rect 45054 599160 45122 599216
rect 45178 599160 45246 599216
rect 45302 599160 62874 599216
rect 62930 599160 62998 599216
rect 63054 599160 63122 599216
rect 63178 599160 63246 599216
rect 63302 599160 80874 599216
rect 80930 599160 80998 599216
rect 81054 599160 81122 599216
rect 81178 599160 81246 599216
rect 81302 599160 98874 599216
rect 98930 599160 98998 599216
rect 99054 599160 99122 599216
rect 99178 599160 99246 599216
rect 99302 599160 116874 599216
rect 116930 599160 116998 599216
rect 117054 599160 117122 599216
rect 117178 599160 117246 599216
rect 117302 599160 134874 599216
rect 134930 599160 134998 599216
rect 135054 599160 135122 599216
rect 135178 599160 135246 599216
rect 135302 599160 152874 599216
rect 152930 599160 152998 599216
rect 153054 599160 153122 599216
rect 153178 599160 153246 599216
rect 153302 599160 170874 599216
rect 170930 599160 170998 599216
rect 171054 599160 171122 599216
rect 171178 599160 171246 599216
rect 171302 599160 188874 599216
rect 188930 599160 188998 599216
rect 189054 599160 189122 599216
rect 189178 599160 189246 599216
rect 189302 599160 206874 599216
rect 206930 599160 206998 599216
rect 207054 599160 207122 599216
rect 207178 599160 207246 599216
rect 207302 599160 224874 599216
rect 224930 599160 224998 599216
rect 225054 599160 225122 599216
rect 225178 599160 225246 599216
rect 225302 599160 242874 599216
rect 242930 599160 242998 599216
rect 243054 599160 243122 599216
rect 243178 599160 243246 599216
rect 243302 599160 260874 599216
rect 260930 599160 260998 599216
rect 261054 599160 261122 599216
rect 261178 599160 261246 599216
rect 261302 599160 278874 599216
rect 278930 599160 278998 599216
rect 279054 599160 279122 599216
rect 279178 599160 279246 599216
rect 279302 599160 296874 599216
rect 296930 599160 296998 599216
rect 297054 599160 297122 599216
rect 297178 599160 297246 599216
rect 297302 599160 314874 599216
rect 314930 599160 314998 599216
rect 315054 599160 315122 599216
rect 315178 599160 315246 599216
rect 315302 599160 332874 599216
rect 332930 599160 332998 599216
rect 333054 599160 333122 599216
rect 333178 599160 333246 599216
rect 333302 599160 350874 599216
rect 350930 599160 350998 599216
rect 351054 599160 351122 599216
rect 351178 599160 351246 599216
rect 351302 599160 368874 599216
rect 368930 599160 368998 599216
rect 369054 599160 369122 599216
rect 369178 599160 369246 599216
rect 369302 599160 386874 599216
rect 386930 599160 386998 599216
rect 387054 599160 387122 599216
rect 387178 599160 387246 599216
rect 387302 599160 404874 599216
rect 404930 599160 404998 599216
rect 405054 599160 405122 599216
rect 405178 599160 405246 599216
rect 405302 599160 422874 599216
rect 422930 599160 422998 599216
rect 423054 599160 423122 599216
rect 423178 599160 423246 599216
rect 423302 599160 440874 599216
rect 440930 599160 440998 599216
rect 441054 599160 441122 599216
rect 441178 599160 441246 599216
rect 441302 599160 458874 599216
rect 458930 599160 458998 599216
rect 459054 599160 459122 599216
rect 459178 599160 459246 599216
rect 459302 599160 476874 599216
rect 476930 599160 476998 599216
rect 477054 599160 477122 599216
rect 477178 599160 477246 599216
rect 477302 599160 494874 599216
rect 494930 599160 494998 599216
rect 495054 599160 495122 599216
rect 495178 599160 495246 599216
rect 495302 599160 512874 599216
rect 512930 599160 512998 599216
rect 513054 599160 513122 599216
rect 513178 599160 513246 599216
rect 513302 599160 530874 599216
rect 530930 599160 530998 599216
rect 531054 599160 531122 599216
rect 531178 599160 531246 599216
rect 531302 599160 548874 599216
rect 548930 599160 548998 599216
rect 549054 599160 549122 599216
rect 549178 599160 549246 599216
rect 549302 599160 566874 599216
rect 566930 599160 566998 599216
rect 567054 599160 567122 599216
rect 567178 599160 567246 599216
rect 567302 599160 584874 599216
rect 584930 599160 584998 599216
rect 585054 599160 585122 599216
rect 585178 599160 585246 599216
rect 585302 599160 599472 599216
rect 599528 599160 599596 599216
rect 599652 599160 599720 599216
rect 599776 599160 599844 599216
rect 599900 599160 599996 599216
rect -12 599092 599996 599160
rect -12 599036 84 599092
rect 140 599036 208 599092
rect 264 599036 332 599092
rect 388 599036 456 599092
rect 512 599036 8874 599092
rect 8930 599036 8998 599092
rect 9054 599036 9122 599092
rect 9178 599036 9246 599092
rect 9302 599036 26874 599092
rect 26930 599036 26998 599092
rect 27054 599036 27122 599092
rect 27178 599036 27246 599092
rect 27302 599036 44874 599092
rect 44930 599036 44998 599092
rect 45054 599036 45122 599092
rect 45178 599036 45246 599092
rect 45302 599036 62874 599092
rect 62930 599036 62998 599092
rect 63054 599036 63122 599092
rect 63178 599036 63246 599092
rect 63302 599036 80874 599092
rect 80930 599036 80998 599092
rect 81054 599036 81122 599092
rect 81178 599036 81246 599092
rect 81302 599036 98874 599092
rect 98930 599036 98998 599092
rect 99054 599036 99122 599092
rect 99178 599036 99246 599092
rect 99302 599036 116874 599092
rect 116930 599036 116998 599092
rect 117054 599036 117122 599092
rect 117178 599036 117246 599092
rect 117302 599036 134874 599092
rect 134930 599036 134998 599092
rect 135054 599036 135122 599092
rect 135178 599036 135246 599092
rect 135302 599036 152874 599092
rect 152930 599036 152998 599092
rect 153054 599036 153122 599092
rect 153178 599036 153246 599092
rect 153302 599036 170874 599092
rect 170930 599036 170998 599092
rect 171054 599036 171122 599092
rect 171178 599036 171246 599092
rect 171302 599036 188874 599092
rect 188930 599036 188998 599092
rect 189054 599036 189122 599092
rect 189178 599036 189246 599092
rect 189302 599036 206874 599092
rect 206930 599036 206998 599092
rect 207054 599036 207122 599092
rect 207178 599036 207246 599092
rect 207302 599036 224874 599092
rect 224930 599036 224998 599092
rect 225054 599036 225122 599092
rect 225178 599036 225246 599092
rect 225302 599036 242874 599092
rect 242930 599036 242998 599092
rect 243054 599036 243122 599092
rect 243178 599036 243246 599092
rect 243302 599036 260874 599092
rect 260930 599036 260998 599092
rect 261054 599036 261122 599092
rect 261178 599036 261246 599092
rect 261302 599036 278874 599092
rect 278930 599036 278998 599092
rect 279054 599036 279122 599092
rect 279178 599036 279246 599092
rect 279302 599036 296874 599092
rect 296930 599036 296998 599092
rect 297054 599036 297122 599092
rect 297178 599036 297246 599092
rect 297302 599036 314874 599092
rect 314930 599036 314998 599092
rect 315054 599036 315122 599092
rect 315178 599036 315246 599092
rect 315302 599036 332874 599092
rect 332930 599036 332998 599092
rect 333054 599036 333122 599092
rect 333178 599036 333246 599092
rect 333302 599036 350874 599092
rect 350930 599036 350998 599092
rect 351054 599036 351122 599092
rect 351178 599036 351246 599092
rect 351302 599036 368874 599092
rect 368930 599036 368998 599092
rect 369054 599036 369122 599092
rect 369178 599036 369246 599092
rect 369302 599036 386874 599092
rect 386930 599036 386998 599092
rect 387054 599036 387122 599092
rect 387178 599036 387246 599092
rect 387302 599036 404874 599092
rect 404930 599036 404998 599092
rect 405054 599036 405122 599092
rect 405178 599036 405246 599092
rect 405302 599036 422874 599092
rect 422930 599036 422998 599092
rect 423054 599036 423122 599092
rect 423178 599036 423246 599092
rect 423302 599036 440874 599092
rect 440930 599036 440998 599092
rect 441054 599036 441122 599092
rect 441178 599036 441246 599092
rect 441302 599036 458874 599092
rect 458930 599036 458998 599092
rect 459054 599036 459122 599092
rect 459178 599036 459246 599092
rect 459302 599036 476874 599092
rect 476930 599036 476998 599092
rect 477054 599036 477122 599092
rect 477178 599036 477246 599092
rect 477302 599036 494874 599092
rect 494930 599036 494998 599092
rect 495054 599036 495122 599092
rect 495178 599036 495246 599092
rect 495302 599036 512874 599092
rect 512930 599036 512998 599092
rect 513054 599036 513122 599092
rect 513178 599036 513246 599092
rect 513302 599036 530874 599092
rect 530930 599036 530998 599092
rect 531054 599036 531122 599092
rect 531178 599036 531246 599092
rect 531302 599036 548874 599092
rect 548930 599036 548998 599092
rect 549054 599036 549122 599092
rect 549178 599036 549246 599092
rect 549302 599036 566874 599092
rect 566930 599036 566998 599092
rect 567054 599036 567122 599092
rect 567178 599036 567246 599092
rect 567302 599036 584874 599092
rect 584930 599036 584998 599092
rect 585054 599036 585122 599092
rect 585178 599036 585246 599092
rect 585302 599036 599472 599092
rect 599528 599036 599596 599092
rect 599652 599036 599720 599092
rect 599776 599036 599844 599092
rect 599900 599036 599996 599092
rect -12 598968 599996 599036
rect -12 598912 84 598968
rect 140 598912 208 598968
rect 264 598912 332 598968
rect 388 598912 456 598968
rect 512 598912 8874 598968
rect 8930 598912 8998 598968
rect 9054 598912 9122 598968
rect 9178 598912 9246 598968
rect 9302 598912 26874 598968
rect 26930 598912 26998 598968
rect 27054 598912 27122 598968
rect 27178 598912 27246 598968
rect 27302 598912 44874 598968
rect 44930 598912 44998 598968
rect 45054 598912 45122 598968
rect 45178 598912 45246 598968
rect 45302 598912 62874 598968
rect 62930 598912 62998 598968
rect 63054 598912 63122 598968
rect 63178 598912 63246 598968
rect 63302 598912 80874 598968
rect 80930 598912 80998 598968
rect 81054 598912 81122 598968
rect 81178 598912 81246 598968
rect 81302 598912 98874 598968
rect 98930 598912 98998 598968
rect 99054 598912 99122 598968
rect 99178 598912 99246 598968
rect 99302 598912 116874 598968
rect 116930 598912 116998 598968
rect 117054 598912 117122 598968
rect 117178 598912 117246 598968
rect 117302 598912 134874 598968
rect 134930 598912 134998 598968
rect 135054 598912 135122 598968
rect 135178 598912 135246 598968
rect 135302 598912 152874 598968
rect 152930 598912 152998 598968
rect 153054 598912 153122 598968
rect 153178 598912 153246 598968
rect 153302 598912 170874 598968
rect 170930 598912 170998 598968
rect 171054 598912 171122 598968
rect 171178 598912 171246 598968
rect 171302 598912 188874 598968
rect 188930 598912 188998 598968
rect 189054 598912 189122 598968
rect 189178 598912 189246 598968
rect 189302 598912 206874 598968
rect 206930 598912 206998 598968
rect 207054 598912 207122 598968
rect 207178 598912 207246 598968
rect 207302 598912 224874 598968
rect 224930 598912 224998 598968
rect 225054 598912 225122 598968
rect 225178 598912 225246 598968
rect 225302 598912 242874 598968
rect 242930 598912 242998 598968
rect 243054 598912 243122 598968
rect 243178 598912 243246 598968
rect 243302 598912 260874 598968
rect 260930 598912 260998 598968
rect 261054 598912 261122 598968
rect 261178 598912 261246 598968
rect 261302 598912 278874 598968
rect 278930 598912 278998 598968
rect 279054 598912 279122 598968
rect 279178 598912 279246 598968
rect 279302 598912 296874 598968
rect 296930 598912 296998 598968
rect 297054 598912 297122 598968
rect 297178 598912 297246 598968
rect 297302 598912 314874 598968
rect 314930 598912 314998 598968
rect 315054 598912 315122 598968
rect 315178 598912 315246 598968
rect 315302 598912 332874 598968
rect 332930 598912 332998 598968
rect 333054 598912 333122 598968
rect 333178 598912 333246 598968
rect 333302 598912 350874 598968
rect 350930 598912 350998 598968
rect 351054 598912 351122 598968
rect 351178 598912 351246 598968
rect 351302 598912 368874 598968
rect 368930 598912 368998 598968
rect 369054 598912 369122 598968
rect 369178 598912 369246 598968
rect 369302 598912 386874 598968
rect 386930 598912 386998 598968
rect 387054 598912 387122 598968
rect 387178 598912 387246 598968
rect 387302 598912 404874 598968
rect 404930 598912 404998 598968
rect 405054 598912 405122 598968
rect 405178 598912 405246 598968
rect 405302 598912 422874 598968
rect 422930 598912 422998 598968
rect 423054 598912 423122 598968
rect 423178 598912 423246 598968
rect 423302 598912 440874 598968
rect 440930 598912 440998 598968
rect 441054 598912 441122 598968
rect 441178 598912 441246 598968
rect 441302 598912 458874 598968
rect 458930 598912 458998 598968
rect 459054 598912 459122 598968
rect 459178 598912 459246 598968
rect 459302 598912 476874 598968
rect 476930 598912 476998 598968
rect 477054 598912 477122 598968
rect 477178 598912 477246 598968
rect 477302 598912 494874 598968
rect 494930 598912 494998 598968
rect 495054 598912 495122 598968
rect 495178 598912 495246 598968
rect 495302 598912 512874 598968
rect 512930 598912 512998 598968
rect 513054 598912 513122 598968
rect 513178 598912 513246 598968
rect 513302 598912 530874 598968
rect 530930 598912 530998 598968
rect 531054 598912 531122 598968
rect 531178 598912 531246 598968
rect 531302 598912 548874 598968
rect 548930 598912 548998 598968
rect 549054 598912 549122 598968
rect 549178 598912 549246 598968
rect 549302 598912 566874 598968
rect 566930 598912 566998 598968
rect 567054 598912 567122 598968
rect 567178 598912 567246 598968
rect 567302 598912 584874 598968
rect 584930 598912 584998 598968
rect 585054 598912 585122 598968
rect 585178 598912 585246 598968
rect 585302 598912 599472 598968
rect 599528 598912 599596 598968
rect 599652 598912 599720 598968
rect 599776 598912 599844 598968
rect 599900 598912 599996 598968
rect -12 598816 599996 598912
rect 948 598380 599036 598476
rect 948 598324 1044 598380
rect 1100 598324 1168 598380
rect 1224 598324 1292 598380
rect 1348 598324 1416 598380
rect 1472 598324 5154 598380
rect 5210 598324 5278 598380
rect 5334 598324 5402 598380
rect 5458 598324 5526 598380
rect 5582 598324 23154 598380
rect 23210 598324 23278 598380
rect 23334 598324 23402 598380
rect 23458 598324 23526 598380
rect 23582 598324 41154 598380
rect 41210 598324 41278 598380
rect 41334 598324 41402 598380
rect 41458 598324 41526 598380
rect 41582 598324 59154 598380
rect 59210 598324 59278 598380
rect 59334 598324 59402 598380
rect 59458 598324 59526 598380
rect 59582 598324 77154 598380
rect 77210 598324 77278 598380
rect 77334 598324 77402 598380
rect 77458 598324 77526 598380
rect 77582 598324 95154 598380
rect 95210 598324 95278 598380
rect 95334 598324 95402 598380
rect 95458 598324 95526 598380
rect 95582 598324 113154 598380
rect 113210 598324 113278 598380
rect 113334 598324 113402 598380
rect 113458 598324 113526 598380
rect 113582 598324 131154 598380
rect 131210 598324 131278 598380
rect 131334 598324 131402 598380
rect 131458 598324 131526 598380
rect 131582 598324 149154 598380
rect 149210 598324 149278 598380
rect 149334 598324 149402 598380
rect 149458 598324 149526 598380
rect 149582 598324 167154 598380
rect 167210 598324 167278 598380
rect 167334 598324 167402 598380
rect 167458 598324 167526 598380
rect 167582 598324 185154 598380
rect 185210 598324 185278 598380
rect 185334 598324 185402 598380
rect 185458 598324 185526 598380
rect 185582 598324 203154 598380
rect 203210 598324 203278 598380
rect 203334 598324 203402 598380
rect 203458 598324 203526 598380
rect 203582 598324 221154 598380
rect 221210 598324 221278 598380
rect 221334 598324 221402 598380
rect 221458 598324 221526 598380
rect 221582 598324 239154 598380
rect 239210 598324 239278 598380
rect 239334 598324 239402 598380
rect 239458 598324 239526 598380
rect 239582 598324 257154 598380
rect 257210 598324 257278 598380
rect 257334 598324 257402 598380
rect 257458 598324 257526 598380
rect 257582 598324 275154 598380
rect 275210 598324 275278 598380
rect 275334 598324 275402 598380
rect 275458 598324 275526 598380
rect 275582 598324 293154 598380
rect 293210 598324 293278 598380
rect 293334 598324 293402 598380
rect 293458 598324 293526 598380
rect 293582 598324 311154 598380
rect 311210 598324 311278 598380
rect 311334 598324 311402 598380
rect 311458 598324 311526 598380
rect 311582 598324 329154 598380
rect 329210 598324 329278 598380
rect 329334 598324 329402 598380
rect 329458 598324 329526 598380
rect 329582 598324 347154 598380
rect 347210 598324 347278 598380
rect 347334 598324 347402 598380
rect 347458 598324 347526 598380
rect 347582 598324 365154 598380
rect 365210 598324 365278 598380
rect 365334 598324 365402 598380
rect 365458 598324 365526 598380
rect 365582 598324 383154 598380
rect 383210 598324 383278 598380
rect 383334 598324 383402 598380
rect 383458 598324 383526 598380
rect 383582 598324 401154 598380
rect 401210 598324 401278 598380
rect 401334 598324 401402 598380
rect 401458 598324 401526 598380
rect 401582 598324 419154 598380
rect 419210 598324 419278 598380
rect 419334 598324 419402 598380
rect 419458 598324 419526 598380
rect 419582 598324 437154 598380
rect 437210 598324 437278 598380
rect 437334 598324 437402 598380
rect 437458 598324 437526 598380
rect 437582 598324 455154 598380
rect 455210 598324 455278 598380
rect 455334 598324 455402 598380
rect 455458 598324 455526 598380
rect 455582 598324 473154 598380
rect 473210 598324 473278 598380
rect 473334 598324 473402 598380
rect 473458 598324 473526 598380
rect 473582 598324 491154 598380
rect 491210 598324 491278 598380
rect 491334 598324 491402 598380
rect 491458 598324 491526 598380
rect 491582 598324 509154 598380
rect 509210 598324 509278 598380
rect 509334 598324 509402 598380
rect 509458 598324 509526 598380
rect 509582 598324 527154 598380
rect 527210 598324 527278 598380
rect 527334 598324 527402 598380
rect 527458 598324 527526 598380
rect 527582 598324 545154 598380
rect 545210 598324 545278 598380
rect 545334 598324 545402 598380
rect 545458 598324 545526 598380
rect 545582 598324 563154 598380
rect 563210 598324 563278 598380
rect 563334 598324 563402 598380
rect 563458 598324 563526 598380
rect 563582 598324 581154 598380
rect 581210 598324 581278 598380
rect 581334 598324 581402 598380
rect 581458 598324 581526 598380
rect 581582 598324 598512 598380
rect 598568 598324 598636 598380
rect 598692 598324 598760 598380
rect 598816 598324 598884 598380
rect 598940 598324 599036 598380
rect 948 598256 599036 598324
rect 948 598200 1044 598256
rect 1100 598200 1168 598256
rect 1224 598200 1292 598256
rect 1348 598200 1416 598256
rect 1472 598200 5154 598256
rect 5210 598200 5278 598256
rect 5334 598200 5402 598256
rect 5458 598200 5526 598256
rect 5582 598200 23154 598256
rect 23210 598200 23278 598256
rect 23334 598200 23402 598256
rect 23458 598200 23526 598256
rect 23582 598200 41154 598256
rect 41210 598200 41278 598256
rect 41334 598200 41402 598256
rect 41458 598200 41526 598256
rect 41582 598200 59154 598256
rect 59210 598200 59278 598256
rect 59334 598200 59402 598256
rect 59458 598200 59526 598256
rect 59582 598200 77154 598256
rect 77210 598200 77278 598256
rect 77334 598200 77402 598256
rect 77458 598200 77526 598256
rect 77582 598200 95154 598256
rect 95210 598200 95278 598256
rect 95334 598200 95402 598256
rect 95458 598200 95526 598256
rect 95582 598200 113154 598256
rect 113210 598200 113278 598256
rect 113334 598200 113402 598256
rect 113458 598200 113526 598256
rect 113582 598200 131154 598256
rect 131210 598200 131278 598256
rect 131334 598200 131402 598256
rect 131458 598200 131526 598256
rect 131582 598200 149154 598256
rect 149210 598200 149278 598256
rect 149334 598200 149402 598256
rect 149458 598200 149526 598256
rect 149582 598200 167154 598256
rect 167210 598200 167278 598256
rect 167334 598200 167402 598256
rect 167458 598200 167526 598256
rect 167582 598200 185154 598256
rect 185210 598200 185278 598256
rect 185334 598200 185402 598256
rect 185458 598200 185526 598256
rect 185582 598200 203154 598256
rect 203210 598200 203278 598256
rect 203334 598200 203402 598256
rect 203458 598200 203526 598256
rect 203582 598200 221154 598256
rect 221210 598200 221278 598256
rect 221334 598200 221402 598256
rect 221458 598200 221526 598256
rect 221582 598200 239154 598256
rect 239210 598200 239278 598256
rect 239334 598200 239402 598256
rect 239458 598200 239526 598256
rect 239582 598200 257154 598256
rect 257210 598200 257278 598256
rect 257334 598200 257402 598256
rect 257458 598200 257526 598256
rect 257582 598200 275154 598256
rect 275210 598200 275278 598256
rect 275334 598200 275402 598256
rect 275458 598200 275526 598256
rect 275582 598200 293154 598256
rect 293210 598200 293278 598256
rect 293334 598200 293402 598256
rect 293458 598200 293526 598256
rect 293582 598200 311154 598256
rect 311210 598200 311278 598256
rect 311334 598200 311402 598256
rect 311458 598200 311526 598256
rect 311582 598200 329154 598256
rect 329210 598200 329278 598256
rect 329334 598200 329402 598256
rect 329458 598200 329526 598256
rect 329582 598200 347154 598256
rect 347210 598200 347278 598256
rect 347334 598200 347402 598256
rect 347458 598200 347526 598256
rect 347582 598200 365154 598256
rect 365210 598200 365278 598256
rect 365334 598200 365402 598256
rect 365458 598200 365526 598256
rect 365582 598200 383154 598256
rect 383210 598200 383278 598256
rect 383334 598200 383402 598256
rect 383458 598200 383526 598256
rect 383582 598200 401154 598256
rect 401210 598200 401278 598256
rect 401334 598200 401402 598256
rect 401458 598200 401526 598256
rect 401582 598200 419154 598256
rect 419210 598200 419278 598256
rect 419334 598200 419402 598256
rect 419458 598200 419526 598256
rect 419582 598200 437154 598256
rect 437210 598200 437278 598256
rect 437334 598200 437402 598256
rect 437458 598200 437526 598256
rect 437582 598200 455154 598256
rect 455210 598200 455278 598256
rect 455334 598200 455402 598256
rect 455458 598200 455526 598256
rect 455582 598200 473154 598256
rect 473210 598200 473278 598256
rect 473334 598200 473402 598256
rect 473458 598200 473526 598256
rect 473582 598200 491154 598256
rect 491210 598200 491278 598256
rect 491334 598200 491402 598256
rect 491458 598200 491526 598256
rect 491582 598200 509154 598256
rect 509210 598200 509278 598256
rect 509334 598200 509402 598256
rect 509458 598200 509526 598256
rect 509582 598200 527154 598256
rect 527210 598200 527278 598256
rect 527334 598200 527402 598256
rect 527458 598200 527526 598256
rect 527582 598200 545154 598256
rect 545210 598200 545278 598256
rect 545334 598200 545402 598256
rect 545458 598200 545526 598256
rect 545582 598200 563154 598256
rect 563210 598200 563278 598256
rect 563334 598200 563402 598256
rect 563458 598200 563526 598256
rect 563582 598200 581154 598256
rect 581210 598200 581278 598256
rect 581334 598200 581402 598256
rect 581458 598200 581526 598256
rect 581582 598200 598512 598256
rect 598568 598200 598636 598256
rect 598692 598200 598760 598256
rect 598816 598200 598884 598256
rect 598940 598200 599036 598256
rect 948 598132 599036 598200
rect 948 598076 1044 598132
rect 1100 598076 1168 598132
rect 1224 598076 1292 598132
rect 1348 598076 1416 598132
rect 1472 598076 5154 598132
rect 5210 598076 5278 598132
rect 5334 598076 5402 598132
rect 5458 598076 5526 598132
rect 5582 598076 23154 598132
rect 23210 598076 23278 598132
rect 23334 598076 23402 598132
rect 23458 598076 23526 598132
rect 23582 598076 41154 598132
rect 41210 598076 41278 598132
rect 41334 598076 41402 598132
rect 41458 598076 41526 598132
rect 41582 598076 59154 598132
rect 59210 598076 59278 598132
rect 59334 598076 59402 598132
rect 59458 598076 59526 598132
rect 59582 598076 77154 598132
rect 77210 598076 77278 598132
rect 77334 598076 77402 598132
rect 77458 598076 77526 598132
rect 77582 598076 95154 598132
rect 95210 598076 95278 598132
rect 95334 598076 95402 598132
rect 95458 598076 95526 598132
rect 95582 598076 113154 598132
rect 113210 598076 113278 598132
rect 113334 598076 113402 598132
rect 113458 598076 113526 598132
rect 113582 598076 131154 598132
rect 131210 598076 131278 598132
rect 131334 598076 131402 598132
rect 131458 598076 131526 598132
rect 131582 598076 149154 598132
rect 149210 598076 149278 598132
rect 149334 598076 149402 598132
rect 149458 598076 149526 598132
rect 149582 598076 167154 598132
rect 167210 598076 167278 598132
rect 167334 598076 167402 598132
rect 167458 598076 167526 598132
rect 167582 598076 185154 598132
rect 185210 598076 185278 598132
rect 185334 598076 185402 598132
rect 185458 598076 185526 598132
rect 185582 598076 203154 598132
rect 203210 598076 203278 598132
rect 203334 598076 203402 598132
rect 203458 598076 203526 598132
rect 203582 598076 221154 598132
rect 221210 598076 221278 598132
rect 221334 598076 221402 598132
rect 221458 598076 221526 598132
rect 221582 598076 239154 598132
rect 239210 598076 239278 598132
rect 239334 598076 239402 598132
rect 239458 598076 239526 598132
rect 239582 598076 257154 598132
rect 257210 598076 257278 598132
rect 257334 598076 257402 598132
rect 257458 598076 257526 598132
rect 257582 598076 275154 598132
rect 275210 598076 275278 598132
rect 275334 598076 275402 598132
rect 275458 598076 275526 598132
rect 275582 598076 293154 598132
rect 293210 598076 293278 598132
rect 293334 598076 293402 598132
rect 293458 598076 293526 598132
rect 293582 598076 311154 598132
rect 311210 598076 311278 598132
rect 311334 598076 311402 598132
rect 311458 598076 311526 598132
rect 311582 598076 329154 598132
rect 329210 598076 329278 598132
rect 329334 598076 329402 598132
rect 329458 598076 329526 598132
rect 329582 598076 347154 598132
rect 347210 598076 347278 598132
rect 347334 598076 347402 598132
rect 347458 598076 347526 598132
rect 347582 598076 365154 598132
rect 365210 598076 365278 598132
rect 365334 598076 365402 598132
rect 365458 598076 365526 598132
rect 365582 598076 383154 598132
rect 383210 598076 383278 598132
rect 383334 598076 383402 598132
rect 383458 598076 383526 598132
rect 383582 598076 401154 598132
rect 401210 598076 401278 598132
rect 401334 598076 401402 598132
rect 401458 598076 401526 598132
rect 401582 598076 419154 598132
rect 419210 598076 419278 598132
rect 419334 598076 419402 598132
rect 419458 598076 419526 598132
rect 419582 598076 437154 598132
rect 437210 598076 437278 598132
rect 437334 598076 437402 598132
rect 437458 598076 437526 598132
rect 437582 598076 455154 598132
rect 455210 598076 455278 598132
rect 455334 598076 455402 598132
rect 455458 598076 455526 598132
rect 455582 598076 473154 598132
rect 473210 598076 473278 598132
rect 473334 598076 473402 598132
rect 473458 598076 473526 598132
rect 473582 598076 491154 598132
rect 491210 598076 491278 598132
rect 491334 598076 491402 598132
rect 491458 598076 491526 598132
rect 491582 598076 509154 598132
rect 509210 598076 509278 598132
rect 509334 598076 509402 598132
rect 509458 598076 509526 598132
rect 509582 598076 527154 598132
rect 527210 598076 527278 598132
rect 527334 598076 527402 598132
rect 527458 598076 527526 598132
rect 527582 598076 545154 598132
rect 545210 598076 545278 598132
rect 545334 598076 545402 598132
rect 545458 598076 545526 598132
rect 545582 598076 563154 598132
rect 563210 598076 563278 598132
rect 563334 598076 563402 598132
rect 563458 598076 563526 598132
rect 563582 598076 581154 598132
rect 581210 598076 581278 598132
rect 581334 598076 581402 598132
rect 581458 598076 581526 598132
rect 581582 598076 598512 598132
rect 598568 598076 598636 598132
rect 598692 598076 598760 598132
rect 598816 598076 598884 598132
rect 598940 598076 599036 598132
rect 948 598008 599036 598076
rect 948 597952 1044 598008
rect 1100 597952 1168 598008
rect 1224 597952 1292 598008
rect 1348 597952 1416 598008
rect 1472 597952 5154 598008
rect 5210 597952 5278 598008
rect 5334 597952 5402 598008
rect 5458 597952 5526 598008
rect 5582 597952 23154 598008
rect 23210 597952 23278 598008
rect 23334 597952 23402 598008
rect 23458 597952 23526 598008
rect 23582 597952 41154 598008
rect 41210 597952 41278 598008
rect 41334 597952 41402 598008
rect 41458 597952 41526 598008
rect 41582 597952 59154 598008
rect 59210 597952 59278 598008
rect 59334 597952 59402 598008
rect 59458 597952 59526 598008
rect 59582 597952 77154 598008
rect 77210 597952 77278 598008
rect 77334 597952 77402 598008
rect 77458 597952 77526 598008
rect 77582 597952 95154 598008
rect 95210 597952 95278 598008
rect 95334 597952 95402 598008
rect 95458 597952 95526 598008
rect 95582 597952 113154 598008
rect 113210 597952 113278 598008
rect 113334 597952 113402 598008
rect 113458 597952 113526 598008
rect 113582 597952 131154 598008
rect 131210 597952 131278 598008
rect 131334 597952 131402 598008
rect 131458 597952 131526 598008
rect 131582 597952 149154 598008
rect 149210 597952 149278 598008
rect 149334 597952 149402 598008
rect 149458 597952 149526 598008
rect 149582 597952 167154 598008
rect 167210 597952 167278 598008
rect 167334 597952 167402 598008
rect 167458 597952 167526 598008
rect 167582 597952 185154 598008
rect 185210 597952 185278 598008
rect 185334 597952 185402 598008
rect 185458 597952 185526 598008
rect 185582 597952 203154 598008
rect 203210 597952 203278 598008
rect 203334 597952 203402 598008
rect 203458 597952 203526 598008
rect 203582 597952 221154 598008
rect 221210 597952 221278 598008
rect 221334 597952 221402 598008
rect 221458 597952 221526 598008
rect 221582 597952 239154 598008
rect 239210 597952 239278 598008
rect 239334 597952 239402 598008
rect 239458 597952 239526 598008
rect 239582 597952 257154 598008
rect 257210 597952 257278 598008
rect 257334 597952 257402 598008
rect 257458 597952 257526 598008
rect 257582 597952 275154 598008
rect 275210 597952 275278 598008
rect 275334 597952 275402 598008
rect 275458 597952 275526 598008
rect 275582 597952 293154 598008
rect 293210 597952 293278 598008
rect 293334 597952 293402 598008
rect 293458 597952 293526 598008
rect 293582 597952 311154 598008
rect 311210 597952 311278 598008
rect 311334 597952 311402 598008
rect 311458 597952 311526 598008
rect 311582 597952 329154 598008
rect 329210 597952 329278 598008
rect 329334 597952 329402 598008
rect 329458 597952 329526 598008
rect 329582 597952 347154 598008
rect 347210 597952 347278 598008
rect 347334 597952 347402 598008
rect 347458 597952 347526 598008
rect 347582 597952 365154 598008
rect 365210 597952 365278 598008
rect 365334 597952 365402 598008
rect 365458 597952 365526 598008
rect 365582 597952 383154 598008
rect 383210 597952 383278 598008
rect 383334 597952 383402 598008
rect 383458 597952 383526 598008
rect 383582 597952 401154 598008
rect 401210 597952 401278 598008
rect 401334 597952 401402 598008
rect 401458 597952 401526 598008
rect 401582 597952 419154 598008
rect 419210 597952 419278 598008
rect 419334 597952 419402 598008
rect 419458 597952 419526 598008
rect 419582 597952 437154 598008
rect 437210 597952 437278 598008
rect 437334 597952 437402 598008
rect 437458 597952 437526 598008
rect 437582 597952 455154 598008
rect 455210 597952 455278 598008
rect 455334 597952 455402 598008
rect 455458 597952 455526 598008
rect 455582 597952 473154 598008
rect 473210 597952 473278 598008
rect 473334 597952 473402 598008
rect 473458 597952 473526 598008
rect 473582 597952 491154 598008
rect 491210 597952 491278 598008
rect 491334 597952 491402 598008
rect 491458 597952 491526 598008
rect 491582 597952 509154 598008
rect 509210 597952 509278 598008
rect 509334 597952 509402 598008
rect 509458 597952 509526 598008
rect 509582 597952 527154 598008
rect 527210 597952 527278 598008
rect 527334 597952 527402 598008
rect 527458 597952 527526 598008
rect 527582 597952 545154 598008
rect 545210 597952 545278 598008
rect 545334 597952 545402 598008
rect 545458 597952 545526 598008
rect 545582 597952 563154 598008
rect 563210 597952 563278 598008
rect 563334 597952 563402 598008
rect 563458 597952 563526 598008
rect 563582 597952 581154 598008
rect 581210 597952 581278 598008
rect 581334 597952 581402 598008
rect 581458 597952 581526 598008
rect 581582 597952 598512 598008
rect 598568 597952 598636 598008
rect 598692 597952 598760 598008
rect 598816 597952 598884 598008
rect 598940 597952 599036 598008
rect 948 597856 599036 597952
rect -12 587918 6134 588014
rect -12 587862 84 587918
rect 140 587862 208 587918
rect 264 587862 332 587918
rect 388 587862 456 587918
rect 512 587862 6134 587918
rect -12 587794 6134 587862
rect -12 587738 84 587794
rect 140 587738 208 587794
rect 264 587738 332 587794
rect 388 587738 456 587794
rect 512 587738 6134 587794
rect -12 587670 6134 587738
rect -12 587614 84 587670
rect 140 587614 208 587670
rect 264 587614 332 587670
rect 388 587614 456 587670
rect 512 587614 6134 587670
rect -12 587546 6134 587614
rect -12 587490 84 587546
rect 140 587490 208 587546
rect 264 587490 332 587546
rect 388 587490 456 587546
rect 512 587490 6134 587546
rect -12 587394 6134 587490
rect 595211 587918 599996 588014
rect 595211 587862 599472 587918
rect 599528 587862 599596 587918
rect 599652 587862 599720 587918
rect 599776 587862 599844 587918
rect 599900 587862 599996 587918
rect 595211 587794 599996 587862
rect 595211 587738 599472 587794
rect 599528 587738 599596 587794
rect 599652 587738 599720 587794
rect 599776 587738 599844 587794
rect 599900 587738 599996 587794
rect 595211 587670 599996 587738
rect 595211 587614 599472 587670
rect 599528 587614 599596 587670
rect 599652 587614 599720 587670
rect 599776 587614 599844 587670
rect 599900 587614 599996 587670
rect 595211 587546 599996 587614
rect 595211 587490 599472 587546
rect 599528 587490 599596 587546
rect 599652 587490 599720 587546
rect 599776 587490 599844 587546
rect 599900 587490 599996 587546
rect 595211 587394 599996 587490
rect -12 581918 6134 582014
rect -12 581862 1044 581918
rect 1100 581862 1168 581918
rect 1224 581862 1292 581918
rect 1348 581862 1416 581918
rect 1472 581862 5154 581918
rect 5210 581862 5278 581918
rect 5334 581862 5402 581918
rect 5458 581862 5526 581918
rect 5582 581862 6134 581918
rect -12 581794 6134 581862
rect -12 581738 1044 581794
rect 1100 581738 1168 581794
rect 1224 581738 1292 581794
rect 1348 581738 1416 581794
rect 1472 581738 5154 581794
rect 5210 581738 5278 581794
rect 5334 581738 5402 581794
rect 5458 581738 5526 581794
rect 5582 581738 6134 581794
rect -12 581670 6134 581738
rect -12 581614 1044 581670
rect 1100 581614 1168 581670
rect 1224 581614 1292 581670
rect 1348 581614 1416 581670
rect 1472 581614 5154 581670
rect 5210 581614 5278 581670
rect 5334 581614 5402 581670
rect 5458 581614 5526 581670
rect 5582 581614 6134 581670
rect -12 581546 6134 581614
rect -12 581490 1044 581546
rect 1100 581490 1168 581546
rect 1224 581490 1292 581546
rect 1348 581490 1416 581546
rect 1472 581490 5154 581546
rect 5210 581490 5278 581546
rect 5334 581490 5402 581546
rect 5458 581490 5526 581546
rect 5582 581490 6134 581546
rect -12 581394 6134 581490
rect 595211 581918 599996 582014
rect 595211 581862 598512 581918
rect 598568 581862 598636 581918
rect 598692 581862 598760 581918
rect 598816 581862 598884 581918
rect 598940 581862 599996 581918
rect 595211 581794 599996 581862
rect 595211 581738 598512 581794
rect 598568 581738 598636 581794
rect 598692 581738 598760 581794
rect 598816 581738 598884 581794
rect 598940 581738 599996 581794
rect 595211 581670 599996 581738
rect 595211 581614 598512 581670
rect 598568 581614 598636 581670
rect 598692 581614 598760 581670
rect 598816 581614 598884 581670
rect 598940 581614 599996 581670
rect 595211 581546 599996 581614
rect 595211 581490 598512 581546
rect 598568 581490 598636 581546
rect 598692 581490 598760 581546
rect 598816 581490 598884 581546
rect 598940 581490 599996 581546
rect 595211 581394 599996 581490
rect -12 569918 6134 570014
rect -12 569862 84 569918
rect 140 569862 208 569918
rect 264 569862 332 569918
rect 388 569862 456 569918
rect 512 569862 6134 569918
rect -12 569794 6134 569862
rect -12 569738 84 569794
rect 140 569738 208 569794
rect 264 569738 332 569794
rect 388 569738 456 569794
rect 512 569738 6134 569794
rect -12 569670 6134 569738
rect -12 569614 84 569670
rect 140 569614 208 569670
rect 264 569614 332 569670
rect 388 569614 456 569670
rect 512 569614 6134 569670
rect -12 569546 6134 569614
rect -12 569490 84 569546
rect 140 569490 208 569546
rect 264 569490 332 569546
rect 388 569490 456 569546
rect 512 569490 6134 569546
rect -12 569394 6134 569490
rect 595211 569918 599996 570014
rect 595211 569862 599472 569918
rect 599528 569862 599596 569918
rect 599652 569862 599720 569918
rect 599776 569862 599844 569918
rect 599900 569862 599996 569918
rect 595211 569794 599996 569862
rect 595211 569738 599472 569794
rect 599528 569738 599596 569794
rect 599652 569738 599720 569794
rect 599776 569738 599844 569794
rect 599900 569738 599996 569794
rect 595211 569670 599996 569738
rect 595211 569614 599472 569670
rect 599528 569614 599596 569670
rect 599652 569614 599720 569670
rect 599776 569614 599844 569670
rect 599900 569614 599996 569670
rect 595211 569546 599996 569614
rect 595211 569490 599472 569546
rect 599528 569490 599596 569546
rect 599652 569490 599720 569546
rect 599776 569490 599844 569546
rect 599900 569490 599996 569546
rect 595211 569394 599996 569490
rect -12 563918 6134 564014
rect -12 563862 1044 563918
rect 1100 563862 1168 563918
rect 1224 563862 1292 563918
rect 1348 563862 1416 563918
rect 1472 563862 5154 563918
rect 5210 563862 5278 563918
rect 5334 563862 5402 563918
rect 5458 563862 5526 563918
rect 5582 563862 6134 563918
rect -12 563794 6134 563862
rect -12 563738 1044 563794
rect 1100 563738 1168 563794
rect 1224 563738 1292 563794
rect 1348 563738 1416 563794
rect 1472 563738 5154 563794
rect 5210 563738 5278 563794
rect 5334 563738 5402 563794
rect 5458 563738 5526 563794
rect 5582 563738 6134 563794
rect -12 563670 6134 563738
rect -12 563614 1044 563670
rect 1100 563614 1168 563670
rect 1224 563614 1292 563670
rect 1348 563614 1416 563670
rect 1472 563614 5154 563670
rect 5210 563614 5278 563670
rect 5334 563614 5402 563670
rect 5458 563614 5526 563670
rect 5582 563614 6134 563670
rect -12 563546 6134 563614
rect -12 563490 1044 563546
rect 1100 563490 1168 563546
rect 1224 563490 1292 563546
rect 1348 563490 1416 563546
rect 1472 563490 5154 563546
rect 5210 563490 5278 563546
rect 5334 563490 5402 563546
rect 5458 563490 5526 563546
rect 5582 563490 6134 563546
rect -12 563394 6134 563490
rect 595211 563918 599996 564014
rect 595211 563862 598512 563918
rect 598568 563862 598636 563918
rect 598692 563862 598760 563918
rect 598816 563862 598884 563918
rect 598940 563862 599996 563918
rect 595211 563794 599996 563862
rect 595211 563738 598512 563794
rect 598568 563738 598636 563794
rect 598692 563738 598760 563794
rect 598816 563738 598884 563794
rect 598940 563738 599996 563794
rect 595211 563670 599996 563738
rect 595211 563614 598512 563670
rect 598568 563614 598636 563670
rect 598692 563614 598760 563670
rect 598816 563614 598884 563670
rect 598940 563614 599996 563670
rect 595211 563546 599996 563614
rect 595211 563490 598512 563546
rect 598568 563490 598636 563546
rect 598692 563490 598760 563546
rect 598816 563490 598884 563546
rect 598940 563490 599996 563546
rect 595211 563394 599996 563490
rect -12 551918 6134 552014
rect -12 551862 84 551918
rect 140 551862 208 551918
rect 264 551862 332 551918
rect 388 551862 456 551918
rect 512 551862 6134 551918
rect -12 551794 6134 551862
rect -12 551738 84 551794
rect 140 551738 208 551794
rect 264 551738 332 551794
rect 388 551738 456 551794
rect 512 551738 6134 551794
rect -12 551670 6134 551738
rect -12 551614 84 551670
rect 140 551614 208 551670
rect 264 551614 332 551670
rect 388 551614 456 551670
rect 512 551614 6134 551670
rect -12 551546 6134 551614
rect -12 551490 84 551546
rect 140 551490 208 551546
rect 264 551490 332 551546
rect 388 551490 456 551546
rect 512 551490 6134 551546
rect -12 551394 6134 551490
rect 595211 551918 599996 552014
rect 595211 551862 599472 551918
rect 599528 551862 599596 551918
rect 599652 551862 599720 551918
rect 599776 551862 599844 551918
rect 599900 551862 599996 551918
rect 595211 551794 599996 551862
rect 595211 551738 599472 551794
rect 599528 551738 599596 551794
rect 599652 551738 599720 551794
rect 599776 551738 599844 551794
rect 599900 551738 599996 551794
rect 595211 551670 599996 551738
rect 595211 551614 599472 551670
rect 599528 551614 599596 551670
rect 599652 551614 599720 551670
rect 599776 551614 599844 551670
rect 599900 551614 599996 551670
rect 595211 551546 599996 551614
rect 595211 551490 599472 551546
rect 599528 551490 599596 551546
rect 599652 551490 599720 551546
rect 599776 551490 599844 551546
rect 599900 551490 599996 551546
rect 595211 551394 599996 551490
rect -12 545918 6134 546014
rect -12 545862 1044 545918
rect 1100 545862 1168 545918
rect 1224 545862 1292 545918
rect 1348 545862 1416 545918
rect 1472 545862 5154 545918
rect 5210 545862 5278 545918
rect 5334 545862 5402 545918
rect 5458 545862 5526 545918
rect 5582 545862 6134 545918
rect -12 545794 6134 545862
rect -12 545738 1044 545794
rect 1100 545738 1168 545794
rect 1224 545738 1292 545794
rect 1348 545738 1416 545794
rect 1472 545738 5154 545794
rect 5210 545738 5278 545794
rect 5334 545738 5402 545794
rect 5458 545738 5526 545794
rect 5582 545738 6134 545794
rect -12 545670 6134 545738
rect -12 545614 1044 545670
rect 1100 545614 1168 545670
rect 1224 545614 1292 545670
rect 1348 545614 1416 545670
rect 1472 545614 5154 545670
rect 5210 545614 5278 545670
rect 5334 545614 5402 545670
rect 5458 545614 5526 545670
rect 5582 545614 6134 545670
rect -12 545546 6134 545614
rect -12 545490 1044 545546
rect 1100 545490 1168 545546
rect 1224 545490 1292 545546
rect 1348 545490 1416 545546
rect 1472 545490 5154 545546
rect 5210 545490 5278 545546
rect 5334 545490 5402 545546
rect 5458 545490 5526 545546
rect 5582 545490 6134 545546
rect -12 545394 6134 545490
rect 595211 545918 599996 546014
rect 595211 545862 598512 545918
rect 598568 545862 598636 545918
rect 598692 545862 598760 545918
rect 598816 545862 598884 545918
rect 598940 545862 599996 545918
rect 595211 545794 599996 545862
rect 595211 545738 598512 545794
rect 598568 545738 598636 545794
rect 598692 545738 598760 545794
rect 598816 545738 598884 545794
rect 598940 545738 599996 545794
rect 595211 545670 599996 545738
rect 595211 545614 598512 545670
rect 598568 545614 598636 545670
rect 598692 545614 598760 545670
rect 598816 545614 598884 545670
rect 598940 545614 599996 545670
rect 595211 545546 599996 545614
rect 595211 545490 598512 545546
rect 598568 545490 598636 545546
rect 598692 545490 598760 545546
rect 598816 545490 598884 545546
rect 598940 545490 599996 545546
rect 595211 545394 599996 545490
rect -12 533918 6134 534014
rect -12 533862 84 533918
rect 140 533862 208 533918
rect 264 533862 332 533918
rect 388 533862 456 533918
rect 512 533862 6134 533918
rect -12 533794 6134 533862
rect -12 533738 84 533794
rect 140 533738 208 533794
rect 264 533738 332 533794
rect 388 533738 456 533794
rect 512 533738 6134 533794
rect -12 533670 6134 533738
rect -12 533614 84 533670
rect 140 533614 208 533670
rect 264 533614 332 533670
rect 388 533614 456 533670
rect 512 533614 6134 533670
rect -12 533546 6134 533614
rect -12 533490 84 533546
rect 140 533490 208 533546
rect 264 533490 332 533546
rect 388 533490 456 533546
rect 512 533490 6134 533546
rect -12 533394 6134 533490
rect 595211 533918 599996 534014
rect 595211 533862 599472 533918
rect 599528 533862 599596 533918
rect 599652 533862 599720 533918
rect 599776 533862 599844 533918
rect 599900 533862 599996 533918
rect 595211 533794 599996 533862
rect 595211 533738 599472 533794
rect 599528 533738 599596 533794
rect 599652 533738 599720 533794
rect 599776 533738 599844 533794
rect 599900 533738 599996 533794
rect 595211 533670 599996 533738
rect 595211 533614 599472 533670
rect 599528 533614 599596 533670
rect 599652 533614 599720 533670
rect 599776 533614 599844 533670
rect 599900 533614 599996 533670
rect 595211 533546 599996 533614
rect 595211 533490 599472 533546
rect 599528 533490 599596 533546
rect 599652 533490 599720 533546
rect 599776 533490 599844 533546
rect 599900 533490 599996 533546
rect 595211 533394 599996 533490
rect -12 527918 6134 528014
rect -12 527862 1044 527918
rect 1100 527862 1168 527918
rect 1224 527862 1292 527918
rect 1348 527862 1416 527918
rect 1472 527862 5154 527918
rect 5210 527862 5278 527918
rect 5334 527862 5402 527918
rect 5458 527862 5526 527918
rect 5582 527862 6134 527918
rect -12 527794 6134 527862
rect -12 527738 1044 527794
rect 1100 527738 1168 527794
rect 1224 527738 1292 527794
rect 1348 527738 1416 527794
rect 1472 527738 5154 527794
rect 5210 527738 5278 527794
rect 5334 527738 5402 527794
rect 5458 527738 5526 527794
rect 5582 527738 6134 527794
rect -12 527670 6134 527738
rect -12 527614 1044 527670
rect 1100 527614 1168 527670
rect 1224 527614 1292 527670
rect 1348 527614 1416 527670
rect 1472 527614 5154 527670
rect 5210 527614 5278 527670
rect 5334 527614 5402 527670
rect 5458 527614 5526 527670
rect 5582 527614 6134 527670
rect -12 527546 6134 527614
rect -12 527490 1044 527546
rect 1100 527490 1168 527546
rect 1224 527490 1292 527546
rect 1348 527490 1416 527546
rect 1472 527490 5154 527546
rect 5210 527490 5278 527546
rect 5334 527490 5402 527546
rect 5458 527490 5526 527546
rect 5582 527490 6134 527546
rect -12 527394 6134 527490
rect 595211 527918 599996 528014
rect 595211 527862 598512 527918
rect 598568 527862 598636 527918
rect 598692 527862 598760 527918
rect 598816 527862 598884 527918
rect 598940 527862 599996 527918
rect 595211 527794 599996 527862
rect 595211 527738 598512 527794
rect 598568 527738 598636 527794
rect 598692 527738 598760 527794
rect 598816 527738 598884 527794
rect 598940 527738 599996 527794
rect 595211 527670 599996 527738
rect 595211 527614 598512 527670
rect 598568 527614 598636 527670
rect 598692 527614 598760 527670
rect 598816 527614 598884 527670
rect 598940 527614 599996 527670
rect 595211 527546 599996 527614
rect 595211 527490 598512 527546
rect 598568 527490 598636 527546
rect 598692 527490 598760 527546
rect 598816 527490 598884 527546
rect 598940 527490 599996 527546
rect 595211 527394 599996 527490
rect -12 515918 6134 516014
rect -12 515862 84 515918
rect 140 515862 208 515918
rect 264 515862 332 515918
rect 388 515862 456 515918
rect 512 515862 6134 515918
rect -12 515794 6134 515862
rect -12 515738 84 515794
rect 140 515738 208 515794
rect 264 515738 332 515794
rect 388 515738 456 515794
rect 512 515738 6134 515794
rect -12 515670 6134 515738
rect -12 515614 84 515670
rect 140 515614 208 515670
rect 264 515614 332 515670
rect 388 515614 456 515670
rect 512 515614 6134 515670
rect -12 515546 6134 515614
rect -12 515490 84 515546
rect 140 515490 208 515546
rect 264 515490 332 515546
rect 388 515490 456 515546
rect 512 515490 6134 515546
rect -12 515394 6134 515490
rect 595211 515918 599996 516014
rect 595211 515862 599472 515918
rect 599528 515862 599596 515918
rect 599652 515862 599720 515918
rect 599776 515862 599844 515918
rect 599900 515862 599996 515918
rect 595211 515794 599996 515862
rect 595211 515738 599472 515794
rect 599528 515738 599596 515794
rect 599652 515738 599720 515794
rect 599776 515738 599844 515794
rect 599900 515738 599996 515794
rect 595211 515670 599996 515738
rect 595211 515614 599472 515670
rect 599528 515614 599596 515670
rect 599652 515614 599720 515670
rect 599776 515614 599844 515670
rect 599900 515614 599996 515670
rect 595211 515546 599996 515614
rect 595211 515490 599472 515546
rect 599528 515490 599596 515546
rect 599652 515490 599720 515546
rect 599776 515490 599844 515546
rect 599900 515490 599996 515546
rect 595211 515394 599996 515490
rect -12 509918 6134 510014
rect -12 509862 1044 509918
rect 1100 509862 1168 509918
rect 1224 509862 1292 509918
rect 1348 509862 1416 509918
rect 1472 509862 5154 509918
rect 5210 509862 5278 509918
rect 5334 509862 5402 509918
rect 5458 509862 5526 509918
rect 5582 509862 6134 509918
rect -12 509794 6134 509862
rect -12 509738 1044 509794
rect 1100 509738 1168 509794
rect 1224 509738 1292 509794
rect 1348 509738 1416 509794
rect 1472 509738 5154 509794
rect 5210 509738 5278 509794
rect 5334 509738 5402 509794
rect 5458 509738 5526 509794
rect 5582 509738 6134 509794
rect -12 509670 6134 509738
rect -12 509614 1044 509670
rect 1100 509614 1168 509670
rect 1224 509614 1292 509670
rect 1348 509614 1416 509670
rect 1472 509614 5154 509670
rect 5210 509614 5278 509670
rect 5334 509614 5402 509670
rect 5458 509614 5526 509670
rect 5582 509614 6134 509670
rect -12 509546 6134 509614
rect -12 509490 1044 509546
rect 1100 509490 1168 509546
rect 1224 509490 1292 509546
rect 1348 509490 1416 509546
rect 1472 509490 5154 509546
rect 5210 509490 5278 509546
rect 5334 509490 5402 509546
rect 5458 509490 5526 509546
rect 5582 509490 6134 509546
rect -12 509394 6134 509490
rect 595211 509918 599996 510014
rect 595211 509862 598512 509918
rect 598568 509862 598636 509918
rect 598692 509862 598760 509918
rect 598816 509862 598884 509918
rect 598940 509862 599996 509918
rect 595211 509794 599996 509862
rect 595211 509738 598512 509794
rect 598568 509738 598636 509794
rect 598692 509738 598760 509794
rect 598816 509738 598884 509794
rect 598940 509738 599996 509794
rect 595211 509670 599996 509738
rect 595211 509614 598512 509670
rect 598568 509614 598636 509670
rect 598692 509614 598760 509670
rect 598816 509614 598884 509670
rect 598940 509614 599996 509670
rect 595211 509546 599996 509614
rect 595211 509490 598512 509546
rect 598568 509490 598636 509546
rect 598692 509490 598760 509546
rect 598816 509490 598884 509546
rect 598940 509490 599996 509546
rect 595211 509394 599996 509490
rect -12 497918 6134 498014
rect -12 497862 84 497918
rect 140 497862 208 497918
rect 264 497862 332 497918
rect 388 497862 456 497918
rect 512 497862 6134 497918
rect -12 497794 6134 497862
rect -12 497738 84 497794
rect 140 497738 208 497794
rect 264 497738 332 497794
rect 388 497738 456 497794
rect 512 497738 6134 497794
rect -12 497670 6134 497738
rect -12 497614 84 497670
rect 140 497614 208 497670
rect 264 497614 332 497670
rect 388 497614 456 497670
rect 512 497614 6134 497670
rect -12 497546 6134 497614
rect -12 497490 84 497546
rect 140 497490 208 497546
rect 264 497490 332 497546
rect 388 497490 456 497546
rect 512 497490 6134 497546
rect -12 497394 6134 497490
rect 595211 497918 599996 498014
rect 595211 497862 599472 497918
rect 599528 497862 599596 497918
rect 599652 497862 599720 497918
rect 599776 497862 599844 497918
rect 599900 497862 599996 497918
rect 595211 497794 599996 497862
rect 595211 497738 599472 497794
rect 599528 497738 599596 497794
rect 599652 497738 599720 497794
rect 599776 497738 599844 497794
rect 599900 497738 599996 497794
rect 595211 497670 599996 497738
rect 595211 497614 599472 497670
rect 599528 497614 599596 497670
rect 599652 497614 599720 497670
rect 599776 497614 599844 497670
rect 599900 497614 599996 497670
rect 595211 497546 599996 497614
rect 595211 497490 599472 497546
rect 599528 497490 599596 497546
rect 599652 497490 599720 497546
rect 599776 497490 599844 497546
rect 599900 497490 599996 497546
rect 595211 497394 599996 497490
rect -12 491918 6134 492014
rect -12 491862 1044 491918
rect 1100 491862 1168 491918
rect 1224 491862 1292 491918
rect 1348 491862 1416 491918
rect 1472 491862 5154 491918
rect 5210 491862 5278 491918
rect 5334 491862 5402 491918
rect 5458 491862 5526 491918
rect 5582 491862 6134 491918
rect -12 491794 6134 491862
rect -12 491738 1044 491794
rect 1100 491738 1168 491794
rect 1224 491738 1292 491794
rect 1348 491738 1416 491794
rect 1472 491738 5154 491794
rect 5210 491738 5278 491794
rect 5334 491738 5402 491794
rect 5458 491738 5526 491794
rect 5582 491738 6134 491794
rect -12 491670 6134 491738
rect -12 491614 1044 491670
rect 1100 491614 1168 491670
rect 1224 491614 1292 491670
rect 1348 491614 1416 491670
rect 1472 491614 5154 491670
rect 5210 491614 5278 491670
rect 5334 491614 5402 491670
rect 5458 491614 5526 491670
rect 5582 491614 6134 491670
rect -12 491546 6134 491614
rect -12 491490 1044 491546
rect 1100 491490 1168 491546
rect 1224 491490 1292 491546
rect 1348 491490 1416 491546
rect 1472 491490 5154 491546
rect 5210 491490 5278 491546
rect 5334 491490 5402 491546
rect 5458 491490 5526 491546
rect 5582 491490 6134 491546
rect -12 491394 6134 491490
rect 595211 491918 599996 492014
rect 595211 491862 598512 491918
rect 598568 491862 598636 491918
rect 598692 491862 598760 491918
rect 598816 491862 598884 491918
rect 598940 491862 599996 491918
rect 595211 491794 599996 491862
rect 595211 491738 598512 491794
rect 598568 491738 598636 491794
rect 598692 491738 598760 491794
rect 598816 491738 598884 491794
rect 598940 491738 599996 491794
rect 595211 491670 599996 491738
rect 595211 491614 598512 491670
rect 598568 491614 598636 491670
rect 598692 491614 598760 491670
rect 598816 491614 598884 491670
rect 598940 491614 599996 491670
rect 595211 491546 599996 491614
rect 595211 491490 598512 491546
rect 598568 491490 598636 491546
rect 598692 491490 598760 491546
rect 598816 491490 598884 491546
rect 598940 491490 599996 491546
rect 595211 491394 599996 491490
rect -12 479918 6134 480014
rect -12 479862 84 479918
rect 140 479862 208 479918
rect 264 479862 332 479918
rect 388 479862 456 479918
rect 512 479862 6134 479918
rect -12 479794 6134 479862
rect -12 479738 84 479794
rect 140 479738 208 479794
rect 264 479738 332 479794
rect 388 479738 456 479794
rect 512 479738 6134 479794
rect -12 479670 6134 479738
rect -12 479614 84 479670
rect 140 479614 208 479670
rect 264 479614 332 479670
rect 388 479614 456 479670
rect 512 479614 6134 479670
rect -12 479546 6134 479614
rect -12 479490 84 479546
rect 140 479490 208 479546
rect 264 479490 332 479546
rect 388 479490 456 479546
rect 512 479490 6134 479546
rect -12 479394 6134 479490
rect 595211 479918 599996 480014
rect 595211 479862 599472 479918
rect 599528 479862 599596 479918
rect 599652 479862 599720 479918
rect 599776 479862 599844 479918
rect 599900 479862 599996 479918
rect 595211 479794 599996 479862
rect 595211 479738 599472 479794
rect 599528 479738 599596 479794
rect 599652 479738 599720 479794
rect 599776 479738 599844 479794
rect 599900 479738 599996 479794
rect 595211 479670 599996 479738
rect 595211 479614 599472 479670
rect 599528 479614 599596 479670
rect 599652 479614 599720 479670
rect 599776 479614 599844 479670
rect 599900 479614 599996 479670
rect 595211 479546 599996 479614
rect 595211 479490 599472 479546
rect 599528 479490 599596 479546
rect 599652 479490 599720 479546
rect 599776 479490 599844 479546
rect 599900 479490 599996 479546
rect 595211 479394 599996 479490
rect -12 473918 6134 474014
rect -12 473862 1044 473918
rect 1100 473862 1168 473918
rect 1224 473862 1292 473918
rect 1348 473862 1416 473918
rect 1472 473862 5154 473918
rect 5210 473862 5278 473918
rect 5334 473862 5402 473918
rect 5458 473862 5526 473918
rect 5582 473862 6134 473918
rect -12 473794 6134 473862
rect -12 473738 1044 473794
rect 1100 473738 1168 473794
rect 1224 473738 1292 473794
rect 1348 473738 1416 473794
rect 1472 473738 5154 473794
rect 5210 473738 5278 473794
rect 5334 473738 5402 473794
rect 5458 473738 5526 473794
rect 5582 473738 6134 473794
rect -12 473670 6134 473738
rect -12 473614 1044 473670
rect 1100 473614 1168 473670
rect 1224 473614 1292 473670
rect 1348 473614 1416 473670
rect 1472 473614 5154 473670
rect 5210 473614 5278 473670
rect 5334 473614 5402 473670
rect 5458 473614 5526 473670
rect 5582 473614 6134 473670
rect -12 473546 6134 473614
rect -12 473490 1044 473546
rect 1100 473490 1168 473546
rect 1224 473490 1292 473546
rect 1348 473490 1416 473546
rect 1472 473490 5154 473546
rect 5210 473490 5278 473546
rect 5334 473490 5402 473546
rect 5458 473490 5526 473546
rect 5582 473490 6134 473546
rect -12 473394 6134 473490
rect 595211 473918 599996 474014
rect 595211 473862 598512 473918
rect 598568 473862 598636 473918
rect 598692 473862 598760 473918
rect 598816 473862 598884 473918
rect 598940 473862 599996 473918
rect 595211 473794 599996 473862
rect 595211 473738 598512 473794
rect 598568 473738 598636 473794
rect 598692 473738 598760 473794
rect 598816 473738 598884 473794
rect 598940 473738 599996 473794
rect 595211 473670 599996 473738
rect 595211 473614 598512 473670
rect 598568 473614 598636 473670
rect 598692 473614 598760 473670
rect 598816 473614 598884 473670
rect 598940 473614 599996 473670
rect 595211 473546 599996 473614
rect 595211 473490 598512 473546
rect 598568 473490 598636 473546
rect 598692 473490 598760 473546
rect 598816 473490 598884 473546
rect 598940 473490 599996 473546
rect 595211 473394 599996 473490
rect -12 461918 6134 462014
rect -12 461862 84 461918
rect 140 461862 208 461918
rect 264 461862 332 461918
rect 388 461862 456 461918
rect 512 461862 6134 461918
rect -12 461794 6134 461862
rect -12 461738 84 461794
rect 140 461738 208 461794
rect 264 461738 332 461794
rect 388 461738 456 461794
rect 512 461738 6134 461794
rect -12 461670 6134 461738
rect -12 461614 84 461670
rect 140 461614 208 461670
rect 264 461614 332 461670
rect 388 461614 456 461670
rect 512 461614 6134 461670
rect -12 461546 6134 461614
rect -12 461490 84 461546
rect 140 461490 208 461546
rect 264 461490 332 461546
rect 388 461490 456 461546
rect 512 461490 6134 461546
rect -12 461394 6134 461490
rect 595211 461918 599996 462014
rect 595211 461862 599472 461918
rect 599528 461862 599596 461918
rect 599652 461862 599720 461918
rect 599776 461862 599844 461918
rect 599900 461862 599996 461918
rect 595211 461794 599996 461862
rect 595211 461738 599472 461794
rect 599528 461738 599596 461794
rect 599652 461738 599720 461794
rect 599776 461738 599844 461794
rect 599900 461738 599996 461794
rect 595211 461670 599996 461738
rect 595211 461614 599472 461670
rect 599528 461614 599596 461670
rect 599652 461614 599720 461670
rect 599776 461614 599844 461670
rect 599900 461614 599996 461670
rect 595211 461546 599996 461614
rect 595211 461490 599472 461546
rect 599528 461490 599596 461546
rect 599652 461490 599720 461546
rect 599776 461490 599844 461546
rect 599900 461490 599996 461546
rect 595211 461394 599996 461490
rect -12 455918 6134 456014
rect -12 455862 1044 455918
rect 1100 455862 1168 455918
rect 1224 455862 1292 455918
rect 1348 455862 1416 455918
rect 1472 455862 5154 455918
rect 5210 455862 5278 455918
rect 5334 455862 5402 455918
rect 5458 455862 5526 455918
rect 5582 455862 6134 455918
rect -12 455794 6134 455862
rect -12 455738 1044 455794
rect 1100 455738 1168 455794
rect 1224 455738 1292 455794
rect 1348 455738 1416 455794
rect 1472 455738 5154 455794
rect 5210 455738 5278 455794
rect 5334 455738 5402 455794
rect 5458 455738 5526 455794
rect 5582 455738 6134 455794
rect -12 455670 6134 455738
rect -12 455614 1044 455670
rect 1100 455614 1168 455670
rect 1224 455614 1292 455670
rect 1348 455614 1416 455670
rect 1472 455614 5154 455670
rect 5210 455614 5278 455670
rect 5334 455614 5402 455670
rect 5458 455614 5526 455670
rect 5582 455614 6134 455670
rect -12 455546 6134 455614
rect -12 455490 1044 455546
rect 1100 455490 1168 455546
rect 1224 455490 1292 455546
rect 1348 455490 1416 455546
rect 1472 455490 5154 455546
rect 5210 455490 5278 455546
rect 5334 455490 5402 455546
rect 5458 455490 5526 455546
rect 5582 455490 6134 455546
rect -12 455394 6134 455490
rect 595211 455918 599996 456014
rect 595211 455862 598512 455918
rect 598568 455862 598636 455918
rect 598692 455862 598760 455918
rect 598816 455862 598884 455918
rect 598940 455862 599996 455918
rect 595211 455794 599996 455862
rect 595211 455738 598512 455794
rect 598568 455738 598636 455794
rect 598692 455738 598760 455794
rect 598816 455738 598884 455794
rect 598940 455738 599996 455794
rect 595211 455670 599996 455738
rect 595211 455614 598512 455670
rect 598568 455614 598636 455670
rect 598692 455614 598760 455670
rect 598816 455614 598884 455670
rect 598940 455614 599996 455670
rect 595211 455546 599996 455614
rect 595211 455490 598512 455546
rect 598568 455490 598636 455546
rect 598692 455490 598760 455546
rect 598816 455490 598884 455546
rect 598940 455490 599996 455546
rect 595211 455394 599996 455490
rect -12 443918 6134 444014
rect -12 443862 84 443918
rect 140 443862 208 443918
rect 264 443862 332 443918
rect 388 443862 456 443918
rect 512 443862 6134 443918
rect -12 443794 6134 443862
rect -12 443738 84 443794
rect 140 443738 208 443794
rect 264 443738 332 443794
rect 388 443738 456 443794
rect 512 443738 6134 443794
rect -12 443670 6134 443738
rect -12 443614 84 443670
rect 140 443614 208 443670
rect 264 443614 332 443670
rect 388 443614 456 443670
rect 512 443614 6134 443670
rect -12 443546 6134 443614
rect -12 443490 84 443546
rect 140 443490 208 443546
rect 264 443490 332 443546
rect 388 443490 456 443546
rect 512 443490 6134 443546
rect -12 443394 6134 443490
rect 595211 443918 599996 444014
rect 595211 443862 599472 443918
rect 599528 443862 599596 443918
rect 599652 443862 599720 443918
rect 599776 443862 599844 443918
rect 599900 443862 599996 443918
rect 595211 443794 599996 443862
rect 595211 443738 599472 443794
rect 599528 443738 599596 443794
rect 599652 443738 599720 443794
rect 599776 443738 599844 443794
rect 599900 443738 599996 443794
rect 595211 443670 599996 443738
rect 595211 443614 599472 443670
rect 599528 443614 599596 443670
rect 599652 443614 599720 443670
rect 599776 443614 599844 443670
rect 599900 443614 599996 443670
rect 595211 443546 599996 443614
rect 595211 443490 599472 443546
rect 599528 443490 599596 443546
rect 599652 443490 599720 443546
rect 599776 443490 599844 443546
rect 599900 443490 599996 443546
rect 595211 443394 599996 443490
rect -12 437918 6134 438014
rect -12 437862 1044 437918
rect 1100 437862 1168 437918
rect 1224 437862 1292 437918
rect 1348 437862 1416 437918
rect 1472 437862 5154 437918
rect 5210 437862 5278 437918
rect 5334 437862 5402 437918
rect 5458 437862 5526 437918
rect 5582 437862 6134 437918
rect -12 437794 6134 437862
rect -12 437738 1044 437794
rect 1100 437738 1168 437794
rect 1224 437738 1292 437794
rect 1348 437738 1416 437794
rect 1472 437738 5154 437794
rect 5210 437738 5278 437794
rect 5334 437738 5402 437794
rect 5458 437738 5526 437794
rect 5582 437738 6134 437794
rect -12 437670 6134 437738
rect -12 437614 1044 437670
rect 1100 437614 1168 437670
rect 1224 437614 1292 437670
rect 1348 437614 1416 437670
rect 1472 437614 5154 437670
rect 5210 437614 5278 437670
rect 5334 437614 5402 437670
rect 5458 437614 5526 437670
rect 5582 437614 6134 437670
rect -12 437546 6134 437614
rect -12 437490 1044 437546
rect 1100 437490 1168 437546
rect 1224 437490 1292 437546
rect 1348 437490 1416 437546
rect 1472 437490 5154 437546
rect 5210 437490 5278 437546
rect 5334 437490 5402 437546
rect 5458 437490 5526 437546
rect 5582 437490 6134 437546
rect -12 437394 6134 437490
rect 595211 437918 599996 438014
rect 595211 437862 598512 437918
rect 598568 437862 598636 437918
rect 598692 437862 598760 437918
rect 598816 437862 598884 437918
rect 598940 437862 599996 437918
rect 595211 437794 599996 437862
rect 595211 437738 598512 437794
rect 598568 437738 598636 437794
rect 598692 437738 598760 437794
rect 598816 437738 598884 437794
rect 598940 437738 599996 437794
rect 595211 437670 599996 437738
rect 595211 437614 598512 437670
rect 598568 437614 598636 437670
rect 598692 437614 598760 437670
rect 598816 437614 598884 437670
rect 598940 437614 599996 437670
rect 595211 437546 599996 437614
rect 595211 437490 598512 437546
rect 598568 437490 598636 437546
rect 598692 437490 598760 437546
rect 598816 437490 598884 437546
rect 598940 437490 599996 437546
rect 595211 437394 599996 437490
rect -12 425918 6134 426014
rect -12 425862 84 425918
rect 140 425862 208 425918
rect 264 425862 332 425918
rect 388 425862 456 425918
rect 512 425862 6134 425918
rect -12 425794 6134 425862
rect -12 425738 84 425794
rect 140 425738 208 425794
rect 264 425738 332 425794
rect 388 425738 456 425794
rect 512 425738 6134 425794
rect -12 425670 6134 425738
rect -12 425614 84 425670
rect 140 425614 208 425670
rect 264 425614 332 425670
rect 388 425614 456 425670
rect 512 425614 6134 425670
rect -12 425546 6134 425614
rect -12 425490 84 425546
rect 140 425490 208 425546
rect 264 425490 332 425546
rect 388 425490 456 425546
rect 512 425490 6134 425546
rect -12 425394 6134 425490
rect 595211 425918 599996 426014
rect 595211 425862 599472 425918
rect 599528 425862 599596 425918
rect 599652 425862 599720 425918
rect 599776 425862 599844 425918
rect 599900 425862 599996 425918
rect 595211 425794 599996 425862
rect 595211 425738 599472 425794
rect 599528 425738 599596 425794
rect 599652 425738 599720 425794
rect 599776 425738 599844 425794
rect 599900 425738 599996 425794
rect 595211 425670 599996 425738
rect 595211 425614 599472 425670
rect 599528 425614 599596 425670
rect 599652 425614 599720 425670
rect 599776 425614 599844 425670
rect 599900 425614 599996 425670
rect 595211 425546 599996 425614
rect 595211 425490 599472 425546
rect 599528 425490 599596 425546
rect 599652 425490 599720 425546
rect 599776 425490 599844 425546
rect 599900 425490 599996 425546
rect 595211 425394 599996 425490
rect -12 419918 6134 420014
rect -12 419862 1044 419918
rect 1100 419862 1168 419918
rect 1224 419862 1292 419918
rect 1348 419862 1416 419918
rect 1472 419862 5154 419918
rect 5210 419862 5278 419918
rect 5334 419862 5402 419918
rect 5458 419862 5526 419918
rect 5582 419862 6134 419918
rect -12 419794 6134 419862
rect -12 419738 1044 419794
rect 1100 419738 1168 419794
rect 1224 419738 1292 419794
rect 1348 419738 1416 419794
rect 1472 419738 5154 419794
rect 5210 419738 5278 419794
rect 5334 419738 5402 419794
rect 5458 419738 5526 419794
rect 5582 419738 6134 419794
rect -12 419670 6134 419738
rect -12 419614 1044 419670
rect 1100 419614 1168 419670
rect 1224 419614 1292 419670
rect 1348 419614 1416 419670
rect 1472 419614 5154 419670
rect 5210 419614 5278 419670
rect 5334 419614 5402 419670
rect 5458 419614 5526 419670
rect 5582 419614 6134 419670
rect -12 419546 6134 419614
rect -12 419490 1044 419546
rect 1100 419490 1168 419546
rect 1224 419490 1292 419546
rect 1348 419490 1416 419546
rect 1472 419490 5154 419546
rect 5210 419490 5278 419546
rect 5334 419490 5402 419546
rect 5458 419490 5526 419546
rect 5582 419490 6134 419546
rect -12 419394 6134 419490
rect 595211 419918 599996 420014
rect 595211 419862 598512 419918
rect 598568 419862 598636 419918
rect 598692 419862 598760 419918
rect 598816 419862 598884 419918
rect 598940 419862 599996 419918
rect 595211 419794 599996 419862
rect 595211 419738 598512 419794
rect 598568 419738 598636 419794
rect 598692 419738 598760 419794
rect 598816 419738 598884 419794
rect 598940 419738 599996 419794
rect 595211 419670 599996 419738
rect 595211 419614 598512 419670
rect 598568 419614 598636 419670
rect 598692 419614 598760 419670
rect 598816 419614 598884 419670
rect 598940 419614 599996 419670
rect 595211 419546 599996 419614
rect 595211 419490 598512 419546
rect 598568 419490 598636 419546
rect 598692 419490 598760 419546
rect 598816 419490 598884 419546
rect 598940 419490 599996 419546
rect 595211 419394 599996 419490
rect -12 407918 6134 408014
rect -12 407862 84 407918
rect 140 407862 208 407918
rect 264 407862 332 407918
rect 388 407862 456 407918
rect 512 407862 6134 407918
rect -12 407794 6134 407862
rect -12 407738 84 407794
rect 140 407738 208 407794
rect 264 407738 332 407794
rect 388 407738 456 407794
rect 512 407738 6134 407794
rect -12 407670 6134 407738
rect -12 407614 84 407670
rect 140 407614 208 407670
rect 264 407614 332 407670
rect 388 407614 456 407670
rect 512 407614 6134 407670
rect -12 407546 6134 407614
rect -12 407490 84 407546
rect 140 407490 208 407546
rect 264 407490 332 407546
rect 388 407490 456 407546
rect 512 407490 6134 407546
rect -12 407394 6134 407490
rect 595211 407918 599996 408014
rect 595211 407862 599472 407918
rect 599528 407862 599596 407918
rect 599652 407862 599720 407918
rect 599776 407862 599844 407918
rect 599900 407862 599996 407918
rect 595211 407794 599996 407862
rect 595211 407738 599472 407794
rect 599528 407738 599596 407794
rect 599652 407738 599720 407794
rect 599776 407738 599844 407794
rect 599900 407738 599996 407794
rect 595211 407670 599996 407738
rect 595211 407614 599472 407670
rect 599528 407614 599596 407670
rect 599652 407614 599720 407670
rect 599776 407614 599844 407670
rect 599900 407614 599996 407670
rect 595211 407546 599996 407614
rect 595211 407490 599472 407546
rect 599528 407490 599596 407546
rect 599652 407490 599720 407546
rect 599776 407490 599844 407546
rect 599900 407490 599996 407546
rect 595211 407394 599996 407490
rect -12 401918 6134 402014
rect -12 401862 1044 401918
rect 1100 401862 1168 401918
rect 1224 401862 1292 401918
rect 1348 401862 1416 401918
rect 1472 401862 5154 401918
rect 5210 401862 5278 401918
rect 5334 401862 5402 401918
rect 5458 401862 5526 401918
rect 5582 401862 6134 401918
rect -12 401794 6134 401862
rect -12 401738 1044 401794
rect 1100 401738 1168 401794
rect 1224 401738 1292 401794
rect 1348 401738 1416 401794
rect 1472 401738 5154 401794
rect 5210 401738 5278 401794
rect 5334 401738 5402 401794
rect 5458 401738 5526 401794
rect 5582 401738 6134 401794
rect -12 401670 6134 401738
rect -12 401614 1044 401670
rect 1100 401614 1168 401670
rect 1224 401614 1292 401670
rect 1348 401614 1416 401670
rect 1472 401614 5154 401670
rect 5210 401614 5278 401670
rect 5334 401614 5402 401670
rect 5458 401614 5526 401670
rect 5582 401614 6134 401670
rect -12 401546 6134 401614
rect -12 401490 1044 401546
rect 1100 401490 1168 401546
rect 1224 401490 1292 401546
rect 1348 401490 1416 401546
rect 1472 401490 5154 401546
rect 5210 401490 5278 401546
rect 5334 401490 5402 401546
rect 5458 401490 5526 401546
rect 5582 401490 6134 401546
rect -12 401394 6134 401490
rect 595211 401918 599996 402014
rect 595211 401862 598512 401918
rect 598568 401862 598636 401918
rect 598692 401862 598760 401918
rect 598816 401862 598884 401918
rect 598940 401862 599996 401918
rect 595211 401794 599996 401862
rect 595211 401738 598512 401794
rect 598568 401738 598636 401794
rect 598692 401738 598760 401794
rect 598816 401738 598884 401794
rect 598940 401738 599996 401794
rect 595211 401670 599996 401738
rect 595211 401614 598512 401670
rect 598568 401614 598636 401670
rect 598692 401614 598760 401670
rect 598816 401614 598884 401670
rect 598940 401614 599996 401670
rect 595211 401546 599996 401614
rect 595211 401490 598512 401546
rect 598568 401490 598636 401546
rect 598692 401490 598760 401546
rect 598816 401490 598884 401546
rect 598940 401490 599996 401546
rect 595211 401394 599996 401490
rect -12 389918 6134 390014
rect -12 389862 84 389918
rect 140 389862 208 389918
rect 264 389862 332 389918
rect 388 389862 456 389918
rect 512 389862 6134 389918
rect -12 389794 6134 389862
rect -12 389738 84 389794
rect 140 389738 208 389794
rect 264 389738 332 389794
rect 388 389738 456 389794
rect 512 389738 6134 389794
rect -12 389670 6134 389738
rect -12 389614 84 389670
rect 140 389614 208 389670
rect 264 389614 332 389670
rect 388 389614 456 389670
rect 512 389614 6134 389670
rect -12 389546 6134 389614
rect -12 389490 84 389546
rect 140 389490 208 389546
rect 264 389490 332 389546
rect 388 389490 456 389546
rect 512 389490 6134 389546
rect -12 389394 6134 389490
rect 595211 389918 599996 390014
rect 595211 389862 599472 389918
rect 599528 389862 599596 389918
rect 599652 389862 599720 389918
rect 599776 389862 599844 389918
rect 599900 389862 599996 389918
rect 595211 389794 599996 389862
rect 595211 389738 599472 389794
rect 599528 389738 599596 389794
rect 599652 389738 599720 389794
rect 599776 389738 599844 389794
rect 599900 389738 599996 389794
rect 595211 389670 599996 389738
rect 595211 389614 599472 389670
rect 599528 389614 599596 389670
rect 599652 389614 599720 389670
rect 599776 389614 599844 389670
rect 599900 389614 599996 389670
rect 595211 389546 599996 389614
rect 595211 389490 599472 389546
rect 599528 389490 599596 389546
rect 599652 389490 599720 389546
rect 599776 389490 599844 389546
rect 599900 389490 599996 389546
rect 595211 389394 599996 389490
rect -12 383918 6134 384014
rect -12 383862 1044 383918
rect 1100 383862 1168 383918
rect 1224 383862 1292 383918
rect 1348 383862 1416 383918
rect 1472 383862 5154 383918
rect 5210 383862 5278 383918
rect 5334 383862 5402 383918
rect 5458 383862 5526 383918
rect 5582 383862 6134 383918
rect -12 383794 6134 383862
rect -12 383738 1044 383794
rect 1100 383738 1168 383794
rect 1224 383738 1292 383794
rect 1348 383738 1416 383794
rect 1472 383738 5154 383794
rect 5210 383738 5278 383794
rect 5334 383738 5402 383794
rect 5458 383738 5526 383794
rect 5582 383738 6134 383794
rect -12 383670 6134 383738
rect -12 383614 1044 383670
rect 1100 383614 1168 383670
rect 1224 383614 1292 383670
rect 1348 383614 1416 383670
rect 1472 383614 5154 383670
rect 5210 383614 5278 383670
rect 5334 383614 5402 383670
rect 5458 383614 5526 383670
rect 5582 383614 6134 383670
rect -12 383546 6134 383614
rect -12 383490 1044 383546
rect 1100 383490 1168 383546
rect 1224 383490 1292 383546
rect 1348 383490 1416 383546
rect 1472 383490 5154 383546
rect 5210 383490 5278 383546
rect 5334 383490 5402 383546
rect 5458 383490 5526 383546
rect 5582 383490 6134 383546
rect -12 383394 6134 383490
rect 595211 383918 599996 384014
rect 595211 383862 598512 383918
rect 598568 383862 598636 383918
rect 598692 383862 598760 383918
rect 598816 383862 598884 383918
rect 598940 383862 599996 383918
rect 595211 383794 599996 383862
rect 595211 383738 598512 383794
rect 598568 383738 598636 383794
rect 598692 383738 598760 383794
rect 598816 383738 598884 383794
rect 598940 383738 599996 383794
rect 595211 383670 599996 383738
rect 595211 383614 598512 383670
rect 598568 383614 598636 383670
rect 598692 383614 598760 383670
rect 598816 383614 598884 383670
rect 598940 383614 599996 383670
rect 595211 383546 599996 383614
rect 595211 383490 598512 383546
rect 598568 383490 598636 383546
rect 598692 383490 598760 383546
rect 598816 383490 598884 383546
rect 598940 383490 599996 383546
rect 595211 383394 599996 383490
rect -12 371918 6134 372014
rect -12 371862 84 371918
rect 140 371862 208 371918
rect 264 371862 332 371918
rect 388 371862 456 371918
rect 512 371862 6134 371918
rect -12 371794 6134 371862
rect -12 371738 84 371794
rect 140 371738 208 371794
rect 264 371738 332 371794
rect 388 371738 456 371794
rect 512 371738 6134 371794
rect -12 371670 6134 371738
rect -12 371614 84 371670
rect 140 371614 208 371670
rect 264 371614 332 371670
rect 388 371614 456 371670
rect 512 371614 6134 371670
rect -12 371546 6134 371614
rect -12 371490 84 371546
rect 140 371490 208 371546
rect 264 371490 332 371546
rect 388 371490 456 371546
rect 512 371490 6134 371546
rect -12 371394 6134 371490
rect 595211 371918 599996 372014
rect 595211 371862 599472 371918
rect 599528 371862 599596 371918
rect 599652 371862 599720 371918
rect 599776 371862 599844 371918
rect 599900 371862 599996 371918
rect 595211 371794 599996 371862
rect 595211 371738 599472 371794
rect 599528 371738 599596 371794
rect 599652 371738 599720 371794
rect 599776 371738 599844 371794
rect 599900 371738 599996 371794
rect 595211 371670 599996 371738
rect 595211 371614 599472 371670
rect 599528 371614 599596 371670
rect 599652 371614 599720 371670
rect 599776 371614 599844 371670
rect 599900 371614 599996 371670
rect 595211 371546 599996 371614
rect 595211 371490 599472 371546
rect 599528 371490 599596 371546
rect 599652 371490 599720 371546
rect 599776 371490 599844 371546
rect 599900 371490 599996 371546
rect 595211 371394 599996 371490
rect -12 365918 6134 366014
rect -12 365862 1044 365918
rect 1100 365862 1168 365918
rect 1224 365862 1292 365918
rect 1348 365862 1416 365918
rect 1472 365862 5154 365918
rect 5210 365862 5278 365918
rect 5334 365862 5402 365918
rect 5458 365862 5526 365918
rect 5582 365862 6134 365918
rect -12 365794 6134 365862
rect -12 365738 1044 365794
rect 1100 365738 1168 365794
rect 1224 365738 1292 365794
rect 1348 365738 1416 365794
rect 1472 365738 5154 365794
rect 5210 365738 5278 365794
rect 5334 365738 5402 365794
rect 5458 365738 5526 365794
rect 5582 365738 6134 365794
rect -12 365670 6134 365738
rect -12 365614 1044 365670
rect 1100 365614 1168 365670
rect 1224 365614 1292 365670
rect 1348 365614 1416 365670
rect 1472 365614 5154 365670
rect 5210 365614 5278 365670
rect 5334 365614 5402 365670
rect 5458 365614 5526 365670
rect 5582 365614 6134 365670
rect -12 365546 6134 365614
rect -12 365490 1044 365546
rect 1100 365490 1168 365546
rect 1224 365490 1292 365546
rect 1348 365490 1416 365546
rect 1472 365490 5154 365546
rect 5210 365490 5278 365546
rect 5334 365490 5402 365546
rect 5458 365490 5526 365546
rect 5582 365490 6134 365546
rect -12 365394 6134 365490
rect 595211 365918 599996 366014
rect 595211 365862 598512 365918
rect 598568 365862 598636 365918
rect 598692 365862 598760 365918
rect 598816 365862 598884 365918
rect 598940 365862 599996 365918
rect 595211 365794 599996 365862
rect 595211 365738 598512 365794
rect 598568 365738 598636 365794
rect 598692 365738 598760 365794
rect 598816 365738 598884 365794
rect 598940 365738 599996 365794
rect 595211 365670 599996 365738
rect 595211 365614 598512 365670
rect 598568 365614 598636 365670
rect 598692 365614 598760 365670
rect 598816 365614 598884 365670
rect 598940 365614 599996 365670
rect 595211 365546 599996 365614
rect 595211 365490 598512 365546
rect 598568 365490 598636 365546
rect 598692 365490 598760 365546
rect 598816 365490 598884 365546
rect 598940 365490 599996 365546
rect 595211 365394 599996 365490
rect -12 353918 6134 354014
rect -12 353862 84 353918
rect 140 353862 208 353918
rect 264 353862 332 353918
rect 388 353862 456 353918
rect 512 353862 6134 353918
rect -12 353794 6134 353862
rect -12 353738 84 353794
rect 140 353738 208 353794
rect 264 353738 332 353794
rect 388 353738 456 353794
rect 512 353738 6134 353794
rect -12 353670 6134 353738
rect -12 353614 84 353670
rect 140 353614 208 353670
rect 264 353614 332 353670
rect 388 353614 456 353670
rect 512 353614 6134 353670
rect -12 353546 6134 353614
rect -12 353490 84 353546
rect 140 353490 208 353546
rect 264 353490 332 353546
rect 388 353490 456 353546
rect 512 353490 6134 353546
rect -12 353394 6134 353490
rect 595211 353918 599996 354014
rect 595211 353862 599472 353918
rect 599528 353862 599596 353918
rect 599652 353862 599720 353918
rect 599776 353862 599844 353918
rect 599900 353862 599996 353918
rect 595211 353794 599996 353862
rect 595211 353738 599472 353794
rect 599528 353738 599596 353794
rect 599652 353738 599720 353794
rect 599776 353738 599844 353794
rect 599900 353738 599996 353794
rect 595211 353670 599996 353738
rect 595211 353614 599472 353670
rect 599528 353614 599596 353670
rect 599652 353614 599720 353670
rect 599776 353614 599844 353670
rect 599900 353614 599996 353670
rect 595211 353546 599996 353614
rect 595211 353490 599472 353546
rect 599528 353490 599596 353546
rect 599652 353490 599720 353546
rect 599776 353490 599844 353546
rect 599900 353490 599996 353546
rect 595211 353394 599996 353490
rect -12 347918 6134 348014
rect -12 347862 1044 347918
rect 1100 347862 1168 347918
rect 1224 347862 1292 347918
rect 1348 347862 1416 347918
rect 1472 347862 5154 347918
rect 5210 347862 5278 347918
rect 5334 347862 5402 347918
rect 5458 347862 5526 347918
rect 5582 347862 6134 347918
rect -12 347794 6134 347862
rect -12 347738 1044 347794
rect 1100 347738 1168 347794
rect 1224 347738 1292 347794
rect 1348 347738 1416 347794
rect 1472 347738 5154 347794
rect 5210 347738 5278 347794
rect 5334 347738 5402 347794
rect 5458 347738 5526 347794
rect 5582 347738 6134 347794
rect -12 347670 6134 347738
rect -12 347614 1044 347670
rect 1100 347614 1168 347670
rect 1224 347614 1292 347670
rect 1348 347614 1416 347670
rect 1472 347614 5154 347670
rect 5210 347614 5278 347670
rect 5334 347614 5402 347670
rect 5458 347614 5526 347670
rect 5582 347614 6134 347670
rect -12 347546 6134 347614
rect -12 347490 1044 347546
rect 1100 347490 1168 347546
rect 1224 347490 1292 347546
rect 1348 347490 1416 347546
rect 1472 347490 5154 347546
rect 5210 347490 5278 347546
rect 5334 347490 5402 347546
rect 5458 347490 5526 347546
rect 5582 347490 6134 347546
rect -12 347394 6134 347490
rect 595211 347918 599996 348014
rect 595211 347862 598512 347918
rect 598568 347862 598636 347918
rect 598692 347862 598760 347918
rect 598816 347862 598884 347918
rect 598940 347862 599996 347918
rect 595211 347794 599996 347862
rect 595211 347738 598512 347794
rect 598568 347738 598636 347794
rect 598692 347738 598760 347794
rect 598816 347738 598884 347794
rect 598940 347738 599996 347794
rect 595211 347670 599996 347738
rect 595211 347614 598512 347670
rect 598568 347614 598636 347670
rect 598692 347614 598760 347670
rect 598816 347614 598884 347670
rect 598940 347614 599996 347670
rect 595211 347546 599996 347614
rect 595211 347490 598512 347546
rect 598568 347490 598636 347546
rect 598692 347490 598760 347546
rect 598816 347490 598884 347546
rect 598940 347490 599996 347546
rect 595211 347394 599996 347490
rect -12 335918 6134 336014
rect -12 335862 84 335918
rect 140 335862 208 335918
rect 264 335862 332 335918
rect 388 335862 456 335918
rect 512 335862 6134 335918
rect -12 335794 6134 335862
rect -12 335738 84 335794
rect 140 335738 208 335794
rect 264 335738 332 335794
rect 388 335738 456 335794
rect 512 335738 6134 335794
rect -12 335670 6134 335738
rect -12 335614 84 335670
rect 140 335614 208 335670
rect 264 335614 332 335670
rect 388 335614 456 335670
rect 512 335614 6134 335670
rect -12 335546 6134 335614
rect -12 335490 84 335546
rect 140 335490 208 335546
rect 264 335490 332 335546
rect 388 335490 456 335546
rect 512 335490 6134 335546
rect -12 335394 6134 335490
rect 595211 335918 599996 336014
rect 595211 335862 599472 335918
rect 599528 335862 599596 335918
rect 599652 335862 599720 335918
rect 599776 335862 599844 335918
rect 599900 335862 599996 335918
rect 595211 335794 599996 335862
rect 595211 335738 599472 335794
rect 599528 335738 599596 335794
rect 599652 335738 599720 335794
rect 599776 335738 599844 335794
rect 599900 335738 599996 335794
rect 595211 335670 599996 335738
rect 595211 335614 599472 335670
rect 599528 335614 599596 335670
rect 599652 335614 599720 335670
rect 599776 335614 599844 335670
rect 599900 335614 599996 335670
rect 595211 335546 599996 335614
rect 595211 335490 599472 335546
rect 599528 335490 599596 335546
rect 599652 335490 599720 335546
rect 599776 335490 599844 335546
rect 599900 335490 599996 335546
rect 595211 335394 599996 335490
rect -12 329918 6134 330014
rect -12 329862 1044 329918
rect 1100 329862 1168 329918
rect 1224 329862 1292 329918
rect 1348 329862 1416 329918
rect 1472 329862 5154 329918
rect 5210 329862 5278 329918
rect 5334 329862 5402 329918
rect 5458 329862 5526 329918
rect 5582 329862 6134 329918
rect -12 329794 6134 329862
rect -12 329738 1044 329794
rect 1100 329738 1168 329794
rect 1224 329738 1292 329794
rect 1348 329738 1416 329794
rect 1472 329738 5154 329794
rect 5210 329738 5278 329794
rect 5334 329738 5402 329794
rect 5458 329738 5526 329794
rect 5582 329738 6134 329794
rect -12 329670 6134 329738
rect -12 329614 1044 329670
rect 1100 329614 1168 329670
rect 1224 329614 1292 329670
rect 1348 329614 1416 329670
rect 1472 329614 5154 329670
rect 5210 329614 5278 329670
rect 5334 329614 5402 329670
rect 5458 329614 5526 329670
rect 5582 329614 6134 329670
rect -12 329546 6134 329614
rect -12 329490 1044 329546
rect 1100 329490 1168 329546
rect 1224 329490 1292 329546
rect 1348 329490 1416 329546
rect 1472 329490 5154 329546
rect 5210 329490 5278 329546
rect 5334 329490 5402 329546
rect 5458 329490 5526 329546
rect 5582 329490 6134 329546
rect -12 329394 6134 329490
rect 595211 329918 599996 330014
rect 595211 329862 598512 329918
rect 598568 329862 598636 329918
rect 598692 329862 598760 329918
rect 598816 329862 598884 329918
rect 598940 329862 599996 329918
rect 595211 329794 599996 329862
rect 595211 329738 598512 329794
rect 598568 329738 598636 329794
rect 598692 329738 598760 329794
rect 598816 329738 598884 329794
rect 598940 329738 599996 329794
rect 595211 329670 599996 329738
rect 595211 329614 598512 329670
rect 598568 329614 598636 329670
rect 598692 329614 598760 329670
rect 598816 329614 598884 329670
rect 598940 329614 599996 329670
rect 595211 329546 599996 329614
rect 595211 329490 598512 329546
rect 598568 329490 598636 329546
rect 598692 329490 598760 329546
rect 598816 329490 598884 329546
rect 598940 329490 599996 329546
rect 595211 329394 599996 329490
rect -12 317918 6134 318014
rect -12 317862 84 317918
rect 140 317862 208 317918
rect 264 317862 332 317918
rect 388 317862 456 317918
rect 512 317862 6134 317918
rect -12 317794 6134 317862
rect -12 317738 84 317794
rect 140 317738 208 317794
rect 264 317738 332 317794
rect 388 317738 456 317794
rect 512 317738 6134 317794
rect -12 317670 6134 317738
rect -12 317614 84 317670
rect 140 317614 208 317670
rect 264 317614 332 317670
rect 388 317614 456 317670
rect 512 317614 6134 317670
rect -12 317546 6134 317614
rect -12 317490 84 317546
rect 140 317490 208 317546
rect 264 317490 332 317546
rect 388 317490 456 317546
rect 512 317490 6134 317546
rect -12 317394 6134 317490
rect 595211 317918 599996 318014
rect 595211 317862 599472 317918
rect 599528 317862 599596 317918
rect 599652 317862 599720 317918
rect 599776 317862 599844 317918
rect 599900 317862 599996 317918
rect 595211 317794 599996 317862
rect 595211 317738 599472 317794
rect 599528 317738 599596 317794
rect 599652 317738 599720 317794
rect 599776 317738 599844 317794
rect 599900 317738 599996 317794
rect 595211 317670 599996 317738
rect 595211 317614 599472 317670
rect 599528 317614 599596 317670
rect 599652 317614 599720 317670
rect 599776 317614 599844 317670
rect 599900 317614 599996 317670
rect 595211 317546 599996 317614
rect 595211 317490 599472 317546
rect 599528 317490 599596 317546
rect 599652 317490 599720 317546
rect 599776 317490 599844 317546
rect 599900 317490 599996 317546
rect 595211 317394 599996 317490
rect -12 311918 6134 312014
rect -12 311862 1044 311918
rect 1100 311862 1168 311918
rect 1224 311862 1292 311918
rect 1348 311862 1416 311918
rect 1472 311862 5154 311918
rect 5210 311862 5278 311918
rect 5334 311862 5402 311918
rect 5458 311862 5526 311918
rect 5582 311862 6134 311918
rect -12 311794 6134 311862
rect -12 311738 1044 311794
rect 1100 311738 1168 311794
rect 1224 311738 1292 311794
rect 1348 311738 1416 311794
rect 1472 311738 5154 311794
rect 5210 311738 5278 311794
rect 5334 311738 5402 311794
rect 5458 311738 5526 311794
rect 5582 311738 6134 311794
rect -12 311670 6134 311738
rect -12 311614 1044 311670
rect 1100 311614 1168 311670
rect 1224 311614 1292 311670
rect 1348 311614 1416 311670
rect 1472 311614 5154 311670
rect 5210 311614 5278 311670
rect 5334 311614 5402 311670
rect 5458 311614 5526 311670
rect 5582 311614 6134 311670
rect -12 311546 6134 311614
rect -12 311490 1044 311546
rect 1100 311490 1168 311546
rect 1224 311490 1292 311546
rect 1348 311490 1416 311546
rect 1472 311490 5154 311546
rect 5210 311490 5278 311546
rect 5334 311490 5402 311546
rect 5458 311490 5526 311546
rect 5582 311490 6134 311546
rect -12 311394 6134 311490
rect 595211 311918 599996 312014
rect 595211 311862 598512 311918
rect 598568 311862 598636 311918
rect 598692 311862 598760 311918
rect 598816 311862 598884 311918
rect 598940 311862 599996 311918
rect 595211 311794 599996 311862
rect 595211 311738 598512 311794
rect 598568 311738 598636 311794
rect 598692 311738 598760 311794
rect 598816 311738 598884 311794
rect 598940 311738 599996 311794
rect 595211 311670 599996 311738
rect 595211 311614 598512 311670
rect 598568 311614 598636 311670
rect 598692 311614 598760 311670
rect 598816 311614 598884 311670
rect 598940 311614 599996 311670
rect 595211 311546 599996 311614
rect 595211 311490 598512 311546
rect 598568 311490 598636 311546
rect 598692 311490 598760 311546
rect 598816 311490 598884 311546
rect 598940 311490 599996 311546
rect 595211 311394 599996 311490
rect -12 299918 6134 300014
rect -12 299862 84 299918
rect 140 299862 208 299918
rect 264 299862 332 299918
rect 388 299862 456 299918
rect 512 299862 6134 299918
rect -12 299794 6134 299862
rect -12 299738 84 299794
rect 140 299738 208 299794
rect 264 299738 332 299794
rect 388 299738 456 299794
rect 512 299738 6134 299794
rect -12 299670 6134 299738
rect -12 299614 84 299670
rect 140 299614 208 299670
rect 264 299614 332 299670
rect 388 299614 456 299670
rect 512 299614 6134 299670
rect -12 299546 6134 299614
rect -12 299490 84 299546
rect 140 299490 208 299546
rect 264 299490 332 299546
rect 388 299490 456 299546
rect 512 299490 6134 299546
rect -12 299394 6134 299490
rect 595211 299918 599996 300014
rect 595211 299862 599472 299918
rect 599528 299862 599596 299918
rect 599652 299862 599720 299918
rect 599776 299862 599844 299918
rect 599900 299862 599996 299918
rect 595211 299794 599996 299862
rect 595211 299738 599472 299794
rect 599528 299738 599596 299794
rect 599652 299738 599720 299794
rect 599776 299738 599844 299794
rect 599900 299738 599996 299794
rect 595211 299670 599996 299738
rect 595211 299614 599472 299670
rect 599528 299614 599596 299670
rect 599652 299614 599720 299670
rect 599776 299614 599844 299670
rect 599900 299614 599996 299670
rect 595211 299546 599996 299614
rect 595211 299490 599472 299546
rect 599528 299490 599596 299546
rect 599652 299490 599720 299546
rect 599776 299490 599844 299546
rect 599900 299490 599996 299546
rect 595211 299394 599996 299490
rect -12 293918 6134 294014
rect -12 293862 1044 293918
rect 1100 293862 1168 293918
rect 1224 293862 1292 293918
rect 1348 293862 1416 293918
rect 1472 293862 5154 293918
rect 5210 293862 5278 293918
rect 5334 293862 5402 293918
rect 5458 293862 5526 293918
rect 5582 293862 6134 293918
rect -12 293794 6134 293862
rect -12 293738 1044 293794
rect 1100 293738 1168 293794
rect 1224 293738 1292 293794
rect 1348 293738 1416 293794
rect 1472 293738 5154 293794
rect 5210 293738 5278 293794
rect 5334 293738 5402 293794
rect 5458 293738 5526 293794
rect 5582 293738 6134 293794
rect -12 293670 6134 293738
rect -12 293614 1044 293670
rect 1100 293614 1168 293670
rect 1224 293614 1292 293670
rect 1348 293614 1416 293670
rect 1472 293614 5154 293670
rect 5210 293614 5278 293670
rect 5334 293614 5402 293670
rect 5458 293614 5526 293670
rect 5582 293614 6134 293670
rect -12 293546 6134 293614
rect -12 293490 1044 293546
rect 1100 293490 1168 293546
rect 1224 293490 1292 293546
rect 1348 293490 1416 293546
rect 1472 293490 5154 293546
rect 5210 293490 5278 293546
rect 5334 293490 5402 293546
rect 5458 293490 5526 293546
rect 5582 293490 6134 293546
rect -12 293394 6134 293490
rect 595211 293918 599996 294014
rect 595211 293862 598512 293918
rect 598568 293862 598636 293918
rect 598692 293862 598760 293918
rect 598816 293862 598884 293918
rect 598940 293862 599996 293918
rect 595211 293794 599996 293862
rect 595211 293738 598512 293794
rect 598568 293738 598636 293794
rect 598692 293738 598760 293794
rect 598816 293738 598884 293794
rect 598940 293738 599996 293794
rect 595211 293670 599996 293738
rect 595211 293614 598512 293670
rect 598568 293614 598636 293670
rect 598692 293614 598760 293670
rect 598816 293614 598884 293670
rect 598940 293614 599996 293670
rect 595211 293546 599996 293614
rect 595211 293490 598512 293546
rect 598568 293490 598636 293546
rect 598692 293490 598760 293546
rect 598816 293490 598884 293546
rect 598940 293490 599996 293546
rect 595211 293394 599996 293490
rect -12 281918 6134 282014
rect -12 281862 84 281918
rect 140 281862 208 281918
rect 264 281862 332 281918
rect 388 281862 456 281918
rect 512 281862 6134 281918
rect -12 281794 6134 281862
rect -12 281738 84 281794
rect 140 281738 208 281794
rect 264 281738 332 281794
rect 388 281738 456 281794
rect 512 281738 6134 281794
rect -12 281670 6134 281738
rect -12 281614 84 281670
rect 140 281614 208 281670
rect 264 281614 332 281670
rect 388 281614 456 281670
rect 512 281614 6134 281670
rect -12 281546 6134 281614
rect -12 281490 84 281546
rect 140 281490 208 281546
rect 264 281490 332 281546
rect 388 281490 456 281546
rect 512 281490 6134 281546
rect -12 281394 6134 281490
rect 595211 281918 599996 282014
rect 595211 281862 599472 281918
rect 599528 281862 599596 281918
rect 599652 281862 599720 281918
rect 599776 281862 599844 281918
rect 599900 281862 599996 281918
rect 595211 281794 599996 281862
rect 595211 281738 599472 281794
rect 599528 281738 599596 281794
rect 599652 281738 599720 281794
rect 599776 281738 599844 281794
rect 599900 281738 599996 281794
rect 595211 281670 599996 281738
rect 595211 281614 599472 281670
rect 599528 281614 599596 281670
rect 599652 281614 599720 281670
rect 599776 281614 599844 281670
rect 599900 281614 599996 281670
rect 595211 281546 599996 281614
rect 595211 281490 599472 281546
rect 599528 281490 599596 281546
rect 599652 281490 599720 281546
rect 599776 281490 599844 281546
rect 599900 281490 599996 281546
rect 595211 281394 599996 281490
rect -12 275918 6134 276014
rect -12 275862 1044 275918
rect 1100 275862 1168 275918
rect 1224 275862 1292 275918
rect 1348 275862 1416 275918
rect 1472 275862 5154 275918
rect 5210 275862 5278 275918
rect 5334 275862 5402 275918
rect 5458 275862 5526 275918
rect 5582 275862 6134 275918
rect -12 275794 6134 275862
rect -12 275738 1044 275794
rect 1100 275738 1168 275794
rect 1224 275738 1292 275794
rect 1348 275738 1416 275794
rect 1472 275738 5154 275794
rect 5210 275738 5278 275794
rect 5334 275738 5402 275794
rect 5458 275738 5526 275794
rect 5582 275738 6134 275794
rect -12 275670 6134 275738
rect -12 275614 1044 275670
rect 1100 275614 1168 275670
rect 1224 275614 1292 275670
rect 1348 275614 1416 275670
rect 1472 275614 5154 275670
rect 5210 275614 5278 275670
rect 5334 275614 5402 275670
rect 5458 275614 5526 275670
rect 5582 275614 6134 275670
rect -12 275546 6134 275614
rect -12 275490 1044 275546
rect 1100 275490 1168 275546
rect 1224 275490 1292 275546
rect 1348 275490 1416 275546
rect 1472 275490 5154 275546
rect 5210 275490 5278 275546
rect 5334 275490 5402 275546
rect 5458 275490 5526 275546
rect 5582 275490 6134 275546
rect -12 275394 6134 275490
rect 595211 275918 599996 276014
rect 595211 275862 598512 275918
rect 598568 275862 598636 275918
rect 598692 275862 598760 275918
rect 598816 275862 598884 275918
rect 598940 275862 599996 275918
rect 595211 275794 599996 275862
rect 595211 275738 598512 275794
rect 598568 275738 598636 275794
rect 598692 275738 598760 275794
rect 598816 275738 598884 275794
rect 598940 275738 599996 275794
rect 595211 275670 599996 275738
rect 595211 275614 598512 275670
rect 598568 275614 598636 275670
rect 598692 275614 598760 275670
rect 598816 275614 598884 275670
rect 598940 275614 599996 275670
rect 595211 275546 599996 275614
rect 595211 275490 598512 275546
rect 598568 275490 598636 275546
rect 598692 275490 598760 275546
rect 598816 275490 598884 275546
rect 598940 275490 599996 275546
rect 595211 275394 599996 275490
rect -12 263918 6134 264014
rect -12 263862 84 263918
rect 140 263862 208 263918
rect 264 263862 332 263918
rect 388 263862 456 263918
rect 512 263862 6134 263918
rect -12 263794 6134 263862
rect -12 263738 84 263794
rect 140 263738 208 263794
rect 264 263738 332 263794
rect 388 263738 456 263794
rect 512 263738 6134 263794
rect -12 263670 6134 263738
rect -12 263614 84 263670
rect 140 263614 208 263670
rect 264 263614 332 263670
rect 388 263614 456 263670
rect 512 263614 6134 263670
rect -12 263546 6134 263614
rect -12 263490 84 263546
rect 140 263490 208 263546
rect 264 263490 332 263546
rect 388 263490 456 263546
rect 512 263490 6134 263546
rect -12 263394 6134 263490
rect 595211 263918 599996 264014
rect 595211 263862 599472 263918
rect 599528 263862 599596 263918
rect 599652 263862 599720 263918
rect 599776 263862 599844 263918
rect 599900 263862 599996 263918
rect 595211 263794 599996 263862
rect 595211 263738 599472 263794
rect 599528 263738 599596 263794
rect 599652 263738 599720 263794
rect 599776 263738 599844 263794
rect 599900 263738 599996 263794
rect 595211 263670 599996 263738
rect 595211 263614 599472 263670
rect 599528 263614 599596 263670
rect 599652 263614 599720 263670
rect 599776 263614 599844 263670
rect 599900 263614 599996 263670
rect 595211 263546 599996 263614
rect 595211 263490 599472 263546
rect 599528 263490 599596 263546
rect 599652 263490 599720 263546
rect 599776 263490 599844 263546
rect 599900 263490 599996 263546
rect 595211 263394 599996 263490
rect -12 257918 6134 258014
rect -12 257862 1044 257918
rect 1100 257862 1168 257918
rect 1224 257862 1292 257918
rect 1348 257862 1416 257918
rect 1472 257862 5154 257918
rect 5210 257862 5278 257918
rect 5334 257862 5402 257918
rect 5458 257862 5526 257918
rect 5582 257862 6134 257918
rect -12 257794 6134 257862
rect -12 257738 1044 257794
rect 1100 257738 1168 257794
rect 1224 257738 1292 257794
rect 1348 257738 1416 257794
rect 1472 257738 5154 257794
rect 5210 257738 5278 257794
rect 5334 257738 5402 257794
rect 5458 257738 5526 257794
rect 5582 257738 6134 257794
rect -12 257670 6134 257738
rect -12 257614 1044 257670
rect 1100 257614 1168 257670
rect 1224 257614 1292 257670
rect 1348 257614 1416 257670
rect 1472 257614 5154 257670
rect 5210 257614 5278 257670
rect 5334 257614 5402 257670
rect 5458 257614 5526 257670
rect 5582 257614 6134 257670
rect -12 257546 6134 257614
rect -12 257490 1044 257546
rect 1100 257490 1168 257546
rect 1224 257490 1292 257546
rect 1348 257490 1416 257546
rect 1472 257490 5154 257546
rect 5210 257490 5278 257546
rect 5334 257490 5402 257546
rect 5458 257490 5526 257546
rect 5582 257490 6134 257546
rect -12 257394 6134 257490
rect 595211 257918 599996 258014
rect 595211 257862 598512 257918
rect 598568 257862 598636 257918
rect 598692 257862 598760 257918
rect 598816 257862 598884 257918
rect 598940 257862 599996 257918
rect 595211 257794 599996 257862
rect 595211 257738 598512 257794
rect 598568 257738 598636 257794
rect 598692 257738 598760 257794
rect 598816 257738 598884 257794
rect 598940 257738 599996 257794
rect 595211 257670 599996 257738
rect 595211 257614 598512 257670
rect 598568 257614 598636 257670
rect 598692 257614 598760 257670
rect 598816 257614 598884 257670
rect 598940 257614 599996 257670
rect 595211 257546 599996 257614
rect 595211 257490 598512 257546
rect 598568 257490 598636 257546
rect 598692 257490 598760 257546
rect 598816 257490 598884 257546
rect 598940 257490 599996 257546
rect 595211 257394 599996 257490
rect -12 245918 6134 246014
rect -12 245862 84 245918
rect 140 245862 208 245918
rect 264 245862 332 245918
rect 388 245862 456 245918
rect 512 245862 6134 245918
rect -12 245794 6134 245862
rect -12 245738 84 245794
rect 140 245738 208 245794
rect 264 245738 332 245794
rect 388 245738 456 245794
rect 512 245738 6134 245794
rect -12 245670 6134 245738
rect -12 245614 84 245670
rect 140 245614 208 245670
rect 264 245614 332 245670
rect 388 245614 456 245670
rect 512 245614 6134 245670
rect -12 245546 6134 245614
rect -12 245490 84 245546
rect 140 245490 208 245546
rect 264 245490 332 245546
rect 388 245490 456 245546
rect 512 245490 6134 245546
rect -12 245394 6134 245490
rect 595211 245918 599996 246014
rect 595211 245862 599472 245918
rect 599528 245862 599596 245918
rect 599652 245862 599720 245918
rect 599776 245862 599844 245918
rect 599900 245862 599996 245918
rect 595211 245794 599996 245862
rect 595211 245738 599472 245794
rect 599528 245738 599596 245794
rect 599652 245738 599720 245794
rect 599776 245738 599844 245794
rect 599900 245738 599996 245794
rect 595211 245670 599996 245738
rect 595211 245614 599472 245670
rect 599528 245614 599596 245670
rect 599652 245614 599720 245670
rect 599776 245614 599844 245670
rect 599900 245614 599996 245670
rect 595211 245546 599996 245614
rect 595211 245490 599472 245546
rect 599528 245490 599596 245546
rect 599652 245490 599720 245546
rect 599776 245490 599844 245546
rect 599900 245490 599996 245546
rect 595211 245394 599996 245490
rect -12 239918 6134 240014
rect -12 239862 1044 239918
rect 1100 239862 1168 239918
rect 1224 239862 1292 239918
rect 1348 239862 1416 239918
rect 1472 239862 5154 239918
rect 5210 239862 5278 239918
rect 5334 239862 5402 239918
rect 5458 239862 5526 239918
rect 5582 239862 6134 239918
rect -12 239794 6134 239862
rect -12 239738 1044 239794
rect 1100 239738 1168 239794
rect 1224 239738 1292 239794
rect 1348 239738 1416 239794
rect 1472 239738 5154 239794
rect 5210 239738 5278 239794
rect 5334 239738 5402 239794
rect 5458 239738 5526 239794
rect 5582 239738 6134 239794
rect -12 239670 6134 239738
rect -12 239614 1044 239670
rect 1100 239614 1168 239670
rect 1224 239614 1292 239670
rect 1348 239614 1416 239670
rect 1472 239614 5154 239670
rect 5210 239614 5278 239670
rect 5334 239614 5402 239670
rect 5458 239614 5526 239670
rect 5582 239614 6134 239670
rect -12 239546 6134 239614
rect -12 239490 1044 239546
rect 1100 239490 1168 239546
rect 1224 239490 1292 239546
rect 1348 239490 1416 239546
rect 1472 239490 5154 239546
rect 5210 239490 5278 239546
rect 5334 239490 5402 239546
rect 5458 239490 5526 239546
rect 5582 239490 6134 239546
rect -12 239394 6134 239490
rect 595211 239918 599996 240014
rect 595211 239862 598512 239918
rect 598568 239862 598636 239918
rect 598692 239862 598760 239918
rect 598816 239862 598884 239918
rect 598940 239862 599996 239918
rect 595211 239794 599996 239862
rect 595211 239738 598512 239794
rect 598568 239738 598636 239794
rect 598692 239738 598760 239794
rect 598816 239738 598884 239794
rect 598940 239738 599996 239794
rect 595211 239670 599996 239738
rect 595211 239614 598512 239670
rect 598568 239614 598636 239670
rect 598692 239614 598760 239670
rect 598816 239614 598884 239670
rect 598940 239614 599996 239670
rect 595211 239546 599996 239614
rect 595211 239490 598512 239546
rect 598568 239490 598636 239546
rect 598692 239490 598760 239546
rect 598816 239490 598884 239546
rect 598940 239490 599996 239546
rect 595211 239394 599996 239490
rect -12 227918 6134 228014
rect -12 227862 84 227918
rect 140 227862 208 227918
rect 264 227862 332 227918
rect 388 227862 456 227918
rect 512 227862 6134 227918
rect -12 227794 6134 227862
rect -12 227738 84 227794
rect 140 227738 208 227794
rect 264 227738 332 227794
rect 388 227738 456 227794
rect 512 227738 6134 227794
rect -12 227670 6134 227738
rect -12 227614 84 227670
rect 140 227614 208 227670
rect 264 227614 332 227670
rect 388 227614 456 227670
rect 512 227614 6134 227670
rect -12 227546 6134 227614
rect -12 227490 84 227546
rect 140 227490 208 227546
rect 264 227490 332 227546
rect 388 227490 456 227546
rect 512 227490 6134 227546
rect -12 227394 6134 227490
rect 595211 227918 599996 228014
rect 595211 227862 599472 227918
rect 599528 227862 599596 227918
rect 599652 227862 599720 227918
rect 599776 227862 599844 227918
rect 599900 227862 599996 227918
rect 595211 227794 599996 227862
rect 595211 227738 599472 227794
rect 599528 227738 599596 227794
rect 599652 227738 599720 227794
rect 599776 227738 599844 227794
rect 599900 227738 599996 227794
rect 595211 227670 599996 227738
rect 595211 227614 599472 227670
rect 599528 227614 599596 227670
rect 599652 227614 599720 227670
rect 599776 227614 599844 227670
rect 599900 227614 599996 227670
rect 595211 227546 599996 227614
rect 595211 227490 599472 227546
rect 599528 227490 599596 227546
rect 599652 227490 599720 227546
rect 599776 227490 599844 227546
rect 599900 227490 599996 227546
rect 595211 227394 599996 227490
rect -12 221918 6134 222014
rect -12 221862 1044 221918
rect 1100 221862 1168 221918
rect 1224 221862 1292 221918
rect 1348 221862 1416 221918
rect 1472 221862 5154 221918
rect 5210 221862 5278 221918
rect 5334 221862 5402 221918
rect 5458 221862 5526 221918
rect 5582 221862 6134 221918
rect -12 221794 6134 221862
rect -12 221738 1044 221794
rect 1100 221738 1168 221794
rect 1224 221738 1292 221794
rect 1348 221738 1416 221794
rect 1472 221738 5154 221794
rect 5210 221738 5278 221794
rect 5334 221738 5402 221794
rect 5458 221738 5526 221794
rect 5582 221738 6134 221794
rect -12 221670 6134 221738
rect -12 221614 1044 221670
rect 1100 221614 1168 221670
rect 1224 221614 1292 221670
rect 1348 221614 1416 221670
rect 1472 221614 5154 221670
rect 5210 221614 5278 221670
rect 5334 221614 5402 221670
rect 5458 221614 5526 221670
rect 5582 221614 6134 221670
rect -12 221546 6134 221614
rect -12 221490 1044 221546
rect 1100 221490 1168 221546
rect 1224 221490 1292 221546
rect 1348 221490 1416 221546
rect 1472 221490 5154 221546
rect 5210 221490 5278 221546
rect 5334 221490 5402 221546
rect 5458 221490 5526 221546
rect 5582 221490 6134 221546
rect -12 221394 6134 221490
rect 595211 221918 599996 222014
rect 595211 221862 598512 221918
rect 598568 221862 598636 221918
rect 598692 221862 598760 221918
rect 598816 221862 598884 221918
rect 598940 221862 599996 221918
rect 595211 221794 599996 221862
rect 595211 221738 598512 221794
rect 598568 221738 598636 221794
rect 598692 221738 598760 221794
rect 598816 221738 598884 221794
rect 598940 221738 599996 221794
rect 595211 221670 599996 221738
rect 595211 221614 598512 221670
rect 598568 221614 598636 221670
rect 598692 221614 598760 221670
rect 598816 221614 598884 221670
rect 598940 221614 599996 221670
rect 595211 221546 599996 221614
rect 595211 221490 598512 221546
rect 598568 221490 598636 221546
rect 598692 221490 598760 221546
rect 598816 221490 598884 221546
rect 598940 221490 599996 221546
rect 595211 221394 599996 221490
rect -12 209918 6134 210014
rect -12 209862 84 209918
rect 140 209862 208 209918
rect 264 209862 332 209918
rect 388 209862 456 209918
rect 512 209862 6134 209918
rect -12 209794 6134 209862
rect -12 209738 84 209794
rect 140 209738 208 209794
rect 264 209738 332 209794
rect 388 209738 456 209794
rect 512 209738 6134 209794
rect -12 209670 6134 209738
rect -12 209614 84 209670
rect 140 209614 208 209670
rect 264 209614 332 209670
rect 388 209614 456 209670
rect 512 209614 6134 209670
rect -12 209546 6134 209614
rect -12 209490 84 209546
rect 140 209490 208 209546
rect 264 209490 332 209546
rect 388 209490 456 209546
rect 512 209490 6134 209546
rect -12 209394 6134 209490
rect 595211 209918 599996 210014
rect 595211 209862 599472 209918
rect 599528 209862 599596 209918
rect 599652 209862 599720 209918
rect 599776 209862 599844 209918
rect 599900 209862 599996 209918
rect 595211 209794 599996 209862
rect 595211 209738 599472 209794
rect 599528 209738 599596 209794
rect 599652 209738 599720 209794
rect 599776 209738 599844 209794
rect 599900 209738 599996 209794
rect 595211 209670 599996 209738
rect 595211 209614 599472 209670
rect 599528 209614 599596 209670
rect 599652 209614 599720 209670
rect 599776 209614 599844 209670
rect 599900 209614 599996 209670
rect 595211 209546 599996 209614
rect 595211 209490 599472 209546
rect 599528 209490 599596 209546
rect 599652 209490 599720 209546
rect 599776 209490 599844 209546
rect 599900 209490 599996 209546
rect 595211 209394 599996 209490
rect -12 203918 6134 204014
rect -12 203862 1044 203918
rect 1100 203862 1168 203918
rect 1224 203862 1292 203918
rect 1348 203862 1416 203918
rect 1472 203862 5154 203918
rect 5210 203862 5278 203918
rect 5334 203862 5402 203918
rect 5458 203862 5526 203918
rect 5582 203862 6134 203918
rect -12 203794 6134 203862
rect -12 203738 1044 203794
rect 1100 203738 1168 203794
rect 1224 203738 1292 203794
rect 1348 203738 1416 203794
rect 1472 203738 5154 203794
rect 5210 203738 5278 203794
rect 5334 203738 5402 203794
rect 5458 203738 5526 203794
rect 5582 203738 6134 203794
rect -12 203670 6134 203738
rect -12 203614 1044 203670
rect 1100 203614 1168 203670
rect 1224 203614 1292 203670
rect 1348 203614 1416 203670
rect 1472 203614 5154 203670
rect 5210 203614 5278 203670
rect 5334 203614 5402 203670
rect 5458 203614 5526 203670
rect 5582 203614 6134 203670
rect -12 203546 6134 203614
rect -12 203490 1044 203546
rect 1100 203490 1168 203546
rect 1224 203490 1292 203546
rect 1348 203490 1416 203546
rect 1472 203490 5154 203546
rect 5210 203490 5278 203546
rect 5334 203490 5402 203546
rect 5458 203490 5526 203546
rect 5582 203490 6134 203546
rect -12 203394 6134 203490
rect 595211 203918 599996 204014
rect 595211 203862 598512 203918
rect 598568 203862 598636 203918
rect 598692 203862 598760 203918
rect 598816 203862 598884 203918
rect 598940 203862 599996 203918
rect 595211 203794 599996 203862
rect 595211 203738 598512 203794
rect 598568 203738 598636 203794
rect 598692 203738 598760 203794
rect 598816 203738 598884 203794
rect 598940 203738 599996 203794
rect 595211 203670 599996 203738
rect 595211 203614 598512 203670
rect 598568 203614 598636 203670
rect 598692 203614 598760 203670
rect 598816 203614 598884 203670
rect 598940 203614 599996 203670
rect 595211 203546 599996 203614
rect 595211 203490 598512 203546
rect 598568 203490 598636 203546
rect 598692 203490 598760 203546
rect 598816 203490 598884 203546
rect 598940 203490 599996 203546
rect 595211 203394 599996 203490
rect -12 191918 6134 192014
rect -12 191862 84 191918
rect 140 191862 208 191918
rect 264 191862 332 191918
rect 388 191862 456 191918
rect 512 191862 6134 191918
rect -12 191794 6134 191862
rect -12 191738 84 191794
rect 140 191738 208 191794
rect 264 191738 332 191794
rect 388 191738 456 191794
rect 512 191738 6134 191794
rect -12 191670 6134 191738
rect -12 191614 84 191670
rect 140 191614 208 191670
rect 264 191614 332 191670
rect 388 191614 456 191670
rect 512 191614 6134 191670
rect -12 191546 6134 191614
rect -12 191490 84 191546
rect 140 191490 208 191546
rect 264 191490 332 191546
rect 388 191490 456 191546
rect 512 191490 6134 191546
rect -12 191394 6134 191490
rect 595211 191918 599996 192014
rect 595211 191862 599472 191918
rect 599528 191862 599596 191918
rect 599652 191862 599720 191918
rect 599776 191862 599844 191918
rect 599900 191862 599996 191918
rect 595211 191794 599996 191862
rect 595211 191738 599472 191794
rect 599528 191738 599596 191794
rect 599652 191738 599720 191794
rect 599776 191738 599844 191794
rect 599900 191738 599996 191794
rect 595211 191670 599996 191738
rect 595211 191614 599472 191670
rect 599528 191614 599596 191670
rect 599652 191614 599720 191670
rect 599776 191614 599844 191670
rect 599900 191614 599996 191670
rect 595211 191546 599996 191614
rect 595211 191490 599472 191546
rect 599528 191490 599596 191546
rect 599652 191490 599720 191546
rect 599776 191490 599844 191546
rect 599900 191490 599996 191546
rect 595211 191394 599996 191490
rect -12 185918 6134 186014
rect -12 185862 1044 185918
rect 1100 185862 1168 185918
rect 1224 185862 1292 185918
rect 1348 185862 1416 185918
rect 1472 185862 5154 185918
rect 5210 185862 5278 185918
rect 5334 185862 5402 185918
rect 5458 185862 5526 185918
rect 5582 185862 6134 185918
rect -12 185794 6134 185862
rect -12 185738 1044 185794
rect 1100 185738 1168 185794
rect 1224 185738 1292 185794
rect 1348 185738 1416 185794
rect 1472 185738 5154 185794
rect 5210 185738 5278 185794
rect 5334 185738 5402 185794
rect 5458 185738 5526 185794
rect 5582 185738 6134 185794
rect -12 185670 6134 185738
rect -12 185614 1044 185670
rect 1100 185614 1168 185670
rect 1224 185614 1292 185670
rect 1348 185614 1416 185670
rect 1472 185614 5154 185670
rect 5210 185614 5278 185670
rect 5334 185614 5402 185670
rect 5458 185614 5526 185670
rect 5582 185614 6134 185670
rect -12 185546 6134 185614
rect -12 185490 1044 185546
rect 1100 185490 1168 185546
rect 1224 185490 1292 185546
rect 1348 185490 1416 185546
rect 1472 185490 5154 185546
rect 5210 185490 5278 185546
rect 5334 185490 5402 185546
rect 5458 185490 5526 185546
rect 5582 185490 6134 185546
rect -12 185394 6134 185490
rect 595211 185918 599996 186014
rect 595211 185862 598512 185918
rect 598568 185862 598636 185918
rect 598692 185862 598760 185918
rect 598816 185862 598884 185918
rect 598940 185862 599996 185918
rect 595211 185794 599996 185862
rect 595211 185738 598512 185794
rect 598568 185738 598636 185794
rect 598692 185738 598760 185794
rect 598816 185738 598884 185794
rect 598940 185738 599996 185794
rect 595211 185670 599996 185738
rect 595211 185614 598512 185670
rect 598568 185614 598636 185670
rect 598692 185614 598760 185670
rect 598816 185614 598884 185670
rect 598940 185614 599996 185670
rect 595211 185546 599996 185614
rect 595211 185490 598512 185546
rect 598568 185490 598636 185546
rect 598692 185490 598760 185546
rect 598816 185490 598884 185546
rect 598940 185490 599996 185546
rect 595211 185394 599996 185490
rect -12 173918 6134 174014
rect -12 173862 84 173918
rect 140 173862 208 173918
rect 264 173862 332 173918
rect 388 173862 456 173918
rect 512 173862 6134 173918
rect -12 173794 6134 173862
rect -12 173738 84 173794
rect 140 173738 208 173794
rect 264 173738 332 173794
rect 388 173738 456 173794
rect 512 173738 6134 173794
rect -12 173670 6134 173738
rect -12 173614 84 173670
rect 140 173614 208 173670
rect 264 173614 332 173670
rect 388 173614 456 173670
rect 512 173614 6134 173670
rect -12 173546 6134 173614
rect -12 173490 84 173546
rect 140 173490 208 173546
rect 264 173490 332 173546
rect 388 173490 456 173546
rect 512 173490 6134 173546
rect -12 173394 6134 173490
rect 595211 173918 599996 174014
rect 595211 173862 599472 173918
rect 599528 173862 599596 173918
rect 599652 173862 599720 173918
rect 599776 173862 599844 173918
rect 599900 173862 599996 173918
rect 595211 173794 599996 173862
rect 595211 173738 599472 173794
rect 599528 173738 599596 173794
rect 599652 173738 599720 173794
rect 599776 173738 599844 173794
rect 599900 173738 599996 173794
rect 595211 173670 599996 173738
rect 595211 173614 599472 173670
rect 599528 173614 599596 173670
rect 599652 173614 599720 173670
rect 599776 173614 599844 173670
rect 599900 173614 599996 173670
rect 595211 173546 599996 173614
rect 595211 173490 599472 173546
rect 599528 173490 599596 173546
rect 599652 173490 599720 173546
rect 599776 173490 599844 173546
rect 599900 173490 599996 173546
rect 595211 173394 599996 173490
rect -12 167918 6134 168014
rect -12 167862 1044 167918
rect 1100 167862 1168 167918
rect 1224 167862 1292 167918
rect 1348 167862 1416 167918
rect 1472 167862 5154 167918
rect 5210 167862 5278 167918
rect 5334 167862 5402 167918
rect 5458 167862 5526 167918
rect 5582 167862 6134 167918
rect -12 167794 6134 167862
rect -12 167738 1044 167794
rect 1100 167738 1168 167794
rect 1224 167738 1292 167794
rect 1348 167738 1416 167794
rect 1472 167738 5154 167794
rect 5210 167738 5278 167794
rect 5334 167738 5402 167794
rect 5458 167738 5526 167794
rect 5582 167738 6134 167794
rect -12 167670 6134 167738
rect -12 167614 1044 167670
rect 1100 167614 1168 167670
rect 1224 167614 1292 167670
rect 1348 167614 1416 167670
rect 1472 167614 5154 167670
rect 5210 167614 5278 167670
rect 5334 167614 5402 167670
rect 5458 167614 5526 167670
rect 5582 167614 6134 167670
rect -12 167546 6134 167614
rect -12 167490 1044 167546
rect 1100 167490 1168 167546
rect 1224 167490 1292 167546
rect 1348 167490 1416 167546
rect 1472 167490 5154 167546
rect 5210 167490 5278 167546
rect 5334 167490 5402 167546
rect 5458 167490 5526 167546
rect 5582 167490 6134 167546
rect -12 167394 6134 167490
rect 595211 167918 599996 168014
rect 595211 167862 598512 167918
rect 598568 167862 598636 167918
rect 598692 167862 598760 167918
rect 598816 167862 598884 167918
rect 598940 167862 599996 167918
rect 595211 167794 599996 167862
rect 595211 167738 598512 167794
rect 598568 167738 598636 167794
rect 598692 167738 598760 167794
rect 598816 167738 598884 167794
rect 598940 167738 599996 167794
rect 595211 167670 599996 167738
rect 595211 167614 598512 167670
rect 598568 167614 598636 167670
rect 598692 167614 598760 167670
rect 598816 167614 598884 167670
rect 598940 167614 599996 167670
rect 595211 167546 599996 167614
rect 595211 167490 598512 167546
rect 598568 167490 598636 167546
rect 598692 167490 598760 167546
rect 598816 167490 598884 167546
rect 598940 167490 599996 167546
rect 595211 167394 599996 167490
rect -12 155918 6134 156014
rect -12 155862 84 155918
rect 140 155862 208 155918
rect 264 155862 332 155918
rect 388 155862 456 155918
rect 512 155862 6134 155918
rect -12 155794 6134 155862
rect -12 155738 84 155794
rect 140 155738 208 155794
rect 264 155738 332 155794
rect 388 155738 456 155794
rect 512 155738 6134 155794
rect -12 155670 6134 155738
rect -12 155614 84 155670
rect 140 155614 208 155670
rect 264 155614 332 155670
rect 388 155614 456 155670
rect 512 155614 6134 155670
rect -12 155546 6134 155614
rect -12 155490 84 155546
rect 140 155490 208 155546
rect 264 155490 332 155546
rect 388 155490 456 155546
rect 512 155490 6134 155546
rect -12 155394 6134 155490
rect 595211 155918 599996 156014
rect 595211 155862 599472 155918
rect 599528 155862 599596 155918
rect 599652 155862 599720 155918
rect 599776 155862 599844 155918
rect 599900 155862 599996 155918
rect 595211 155794 599996 155862
rect 595211 155738 599472 155794
rect 599528 155738 599596 155794
rect 599652 155738 599720 155794
rect 599776 155738 599844 155794
rect 599900 155738 599996 155794
rect 595211 155670 599996 155738
rect 595211 155614 599472 155670
rect 599528 155614 599596 155670
rect 599652 155614 599720 155670
rect 599776 155614 599844 155670
rect 599900 155614 599996 155670
rect 595211 155546 599996 155614
rect 595211 155490 599472 155546
rect 599528 155490 599596 155546
rect 599652 155490 599720 155546
rect 599776 155490 599844 155546
rect 599900 155490 599996 155546
rect 595211 155394 599996 155490
rect -12 149918 6134 150014
rect -12 149862 1044 149918
rect 1100 149862 1168 149918
rect 1224 149862 1292 149918
rect 1348 149862 1416 149918
rect 1472 149862 5154 149918
rect 5210 149862 5278 149918
rect 5334 149862 5402 149918
rect 5458 149862 5526 149918
rect 5582 149862 6134 149918
rect -12 149794 6134 149862
rect -12 149738 1044 149794
rect 1100 149738 1168 149794
rect 1224 149738 1292 149794
rect 1348 149738 1416 149794
rect 1472 149738 5154 149794
rect 5210 149738 5278 149794
rect 5334 149738 5402 149794
rect 5458 149738 5526 149794
rect 5582 149738 6134 149794
rect -12 149670 6134 149738
rect -12 149614 1044 149670
rect 1100 149614 1168 149670
rect 1224 149614 1292 149670
rect 1348 149614 1416 149670
rect 1472 149614 5154 149670
rect 5210 149614 5278 149670
rect 5334 149614 5402 149670
rect 5458 149614 5526 149670
rect 5582 149614 6134 149670
rect -12 149546 6134 149614
rect -12 149490 1044 149546
rect 1100 149490 1168 149546
rect 1224 149490 1292 149546
rect 1348 149490 1416 149546
rect 1472 149490 5154 149546
rect 5210 149490 5278 149546
rect 5334 149490 5402 149546
rect 5458 149490 5526 149546
rect 5582 149490 6134 149546
rect -12 149394 6134 149490
rect 595211 149918 599996 150014
rect 595211 149862 598512 149918
rect 598568 149862 598636 149918
rect 598692 149862 598760 149918
rect 598816 149862 598884 149918
rect 598940 149862 599996 149918
rect 595211 149794 599996 149862
rect 595211 149738 598512 149794
rect 598568 149738 598636 149794
rect 598692 149738 598760 149794
rect 598816 149738 598884 149794
rect 598940 149738 599996 149794
rect 595211 149670 599996 149738
rect 595211 149614 598512 149670
rect 598568 149614 598636 149670
rect 598692 149614 598760 149670
rect 598816 149614 598884 149670
rect 598940 149614 599996 149670
rect 595211 149546 599996 149614
rect 595211 149490 598512 149546
rect 598568 149490 598636 149546
rect 598692 149490 598760 149546
rect 598816 149490 598884 149546
rect 598940 149490 599996 149546
rect 595211 149394 599996 149490
rect -12 137918 6134 138014
rect -12 137862 84 137918
rect 140 137862 208 137918
rect 264 137862 332 137918
rect 388 137862 456 137918
rect 512 137862 6134 137918
rect -12 137794 6134 137862
rect -12 137738 84 137794
rect 140 137738 208 137794
rect 264 137738 332 137794
rect 388 137738 456 137794
rect 512 137738 6134 137794
rect -12 137670 6134 137738
rect -12 137614 84 137670
rect 140 137614 208 137670
rect 264 137614 332 137670
rect 388 137614 456 137670
rect 512 137614 6134 137670
rect -12 137546 6134 137614
rect -12 137490 84 137546
rect 140 137490 208 137546
rect 264 137490 332 137546
rect 388 137490 456 137546
rect 512 137490 6134 137546
rect -12 137394 6134 137490
rect 595211 137918 599996 138014
rect 595211 137862 599472 137918
rect 599528 137862 599596 137918
rect 599652 137862 599720 137918
rect 599776 137862 599844 137918
rect 599900 137862 599996 137918
rect 595211 137794 599996 137862
rect 595211 137738 599472 137794
rect 599528 137738 599596 137794
rect 599652 137738 599720 137794
rect 599776 137738 599844 137794
rect 599900 137738 599996 137794
rect 595211 137670 599996 137738
rect 595211 137614 599472 137670
rect 599528 137614 599596 137670
rect 599652 137614 599720 137670
rect 599776 137614 599844 137670
rect 599900 137614 599996 137670
rect 595211 137546 599996 137614
rect 595211 137490 599472 137546
rect 599528 137490 599596 137546
rect 599652 137490 599720 137546
rect 599776 137490 599844 137546
rect 599900 137490 599996 137546
rect 595211 137394 599996 137490
rect -12 131918 6134 132014
rect -12 131862 1044 131918
rect 1100 131862 1168 131918
rect 1224 131862 1292 131918
rect 1348 131862 1416 131918
rect 1472 131862 5154 131918
rect 5210 131862 5278 131918
rect 5334 131862 5402 131918
rect 5458 131862 5526 131918
rect 5582 131862 6134 131918
rect -12 131794 6134 131862
rect -12 131738 1044 131794
rect 1100 131738 1168 131794
rect 1224 131738 1292 131794
rect 1348 131738 1416 131794
rect 1472 131738 5154 131794
rect 5210 131738 5278 131794
rect 5334 131738 5402 131794
rect 5458 131738 5526 131794
rect 5582 131738 6134 131794
rect -12 131670 6134 131738
rect -12 131614 1044 131670
rect 1100 131614 1168 131670
rect 1224 131614 1292 131670
rect 1348 131614 1416 131670
rect 1472 131614 5154 131670
rect 5210 131614 5278 131670
rect 5334 131614 5402 131670
rect 5458 131614 5526 131670
rect 5582 131614 6134 131670
rect -12 131546 6134 131614
rect -12 131490 1044 131546
rect 1100 131490 1168 131546
rect 1224 131490 1292 131546
rect 1348 131490 1416 131546
rect 1472 131490 5154 131546
rect 5210 131490 5278 131546
rect 5334 131490 5402 131546
rect 5458 131490 5526 131546
rect 5582 131490 6134 131546
rect -12 131394 6134 131490
rect 595211 131918 599996 132014
rect 595211 131862 598512 131918
rect 598568 131862 598636 131918
rect 598692 131862 598760 131918
rect 598816 131862 598884 131918
rect 598940 131862 599996 131918
rect 595211 131794 599996 131862
rect 595211 131738 598512 131794
rect 598568 131738 598636 131794
rect 598692 131738 598760 131794
rect 598816 131738 598884 131794
rect 598940 131738 599996 131794
rect 595211 131670 599996 131738
rect 595211 131614 598512 131670
rect 598568 131614 598636 131670
rect 598692 131614 598760 131670
rect 598816 131614 598884 131670
rect 598940 131614 599996 131670
rect 595211 131546 599996 131614
rect 595211 131490 598512 131546
rect 598568 131490 598636 131546
rect 598692 131490 598760 131546
rect 598816 131490 598884 131546
rect 598940 131490 599996 131546
rect 595211 131394 599996 131490
rect -12 119918 6134 120014
rect -12 119862 84 119918
rect 140 119862 208 119918
rect 264 119862 332 119918
rect 388 119862 456 119918
rect 512 119862 6134 119918
rect -12 119794 6134 119862
rect -12 119738 84 119794
rect 140 119738 208 119794
rect 264 119738 332 119794
rect 388 119738 456 119794
rect 512 119738 6134 119794
rect -12 119670 6134 119738
rect -12 119614 84 119670
rect 140 119614 208 119670
rect 264 119614 332 119670
rect 388 119614 456 119670
rect 512 119614 6134 119670
rect -12 119546 6134 119614
rect -12 119490 84 119546
rect 140 119490 208 119546
rect 264 119490 332 119546
rect 388 119490 456 119546
rect 512 119490 6134 119546
rect -12 119394 6134 119490
rect 595211 119918 599996 120014
rect 595211 119862 599472 119918
rect 599528 119862 599596 119918
rect 599652 119862 599720 119918
rect 599776 119862 599844 119918
rect 599900 119862 599996 119918
rect 595211 119794 599996 119862
rect 595211 119738 599472 119794
rect 599528 119738 599596 119794
rect 599652 119738 599720 119794
rect 599776 119738 599844 119794
rect 599900 119738 599996 119794
rect 595211 119670 599996 119738
rect 595211 119614 599472 119670
rect 599528 119614 599596 119670
rect 599652 119614 599720 119670
rect 599776 119614 599844 119670
rect 599900 119614 599996 119670
rect 595211 119546 599996 119614
rect 595211 119490 599472 119546
rect 599528 119490 599596 119546
rect 599652 119490 599720 119546
rect 599776 119490 599844 119546
rect 599900 119490 599996 119546
rect 595211 119394 599996 119490
rect -12 113918 6134 114014
rect -12 113862 1044 113918
rect 1100 113862 1168 113918
rect 1224 113862 1292 113918
rect 1348 113862 1416 113918
rect 1472 113862 5154 113918
rect 5210 113862 5278 113918
rect 5334 113862 5402 113918
rect 5458 113862 5526 113918
rect 5582 113862 6134 113918
rect -12 113794 6134 113862
rect -12 113738 1044 113794
rect 1100 113738 1168 113794
rect 1224 113738 1292 113794
rect 1348 113738 1416 113794
rect 1472 113738 5154 113794
rect 5210 113738 5278 113794
rect 5334 113738 5402 113794
rect 5458 113738 5526 113794
rect 5582 113738 6134 113794
rect -12 113670 6134 113738
rect -12 113614 1044 113670
rect 1100 113614 1168 113670
rect 1224 113614 1292 113670
rect 1348 113614 1416 113670
rect 1472 113614 5154 113670
rect 5210 113614 5278 113670
rect 5334 113614 5402 113670
rect 5458 113614 5526 113670
rect 5582 113614 6134 113670
rect -12 113546 6134 113614
rect -12 113490 1044 113546
rect 1100 113490 1168 113546
rect 1224 113490 1292 113546
rect 1348 113490 1416 113546
rect 1472 113490 5154 113546
rect 5210 113490 5278 113546
rect 5334 113490 5402 113546
rect 5458 113490 5526 113546
rect 5582 113490 6134 113546
rect -12 113394 6134 113490
rect 595211 113918 599996 114014
rect 595211 113862 598512 113918
rect 598568 113862 598636 113918
rect 598692 113862 598760 113918
rect 598816 113862 598884 113918
rect 598940 113862 599996 113918
rect 595211 113794 599996 113862
rect 595211 113738 598512 113794
rect 598568 113738 598636 113794
rect 598692 113738 598760 113794
rect 598816 113738 598884 113794
rect 598940 113738 599996 113794
rect 595211 113670 599996 113738
rect 595211 113614 598512 113670
rect 598568 113614 598636 113670
rect 598692 113614 598760 113670
rect 598816 113614 598884 113670
rect 598940 113614 599996 113670
rect 595211 113546 599996 113614
rect 595211 113490 598512 113546
rect 598568 113490 598636 113546
rect 598692 113490 598760 113546
rect 598816 113490 598884 113546
rect 598940 113490 599996 113546
rect 595211 113394 599996 113490
rect -12 101918 6134 102014
rect -12 101862 84 101918
rect 140 101862 208 101918
rect 264 101862 332 101918
rect 388 101862 456 101918
rect 512 101862 6134 101918
rect -12 101794 6134 101862
rect -12 101738 84 101794
rect 140 101738 208 101794
rect 264 101738 332 101794
rect 388 101738 456 101794
rect 512 101738 6134 101794
rect -12 101670 6134 101738
rect -12 101614 84 101670
rect 140 101614 208 101670
rect 264 101614 332 101670
rect 388 101614 456 101670
rect 512 101614 6134 101670
rect -12 101546 6134 101614
rect -12 101490 84 101546
rect 140 101490 208 101546
rect 264 101490 332 101546
rect 388 101490 456 101546
rect 512 101490 6134 101546
rect -12 101394 6134 101490
rect 595211 101918 599996 102014
rect 595211 101862 599472 101918
rect 599528 101862 599596 101918
rect 599652 101862 599720 101918
rect 599776 101862 599844 101918
rect 599900 101862 599996 101918
rect 595211 101794 599996 101862
rect 595211 101738 599472 101794
rect 599528 101738 599596 101794
rect 599652 101738 599720 101794
rect 599776 101738 599844 101794
rect 599900 101738 599996 101794
rect 595211 101670 599996 101738
rect 595211 101614 599472 101670
rect 599528 101614 599596 101670
rect 599652 101614 599720 101670
rect 599776 101614 599844 101670
rect 599900 101614 599996 101670
rect 595211 101546 599996 101614
rect 595211 101490 599472 101546
rect 599528 101490 599596 101546
rect 599652 101490 599720 101546
rect 599776 101490 599844 101546
rect 599900 101490 599996 101546
rect 595211 101394 599996 101490
rect -12 95918 6134 96014
rect -12 95862 1044 95918
rect 1100 95862 1168 95918
rect 1224 95862 1292 95918
rect 1348 95862 1416 95918
rect 1472 95862 5154 95918
rect 5210 95862 5278 95918
rect 5334 95862 5402 95918
rect 5458 95862 5526 95918
rect 5582 95862 6134 95918
rect -12 95794 6134 95862
rect -12 95738 1044 95794
rect 1100 95738 1168 95794
rect 1224 95738 1292 95794
rect 1348 95738 1416 95794
rect 1472 95738 5154 95794
rect 5210 95738 5278 95794
rect 5334 95738 5402 95794
rect 5458 95738 5526 95794
rect 5582 95738 6134 95794
rect -12 95670 6134 95738
rect -12 95614 1044 95670
rect 1100 95614 1168 95670
rect 1224 95614 1292 95670
rect 1348 95614 1416 95670
rect 1472 95614 5154 95670
rect 5210 95614 5278 95670
rect 5334 95614 5402 95670
rect 5458 95614 5526 95670
rect 5582 95614 6134 95670
rect -12 95546 6134 95614
rect -12 95490 1044 95546
rect 1100 95490 1168 95546
rect 1224 95490 1292 95546
rect 1348 95490 1416 95546
rect 1472 95490 5154 95546
rect 5210 95490 5278 95546
rect 5334 95490 5402 95546
rect 5458 95490 5526 95546
rect 5582 95490 6134 95546
rect -12 95394 6134 95490
rect 595211 95918 599996 96014
rect 595211 95862 598512 95918
rect 598568 95862 598636 95918
rect 598692 95862 598760 95918
rect 598816 95862 598884 95918
rect 598940 95862 599996 95918
rect 595211 95794 599996 95862
rect 595211 95738 598512 95794
rect 598568 95738 598636 95794
rect 598692 95738 598760 95794
rect 598816 95738 598884 95794
rect 598940 95738 599996 95794
rect 595211 95670 599996 95738
rect 595211 95614 598512 95670
rect 598568 95614 598636 95670
rect 598692 95614 598760 95670
rect 598816 95614 598884 95670
rect 598940 95614 599996 95670
rect 595211 95546 599996 95614
rect 595211 95490 598512 95546
rect 598568 95490 598636 95546
rect 598692 95490 598760 95546
rect 598816 95490 598884 95546
rect 598940 95490 599996 95546
rect 595211 95394 599996 95490
rect -12 83918 6134 84014
rect -12 83862 84 83918
rect 140 83862 208 83918
rect 264 83862 332 83918
rect 388 83862 456 83918
rect 512 83862 6134 83918
rect -12 83794 6134 83862
rect -12 83738 84 83794
rect 140 83738 208 83794
rect 264 83738 332 83794
rect 388 83738 456 83794
rect 512 83738 6134 83794
rect -12 83670 6134 83738
rect -12 83614 84 83670
rect 140 83614 208 83670
rect 264 83614 332 83670
rect 388 83614 456 83670
rect 512 83614 6134 83670
rect -12 83546 6134 83614
rect -12 83490 84 83546
rect 140 83490 208 83546
rect 264 83490 332 83546
rect 388 83490 456 83546
rect 512 83490 6134 83546
rect -12 83394 6134 83490
rect 595211 83918 599996 84014
rect 595211 83862 599472 83918
rect 599528 83862 599596 83918
rect 599652 83862 599720 83918
rect 599776 83862 599844 83918
rect 599900 83862 599996 83918
rect 595211 83794 599996 83862
rect 595211 83738 599472 83794
rect 599528 83738 599596 83794
rect 599652 83738 599720 83794
rect 599776 83738 599844 83794
rect 599900 83738 599996 83794
rect 595211 83670 599996 83738
rect 595211 83614 599472 83670
rect 599528 83614 599596 83670
rect 599652 83614 599720 83670
rect 599776 83614 599844 83670
rect 599900 83614 599996 83670
rect 595211 83546 599996 83614
rect 595211 83490 599472 83546
rect 599528 83490 599596 83546
rect 599652 83490 599720 83546
rect 599776 83490 599844 83546
rect 599900 83490 599996 83546
rect 595211 83394 599996 83490
rect -12 77918 6134 78014
rect -12 77862 1044 77918
rect 1100 77862 1168 77918
rect 1224 77862 1292 77918
rect 1348 77862 1416 77918
rect 1472 77862 5154 77918
rect 5210 77862 5278 77918
rect 5334 77862 5402 77918
rect 5458 77862 5526 77918
rect 5582 77862 6134 77918
rect -12 77794 6134 77862
rect -12 77738 1044 77794
rect 1100 77738 1168 77794
rect 1224 77738 1292 77794
rect 1348 77738 1416 77794
rect 1472 77738 5154 77794
rect 5210 77738 5278 77794
rect 5334 77738 5402 77794
rect 5458 77738 5526 77794
rect 5582 77738 6134 77794
rect -12 77670 6134 77738
rect -12 77614 1044 77670
rect 1100 77614 1168 77670
rect 1224 77614 1292 77670
rect 1348 77614 1416 77670
rect 1472 77614 5154 77670
rect 5210 77614 5278 77670
rect 5334 77614 5402 77670
rect 5458 77614 5526 77670
rect 5582 77614 6134 77670
rect -12 77546 6134 77614
rect -12 77490 1044 77546
rect 1100 77490 1168 77546
rect 1224 77490 1292 77546
rect 1348 77490 1416 77546
rect 1472 77490 5154 77546
rect 5210 77490 5278 77546
rect 5334 77490 5402 77546
rect 5458 77490 5526 77546
rect 5582 77490 6134 77546
rect -12 77394 6134 77490
rect 595211 77918 599996 78014
rect 595211 77862 598512 77918
rect 598568 77862 598636 77918
rect 598692 77862 598760 77918
rect 598816 77862 598884 77918
rect 598940 77862 599996 77918
rect 595211 77794 599996 77862
rect 595211 77738 598512 77794
rect 598568 77738 598636 77794
rect 598692 77738 598760 77794
rect 598816 77738 598884 77794
rect 598940 77738 599996 77794
rect 595211 77670 599996 77738
rect 595211 77614 598512 77670
rect 598568 77614 598636 77670
rect 598692 77614 598760 77670
rect 598816 77614 598884 77670
rect 598940 77614 599996 77670
rect 595211 77546 599996 77614
rect 595211 77490 598512 77546
rect 598568 77490 598636 77546
rect 598692 77490 598760 77546
rect 598816 77490 598884 77546
rect 598940 77490 599996 77546
rect 595211 77394 599996 77490
rect -12 65918 6134 66014
rect -12 65862 84 65918
rect 140 65862 208 65918
rect 264 65862 332 65918
rect 388 65862 456 65918
rect 512 65862 6134 65918
rect -12 65794 6134 65862
rect -12 65738 84 65794
rect 140 65738 208 65794
rect 264 65738 332 65794
rect 388 65738 456 65794
rect 512 65738 6134 65794
rect -12 65670 6134 65738
rect -12 65614 84 65670
rect 140 65614 208 65670
rect 264 65614 332 65670
rect 388 65614 456 65670
rect 512 65614 6134 65670
rect -12 65546 6134 65614
rect -12 65490 84 65546
rect 140 65490 208 65546
rect 264 65490 332 65546
rect 388 65490 456 65546
rect 512 65490 6134 65546
rect -12 65394 6134 65490
rect 595211 65918 599996 66014
rect 595211 65862 599472 65918
rect 599528 65862 599596 65918
rect 599652 65862 599720 65918
rect 599776 65862 599844 65918
rect 599900 65862 599996 65918
rect 595211 65794 599996 65862
rect 595211 65738 599472 65794
rect 599528 65738 599596 65794
rect 599652 65738 599720 65794
rect 599776 65738 599844 65794
rect 599900 65738 599996 65794
rect 595211 65670 599996 65738
rect 595211 65614 599472 65670
rect 599528 65614 599596 65670
rect 599652 65614 599720 65670
rect 599776 65614 599844 65670
rect 599900 65614 599996 65670
rect 595211 65546 599996 65614
rect 595211 65490 599472 65546
rect 599528 65490 599596 65546
rect 599652 65490 599720 65546
rect 599776 65490 599844 65546
rect 599900 65490 599996 65546
rect 595211 65394 599996 65490
rect -12 59918 6134 60014
rect -12 59862 1044 59918
rect 1100 59862 1168 59918
rect 1224 59862 1292 59918
rect 1348 59862 1416 59918
rect 1472 59862 5154 59918
rect 5210 59862 5278 59918
rect 5334 59862 5402 59918
rect 5458 59862 5526 59918
rect 5582 59862 6134 59918
rect -12 59794 6134 59862
rect -12 59738 1044 59794
rect 1100 59738 1168 59794
rect 1224 59738 1292 59794
rect 1348 59738 1416 59794
rect 1472 59738 5154 59794
rect 5210 59738 5278 59794
rect 5334 59738 5402 59794
rect 5458 59738 5526 59794
rect 5582 59738 6134 59794
rect -12 59670 6134 59738
rect -12 59614 1044 59670
rect 1100 59614 1168 59670
rect 1224 59614 1292 59670
rect 1348 59614 1416 59670
rect 1472 59614 5154 59670
rect 5210 59614 5278 59670
rect 5334 59614 5402 59670
rect 5458 59614 5526 59670
rect 5582 59614 6134 59670
rect -12 59546 6134 59614
rect -12 59490 1044 59546
rect 1100 59490 1168 59546
rect 1224 59490 1292 59546
rect 1348 59490 1416 59546
rect 1472 59490 5154 59546
rect 5210 59490 5278 59546
rect 5334 59490 5402 59546
rect 5458 59490 5526 59546
rect 5582 59490 6134 59546
rect -12 59394 6134 59490
rect 595211 59918 599996 60014
rect 595211 59862 598512 59918
rect 598568 59862 598636 59918
rect 598692 59862 598760 59918
rect 598816 59862 598884 59918
rect 598940 59862 599996 59918
rect 595211 59794 599996 59862
rect 595211 59738 598512 59794
rect 598568 59738 598636 59794
rect 598692 59738 598760 59794
rect 598816 59738 598884 59794
rect 598940 59738 599996 59794
rect 595211 59670 599996 59738
rect 595211 59614 598512 59670
rect 598568 59614 598636 59670
rect 598692 59614 598760 59670
rect 598816 59614 598884 59670
rect 598940 59614 599996 59670
rect 595211 59546 599996 59614
rect 595211 59490 598512 59546
rect 598568 59490 598636 59546
rect 598692 59490 598760 59546
rect 598816 59490 598884 59546
rect 598940 59490 599996 59546
rect 595211 59394 599996 59490
rect -12 47918 6134 48014
rect -12 47862 84 47918
rect 140 47862 208 47918
rect 264 47862 332 47918
rect 388 47862 456 47918
rect 512 47862 6134 47918
rect -12 47794 6134 47862
rect -12 47738 84 47794
rect 140 47738 208 47794
rect 264 47738 332 47794
rect 388 47738 456 47794
rect 512 47738 6134 47794
rect -12 47670 6134 47738
rect -12 47614 84 47670
rect 140 47614 208 47670
rect 264 47614 332 47670
rect 388 47614 456 47670
rect 512 47614 6134 47670
rect -12 47546 6134 47614
rect -12 47490 84 47546
rect 140 47490 208 47546
rect 264 47490 332 47546
rect 388 47490 456 47546
rect 512 47490 6134 47546
rect -12 47394 6134 47490
rect 595211 47918 599996 48014
rect 595211 47862 599472 47918
rect 599528 47862 599596 47918
rect 599652 47862 599720 47918
rect 599776 47862 599844 47918
rect 599900 47862 599996 47918
rect 595211 47794 599996 47862
rect 595211 47738 599472 47794
rect 599528 47738 599596 47794
rect 599652 47738 599720 47794
rect 599776 47738 599844 47794
rect 599900 47738 599996 47794
rect 595211 47670 599996 47738
rect 595211 47614 599472 47670
rect 599528 47614 599596 47670
rect 599652 47614 599720 47670
rect 599776 47614 599844 47670
rect 599900 47614 599996 47670
rect 595211 47546 599996 47614
rect 595211 47490 599472 47546
rect 599528 47490 599596 47546
rect 599652 47490 599720 47546
rect 599776 47490 599844 47546
rect 599900 47490 599996 47546
rect 595211 47394 599996 47490
rect -12 41918 6134 42014
rect -12 41862 1044 41918
rect 1100 41862 1168 41918
rect 1224 41862 1292 41918
rect 1348 41862 1416 41918
rect 1472 41862 5154 41918
rect 5210 41862 5278 41918
rect 5334 41862 5402 41918
rect 5458 41862 5526 41918
rect 5582 41862 6134 41918
rect -12 41794 6134 41862
rect -12 41738 1044 41794
rect 1100 41738 1168 41794
rect 1224 41738 1292 41794
rect 1348 41738 1416 41794
rect 1472 41738 5154 41794
rect 5210 41738 5278 41794
rect 5334 41738 5402 41794
rect 5458 41738 5526 41794
rect 5582 41738 6134 41794
rect -12 41670 6134 41738
rect -12 41614 1044 41670
rect 1100 41614 1168 41670
rect 1224 41614 1292 41670
rect 1348 41614 1416 41670
rect 1472 41614 5154 41670
rect 5210 41614 5278 41670
rect 5334 41614 5402 41670
rect 5458 41614 5526 41670
rect 5582 41614 6134 41670
rect -12 41546 6134 41614
rect -12 41490 1044 41546
rect 1100 41490 1168 41546
rect 1224 41490 1292 41546
rect 1348 41490 1416 41546
rect 1472 41490 5154 41546
rect 5210 41490 5278 41546
rect 5334 41490 5402 41546
rect 5458 41490 5526 41546
rect 5582 41490 6134 41546
rect -12 41394 6134 41490
rect 595211 41918 599996 42014
rect 595211 41862 598512 41918
rect 598568 41862 598636 41918
rect 598692 41862 598760 41918
rect 598816 41862 598884 41918
rect 598940 41862 599996 41918
rect 595211 41794 599996 41862
rect 595211 41738 598512 41794
rect 598568 41738 598636 41794
rect 598692 41738 598760 41794
rect 598816 41738 598884 41794
rect 598940 41738 599996 41794
rect 595211 41670 599996 41738
rect 595211 41614 598512 41670
rect 598568 41614 598636 41670
rect 598692 41614 598760 41670
rect 598816 41614 598884 41670
rect 598940 41614 599996 41670
rect 595211 41546 599996 41614
rect 595211 41490 598512 41546
rect 598568 41490 598636 41546
rect 598692 41490 598760 41546
rect 598816 41490 598884 41546
rect 598940 41490 599996 41546
rect 595211 41394 599996 41490
rect -12 29918 6134 30014
rect -12 29862 84 29918
rect 140 29862 208 29918
rect 264 29862 332 29918
rect 388 29862 456 29918
rect 512 29862 6134 29918
rect -12 29794 6134 29862
rect -12 29738 84 29794
rect 140 29738 208 29794
rect 264 29738 332 29794
rect 388 29738 456 29794
rect 512 29738 6134 29794
rect -12 29670 6134 29738
rect -12 29614 84 29670
rect 140 29614 208 29670
rect 264 29614 332 29670
rect 388 29614 456 29670
rect 512 29614 6134 29670
rect -12 29546 6134 29614
rect -12 29490 84 29546
rect 140 29490 208 29546
rect 264 29490 332 29546
rect 388 29490 456 29546
rect 512 29490 6134 29546
rect -12 29394 6134 29490
rect 595211 29918 599996 30014
rect 595211 29862 599472 29918
rect 599528 29862 599596 29918
rect 599652 29862 599720 29918
rect 599776 29862 599844 29918
rect 599900 29862 599996 29918
rect 595211 29794 599996 29862
rect 595211 29738 599472 29794
rect 599528 29738 599596 29794
rect 599652 29738 599720 29794
rect 599776 29738 599844 29794
rect 599900 29738 599996 29794
rect 595211 29670 599996 29738
rect 595211 29614 599472 29670
rect 599528 29614 599596 29670
rect 599652 29614 599720 29670
rect 599776 29614 599844 29670
rect 599900 29614 599996 29670
rect 595211 29546 599996 29614
rect 595211 29490 599472 29546
rect 599528 29490 599596 29546
rect 599652 29490 599720 29546
rect 599776 29490 599844 29546
rect 599900 29490 599996 29546
rect 595211 29394 599996 29490
rect -12 23918 6134 24014
rect -12 23862 1044 23918
rect 1100 23862 1168 23918
rect 1224 23862 1292 23918
rect 1348 23862 1416 23918
rect 1472 23862 5154 23918
rect 5210 23862 5278 23918
rect 5334 23862 5402 23918
rect 5458 23862 5526 23918
rect 5582 23862 6134 23918
rect -12 23794 6134 23862
rect -12 23738 1044 23794
rect 1100 23738 1168 23794
rect 1224 23738 1292 23794
rect 1348 23738 1416 23794
rect 1472 23738 5154 23794
rect 5210 23738 5278 23794
rect 5334 23738 5402 23794
rect 5458 23738 5526 23794
rect 5582 23738 6134 23794
rect -12 23670 6134 23738
rect -12 23614 1044 23670
rect 1100 23614 1168 23670
rect 1224 23614 1292 23670
rect 1348 23614 1416 23670
rect 1472 23614 5154 23670
rect 5210 23614 5278 23670
rect 5334 23614 5402 23670
rect 5458 23614 5526 23670
rect 5582 23614 6134 23670
rect -12 23546 6134 23614
rect -12 23490 1044 23546
rect 1100 23490 1168 23546
rect 1224 23490 1292 23546
rect 1348 23490 1416 23546
rect 1472 23490 5154 23546
rect 5210 23490 5278 23546
rect 5334 23490 5402 23546
rect 5458 23490 5526 23546
rect 5582 23490 6134 23546
rect -12 23394 6134 23490
rect 595211 23918 599996 24014
rect 595211 23862 598512 23918
rect 598568 23862 598636 23918
rect 598692 23862 598760 23918
rect 598816 23862 598884 23918
rect 598940 23862 599996 23918
rect 595211 23794 599996 23862
rect 595211 23738 598512 23794
rect 598568 23738 598636 23794
rect 598692 23738 598760 23794
rect 598816 23738 598884 23794
rect 598940 23738 599996 23794
rect 595211 23670 599996 23738
rect 595211 23614 598512 23670
rect 598568 23614 598636 23670
rect 598692 23614 598760 23670
rect 598816 23614 598884 23670
rect 598940 23614 599996 23670
rect 595211 23546 599996 23614
rect 595211 23490 598512 23546
rect 598568 23490 598636 23546
rect 598692 23490 598760 23546
rect 598816 23490 598884 23546
rect 598940 23490 599996 23546
rect 595211 23394 599996 23490
rect -12 11918 6134 12014
rect -12 11862 84 11918
rect 140 11862 208 11918
rect 264 11862 332 11918
rect 388 11862 456 11918
rect 512 11862 6134 11918
rect -12 11794 6134 11862
rect -12 11738 84 11794
rect 140 11738 208 11794
rect 264 11738 332 11794
rect 388 11738 456 11794
rect 512 11738 6134 11794
rect -12 11670 6134 11738
rect -12 11614 84 11670
rect 140 11614 208 11670
rect 264 11614 332 11670
rect 388 11614 456 11670
rect 512 11614 6134 11670
rect -12 11546 6134 11614
rect -12 11490 84 11546
rect 140 11490 208 11546
rect 264 11490 332 11546
rect 388 11490 456 11546
rect 512 11490 6134 11546
rect -12 11394 6134 11490
rect 595211 11918 599996 12014
rect 595211 11862 599472 11918
rect 599528 11862 599596 11918
rect 599652 11862 599720 11918
rect 599776 11862 599844 11918
rect 599900 11862 599996 11918
rect 595211 11794 599996 11862
rect 595211 11738 599472 11794
rect 599528 11738 599596 11794
rect 599652 11738 599720 11794
rect 599776 11738 599844 11794
rect 599900 11738 599996 11794
rect 595211 11670 599996 11738
rect 595211 11614 599472 11670
rect 599528 11614 599596 11670
rect 599652 11614 599720 11670
rect 599776 11614 599844 11670
rect 599900 11614 599996 11670
rect 595211 11546 599996 11614
rect 595211 11490 599472 11546
rect 599528 11490 599596 11546
rect 599652 11490 599720 11546
rect 599776 11490 599844 11546
rect 599900 11490 599996 11546
rect 595211 11394 599996 11490
rect -12 5918 6134 6014
rect -12 5862 1044 5918
rect 1100 5862 1168 5918
rect 1224 5862 1292 5918
rect 1348 5862 1416 5918
rect 1472 5862 5154 5918
rect 5210 5862 5278 5918
rect 5334 5862 5402 5918
rect 5458 5862 5526 5918
rect 5582 5862 6134 5918
rect -12 5794 6134 5862
rect -12 5738 1044 5794
rect 1100 5738 1168 5794
rect 1224 5738 1292 5794
rect 1348 5738 1416 5794
rect 1472 5738 5154 5794
rect 5210 5738 5278 5794
rect 5334 5738 5402 5794
rect 5458 5738 5526 5794
rect 5582 5738 6134 5794
rect -12 5670 6134 5738
rect -12 5614 1044 5670
rect 1100 5614 1168 5670
rect 1224 5614 1292 5670
rect 1348 5614 1416 5670
rect 1472 5614 5154 5670
rect 5210 5614 5278 5670
rect 5334 5614 5402 5670
rect 5458 5614 5526 5670
rect 5582 5614 6134 5670
rect -12 5546 6134 5614
rect -12 5490 1044 5546
rect 1100 5490 1168 5546
rect 1224 5490 1292 5546
rect 1348 5490 1416 5546
rect 1472 5490 5154 5546
rect 5210 5490 5278 5546
rect 5334 5490 5402 5546
rect 5458 5490 5526 5546
rect 5582 5490 6134 5546
rect -12 5394 6134 5490
rect 595211 5918 599996 6014
rect 595211 5862 598512 5918
rect 598568 5862 598636 5918
rect 598692 5862 598760 5918
rect 598816 5862 598884 5918
rect 598940 5862 599996 5918
rect 595211 5794 599996 5862
rect 595211 5738 598512 5794
rect 598568 5738 598636 5794
rect 598692 5738 598760 5794
rect 598816 5738 598884 5794
rect 598940 5738 599996 5794
rect 595211 5670 599996 5738
rect 595211 5614 598512 5670
rect 598568 5614 598636 5670
rect 598692 5614 598760 5670
rect 598816 5614 598884 5670
rect 598940 5614 599996 5670
rect 595211 5546 599996 5614
rect 595211 5490 598512 5546
rect 598568 5490 598636 5546
rect 598692 5490 598760 5546
rect 598816 5490 598884 5546
rect 598940 5490 599996 5546
rect 595211 5394 599996 5490
rect 948 1808 599036 1904
rect 948 1752 1044 1808
rect 1100 1752 1168 1808
rect 1224 1752 1292 1808
rect 1348 1752 1416 1808
rect 1472 1752 5154 1808
rect 5210 1752 5278 1808
rect 5334 1752 5402 1808
rect 5458 1752 5526 1808
rect 5582 1752 23154 1808
rect 23210 1752 23278 1808
rect 23334 1752 23402 1808
rect 23458 1752 23526 1808
rect 23582 1752 41154 1808
rect 41210 1752 41278 1808
rect 41334 1752 41402 1808
rect 41458 1752 41526 1808
rect 41582 1752 59154 1808
rect 59210 1752 59278 1808
rect 59334 1752 59402 1808
rect 59458 1752 59526 1808
rect 59582 1752 77154 1808
rect 77210 1752 77278 1808
rect 77334 1752 77402 1808
rect 77458 1752 77526 1808
rect 77582 1752 95154 1808
rect 95210 1752 95278 1808
rect 95334 1752 95402 1808
rect 95458 1752 95526 1808
rect 95582 1752 113154 1808
rect 113210 1752 113278 1808
rect 113334 1752 113402 1808
rect 113458 1752 113526 1808
rect 113582 1752 131154 1808
rect 131210 1752 131278 1808
rect 131334 1752 131402 1808
rect 131458 1752 131526 1808
rect 131582 1752 149154 1808
rect 149210 1752 149278 1808
rect 149334 1752 149402 1808
rect 149458 1752 149526 1808
rect 149582 1752 167154 1808
rect 167210 1752 167278 1808
rect 167334 1752 167402 1808
rect 167458 1752 167526 1808
rect 167582 1752 185154 1808
rect 185210 1752 185278 1808
rect 185334 1752 185402 1808
rect 185458 1752 185526 1808
rect 185582 1752 203154 1808
rect 203210 1752 203278 1808
rect 203334 1752 203402 1808
rect 203458 1752 203526 1808
rect 203582 1752 221154 1808
rect 221210 1752 221278 1808
rect 221334 1752 221402 1808
rect 221458 1752 221526 1808
rect 221582 1752 239154 1808
rect 239210 1752 239278 1808
rect 239334 1752 239402 1808
rect 239458 1752 239526 1808
rect 239582 1752 257154 1808
rect 257210 1752 257278 1808
rect 257334 1752 257402 1808
rect 257458 1752 257526 1808
rect 257582 1752 275154 1808
rect 275210 1752 275278 1808
rect 275334 1752 275402 1808
rect 275458 1752 275526 1808
rect 275582 1752 293154 1808
rect 293210 1752 293278 1808
rect 293334 1752 293402 1808
rect 293458 1752 293526 1808
rect 293582 1752 311154 1808
rect 311210 1752 311278 1808
rect 311334 1752 311402 1808
rect 311458 1752 311526 1808
rect 311582 1752 329154 1808
rect 329210 1752 329278 1808
rect 329334 1752 329402 1808
rect 329458 1752 329526 1808
rect 329582 1752 347154 1808
rect 347210 1752 347278 1808
rect 347334 1752 347402 1808
rect 347458 1752 347526 1808
rect 347582 1752 365154 1808
rect 365210 1752 365278 1808
rect 365334 1752 365402 1808
rect 365458 1752 365526 1808
rect 365582 1752 383154 1808
rect 383210 1752 383278 1808
rect 383334 1752 383402 1808
rect 383458 1752 383526 1808
rect 383582 1752 401154 1808
rect 401210 1752 401278 1808
rect 401334 1752 401402 1808
rect 401458 1752 401526 1808
rect 401582 1752 419154 1808
rect 419210 1752 419278 1808
rect 419334 1752 419402 1808
rect 419458 1752 419526 1808
rect 419582 1752 437154 1808
rect 437210 1752 437278 1808
rect 437334 1752 437402 1808
rect 437458 1752 437526 1808
rect 437582 1752 455154 1808
rect 455210 1752 455278 1808
rect 455334 1752 455402 1808
rect 455458 1752 455526 1808
rect 455582 1752 473154 1808
rect 473210 1752 473278 1808
rect 473334 1752 473402 1808
rect 473458 1752 473526 1808
rect 473582 1752 491154 1808
rect 491210 1752 491278 1808
rect 491334 1752 491402 1808
rect 491458 1752 491526 1808
rect 491582 1752 509154 1808
rect 509210 1752 509278 1808
rect 509334 1752 509402 1808
rect 509458 1752 509526 1808
rect 509582 1752 527154 1808
rect 527210 1752 527278 1808
rect 527334 1752 527402 1808
rect 527458 1752 527526 1808
rect 527582 1752 545154 1808
rect 545210 1752 545278 1808
rect 545334 1752 545402 1808
rect 545458 1752 545526 1808
rect 545582 1752 563154 1808
rect 563210 1752 563278 1808
rect 563334 1752 563402 1808
rect 563458 1752 563526 1808
rect 563582 1752 581154 1808
rect 581210 1752 581278 1808
rect 581334 1752 581402 1808
rect 581458 1752 581526 1808
rect 581582 1752 598512 1808
rect 598568 1752 598636 1808
rect 598692 1752 598760 1808
rect 598816 1752 598884 1808
rect 598940 1752 599036 1808
rect 948 1684 599036 1752
rect 948 1628 1044 1684
rect 1100 1628 1168 1684
rect 1224 1628 1292 1684
rect 1348 1628 1416 1684
rect 1472 1628 5154 1684
rect 5210 1628 5278 1684
rect 5334 1628 5402 1684
rect 5458 1628 5526 1684
rect 5582 1628 23154 1684
rect 23210 1628 23278 1684
rect 23334 1628 23402 1684
rect 23458 1628 23526 1684
rect 23582 1628 41154 1684
rect 41210 1628 41278 1684
rect 41334 1628 41402 1684
rect 41458 1628 41526 1684
rect 41582 1628 59154 1684
rect 59210 1628 59278 1684
rect 59334 1628 59402 1684
rect 59458 1628 59526 1684
rect 59582 1628 77154 1684
rect 77210 1628 77278 1684
rect 77334 1628 77402 1684
rect 77458 1628 77526 1684
rect 77582 1628 95154 1684
rect 95210 1628 95278 1684
rect 95334 1628 95402 1684
rect 95458 1628 95526 1684
rect 95582 1628 113154 1684
rect 113210 1628 113278 1684
rect 113334 1628 113402 1684
rect 113458 1628 113526 1684
rect 113582 1628 131154 1684
rect 131210 1628 131278 1684
rect 131334 1628 131402 1684
rect 131458 1628 131526 1684
rect 131582 1628 149154 1684
rect 149210 1628 149278 1684
rect 149334 1628 149402 1684
rect 149458 1628 149526 1684
rect 149582 1628 167154 1684
rect 167210 1628 167278 1684
rect 167334 1628 167402 1684
rect 167458 1628 167526 1684
rect 167582 1628 185154 1684
rect 185210 1628 185278 1684
rect 185334 1628 185402 1684
rect 185458 1628 185526 1684
rect 185582 1628 203154 1684
rect 203210 1628 203278 1684
rect 203334 1628 203402 1684
rect 203458 1628 203526 1684
rect 203582 1628 221154 1684
rect 221210 1628 221278 1684
rect 221334 1628 221402 1684
rect 221458 1628 221526 1684
rect 221582 1628 239154 1684
rect 239210 1628 239278 1684
rect 239334 1628 239402 1684
rect 239458 1628 239526 1684
rect 239582 1628 257154 1684
rect 257210 1628 257278 1684
rect 257334 1628 257402 1684
rect 257458 1628 257526 1684
rect 257582 1628 275154 1684
rect 275210 1628 275278 1684
rect 275334 1628 275402 1684
rect 275458 1628 275526 1684
rect 275582 1628 293154 1684
rect 293210 1628 293278 1684
rect 293334 1628 293402 1684
rect 293458 1628 293526 1684
rect 293582 1628 311154 1684
rect 311210 1628 311278 1684
rect 311334 1628 311402 1684
rect 311458 1628 311526 1684
rect 311582 1628 329154 1684
rect 329210 1628 329278 1684
rect 329334 1628 329402 1684
rect 329458 1628 329526 1684
rect 329582 1628 347154 1684
rect 347210 1628 347278 1684
rect 347334 1628 347402 1684
rect 347458 1628 347526 1684
rect 347582 1628 365154 1684
rect 365210 1628 365278 1684
rect 365334 1628 365402 1684
rect 365458 1628 365526 1684
rect 365582 1628 383154 1684
rect 383210 1628 383278 1684
rect 383334 1628 383402 1684
rect 383458 1628 383526 1684
rect 383582 1628 401154 1684
rect 401210 1628 401278 1684
rect 401334 1628 401402 1684
rect 401458 1628 401526 1684
rect 401582 1628 419154 1684
rect 419210 1628 419278 1684
rect 419334 1628 419402 1684
rect 419458 1628 419526 1684
rect 419582 1628 437154 1684
rect 437210 1628 437278 1684
rect 437334 1628 437402 1684
rect 437458 1628 437526 1684
rect 437582 1628 455154 1684
rect 455210 1628 455278 1684
rect 455334 1628 455402 1684
rect 455458 1628 455526 1684
rect 455582 1628 473154 1684
rect 473210 1628 473278 1684
rect 473334 1628 473402 1684
rect 473458 1628 473526 1684
rect 473582 1628 491154 1684
rect 491210 1628 491278 1684
rect 491334 1628 491402 1684
rect 491458 1628 491526 1684
rect 491582 1628 509154 1684
rect 509210 1628 509278 1684
rect 509334 1628 509402 1684
rect 509458 1628 509526 1684
rect 509582 1628 527154 1684
rect 527210 1628 527278 1684
rect 527334 1628 527402 1684
rect 527458 1628 527526 1684
rect 527582 1628 545154 1684
rect 545210 1628 545278 1684
rect 545334 1628 545402 1684
rect 545458 1628 545526 1684
rect 545582 1628 563154 1684
rect 563210 1628 563278 1684
rect 563334 1628 563402 1684
rect 563458 1628 563526 1684
rect 563582 1628 581154 1684
rect 581210 1628 581278 1684
rect 581334 1628 581402 1684
rect 581458 1628 581526 1684
rect 581582 1628 598512 1684
rect 598568 1628 598636 1684
rect 598692 1628 598760 1684
rect 598816 1628 598884 1684
rect 598940 1628 599036 1684
rect 948 1560 599036 1628
rect 948 1504 1044 1560
rect 1100 1504 1168 1560
rect 1224 1504 1292 1560
rect 1348 1504 1416 1560
rect 1472 1504 5154 1560
rect 5210 1504 5278 1560
rect 5334 1504 5402 1560
rect 5458 1504 5526 1560
rect 5582 1504 23154 1560
rect 23210 1504 23278 1560
rect 23334 1504 23402 1560
rect 23458 1504 23526 1560
rect 23582 1504 41154 1560
rect 41210 1504 41278 1560
rect 41334 1504 41402 1560
rect 41458 1504 41526 1560
rect 41582 1504 59154 1560
rect 59210 1504 59278 1560
rect 59334 1504 59402 1560
rect 59458 1504 59526 1560
rect 59582 1504 77154 1560
rect 77210 1504 77278 1560
rect 77334 1504 77402 1560
rect 77458 1504 77526 1560
rect 77582 1504 95154 1560
rect 95210 1504 95278 1560
rect 95334 1504 95402 1560
rect 95458 1504 95526 1560
rect 95582 1504 113154 1560
rect 113210 1504 113278 1560
rect 113334 1504 113402 1560
rect 113458 1504 113526 1560
rect 113582 1504 131154 1560
rect 131210 1504 131278 1560
rect 131334 1504 131402 1560
rect 131458 1504 131526 1560
rect 131582 1504 149154 1560
rect 149210 1504 149278 1560
rect 149334 1504 149402 1560
rect 149458 1504 149526 1560
rect 149582 1504 167154 1560
rect 167210 1504 167278 1560
rect 167334 1504 167402 1560
rect 167458 1504 167526 1560
rect 167582 1504 185154 1560
rect 185210 1504 185278 1560
rect 185334 1504 185402 1560
rect 185458 1504 185526 1560
rect 185582 1504 203154 1560
rect 203210 1504 203278 1560
rect 203334 1504 203402 1560
rect 203458 1504 203526 1560
rect 203582 1504 221154 1560
rect 221210 1504 221278 1560
rect 221334 1504 221402 1560
rect 221458 1504 221526 1560
rect 221582 1504 239154 1560
rect 239210 1504 239278 1560
rect 239334 1504 239402 1560
rect 239458 1504 239526 1560
rect 239582 1504 257154 1560
rect 257210 1504 257278 1560
rect 257334 1504 257402 1560
rect 257458 1504 257526 1560
rect 257582 1504 275154 1560
rect 275210 1504 275278 1560
rect 275334 1504 275402 1560
rect 275458 1504 275526 1560
rect 275582 1504 293154 1560
rect 293210 1504 293278 1560
rect 293334 1504 293402 1560
rect 293458 1504 293526 1560
rect 293582 1504 311154 1560
rect 311210 1504 311278 1560
rect 311334 1504 311402 1560
rect 311458 1504 311526 1560
rect 311582 1504 329154 1560
rect 329210 1504 329278 1560
rect 329334 1504 329402 1560
rect 329458 1504 329526 1560
rect 329582 1504 347154 1560
rect 347210 1504 347278 1560
rect 347334 1504 347402 1560
rect 347458 1504 347526 1560
rect 347582 1504 365154 1560
rect 365210 1504 365278 1560
rect 365334 1504 365402 1560
rect 365458 1504 365526 1560
rect 365582 1504 383154 1560
rect 383210 1504 383278 1560
rect 383334 1504 383402 1560
rect 383458 1504 383526 1560
rect 383582 1504 401154 1560
rect 401210 1504 401278 1560
rect 401334 1504 401402 1560
rect 401458 1504 401526 1560
rect 401582 1504 419154 1560
rect 419210 1504 419278 1560
rect 419334 1504 419402 1560
rect 419458 1504 419526 1560
rect 419582 1504 437154 1560
rect 437210 1504 437278 1560
rect 437334 1504 437402 1560
rect 437458 1504 437526 1560
rect 437582 1504 455154 1560
rect 455210 1504 455278 1560
rect 455334 1504 455402 1560
rect 455458 1504 455526 1560
rect 455582 1504 473154 1560
rect 473210 1504 473278 1560
rect 473334 1504 473402 1560
rect 473458 1504 473526 1560
rect 473582 1504 491154 1560
rect 491210 1504 491278 1560
rect 491334 1504 491402 1560
rect 491458 1504 491526 1560
rect 491582 1504 509154 1560
rect 509210 1504 509278 1560
rect 509334 1504 509402 1560
rect 509458 1504 509526 1560
rect 509582 1504 527154 1560
rect 527210 1504 527278 1560
rect 527334 1504 527402 1560
rect 527458 1504 527526 1560
rect 527582 1504 545154 1560
rect 545210 1504 545278 1560
rect 545334 1504 545402 1560
rect 545458 1504 545526 1560
rect 545582 1504 563154 1560
rect 563210 1504 563278 1560
rect 563334 1504 563402 1560
rect 563458 1504 563526 1560
rect 563582 1504 581154 1560
rect 581210 1504 581278 1560
rect 581334 1504 581402 1560
rect 581458 1504 581526 1560
rect 581582 1504 598512 1560
rect 598568 1504 598636 1560
rect 598692 1504 598760 1560
rect 598816 1504 598884 1560
rect 598940 1504 599036 1560
rect 948 1436 599036 1504
rect 948 1380 1044 1436
rect 1100 1380 1168 1436
rect 1224 1380 1292 1436
rect 1348 1380 1416 1436
rect 1472 1380 5154 1436
rect 5210 1380 5278 1436
rect 5334 1380 5402 1436
rect 5458 1380 5526 1436
rect 5582 1380 23154 1436
rect 23210 1380 23278 1436
rect 23334 1380 23402 1436
rect 23458 1380 23526 1436
rect 23582 1380 41154 1436
rect 41210 1380 41278 1436
rect 41334 1380 41402 1436
rect 41458 1380 41526 1436
rect 41582 1380 59154 1436
rect 59210 1380 59278 1436
rect 59334 1380 59402 1436
rect 59458 1380 59526 1436
rect 59582 1380 77154 1436
rect 77210 1380 77278 1436
rect 77334 1380 77402 1436
rect 77458 1380 77526 1436
rect 77582 1380 95154 1436
rect 95210 1380 95278 1436
rect 95334 1380 95402 1436
rect 95458 1380 95526 1436
rect 95582 1380 113154 1436
rect 113210 1380 113278 1436
rect 113334 1380 113402 1436
rect 113458 1380 113526 1436
rect 113582 1380 131154 1436
rect 131210 1380 131278 1436
rect 131334 1380 131402 1436
rect 131458 1380 131526 1436
rect 131582 1380 149154 1436
rect 149210 1380 149278 1436
rect 149334 1380 149402 1436
rect 149458 1380 149526 1436
rect 149582 1380 167154 1436
rect 167210 1380 167278 1436
rect 167334 1380 167402 1436
rect 167458 1380 167526 1436
rect 167582 1380 185154 1436
rect 185210 1380 185278 1436
rect 185334 1380 185402 1436
rect 185458 1380 185526 1436
rect 185582 1380 203154 1436
rect 203210 1380 203278 1436
rect 203334 1380 203402 1436
rect 203458 1380 203526 1436
rect 203582 1380 221154 1436
rect 221210 1380 221278 1436
rect 221334 1380 221402 1436
rect 221458 1380 221526 1436
rect 221582 1380 239154 1436
rect 239210 1380 239278 1436
rect 239334 1380 239402 1436
rect 239458 1380 239526 1436
rect 239582 1380 257154 1436
rect 257210 1380 257278 1436
rect 257334 1380 257402 1436
rect 257458 1380 257526 1436
rect 257582 1380 275154 1436
rect 275210 1380 275278 1436
rect 275334 1380 275402 1436
rect 275458 1380 275526 1436
rect 275582 1380 293154 1436
rect 293210 1380 293278 1436
rect 293334 1380 293402 1436
rect 293458 1380 293526 1436
rect 293582 1380 311154 1436
rect 311210 1380 311278 1436
rect 311334 1380 311402 1436
rect 311458 1380 311526 1436
rect 311582 1380 329154 1436
rect 329210 1380 329278 1436
rect 329334 1380 329402 1436
rect 329458 1380 329526 1436
rect 329582 1380 347154 1436
rect 347210 1380 347278 1436
rect 347334 1380 347402 1436
rect 347458 1380 347526 1436
rect 347582 1380 365154 1436
rect 365210 1380 365278 1436
rect 365334 1380 365402 1436
rect 365458 1380 365526 1436
rect 365582 1380 383154 1436
rect 383210 1380 383278 1436
rect 383334 1380 383402 1436
rect 383458 1380 383526 1436
rect 383582 1380 401154 1436
rect 401210 1380 401278 1436
rect 401334 1380 401402 1436
rect 401458 1380 401526 1436
rect 401582 1380 419154 1436
rect 419210 1380 419278 1436
rect 419334 1380 419402 1436
rect 419458 1380 419526 1436
rect 419582 1380 437154 1436
rect 437210 1380 437278 1436
rect 437334 1380 437402 1436
rect 437458 1380 437526 1436
rect 437582 1380 455154 1436
rect 455210 1380 455278 1436
rect 455334 1380 455402 1436
rect 455458 1380 455526 1436
rect 455582 1380 473154 1436
rect 473210 1380 473278 1436
rect 473334 1380 473402 1436
rect 473458 1380 473526 1436
rect 473582 1380 491154 1436
rect 491210 1380 491278 1436
rect 491334 1380 491402 1436
rect 491458 1380 491526 1436
rect 491582 1380 509154 1436
rect 509210 1380 509278 1436
rect 509334 1380 509402 1436
rect 509458 1380 509526 1436
rect 509582 1380 527154 1436
rect 527210 1380 527278 1436
rect 527334 1380 527402 1436
rect 527458 1380 527526 1436
rect 527582 1380 545154 1436
rect 545210 1380 545278 1436
rect 545334 1380 545402 1436
rect 545458 1380 545526 1436
rect 545582 1380 563154 1436
rect 563210 1380 563278 1436
rect 563334 1380 563402 1436
rect 563458 1380 563526 1436
rect 563582 1380 581154 1436
rect 581210 1380 581278 1436
rect 581334 1380 581402 1436
rect 581458 1380 581526 1436
rect 581582 1380 598512 1436
rect 598568 1380 598636 1436
rect 598692 1380 598760 1436
rect 598816 1380 598884 1436
rect 598940 1380 599036 1436
rect 948 1284 599036 1380
rect -12 848 599996 944
rect -12 792 84 848
rect 140 792 208 848
rect 264 792 332 848
rect 388 792 456 848
rect 512 792 8874 848
rect 8930 792 8998 848
rect 9054 792 9122 848
rect 9178 792 9246 848
rect 9302 792 26874 848
rect 26930 792 26998 848
rect 27054 792 27122 848
rect 27178 792 27246 848
rect 27302 792 44874 848
rect 44930 792 44998 848
rect 45054 792 45122 848
rect 45178 792 45246 848
rect 45302 792 62874 848
rect 62930 792 62998 848
rect 63054 792 63122 848
rect 63178 792 63246 848
rect 63302 792 80874 848
rect 80930 792 80998 848
rect 81054 792 81122 848
rect 81178 792 81246 848
rect 81302 792 98874 848
rect 98930 792 98998 848
rect 99054 792 99122 848
rect 99178 792 99246 848
rect 99302 792 116874 848
rect 116930 792 116998 848
rect 117054 792 117122 848
rect 117178 792 117246 848
rect 117302 792 134874 848
rect 134930 792 134998 848
rect 135054 792 135122 848
rect 135178 792 135246 848
rect 135302 792 152874 848
rect 152930 792 152998 848
rect 153054 792 153122 848
rect 153178 792 153246 848
rect 153302 792 170874 848
rect 170930 792 170998 848
rect 171054 792 171122 848
rect 171178 792 171246 848
rect 171302 792 188874 848
rect 188930 792 188998 848
rect 189054 792 189122 848
rect 189178 792 189246 848
rect 189302 792 206874 848
rect 206930 792 206998 848
rect 207054 792 207122 848
rect 207178 792 207246 848
rect 207302 792 224874 848
rect 224930 792 224998 848
rect 225054 792 225122 848
rect 225178 792 225246 848
rect 225302 792 242874 848
rect 242930 792 242998 848
rect 243054 792 243122 848
rect 243178 792 243246 848
rect 243302 792 260874 848
rect 260930 792 260998 848
rect 261054 792 261122 848
rect 261178 792 261246 848
rect 261302 792 278874 848
rect 278930 792 278998 848
rect 279054 792 279122 848
rect 279178 792 279246 848
rect 279302 792 296874 848
rect 296930 792 296998 848
rect 297054 792 297122 848
rect 297178 792 297246 848
rect 297302 792 314874 848
rect 314930 792 314998 848
rect 315054 792 315122 848
rect 315178 792 315246 848
rect 315302 792 332874 848
rect 332930 792 332998 848
rect 333054 792 333122 848
rect 333178 792 333246 848
rect 333302 792 350874 848
rect 350930 792 350998 848
rect 351054 792 351122 848
rect 351178 792 351246 848
rect 351302 792 368874 848
rect 368930 792 368998 848
rect 369054 792 369122 848
rect 369178 792 369246 848
rect 369302 792 386874 848
rect 386930 792 386998 848
rect 387054 792 387122 848
rect 387178 792 387246 848
rect 387302 792 404874 848
rect 404930 792 404998 848
rect 405054 792 405122 848
rect 405178 792 405246 848
rect 405302 792 422874 848
rect 422930 792 422998 848
rect 423054 792 423122 848
rect 423178 792 423246 848
rect 423302 792 440874 848
rect 440930 792 440998 848
rect 441054 792 441122 848
rect 441178 792 441246 848
rect 441302 792 458874 848
rect 458930 792 458998 848
rect 459054 792 459122 848
rect 459178 792 459246 848
rect 459302 792 476874 848
rect 476930 792 476998 848
rect 477054 792 477122 848
rect 477178 792 477246 848
rect 477302 792 494874 848
rect 494930 792 494998 848
rect 495054 792 495122 848
rect 495178 792 495246 848
rect 495302 792 512874 848
rect 512930 792 512998 848
rect 513054 792 513122 848
rect 513178 792 513246 848
rect 513302 792 530874 848
rect 530930 792 530998 848
rect 531054 792 531122 848
rect 531178 792 531246 848
rect 531302 792 548874 848
rect 548930 792 548998 848
rect 549054 792 549122 848
rect 549178 792 549246 848
rect 549302 792 566874 848
rect 566930 792 566998 848
rect 567054 792 567122 848
rect 567178 792 567246 848
rect 567302 792 584874 848
rect 584930 792 584998 848
rect 585054 792 585122 848
rect 585178 792 585246 848
rect 585302 792 599472 848
rect 599528 792 599596 848
rect 599652 792 599720 848
rect 599776 792 599844 848
rect 599900 792 599996 848
rect -12 724 599996 792
rect -12 668 84 724
rect 140 668 208 724
rect 264 668 332 724
rect 388 668 456 724
rect 512 668 8874 724
rect 8930 668 8998 724
rect 9054 668 9122 724
rect 9178 668 9246 724
rect 9302 668 26874 724
rect 26930 668 26998 724
rect 27054 668 27122 724
rect 27178 668 27246 724
rect 27302 668 44874 724
rect 44930 668 44998 724
rect 45054 668 45122 724
rect 45178 668 45246 724
rect 45302 668 62874 724
rect 62930 668 62998 724
rect 63054 668 63122 724
rect 63178 668 63246 724
rect 63302 668 80874 724
rect 80930 668 80998 724
rect 81054 668 81122 724
rect 81178 668 81246 724
rect 81302 668 98874 724
rect 98930 668 98998 724
rect 99054 668 99122 724
rect 99178 668 99246 724
rect 99302 668 116874 724
rect 116930 668 116998 724
rect 117054 668 117122 724
rect 117178 668 117246 724
rect 117302 668 134874 724
rect 134930 668 134998 724
rect 135054 668 135122 724
rect 135178 668 135246 724
rect 135302 668 152874 724
rect 152930 668 152998 724
rect 153054 668 153122 724
rect 153178 668 153246 724
rect 153302 668 170874 724
rect 170930 668 170998 724
rect 171054 668 171122 724
rect 171178 668 171246 724
rect 171302 668 188874 724
rect 188930 668 188998 724
rect 189054 668 189122 724
rect 189178 668 189246 724
rect 189302 668 206874 724
rect 206930 668 206998 724
rect 207054 668 207122 724
rect 207178 668 207246 724
rect 207302 668 224874 724
rect 224930 668 224998 724
rect 225054 668 225122 724
rect 225178 668 225246 724
rect 225302 668 242874 724
rect 242930 668 242998 724
rect 243054 668 243122 724
rect 243178 668 243246 724
rect 243302 668 260874 724
rect 260930 668 260998 724
rect 261054 668 261122 724
rect 261178 668 261246 724
rect 261302 668 278874 724
rect 278930 668 278998 724
rect 279054 668 279122 724
rect 279178 668 279246 724
rect 279302 668 296874 724
rect 296930 668 296998 724
rect 297054 668 297122 724
rect 297178 668 297246 724
rect 297302 668 314874 724
rect 314930 668 314998 724
rect 315054 668 315122 724
rect 315178 668 315246 724
rect 315302 668 332874 724
rect 332930 668 332998 724
rect 333054 668 333122 724
rect 333178 668 333246 724
rect 333302 668 350874 724
rect 350930 668 350998 724
rect 351054 668 351122 724
rect 351178 668 351246 724
rect 351302 668 368874 724
rect 368930 668 368998 724
rect 369054 668 369122 724
rect 369178 668 369246 724
rect 369302 668 386874 724
rect 386930 668 386998 724
rect 387054 668 387122 724
rect 387178 668 387246 724
rect 387302 668 404874 724
rect 404930 668 404998 724
rect 405054 668 405122 724
rect 405178 668 405246 724
rect 405302 668 422874 724
rect 422930 668 422998 724
rect 423054 668 423122 724
rect 423178 668 423246 724
rect 423302 668 440874 724
rect 440930 668 440998 724
rect 441054 668 441122 724
rect 441178 668 441246 724
rect 441302 668 458874 724
rect 458930 668 458998 724
rect 459054 668 459122 724
rect 459178 668 459246 724
rect 459302 668 476874 724
rect 476930 668 476998 724
rect 477054 668 477122 724
rect 477178 668 477246 724
rect 477302 668 494874 724
rect 494930 668 494998 724
rect 495054 668 495122 724
rect 495178 668 495246 724
rect 495302 668 512874 724
rect 512930 668 512998 724
rect 513054 668 513122 724
rect 513178 668 513246 724
rect 513302 668 530874 724
rect 530930 668 530998 724
rect 531054 668 531122 724
rect 531178 668 531246 724
rect 531302 668 548874 724
rect 548930 668 548998 724
rect 549054 668 549122 724
rect 549178 668 549246 724
rect 549302 668 566874 724
rect 566930 668 566998 724
rect 567054 668 567122 724
rect 567178 668 567246 724
rect 567302 668 584874 724
rect 584930 668 584998 724
rect 585054 668 585122 724
rect 585178 668 585246 724
rect 585302 668 599472 724
rect 599528 668 599596 724
rect 599652 668 599720 724
rect 599776 668 599844 724
rect 599900 668 599996 724
rect -12 600 599996 668
rect -12 544 84 600
rect 140 544 208 600
rect 264 544 332 600
rect 388 544 456 600
rect 512 544 8874 600
rect 8930 544 8998 600
rect 9054 544 9122 600
rect 9178 544 9246 600
rect 9302 544 26874 600
rect 26930 544 26998 600
rect 27054 544 27122 600
rect 27178 544 27246 600
rect 27302 544 44874 600
rect 44930 544 44998 600
rect 45054 544 45122 600
rect 45178 544 45246 600
rect 45302 544 62874 600
rect 62930 544 62998 600
rect 63054 544 63122 600
rect 63178 544 63246 600
rect 63302 544 80874 600
rect 80930 544 80998 600
rect 81054 544 81122 600
rect 81178 544 81246 600
rect 81302 544 98874 600
rect 98930 544 98998 600
rect 99054 544 99122 600
rect 99178 544 99246 600
rect 99302 544 116874 600
rect 116930 544 116998 600
rect 117054 544 117122 600
rect 117178 544 117246 600
rect 117302 544 134874 600
rect 134930 544 134998 600
rect 135054 544 135122 600
rect 135178 544 135246 600
rect 135302 544 152874 600
rect 152930 544 152998 600
rect 153054 544 153122 600
rect 153178 544 153246 600
rect 153302 544 170874 600
rect 170930 544 170998 600
rect 171054 544 171122 600
rect 171178 544 171246 600
rect 171302 544 188874 600
rect 188930 544 188998 600
rect 189054 544 189122 600
rect 189178 544 189246 600
rect 189302 544 206874 600
rect 206930 544 206998 600
rect 207054 544 207122 600
rect 207178 544 207246 600
rect 207302 544 224874 600
rect 224930 544 224998 600
rect 225054 544 225122 600
rect 225178 544 225246 600
rect 225302 544 242874 600
rect 242930 544 242998 600
rect 243054 544 243122 600
rect 243178 544 243246 600
rect 243302 544 260874 600
rect 260930 544 260998 600
rect 261054 544 261122 600
rect 261178 544 261246 600
rect 261302 544 278874 600
rect 278930 544 278998 600
rect 279054 544 279122 600
rect 279178 544 279246 600
rect 279302 544 296874 600
rect 296930 544 296998 600
rect 297054 544 297122 600
rect 297178 544 297246 600
rect 297302 544 314874 600
rect 314930 544 314998 600
rect 315054 544 315122 600
rect 315178 544 315246 600
rect 315302 544 332874 600
rect 332930 544 332998 600
rect 333054 544 333122 600
rect 333178 544 333246 600
rect 333302 544 350874 600
rect 350930 544 350998 600
rect 351054 544 351122 600
rect 351178 544 351246 600
rect 351302 544 368874 600
rect 368930 544 368998 600
rect 369054 544 369122 600
rect 369178 544 369246 600
rect 369302 544 386874 600
rect 386930 544 386998 600
rect 387054 544 387122 600
rect 387178 544 387246 600
rect 387302 544 404874 600
rect 404930 544 404998 600
rect 405054 544 405122 600
rect 405178 544 405246 600
rect 405302 544 422874 600
rect 422930 544 422998 600
rect 423054 544 423122 600
rect 423178 544 423246 600
rect 423302 544 440874 600
rect 440930 544 440998 600
rect 441054 544 441122 600
rect 441178 544 441246 600
rect 441302 544 458874 600
rect 458930 544 458998 600
rect 459054 544 459122 600
rect 459178 544 459246 600
rect 459302 544 476874 600
rect 476930 544 476998 600
rect 477054 544 477122 600
rect 477178 544 477246 600
rect 477302 544 494874 600
rect 494930 544 494998 600
rect 495054 544 495122 600
rect 495178 544 495246 600
rect 495302 544 512874 600
rect 512930 544 512998 600
rect 513054 544 513122 600
rect 513178 544 513246 600
rect 513302 544 530874 600
rect 530930 544 530998 600
rect 531054 544 531122 600
rect 531178 544 531246 600
rect 531302 544 548874 600
rect 548930 544 548998 600
rect 549054 544 549122 600
rect 549178 544 549246 600
rect 549302 544 566874 600
rect 566930 544 566998 600
rect 567054 544 567122 600
rect 567178 544 567246 600
rect 567302 544 584874 600
rect 584930 544 584998 600
rect 585054 544 585122 600
rect 585178 544 585246 600
rect 585302 544 599472 600
rect 599528 544 599596 600
rect 599652 544 599720 600
rect 599776 544 599844 600
rect 599900 544 599996 600
rect -12 476 599996 544
rect -12 420 84 476
rect 140 420 208 476
rect 264 420 332 476
rect 388 420 456 476
rect 512 420 8874 476
rect 8930 420 8998 476
rect 9054 420 9122 476
rect 9178 420 9246 476
rect 9302 420 26874 476
rect 26930 420 26998 476
rect 27054 420 27122 476
rect 27178 420 27246 476
rect 27302 420 44874 476
rect 44930 420 44998 476
rect 45054 420 45122 476
rect 45178 420 45246 476
rect 45302 420 62874 476
rect 62930 420 62998 476
rect 63054 420 63122 476
rect 63178 420 63246 476
rect 63302 420 80874 476
rect 80930 420 80998 476
rect 81054 420 81122 476
rect 81178 420 81246 476
rect 81302 420 98874 476
rect 98930 420 98998 476
rect 99054 420 99122 476
rect 99178 420 99246 476
rect 99302 420 116874 476
rect 116930 420 116998 476
rect 117054 420 117122 476
rect 117178 420 117246 476
rect 117302 420 134874 476
rect 134930 420 134998 476
rect 135054 420 135122 476
rect 135178 420 135246 476
rect 135302 420 152874 476
rect 152930 420 152998 476
rect 153054 420 153122 476
rect 153178 420 153246 476
rect 153302 420 170874 476
rect 170930 420 170998 476
rect 171054 420 171122 476
rect 171178 420 171246 476
rect 171302 420 188874 476
rect 188930 420 188998 476
rect 189054 420 189122 476
rect 189178 420 189246 476
rect 189302 420 206874 476
rect 206930 420 206998 476
rect 207054 420 207122 476
rect 207178 420 207246 476
rect 207302 420 224874 476
rect 224930 420 224998 476
rect 225054 420 225122 476
rect 225178 420 225246 476
rect 225302 420 242874 476
rect 242930 420 242998 476
rect 243054 420 243122 476
rect 243178 420 243246 476
rect 243302 420 260874 476
rect 260930 420 260998 476
rect 261054 420 261122 476
rect 261178 420 261246 476
rect 261302 420 278874 476
rect 278930 420 278998 476
rect 279054 420 279122 476
rect 279178 420 279246 476
rect 279302 420 296874 476
rect 296930 420 296998 476
rect 297054 420 297122 476
rect 297178 420 297246 476
rect 297302 420 314874 476
rect 314930 420 314998 476
rect 315054 420 315122 476
rect 315178 420 315246 476
rect 315302 420 332874 476
rect 332930 420 332998 476
rect 333054 420 333122 476
rect 333178 420 333246 476
rect 333302 420 350874 476
rect 350930 420 350998 476
rect 351054 420 351122 476
rect 351178 420 351246 476
rect 351302 420 368874 476
rect 368930 420 368998 476
rect 369054 420 369122 476
rect 369178 420 369246 476
rect 369302 420 386874 476
rect 386930 420 386998 476
rect 387054 420 387122 476
rect 387178 420 387246 476
rect 387302 420 404874 476
rect 404930 420 404998 476
rect 405054 420 405122 476
rect 405178 420 405246 476
rect 405302 420 422874 476
rect 422930 420 422998 476
rect 423054 420 423122 476
rect 423178 420 423246 476
rect 423302 420 440874 476
rect 440930 420 440998 476
rect 441054 420 441122 476
rect 441178 420 441246 476
rect 441302 420 458874 476
rect 458930 420 458998 476
rect 459054 420 459122 476
rect 459178 420 459246 476
rect 459302 420 476874 476
rect 476930 420 476998 476
rect 477054 420 477122 476
rect 477178 420 477246 476
rect 477302 420 494874 476
rect 494930 420 494998 476
rect 495054 420 495122 476
rect 495178 420 495246 476
rect 495302 420 512874 476
rect 512930 420 512998 476
rect 513054 420 513122 476
rect 513178 420 513246 476
rect 513302 420 530874 476
rect 530930 420 530998 476
rect 531054 420 531122 476
rect 531178 420 531246 476
rect 531302 420 548874 476
rect 548930 420 548998 476
rect 549054 420 549122 476
rect 549178 420 549246 476
rect 549302 420 566874 476
rect 566930 420 566998 476
rect 567054 420 567122 476
rect 567178 420 567246 476
rect 567302 420 584874 476
rect 584930 420 584998 476
rect 585054 420 585122 476
rect 585178 420 585246 476
rect 585302 420 599472 476
rect 599528 420 599596 476
rect 599652 420 599720 476
rect 599776 420 599844 476
rect 599900 420 599996 476
rect -12 324 599996 420
<< labels >>
flabel metal3 s 599520 6664 600960 6888 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 599520 406504 600960 406728 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 599520 446488 600960 446712 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 599520 486472 600960 486696 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 599520 526456 600960 526680 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 599520 566440 600960 566664 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 588168 599520 588392 600960 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 521640 599520 521864 600960 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 455112 599520 455336 600960 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 388584 599520 388808 600960 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 322056 599520 322280 600960 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 599520 46648 600960 46872 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 255528 599520 255752 600960 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 189000 599520 189224 600960 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 122472 599520 122696 600960 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55944 599520 56168 600960 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 591416 480 591640 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 548744 480 548968 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 506072 480 506296 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 463400 480 463624 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 420728 480 420952 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 378056 480 378280 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 599520 86632 600960 86856 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 335384 480 335608 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 292712 480 292936 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 250040 480 250264 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 207368 480 207592 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 164696 480 164920 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 122024 480 122248 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79352 480 79576 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36680 480 36904 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 599520 126616 600960 126840 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 599520 166600 600960 166824 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 599520 206584 600960 206808 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 599520 246568 600960 246792 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 599520 286552 600960 286776 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 599520 326536 600960 326760 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 599520 366520 600960 366744 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 599520 33320 600960 33544 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 599520 433160 600960 433384 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 599520 473144 600960 473368 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 599520 513128 600960 513352 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 599520 553112 600960 553336 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 599520 593096 600960 593320 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 543816 599520 544040 600960 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 477288 599520 477512 600960 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 410760 599520 410984 600960 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 344232 599520 344456 600960 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 277704 599520 277928 600960 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 599520 73304 600960 73528 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 211176 599520 211400 600960 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 144648 599520 144872 600960 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 78120 599520 78344 600960 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11592 599520 11816 600960 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 562968 480 563192 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 520296 480 520520 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 477624 480 477848 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 434952 480 435176 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 392280 480 392504 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 349608 480 349832 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 599520 113288 600960 113512 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 306936 480 307160 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 264264 480 264488 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 221592 480 221816 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 178920 480 179144 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 136248 480 136472 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93576 480 93800 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8232 480 8456 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 599520 153272 600960 153496 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 599520 193256 600960 193480 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 599520 233240 600960 233464 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 599520 273224 600960 273448 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 599520 313208 600960 313432 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 599520 353192 600960 353416 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 599520 393176 600960 393400 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 599520 19992 600960 20216 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 599520 419832 600960 420056 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 599520 459816 600960 460040 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 599520 499800 600960 500024 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 599520 539784 600960 540008 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 599520 579768 600960 579992 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 565992 599520 566216 600960 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 499464 599520 499688 600960 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 432936 599520 433160 600960 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 366408 599520 366632 600960 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 299880 599520 300104 600960 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 599520 59976 600960 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 233352 599520 233576 600960 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 166824 599520 167048 600960 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 100296 599520 100520 600960 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33768 599520 33992 600960 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 577192 480 577416 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 534520 480 534744 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 491848 480 492072 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 449176 480 449400 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 406504 480 406728 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 363832 480 364056 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 599520 99960 600960 100184 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 321160 480 321384 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 278488 480 278712 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 235816 480 236040 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 193144 480 193368 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 150472 480 150696 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107800 480 108024 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65128 480 65352 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22456 480 22680 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 599520 139944 600960 140168 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 599520 179928 600960 180152 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 599520 219912 600960 220136 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 599520 259896 600960 260120 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 599520 299880 600960 300104 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 599520 339864 600960 340088 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 599520 379848 600960 380072 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 586376 -960 586600 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s 948 1284 1568 598476 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 948 1284 599036 1904 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 948 597856 599036 598476 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 598416 1284 599036 598476 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5058 324 5678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 23058 324 23678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 41058 324 41678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 59058 324 59678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 77058 324 77678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 95058 324 95678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 113058 324 113678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 131058 324 131678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 149058 324 149678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 167058 324 167678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 185058 324 185678 169874 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 185058 287294 185678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 203058 324 203678 169874 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 203058 287294 203678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 221058 324 221678 169874 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 221058 287294 221678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 239058 324 239678 169874 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 239058 287294 239678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 257058 324 257678 169874 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 257058 287294 257678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 275058 324 275678 170020 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 275058 287932 275678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 293058 324 293678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 311058 324 311678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 329058 324 329678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 347058 324 347678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 365058 324 365678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 383058 324 383678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 401058 324 401678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 419058 324 419678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 437058 324 437678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 455058 324 455678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 473058 324 473678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 491058 324 491678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 509058 324 509678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527058 324 527678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 545058 324 545678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 563058 324 563678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 581058 324 581678 599436 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 5394 599996 6014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 23394 599996 24014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 41394 599996 42014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 59394 599996 60014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 77394 599996 78014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 95394 599996 96014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 113394 599996 114014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 131394 599996 132014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 149394 599996 150014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 167394 599996 168014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 185394 599996 186014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 203394 599996 204014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 221394 599996 222014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 239394 599996 240014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 257394 599996 258014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 275394 599996 276014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 293394 599996 294014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 311394 599996 312014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 329394 599996 330014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 347394 599996 348014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 365394 599996 366014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 383394 599996 384014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 401394 599996 402014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 419394 599996 420014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 437394 599996 438014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 455394 599996 456014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 473394 599996 474014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 491394 599996 492014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 509394 599996 510014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 527394 599996 528014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 545394 599996 546014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 563394 599996 564014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -12 581394 599996 582014 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -12 324 608 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 324 599996 944 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 598816 599996 599436 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 599376 324 599996 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 8778 324 9398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 26778 324 27398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 44778 324 45398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 62778 324 63398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 80778 324 81398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 98778 324 99398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 116778 324 117398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 134778 324 135398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 152778 324 153398 170020 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 152778 287932 153398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 170778 324 171398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188778 324 189398 169874 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 188778 287294 189398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 206778 324 207398 169874 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 206778 287294 207398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224778 324 225398 169874 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224778 287294 225398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 242778 324 243398 169874 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 242778 287294 243398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 260778 324 261398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 278778 324 279398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 296778 324 297398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 314778 324 315398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 332778 324 333398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 350778 324 351398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 368778 324 369398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 386778 324 387398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 404778 324 405398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 422778 324 423398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 440778 324 441398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 458778 324 459398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 476778 324 477398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 494778 324 495398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 512778 324 513398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 530778 324 531398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 548778 324 549398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 566778 324 567398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 584778 324 585398 599436 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 11394 599996 12014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 29394 599996 30014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 47394 599996 48014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 65394 599996 66014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 83394 599996 84014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 101394 599996 102014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 119394 599996 120014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 137394 599996 138014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 155394 599996 156014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 173394 599996 174014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 191394 599996 192014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 209394 599996 210014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 227394 599996 228014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 245394 599996 246014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 263394 599996 264014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 281394 599996 282014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 299394 599996 300014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 317394 599996 318014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 335394 599996 336014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 353394 599996 354014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 371394 599996 372014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 389394 599996 390014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 407394 599996 408014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 425394 599996 426014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 443394 599996 444014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 461394 599996 462014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 479394 599996 480014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 497394 599996 498014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 515394 599996 516014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 533394 599996 534014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 551394 599996 552014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 569394 599996 570014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -12 587394 599996 588014 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel metal2 454328 599592 454328 599592 0 io_in[17]
rlabel metal2 121688 599592 121688 599592 0 io_in[22]
rlabel metal3 3990 591416 3990 591416 0 io_in[24]
rlabel metal3 392 548184 392 548184 0 io_in[25]
rlabel metal3 392 462672 392 462672 0 io_in[27]
rlabel metal3 392 420336 392 420336 0 io_in[28]
rlabel metal3 392 334824 392 334824 0 io_in[30]
rlabel metal3 392 292488 392 292488 0 io_in[31]
rlabel metal3 392 249312 392 249312 0 io_in[32]
rlabel metal3 392 206976 392 206976 0 io_in[33]
rlabel metal3 392 121464 392 121464 0 io_in[35]
rlabel metal3 392 35952 392 35952 0 io_in[37]
rlabel metal2 595560 217168 595560 217168 0 io_in[3]
rlabel metal2 78344 597562 78344 597562 0 io_oeb[22]
rlabel metal2 10808 599592 10808 599592 0 io_oeb[23]
rlabel metal3 392 519680 392 519680 0 io_oeb[25]
rlabel metal3 2422 477624 2422 477624 0 io_oeb[26]
rlabel metal3 2366 434952 2366 434952 0 io_oeb[27]
rlabel metal3 392 391832 392 391832 0 io_oeb[28]
rlabel metal3 2646 306936 2646 306936 0 io_oeb[30]
rlabel metal3 392 263984 392 263984 0 io_oeb[31]
rlabel metal3 3990 221704 3990 221704 0 io_oeb[32]
rlabel metal3 392 178472 392 178472 0 io_oeb[33]
rlabel metal3 392 92960 392 92960 0 io_oeb[35]
rlabel metal3 392 50624 392 50624 0 io_oeb[36]
rlabel metal3 5670 8344 5670 8344 0 io_oeb[37]
rlabel metal2 595672 233016 595672 233016 0 io_oeb[3]
rlabel metal2 596120 302344 596120 302344 0 io_oeb[7]
rlabel metal3 599592 352968 599592 352968 0 io_oeb[8]
rlabel metal3 599592 539504 599592 539504 0 io_out[13]
rlabel metal2 499184 599592 499184 599592 0 io_out[16]
rlabel metal2 166544 599592 166544 599592 0 io_out[21]
rlabel metal3 2310 534520 2310 534520 0 io_out[25]
rlabel metal3 392 491176 392 491176 0 io_out[26]
rlabel metal3 392 448840 392 448840 0 io_out[27]
rlabel metal3 2534 363832 2534 363832 0 io_out[29]
rlabel metal3 392 277816 392 277816 0 io_out[31]
rlabel metal3 392 235480 392 235480 0 io_out[32]
rlabel metal3 2310 65352 2310 65352 0 io_out[36]
rlabel metal3 392 22120 392 22120 0 io_out[37]
rlabel metal3 599592 139664 599592 139664 0 io_out[3]
rlabel metal2 596008 287168 596008 287168 0 io_out[6]
rlabel metal2 282912 392 282912 392 0 la_data_in[12]
rlabel metal2 346248 392 346248 392 0 la_data_in[23]
rlabel metal2 351624 392 351624 392 0 la_data_in[24]
rlabel metal2 369320 1470 369320 1470 0 la_data_in[27]
rlabel metal2 374920 280 374920 280 0 la_data_in[28]
rlabel metal2 380184 392 380184 392 0 la_data_in[29]
rlabel metal2 225848 392 225848 392 0 la_data_in[2]
rlabel metal2 391776 392 391776 392 0 la_data_in[31]
rlabel metal2 397152 392 397152 392 0 la_data_in[32]
rlabel metal2 403368 392 403368 392 0 la_data_in[33]
rlabel metal2 408744 392 408744 392 0 la_data_in[34]
rlabel metal2 425712 392 425712 392 0 la_data_in[37]
rlabel metal2 431928 392 431928 392 0 la_data_in[38]
rlabel metal2 448896 392 448896 392 0 la_data_in[41]
rlabel metal2 454272 392 454272 392 0 la_data_in[42]
rlabel metal2 460488 392 460488 392 0 la_data_in[43]
rlabel metal2 465864 392 465864 392 0 la_data_in[44]
rlabel metal2 477456 392 477456 392 0 la_data_in[46]
rlabel metal2 482832 392 482832 392 0 la_data_in[47]
rlabel metal2 237944 1638 237944 1638 0 la_data_in[4]
rlabel metal2 517608 392 517608 392 0 la_data_in[53]
rlabel metal2 522984 392 522984 392 0 la_data_in[54]
rlabel metal2 534576 392 534576 392 0 la_data_in[56]
rlabel metal2 539952 392 539952 392 0 la_data_in[57]
rlabel metal2 546168 392 546168 392 0 la_data_in[58]
rlabel metal2 551544 392 551544 392 0 la_data_in[59]
rlabel metal2 574728 392 574728 392 0 la_data_in[63]
rlabel metal2 265944 392 265944 392 0 la_data_in[9]
rlabel metal2 279384 392 279384 392 0 la_data_out[11]
rlabel metal2 290920 392 290920 392 0 la_data_out[13]
rlabel metal2 296296 392 296296 392 0 la_data_out[14]
rlabel metal2 307888 392 307888 392 0 la_data_out[16]
rlabel metal2 353416 392 353416 392 0 la_data_out[24]
rlabel metal2 376600 392 376600 392 0 la_data_out[28]
rlabel metal2 381976 392 381976 392 0 la_data_out[29]
rlabel metal2 393568 392 393568 392 0 la_data_out[31]
rlabel metal2 422128 392 422128 392 0 la_data_out[36]
rlabel metal2 433720 392 433720 392 0 la_data_out[38]
rlabel metal2 450688 392 450688 392 0 la_data_out[41]
rlabel metal2 462280 392 462280 392 0 la_data_out[43]
rlabel metal2 467656 392 467656 392 0 la_data_out[44]
rlabel metal2 496216 392 496216 392 0 la_data_out[49]
rlabel metal2 239176 392 239176 392 0 la_data_out[4]
rlabel metal2 519400 392 519400 392 0 la_data_out[53]
rlabel metal2 524776 392 524776 392 0 la_data_out[54]
rlabel metal2 536368 392 536368 392 0 la_data_out[56]
rlabel metal2 553336 392 553336 392 0 la_data_out[59]
rlabel metal2 262416 392 262416 392 0 la_data_out[8]
rlabel metal2 218624 392 218624 392 0 la_oenb[0]
rlabel metal2 275744 392 275744 392 0 la_oenb[10]
rlabel metal2 281120 392 281120 392 0 la_oenb[11]
rlabel metal2 292712 392 292712 392 0 la_oenb[13]
rlabel metal2 298088 392 298088 392 0 la_oenb[14]
rlabel metal2 304304 392 304304 392 0 la_oenb[15]
rlabel metal2 309680 392 309680 392 0 la_oenb[16]
rlabel metal2 326648 392 326648 392 0 la_oenb[19]
rlabel metal2 355208 392 355208 392 0 la_oenb[24]
rlabel metal2 378392 392 378392 392 0 la_oenb[28]
rlabel metal2 389984 392 389984 392 0 la_oenb[30]
rlabel metal2 395360 392 395360 392 0 la_oenb[31]
rlabel metal2 406952 392 406952 392 0 la_oenb[33]
rlabel metal2 412328 392 412328 392 0 la_oenb[34]
rlabel metal2 423920 392 423920 392 0 la_oenb[36]
rlabel metal2 235592 392 235592 392 0 la_oenb[3]
rlabel metal2 447104 392 447104 392 0 la_oenb[40]
rlabel metal2 452480 392 452480 392 0 la_oenb[41]
rlabel metal2 464072 392 464072 392 0 la_oenb[43]
rlabel metal2 469448 392 469448 392 0 la_oenb[44]
rlabel metal2 241024 392 241024 392 0 la_oenb[4]
rlabel metal2 521192 392 521192 392 0 la_oenb[53]
rlabel metal2 538160 392 538160 392 0 la_oenb[56]
rlabel metal2 549752 392 549752 392 0 la_oenb[58]
rlabel metal2 555128 392 555128 392 0 la_oenb[59]
rlabel metal2 583688 392 583688 392 0 user_irq[1]
rlabel metal2 24080 392 24080 392 0 wbs_adr_i[0]
rlabel metal2 95368 2254 95368 2254 0 wbs_adr_i[11]
rlabel metal2 106176 392 106176 392 0 wbs_adr_i[13]
rlabel metal2 111552 392 111552 392 0 wbs_adr_i[14]
rlabel metal2 118216 2254 118216 2254 0 wbs_adr_i[15]
rlabel metal2 123144 392 123144 392 0 wbs_adr_i[16]
rlabel metal2 135352 2310 135352 2310 0 wbs_adr_i[18]
rlabel metal2 140112 392 140112 392 0 wbs_adr_i[19]
rlabel metal2 32088 392 32088 392 0 wbs_adr_i[1]
rlabel metal2 146328 392 146328 392 0 wbs_adr_i[20]
rlabel metal2 163464 392 163464 392 0 wbs_adr_i[23]
rlabel metal2 40152 2254 40152 2254 0 wbs_adr_i[2]
rlabel metal2 54432 392 54432 392 0 wbs_adr_i[4]
rlabel metal2 60648 392 60648 392 0 wbs_adr_i[5]
rlabel metal2 82992 392 82992 392 0 wbs_adr_i[9]
rlabel metal2 25872 392 25872 392 0 wbs_dat_i[0]
rlabel metal2 91560 2254 91560 2254 0 wbs_dat_i[10]
rlabel metal2 96376 392 96376 392 0 wbs_dat_i[11]
rlabel metal2 107968 392 107968 392 0 wbs_dat_i[13]
rlabel metal2 125104 392 125104 392 0 wbs_dat_i[16]
rlabel metal2 131544 2254 131544 2254 0 wbs_dat_i[17]
rlabel metal2 33880 392 33880 392 0 wbs_dat_i[1]
rlabel metal2 165088 392 165088 392 0 wbs_dat_i[23]
rlabel metal2 176680 392 176680 392 0 wbs_dat_i[25]
rlabel metal2 194152 2254 194152 2254 0 wbs_dat_i[28]
rlabel metal2 41944 2310 41944 2310 0 wbs_dat_i[2]
rlabel metal2 205240 392 205240 392 0 wbs_dat_i[30]
rlabel metal2 210672 392 210672 392 0 wbs_dat_i[31]
rlabel metal2 49056 392 49056 392 0 wbs_dat_i[3]
rlabel metal2 67816 392 67816 392 0 wbs_dat_i[6]
rlabel metal2 80136 2198 80136 2198 0 wbs_dat_i[8]
rlabel metal2 92792 392 92792 392 0 wbs_dat_o[10]
rlabel metal2 104384 392 104384 392 0 wbs_dat_o[12]
rlabel metal2 109760 392 109760 392 0 wbs_dat_o[13]
rlabel metal2 121352 392 121352 392 0 wbs_dat_o[15]
rlabel metal2 139160 2310 139160 2310 0 wbs_dat_o[18]
rlabel metal2 35672 392 35672 392 0 wbs_dat_o[1]
rlabel metal2 149912 392 149912 392 0 wbs_dat_o[20]
rlabel metal2 155288 392 155288 392 0 wbs_dat_o[21]
rlabel metal2 161504 392 161504 392 0 wbs_dat_o[22]
rlabel metal2 167720 2310 167720 2310 0 wbs_dat_o[23]
rlabel metal2 178528 392 178528 392 0 wbs_dat_o[25]
rlabel metal2 183904 392 183904 392 0 wbs_dat_o[26]
rlabel metal2 195440 392 195440 392 0 wbs_dat_o[28]
rlabel metal2 50848 392 50848 392 0 wbs_dat_o[3]
rlabel metal2 59192 2254 59192 2254 0 wbs_dat_o[4]
rlabel metal2 70504 2254 70504 2254 0 wbs_dat_o[6]
rlabel metal2 82040 2254 82040 2254 0 wbs_dat_o[8]
rlabel metal2 37464 392 37464 392 0 wbs_sel_i[1]
rlabel metal2 45864 2254 45864 2254 0 wbs_sel_i[2]
rlabel metal2 23016 2310 23016 2310 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 600000 600000
<< end >>
