magic
tech gf180mcuC
magscale 1 5
timestamp 1670230241
<< obsm1 >>
rect 672 1538 39312 18454
<< metal2 >>
rect 2520 19600 2576 20000
rect 7504 19600 7560 20000
rect 12488 19600 12544 20000
rect 17472 19600 17528 20000
rect 22456 19600 22512 20000
rect 27440 19600 27496 20000
rect 32424 19600 32480 20000
rect 37408 19600 37464 20000
rect 840 0 896 400
rect 2072 0 2128 400
rect 3304 0 3360 400
rect 4536 0 4592 400
rect 5768 0 5824 400
rect 7000 0 7056 400
rect 8232 0 8288 400
rect 9464 0 9520 400
rect 10696 0 10752 400
rect 11928 0 11984 400
rect 13160 0 13216 400
rect 14392 0 14448 400
rect 15624 0 15680 400
rect 16856 0 16912 400
rect 18088 0 18144 400
rect 19320 0 19376 400
rect 20552 0 20608 400
rect 21784 0 21840 400
rect 23016 0 23072 400
rect 24248 0 24304 400
rect 25480 0 25536 400
rect 26712 0 26768 400
rect 27944 0 28000 400
rect 29176 0 29232 400
rect 30408 0 30464 400
rect 31640 0 31696 400
rect 32872 0 32928 400
rect 34104 0 34160 400
rect 35336 0 35392 400
rect 36568 0 36624 400
rect 37800 0 37856 400
rect 39032 0 39088 400
<< obsm2 >>
rect 854 19570 2490 19642
rect 2606 19570 7474 19642
rect 7590 19570 12458 19642
rect 12574 19570 17442 19642
rect 17558 19570 22426 19642
rect 22542 19570 27410 19642
rect 27526 19570 32394 19642
rect 32510 19570 37378 19642
rect 37494 19570 39130 19642
rect 854 430 39130 19570
rect 926 350 2042 430
rect 2158 350 3274 430
rect 3390 350 4506 430
rect 4622 350 5738 430
rect 5854 350 6970 430
rect 7086 350 8202 430
rect 8318 350 9434 430
rect 9550 350 10666 430
rect 10782 350 11898 430
rect 12014 350 13130 430
rect 13246 350 14362 430
rect 14478 350 15594 430
rect 15710 350 16826 430
rect 16942 350 18058 430
rect 18174 350 19290 430
rect 19406 350 20522 430
rect 20638 350 21754 430
rect 21870 350 22986 430
rect 23102 350 24218 430
rect 24334 350 25450 430
rect 25566 350 26682 430
rect 26798 350 27914 430
rect 28030 350 29146 430
rect 29262 350 30378 430
rect 30494 350 31610 430
rect 31726 350 32842 430
rect 32958 350 34074 430
rect 34190 350 35306 430
rect 35422 350 36538 430
rect 36654 350 37770 430
rect 37886 350 39002 430
rect 39118 350 39130 430
<< obsm3 >>
rect 1185 1554 39135 18438
<< metal4 >>
rect 2054 1538 2554 18454
rect 4554 1538 5054 18454
rect 7054 1538 7554 18454
rect 9554 1538 10054 18454
rect 12054 1538 12554 18454
rect 14554 1538 15054 18454
rect 17054 1538 17554 18454
rect 19554 1538 20054 18454
rect 22054 1538 22554 18454
rect 24554 1538 25054 18454
rect 27054 1538 27554 18454
rect 29554 1538 30054 18454
rect 32054 1538 32554 18454
rect 34554 1538 35054 18454
rect 37054 1538 37554 18454
<< obsm4 >>
rect 31990 2193 32024 4471
rect 32584 2193 34524 4471
rect 35084 2193 36946 4471
<< labels >>
rlabel metal2 s 37408 19600 37464 20000 6 cap_series_gygyn
port 1 nsew signal bidirectional
rlabel metal2 s 32424 19600 32480 20000 6 cap_series_gygyp
port 2 nsew signal bidirectional
rlabel metal2 s 27440 19600 27496 20000 6 cap_series_gyn
port 3 nsew signal bidirectional
rlabel metal2 s 22456 19600 22512 20000 6 cap_series_gyp
port 4 nsew signal bidirectional
rlabel metal2 s 17472 19600 17528 20000 6 cap_shunt_gyn
port 5 nsew signal bidirectional
rlabel metal2 s 12488 19600 12544 20000 6 cap_shunt_gyp
port 6 nsew signal bidirectional
rlabel metal2 s 7504 19600 7560 20000 6 cap_shunt_n
port 7 nsew signal bidirectional
rlabel metal2 s 2520 19600 2576 20000 6 cap_shunt_p
port 8 nsew signal bidirectional
rlabel metal2 s 14392 0 14448 400 6 tune_series_gy[0]
port 9 nsew signal input
rlabel metal2 s 15624 0 15680 400 6 tune_series_gy[1]
port 10 nsew signal input
rlabel metal2 s 16856 0 16912 400 6 tune_series_gy[2]
port 11 nsew signal input
rlabel metal2 s 18088 0 18144 400 6 tune_series_gy[3]
port 12 nsew signal input
rlabel metal2 s 19320 0 19376 400 6 tune_series_gy[4]
port 13 nsew signal input
rlabel metal2 s 20552 0 20608 400 6 tune_series_gy[5]
port 14 nsew signal input
rlabel metal2 s 21784 0 21840 400 6 tune_series_gy[6]
port 15 nsew signal input
rlabel metal2 s 23016 0 23072 400 6 tune_series_gy[7]
port 16 nsew signal input
rlabel metal2 s 24248 0 24304 400 6 tune_series_gygy[0]
port 17 nsew signal input
rlabel metal2 s 25480 0 25536 400 6 tune_series_gygy[1]
port 18 nsew signal input
rlabel metal2 s 26712 0 26768 400 6 tune_series_gygy[2]
port 19 nsew signal input
rlabel metal2 s 27944 0 28000 400 6 tune_series_gygy[3]
port 20 nsew signal input
rlabel metal2 s 29176 0 29232 400 6 tune_series_gygy[4]
port 21 nsew signal input
rlabel metal2 s 30408 0 30464 400 6 tune_series_gygy[5]
port 22 nsew signal input
rlabel metal2 s 31640 0 31696 400 6 tune_series_gygy[6]
port 23 nsew signal input
rlabel metal2 s 32872 0 32928 400 6 tune_series_gygy[7]
port 24 nsew signal input
rlabel metal2 s 840 0 896 400 6 tune_shunt[0]
port 25 nsew signal input
rlabel metal2 s 13160 0 13216 400 6 tune_shunt[10]
port 26 nsew signal input
rlabel metal2 s 2072 0 2128 400 6 tune_shunt[1]
port 27 nsew signal input
rlabel metal2 s 3304 0 3360 400 6 tune_shunt[2]
port 28 nsew signal input
rlabel metal2 s 4536 0 4592 400 6 tune_shunt[3]
port 29 nsew signal input
rlabel metal2 s 5768 0 5824 400 6 tune_shunt[4]
port 30 nsew signal input
rlabel metal2 s 7000 0 7056 400 6 tune_shunt[5]
port 31 nsew signal input
rlabel metal2 s 8232 0 8288 400 6 tune_shunt[6]
port 32 nsew signal input
rlabel metal2 s 9464 0 9520 400 6 tune_shunt[7]
port 33 nsew signal input
rlabel metal2 s 10696 0 10752 400 6 tune_shunt[8]
port 34 nsew signal input
rlabel metal2 s 11928 0 11984 400 6 tune_shunt[9]
port 35 nsew signal input
rlabel metal2 s 34104 0 34160 400 6 tune_shunt_gy[0]
port 36 nsew signal input
rlabel metal2 s 35336 0 35392 400 6 tune_shunt_gy[1]
port 37 nsew signal input
rlabel metal2 s 36568 0 36624 400 6 tune_shunt_gy[2]
port 38 nsew signal input
rlabel metal2 s 37800 0 37856 400 6 tune_shunt_gy[3]
port 39 nsew signal input
rlabel metal2 s 39032 0 39088 400 6 tune_shunt_gy[4]
port 40 nsew signal input
rlabel metal4 s 2054 1538 2554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 7054 1538 7554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 12054 1538 12554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 17054 1538 17554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 22054 1538 22554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 27054 1538 27554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 32054 1538 32554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 37054 1538 37554 18454 6 vdd
port 41 nsew power bidirectional
rlabel metal4 s 4554 1538 5054 18454 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 9554 1538 10054 18454 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 14554 1538 15054 18454 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 19554 1538 20054 18454 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 24554 1538 25054 18454 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 29554 1538 30054 18454 6 vss
port 42 nsew ground bidirectional
rlabel metal4 s 34554 1538 35054 18454 6 vss
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1453588
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/caparray_s2/runs/22_12_05_03_50/results/signoff/caparray_s2.magic.gds
string GDS_START 56750
<< end >>

