magic
tech gf180mcuC
magscale 1 5
timestamp 1670230331
<< metal1 >>
rect 672 18437 39312 18454
rect 672 18411 2074 18437
rect 2100 18411 2136 18437
rect 2162 18411 2198 18437
rect 2224 18411 2260 18437
rect 2286 18411 2322 18437
rect 2348 18411 2384 18437
rect 2410 18411 2446 18437
rect 2472 18411 2508 18437
rect 2534 18411 7074 18437
rect 7100 18411 7136 18437
rect 7162 18411 7198 18437
rect 7224 18411 7260 18437
rect 7286 18411 7322 18437
rect 7348 18411 7384 18437
rect 7410 18411 7446 18437
rect 7472 18411 7508 18437
rect 7534 18411 12074 18437
rect 12100 18411 12136 18437
rect 12162 18411 12198 18437
rect 12224 18411 12260 18437
rect 12286 18411 12322 18437
rect 12348 18411 12384 18437
rect 12410 18411 12446 18437
rect 12472 18411 12508 18437
rect 12534 18411 17074 18437
rect 17100 18411 17136 18437
rect 17162 18411 17198 18437
rect 17224 18411 17260 18437
rect 17286 18411 17322 18437
rect 17348 18411 17384 18437
rect 17410 18411 17446 18437
rect 17472 18411 17508 18437
rect 17534 18411 22074 18437
rect 22100 18411 22136 18437
rect 22162 18411 22198 18437
rect 22224 18411 22260 18437
rect 22286 18411 22322 18437
rect 22348 18411 22384 18437
rect 22410 18411 22446 18437
rect 22472 18411 22508 18437
rect 22534 18411 27074 18437
rect 27100 18411 27136 18437
rect 27162 18411 27198 18437
rect 27224 18411 27260 18437
rect 27286 18411 27322 18437
rect 27348 18411 27384 18437
rect 27410 18411 27446 18437
rect 27472 18411 27508 18437
rect 27534 18411 32074 18437
rect 32100 18411 32136 18437
rect 32162 18411 32198 18437
rect 32224 18411 32260 18437
rect 32286 18411 32322 18437
rect 32348 18411 32384 18437
rect 32410 18411 32446 18437
rect 32472 18411 32508 18437
rect 32534 18411 37074 18437
rect 37100 18411 37136 18437
rect 37162 18411 37198 18437
rect 37224 18411 37260 18437
rect 37286 18411 37322 18437
rect 37348 18411 37384 18437
rect 37410 18411 37446 18437
rect 37472 18411 37508 18437
rect 37534 18411 39312 18437
rect 672 18394 39312 18411
rect 11097 18215 11103 18241
rect 11129 18215 11135 18241
rect 11825 18215 11831 18241
rect 11857 18215 11863 18241
rect 13337 18215 13343 18241
rect 13369 18215 13375 18241
rect 14233 18215 14239 18241
rect 14265 18215 14271 18241
rect 14625 18215 14631 18241
rect 14657 18215 14663 18241
rect 15801 18215 15807 18241
rect 15833 18215 15839 18241
rect 12049 18159 12055 18185
rect 12081 18159 12087 18185
rect 14233 18159 14239 18185
rect 14265 18159 14271 18185
rect 15801 18159 15807 18185
rect 15833 18159 15839 18185
rect 672 18045 39312 18062
rect 672 18019 4574 18045
rect 4600 18019 4636 18045
rect 4662 18019 4698 18045
rect 4724 18019 4760 18045
rect 4786 18019 4822 18045
rect 4848 18019 4884 18045
rect 4910 18019 4946 18045
rect 4972 18019 5008 18045
rect 5034 18019 9574 18045
rect 9600 18019 9636 18045
rect 9662 18019 9698 18045
rect 9724 18019 9760 18045
rect 9786 18019 9822 18045
rect 9848 18019 9884 18045
rect 9910 18019 9946 18045
rect 9972 18019 10008 18045
rect 10034 18019 14574 18045
rect 14600 18019 14636 18045
rect 14662 18019 14698 18045
rect 14724 18019 14760 18045
rect 14786 18019 14822 18045
rect 14848 18019 14884 18045
rect 14910 18019 14946 18045
rect 14972 18019 15008 18045
rect 15034 18019 19574 18045
rect 19600 18019 19636 18045
rect 19662 18019 19698 18045
rect 19724 18019 19760 18045
rect 19786 18019 19822 18045
rect 19848 18019 19884 18045
rect 19910 18019 19946 18045
rect 19972 18019 20008 18045
rect 20034 18019 24574 18045
rect 24600 18019 24636 18045
rect 24662 18019 24698 18045
rect 24724 18019 24760 18045
rect 24786 18019 24822 18045
rect 24848 18019 24884 18045
rect 24910 18019 24946 18045
rect 24972 18019 25008 18045
rect 25034 18019 29574 18045
rect 29600 18019 29636 18045
rect 29662 18019 29698 18045
rect 29724 18019 29760 18045
rect 29786 18019 29822 18045
rect 29848 18019 29884 18045
rect 29910 18019 29946 18045
rect 29972 18019 30008 18045
rect 30034 18019 34574 18045
rect 34600 18019 34636 18045
rect 34662 18019 34698 18045
rect 34724 18019 34760 18045
rect 34786 18019 34822 18045
rect 34848 18019 34884 18045
rect 34910 18019 34946 18045
rect 34972 18019 35008 18045
rect 35034 18019 39312 18045
rect 672 18002 39312 18019
rect 14569 17879 14575 17905
rect 14601 17879 14607 17905
rect 15913 17879 15919 17905
rect 15945 17879 15951 17905
rect 9809 17823 9815 17849
rect 9841 17823 9847 17849
rect 10257 17823 10263 17849
rect 10289 17823 10295 17849
rect 10481 17823 10487 17849
rect 10513 17823 10519 17849
rect 11265 17823 11271 17849
rect 11297 17823 11303 17849
rect 11825 17823 11831 17849
rect 11857 17823 11863 17849
rect 11937 17823 11943 17849
rect 11969 17823 11975 17849
rect 13393 17823 13399 17849
rect 13425 17823 13431 17849
rect 14569 17823 14575 17849
rect 14601 17823 14607 17849
rect 15073 17823 15079 17849
rect 15105 17823 15111 17849
rect 15913 17823 15919 17849
rect 15945 17823 15951 17849
rect 672 17653 39312 17670
rect 672 17627 2074 17653
rect 2100 17627 2136 17653
rect 2162 17627 2198 17653
rect 2224 17627 2260 17653
rect 2286 17627 2322 17653
rect 2348 17627 2384 17653
rect 2410 17627 2446 17653
rect 2472 17627 2508 17653
rect 2534 17627 7074 17653
rect 7100 17627 7136 17653
rect 7162 17627 7198 17653
rect 7224 17627 7260 17653
rect 7286 17627 7322 17653
rect 7348 17627 7384 17653
rect 7410 17627 7446 17653
rect 7472 17627 7508 17653
rect 7534 17627 12074 17653
rect 12100 17627 12136 17653
rect 12162 17627 12198 17653
rect 12224 17627 12260 17653
rect 12286 17627 12322 17653
rect 12348 17627 12384 17653
rect 12410 17627 12446 17653
rect 12472 17627 12508 17653
rect 12534 17627 17074 17653
rect 17100 17627 17136 17653
rect 17162 17627 17198 17653
rect 17224 17627 17260 17653
rect 17286 17627 17322 17653
rect 17348 17627 17384 17653
rect 17410 17627 17446 17653
rect 17472 17627 17508 17653
rect 17534 17627 22074 17653
rect 22100 17627 22136 17653
rect 22162 17627 22198 17653
rect 22224 17627 22260 17653
rect 22286 17627 22322 17653
rect 22348 17627 22384 17653
rect 22410 17627 22446 17653
rect 22472 17627 22508 17653
rect 22534 17627 27074 17653
rect 27100 17627 27136 17653
rect 27162 17627 27198 17653
rect 27224 17627 27260 17653
rect 27286 17627 27322 17653
rect 27348 17627 27384 17653
rect 27410 17627 27446 17653
rect 27472 17627 27508 17653
rect 27534 17627 32074 17653
rect 32100 17627 32136 17653
rect 32162 17627 32198 17653
rect 32224 17627 32260 17653
rect 32286 17627 32322 17653
rect 32348 17627 32384 17653
rect 32410 17627 32446 17653
rect 32472 17627 32508 17653
rect 32534 17627 37074 17653
rect 37100 17627 37136 17653
rect 37162 17627 37198 17653
rect 37224 17627 37260 17653
rect 37286 17627 37322 17653
rect 37348 17627 37384 17653
rect 37410 17627 37446 17653
rect 37472 17627 37508 17653
rect 37534 17627 39312 17653
rect 672 17610 39312 17627
rect 9249 17431 9255 17457
rect 9281 17431 9287 17457
rect 10369 17431 10375 17457
rect 10401 17431 10407 17457
rect 11769 17431 11775 17457
rect 11801 17431 11807 17457
rect 12217 17431 12223 17457
rect 12249 17431 12255 17457
rect 12441 17431 12447 17457
rect 12473 17431 12479 17457
rect 13281 17431 13287 17457
rect 13313 17431 13319 17457
rect 14233 17431 14239 17457
rect 14265 17431 14271 17457
rect 15073 17431 15079 17457
rect 15105 17431 15111 17457
rect 15969 17431 15975 17457
rect 16001 17431 16007 17457
rect 16249 17431 16255 17457
rect 16281 17431 16287 17457
rect 16753 17431 16759 17457
rect 16785 17431 16791 17457
rect 16921 17431 16927 17457
rect 16953 17431 16959 17457
rect 10369 17375 10375 17401
rect 10401 17375 10407 17401
rect 14233 17375 14239 17401
rect 14265 17375 14271 17401
rect 15969 17375 15975 17401
rect 16001 17375 16007 17401
rect 672 17261 39312 17278
rect 672 17235 4574 17261
rect 4600 17235 4636 17261
rect 4662 17235 4698 17261
rect 4724 17235 4760 17261
rect 4786 17235 4822 17261
rect 4848 17235 4884 17261
rect 4910 17235 4946 17261
rect 4972 17235 5008 17261
rect 5034 17235 9574 17261
rect 9600 17235 9636 17261
rect 9662 17235 9698 17261
rect 9724 17235 9760 17261
rect 9786 17235 9822 17261
rect 9848 17235 9884 17261
rect 9910 17235 9946 17261
rect 9972 17235 10008 17261
rect 10034 17235 14574 17261
rect 14600 17235 14636 17261
rect 14662 17235 14698 17261
rect 14724 17235 14760 17261
rect 14786 17235 14822 17261
rect 14848 17235 14884 17261
rect 14910 17235 14946 17261
rect 14972 17235 15008 17261
rect 15034 17235 19574 17261
rect 19600 17235 19636 17261
rect 19662 17235 19698 17261
rect 19724 17235 19760 17261
rect 19786 17235 19822 17261
rect 19848 17235 19884 17261
rect 19910 17235 19946 17261
rect 19972 17235 20008 17261
rect 20034 17235 24574 17261
rect 24600 17235 24636 17261
rect 24662 17235 24698 17261
rect 24724 17235 24760 17261
rect 24786 17235 24822 17261
rect 24848 17235 24884 17261
rect 24910 17235 24946 17261
rect 24972 17235 25008 17261
rect 25034 17235 29574 17261
rect 29600 17235 29636 17261
rect 29662 17235 29698 17261
rect 29724 17235 29760 17261
rect 29786 17235 29822 17261
rect 29848 17235 29884 17261
rect 29910 17235 29946 17261
rect 29972 17235 30008 17261
rect 30034 17235 34574 17261
rect 34600 17235 34636 17261
rect 34662 17235 34698 17261
rect 34724 17235 34760 17261
rect 34786 17235 34822 17261
rect 34848 17235 34884 17261
rect 34910 17235 34946 17261
rect 34972 17235 35008 17261
rect 35034 17235 39312 17261
rect 672 17218 39312 17235
rect 16137 17095 16143 17121
rect 16169 17095 16175 17121
rect 17873 17095 17879 17121
rect 17905 17095 17911 17121
rect 10089 17039 10095 17065
rect 10121 17039 10127 17065
rect 10369 17039 10375 17065
rect 10401 17039 10407 17065
rect 10481 17039 10487 17065
rect 10513 17039 10519 17065
rect 11265 17039 11271 17065
rect 11297 17039 11303 17065
rect 11825 17039 11831 17065
rect 11857 17039 11863 17065
rect 11937 17039 11943 17065
rect 11969 17039 11975 17065
rect 13729 17039 13735 17065
rect 13761 17039 13767 17065
rect 14289 17039 14295 17065
rect 14321 17039 14327 17065
rect 14457 17039 14463 17065
rect 14489 17039 14495 17065
rect 15185 17039 15191 17065
rect 15217 17039 15223 17065
rect 15969 17039 15975 17065
rect 16001 17039 16007 17065
rect 16809 17039 16815 17065
rect 16841 17039 16847 17065
rect 17873 17039 17879 17065
rect 17905 17039 17911 17065
rect 672 16869 39312 16886
rect 672 16843 2074 16869
rect 2100 16843 2136 16869
rect 2162 16843 2198 16869
rect 2224 16843 2260 16869
rect 2286 16843 2322 16869
rect 2348 16843 2384 16869
rect 2410 16843 2446 16869
rect 2472 16843 2508 16869
rect 2534 16843 7074 16869
rect 7100 16843 7136 16869
rect 7162 16843 7198 16869
rect 7224 16843 7260 16869
rect 7286 16843 7322 16869
rect 7348 16843 7384 16869
rect 7410 16843 7446 16869
rect 7472 16843 7508 16869
rect 7534 16843 12074 16869
rect 12100 16843 12136 16869
rect 12162 16843 12198 16869
rect 12224 16843 12260 16869
rect 12286 16843 12322 16869
rect 12348 16843 12384 16869
rect 12410 16843 12446 16869
rect 12472 16843 12508 16869
rect 12534 16843 17074 16869
rect 17100 16843 17136 16869
rect 17162 16843 17198 16869
rect 17224 16843 17260 16869
rect 17286 16843 17322 16869
rect 17348 16843 17384 16869
rect 17410 16843 17446 16869
rect 17472 16843 17508 16869
rect 17534 16843 22074 16869
rect 22100 16843 22136 16869
rect 22162 16843 22198 16869
rect 22224 16843 22260 16869
rect 22286 16843 22322 16869
rect 22348 16843 22384 16869
rect 22410 16843 22446 16869
rect 22472 16843 22508 16869
rect 22534 16843 27074 16869
rect 27100 16843 27136 16869
rect 27162 16843 27198 16869
rect 27224 16843 27260 16869
rect 27286 16843 27322 16869
rect 27348 16843 27384 16869
rect 27410 16843 27446 16869
rect 27472 16843 27508 16869
rect 27534 16843 32074 16869
rect 32100 16843 32136 16869
rect 32162 16843 32198 16869
rect 32224 16843 32260 16869
rect 32286 16843 32322 16869
rect 32348 16843 32384 16869
rect 32410 16843 32446 16869
rect 32472 16843 32508 16869
rect 32534 16843 37074 16869
rect 37100 16843 37136 16869
rect 37162 16843 37198 16869
rect 37224 16843 37260 16869
rect 37286 16843 37322 16869
rect 37348 16843 37384 16869
rect 37410 16843 37446 16869
rect 37472 16843 37508 16869
rect 37534 16843 39312 16869
rect 672 16826 39312 16843
rect 7793 16647 7799 16673
rect 7825 16647 7831 16673
rect 8969 16647 8975 16673
rect 9001 16647 9007 16673
rect 9473 16647 9479 16673
rect 9505 16647 9511 16673
rect 10425 16647 10431 16673
rect 10457 16647 10463 16673
rect 11769 16647 11775 16673
rect 11801 16647 11807 16673
rect 12217 16647 12223 16673
rect 12249 16647 12255 16673
rect 12441 16647 12447 16673
rect 12473 16647 12479 16673
rect 13281 16647 13287 16673
rect 13313 16647 13319 16673
rect 14233 16647 14239 16673
rect 14265 16647 14271 16673
rect 15073 16647 15079 16673
rect 15105 16647 15111 16673
rect 15969 16647 15975 16673
rect 16001 16647 16007 16673
rect 16249 16647 16255 16673
rect 16281 16647 16287 16673
rect 16753 16647 16759 16673
rect 16785 16647 16791 16673
rect 16921 16647 16927 16673
rect 16953 16647 16959 16673
rect 8969 16591 8975 16617
rect 9001 16591 9007 16617
rect 10425 16591 10431 16617
rect 10457 16591 10463 16617
rect 14233 16591 14239 16617
rect 14265 16591 14271 16617
rect 15969 16591 15975 16617
rect 16001 16591 16007 16617
rect 672 16477 39312 16494
rect 672 16451 4574 16477
rect 4600 16451 4636 16477
rect 4662 16451 4698 16477
rect 4724 16451 4760 16477
rect 4786 16451 4822 16477
rect 4848 16451 4884 16477
rect 4910 16451 4946 16477
rect 4972 16451 5008 16477
rect 5034 16451 9574 16477
rect 9600 16451 9636 16477
rect 9662 16451 9698 16477
rect 9724 16451 9760 16477
rect 9786 16451 9822 16477
rect 9848 16451 9884 16477
rect 9910 16451 9946 16477
rect 9972 16451 10008 16477
rect 10034 16451 14574 16477
rect 14600 16451 14636 16477
rect 14662 16451 14698 16477
rect 14724 16451 14760 16477
rect 14786 16451 14822 16477
rect 14848 16451 14884 16477
rect 14910 16451 14946 16477
rect 14972 16451 15008 16477
rect 15034 16451 19574 16477
rect 19600 16451 19636 16477
rect 19662 16451 19698 16477
rect 19724 16451 19760 16477
rect 19786 16451 19822 16477
rect 19848 16451 19884 16477
rect 19910 16451 19946 16477
rect 19972 16451 20008 16477
rect 20034 16451 24574 16477
rect 24600 16451 24636 16477
rect 24662 16451 24698 16477
rect 24724 16451 24760 16477
rect 24786 16451 24822 16477
rect 24848 16451 24884 16477
rect 24910 16451 24946 16477
rect 24972 16451 25008 16477
rect 25034 16451 29574 16477
rect 29600 16451 29636 16477
rect 29662 16451 29698 16477
rect 29724 16451 29760 16477
rect 29786 16451 29822 16477
rect 29848 16451 29884 16477
rect 29910 16451 29946 16477
rect 29972 16451 30008 16477
rect 30034 16451 34574 16477
rect 34600 16451 34636 16477
rect 34662 16451 34698 16477
rect 34724 16451 34760 16477
rect 34786 16451 34822 16477
rect 34848 16451 34884 16477
rect 34910 16451 34946 16477
rect 34972 16451 35008 16477
rect 35034 16451 39312 16477
rect 672 16434 39312 16451
rect 10985 16311 10991 16337
rect 11017 16311 11023 16337
rect 14625 16311 14631 16337
rect 14657 16311 14663 16337
rect 16305 16311 16311 16337
rect 16337 16311 16343 16337
rect 17873 16311 17879 16337
rect 17905 16311 17911 16337
rect 10089 16255 10095 16281
rect 10121 16255 10127 16281
rect 10985 16255 10991 16281
rect 11017 16255 11023 16281
rect 11265 16255 11271 16281
rect 11297 16255 11303 16281
rect 11825 16255 11831 16281
rect 11857 16255 11863 16281
rect 11937 16255 11943 16281
rect 11969 16255 11975 16281
rect 13729 16255 13735 16281
rect 13761 16255 13767 16281
rect 14401 16255 14407 16281
rect 14433 16255 14439 16281
rect 15129 16255 15135 16281
rect 15161 16255 15167 16281
rect 16305 16255 16311 16281
rect 16337 16255 16343 16281
rect 16809 16255 16815 16281
rect 16841 16255 16847 16281
rect 17873 16255 17879 16281
rect 17905 16255 17911 16281
rect 18265 16255 18271 16281
rect 18297 16255 18303 16281
rect 18713 16255 18719 16281
rect 18745 16255 18751 16281
rect 18937 16255 18943 16281
rect 18969 16255 18975 16281
rect 672 16085 39312 16102
rect 672 16059 2074 16085
rect 2100 16059 2136 16085
rect 2162 16059 2198 16085
rect 2224 16059 2260 16085
rect 2286 16059 2322 16085
rect 2348 16059 2384 16085
rect 2410 16059 2446 16085
rect 2472 16059 2508 16085
rect 2534 16059 7074 16085
rect 7100 16059 7136 16085
rect 7162 16059 7198 16085
rect 7224 16059 7260 16085
rect 7286 16059 7322 16085
rect 7348 16059 7384 16085
rect 7410 16059 7446 16085
rect 7472 16059 7508 16085
rect 7534 16059 12074 16085
rect 12100 16059 12136 16085
rect 12162 16059 12198 16085
rect 12224 16059 12260 16085
rect 12286 16059 12322 16085
rect 12348 16059 12384 16085
rect 12410 16059 12446 16085
rect 12472 16059 12508 16085
rect 12534 16059 17074 16085
rect 17100 16059 17136 16085
rect 17162 16059 17198 16085
rect 17224 16059 17260 16085
rect 17286 16059 17322 16085
rect 17348 16059 17384 16085
rect 17410 16059 17446 16085
rect 17472 16059 17508 16085
rect 17534 16059 22074 16085
rect 22100 16059 22136 16085
rect 22162 16059 22198 16085
rect 22224 16059 22260 16085
rect 22286 16059 22322 16085
rect 22348 16059 22384 16085
rect 22410 16059 22446 16085
rect 22472 16059 22508 16085
rect 22534 16059 27074 16085
rect 27100 16059 27136 16085
rect 27162 16059 27198 16085
rect 27224 16059 27260 16085
rect 27286 16059 27322 16085
rect 27348 16059 27384 16085
rect 27410 16059 27446 16085
rect 27472 16059 27508 16085
rect 27534 16059 32074 16085
rect 32100 16059 32136 16085
rect 32162 16059 32198 16085
rect 32224 16059 32260 16085
rect 32286 16059 32322 16085
rect 32348 16059 32384 16085
rect 32410 16059 32446 16085
rect 32472 16059 32508 16085
rect 32534 16059 37074 16085
rect 37100 16059 37136 16085
rect 37162 16059 37198 16085
rect 37224 16059 37260 16085
rect 37286 16059 37322 16085
rect 37348 16059 37384 16085
rect 37410 16059 37446 16085
rect 37472 16059 37508 16085
rect 37534 16059 39312 16085
rect 672 16042 39312 16059
rect 8073 15863 8079 15889
rect 8105 15863 8111 15889
rect 8969 15863 8975 15889
rect 9001 15863 9007 15889
rect 9473 15863 9479 15889
rect 9505 15863 9511 15889
rect 10425 15863 10431 15889
rect 10457 15863 10463 15889
rect 11769 15863 11775 15889
rect 11801 15863 11807 15889
rect 12217 15863 12223 15889
rect 12249 15863 12255 15889
rect 12441 15863 12447 15889
rect 12473 15863 12479 15889
rect 13281 15863 13287 15889
rect 13313 15863 13319 15889
rect 14401 15863 14407 15889
rect 14433 15863 14439 15889
rect 15073 15863 15079 15889
rect 15105 15863 15111 15889
rect 15969 15863 15975 15889
rect 16001 15863 16007 15889
rect 16249 15863 16255 15889
rect 16281 15863 16287 15889
rect 16809 15863 16815 15889
rect 16841 15863 16847 15889
rect 16921 15863 16927 15889
rect 16953 15863 16959 15889
rect 18769 15863 18775 15889
rect 18801 15863 18807 15889
rect 19217 15863 19223 15889
rect 19249 15863 19255 15889
rect 19441 15863 19447 15889
rect 19473 15863 19479 15889
rect 8969 15807 8975 15833
rect 9001 15807 9007 15833
rect 10425 15807 10431 15833
rect 10457 15807 10463 15833
rect 14401 15807 14407 15833
rect 14433 15807 14439 15833
rect 15969 15807 15975 15833
rect 16001 15807 16007 15833
rect 672 15693 39312 15710
rect 672 15667 4574 15693
rect 4600 15667 4636 15693
rect 4662 15667 4698 15693
rect 4724 15667 4760 15693
rect 4786 15667 4822 15693
rect 4848 15667 4884 15693
rect 4910 15667 4946 15693
rect 4972 15667 5008 15693
rect 5034 15667 9574 15693
rect 9600 15667 9636 15693
rect 9662 15667 9698 15693
rect 9724 15667 9760 15693
rect 9786 15667 9822 15693
rect 9848 15667 9884 15693
rect 9910 15667 9946 15693
rect 9972 15667 10008 15693
rect 10034 15667 14574 15693
rect 14600 15667 14636 15693
rect 14662 15667 14698 15693
rect 14724 15667 14760 15693
rect 14786 15667 14822 15693
rect 14848 15667 14884 15693
rect 14910 15667 14946 15693
rect 14972 15667 15008 15693
rect 15034 15667 19574 15693
rect 19600 15667 19636 15693
rect 19662 15667 19698 15693
rect 19724 15667 19760 15693
rect 19786 15667 19822 15693
rect 19848 15667 19884 15693
rect 19910 15667 19946 15693
rect 19972 15667 20008 15693
rect 20034 15667 24574 15693
rect 24600 15667 24636 15693
rect 24662 15667 24698 15693
rect 24724 15667 24760 15693
rect 24786 15667 24822 15693
rect 24848 15667 24884 15693
rect 24910 15667 24946 15693
rect 24972 15667 25008 15693
rect 25034 15667 29574 15693
rect 29600 15667 29636 15693
rect 29662 15667 29698 15693
rect 29724 15667 29760 15693
rect 29786 15667 29822 15693
rect 29848 15667 29884 15693
rect 29910 15667 29946 15693
rect 29972 15667 30008 15693
rect 30034 15667 34574 15693
rect 34600 15667 34636 15693
rect 34662 15667 34698 15693
rect 34724 15667 34760 15693
rect 34786 15667 34822 15693
rect 34848 15667 34884 15693
rect 34910 15667 34946 15693
rect 34972 15667 35008 15693
rect 35034 15667 39312 15693
rect 672 15650 39312 15667
rect 1857 15527 1863 15553
rect 1889 15527 1895 15553
rect 4489 15527 4495 15553
rect 4521 15527 4527 15553
rect 7009 15527 7015 15553
rect 7041 15527 7047 15553
rect 8465 15527 8471 15553
rect 8497 15527 8503 15553
rect 10985 15527 10991 15553
rect 11017 15527 11023 15553
rect 16137 15527 16143 15553
rect 16169 15527 16175 15553
rect 17873 15527 17879 15553
rect 17905 15527 17911 15553
rect 23417 15527 23423 15553
rect 23449 15527 23455 15553
rect 1857 15471 1863 15497
rect 1889 15471 1895 15497
rect 2753 15471 2759 15497
rect 2785 15471 2791 15497
rect 3313 15471 3319 15497
rect 3345 15471 3351 15497
rect 4489 15471 4495 15497
rect 4521 15471 4527 15497
rect 6113 15471 6119 15497
rect 6145 15471 6151 15497
rect 7009 15471 7015 15497
rect 7041 15471 7047 15497
rect 7569 15471 7575 15497
rect 7601 15471 7607 15497
rect 8465 15471 8471 15497
rect 8497 15471 8503 15497
rect 10033 15471 10039 15497
rect 10065 15471 10071 15497
rect 10985 15471 10991 15497
rect 11017 15471 11023 15497
rect 11265 15471 11271 15497
rect 11297 15471 11303 15497
rect 11825 15471 11831 15497
rect 11857 15471 11863 15497
rect 11937 15471 11943 15497
rect 11969 15471 11975 15497
rect 13729 15471 13735 15497
rect 13761 15471 13767 15497
rect 14289 15471 14295 15497
rect 14321 15471 14327 15497
rect 14457 15471 14463 15497
rect 14489 15471 14495 15497
rect 15185 15471 15191 15497
rect 15217 15471 15223 15497
rect 15969 15471 15975 15497
rect 16001 15471 16007 15497
rect 16809 15471 16815 15497
rect 16841 15471 16847 15497
rect 17873 15471 17879 15497
rect 17905 15471 17911 15497
rect 18265 15471 18271 15497
rect 18297 15471 18303 15497
rect 18713 15471 18719 15497
rect 18745 15471 18751 15497
rect 18937 15471 18943 15497
rect 18969 15471 18975 15497
rect 20785 15471 20791 15497
rect 20817 15471 20823 15497
rect 21233 15471 21239 15497
rect 21265 15471 21271 15497
rect 21457 15471 21463 15497
rect 21489 15471 21495 15497
rect 22521 15471 22527 15497
rect 22553 15471 22559 15497
rect 23417 15471 23423 15497
rect 23449 15471 23455 15497
rect 672 15301 39312 15318
rect 672 15275 2074 15301
rect 2100 15275 2136 15301
rect 2162 15275 2198 15301
rect 2224 15275 2260 15301
rect 2286 15275 2322 15301
rect 2348 15275 2384 15301
rect 2410 15275 2446 15301
rect 2472 15275 2508 15301
rect 2534 15275 7074 15301
rect 7100 15275 7136 15301
rect 7162 15275 7198 15301
rect 7224 15275 7260 15301
rect 7286 15275 7322 15301
rect 7348 15275 7384 15301
rect 7410 15275 7446 15301
rect 7472 15275 7508 15301
rect 7534 15275 12074 15301
rect 12100 15275 12136 15301
rect 12162 15275 12198 15301
rect 12224 15275 12260 15301
rect 12286 15275 12322 15301
rect 12348 15275 12384 15301
rect 12410 15275 12446 15301
rect 12472 15275 12508 15301
rect 12534 15275 17074 15301
rect 17100 15275 17136 15301
rect 17162 15275 17198 15301
rect 17224 15275 17260 15301
rect 17286 15275 17322 15301
rect 17348 15275 17384 15301
rect 17410 15275 17446 15301
rect 17472 15275 17508 15301
rect 17534 15275 22074 15301
rect 22100 15275 22136 15301
rect 22162 15275 22198 15301
rect 22224 15275 22260 15301
rect 22286 15275 22322 15301
rect 22348 15275 22384 15301
rect 22410 15275 22446 15301
rect 22472 15275 22508 15301
rect 22534 15275 27074 15301
rect 27100 15275 27136 15301
rect 27162 15275 27198 15301
rect 27224 15275 27260 15301
rect 27286 15275 27322 15301
rect 27348 15275 27384 15301
rect 27410 15275 27446 15301
rect 27472 15275 27508 15301
rect 27534 15275 32074 15301
rect 32100 15275 32136 15301
rect 32162 15275 32198 15301
rect 32224 15275 32260 15301
rect 32286 15275 32322 15301
rect 32348 15275 32384 15301
rect 32410 15275 32446 15301
rect 32472 15275 32508 15301
rect 32534 15275 37074 15301
rect 37100 15275 37136 15301
rect 37162 15275 37198 15301
rect 37224 15275 37260 15301
rect 37286 15275 37322 15301
rect 37348 15275 37384 15301
rect 37410 15275 37446 15301
rect 37472 15275 37508 15301
rect 37534 15275 39312 15301
rect 672 15258 39312 15275
rect 1521 15079 1527 15105
rect 1553 15079 1559 15105
rect 2473 15079 2479 15105
rect 2505 15079 2511 15105
rect 3817 15079 3823 15105
rect 3849 15079 3855 15105
rect 4377 15079 4383 15105
rect 4409 15079 4415 15105
rect 4489 15079 4495 15105
rect 4521 15079 4527 15105
rect 5553 15079 5559 15105
rect 5585 15079 5591 15105
rect 5833 15079 5839 15105
rect 5865 15079 5871 15105
rect 6449 15079 6455 15105
rect 6481 15079 6487 15105
rect 8073 15079 8079 15105
rect 8105 15079 8111 15105
rect 8969 15079 8975 15105
rect 9001 15079 9007 15105
rect 9473 15079 9479 15105
rect 9505 15079 9511 15105
rect 10425 15079 10431 15105
rect 10457 15079 10463 15105
rect 11769 15079 11775 15105
rect 11801 15079 11807 15105
rect 12721 15079 12727 15105
rect 12753 15079 12759 15105
rect 13281 15079 13287 15105
rect 13313 15079 13319 15105
rect 14401 15079 14407 15105
rect 14433 15079 14439 15105
rect 15073 15079 15079 15105
rect 15105 15079 15111 15105
rect 15969 15079 15975 15105
rect 16001 15079 16007 15105
rect 16249 15079 16255 15105
rect 16281 15079 16287 15105
rect 16977 15079 16983 15105
rect 17009 15079 17015 15105
rect 18825 15079 18831 15105
rect 18857 15079 18863 15105
rect 19329 15079 19335 15105
rect 19361 15079 19367 15105
rect 19441 15079 19447 15105
rect 19473 15079 19479 15105
rect 20505 15079 20511 15105
rect 20537 15079 20543 15105
rect 21009 15079 21015 15105
rect 21041 15079 21047 15105
rect 23025 15079 23031 15105
rect 23057 15079 23063 15105
rect 23921 15079 23927 15105
rect 23953 15079 23959 15105
rect 24481 15079 24487 15105
rect 24513 15079 24519 15105
rect 25321 15079 25327 15105
rect 25353 15079 25359 15105
rect 1521 15023 1527 15049
rect 1553 15023 1559 15049
rect 8969 15023 8975 15049
rect 9001 15023 9007 15049
rect 10425 15023 10431 15049
rect 10457 15023 10463 15049
rect 12721 15023 12727 15049
rect 12753 15023 12759 15049
rect 14401 15023 14407 15049
rect 14433 15023 14439 15049
rect 15969 15023 15975 15049
rect 16001 15023 16007 15049
rect 17201 15023 17207 15049
rect 17233 15023 17239 15049
rect 21177 15023 21183 15049
rect 21209 15023 21215 15049
rect 23921 15023 23927 15049
rect 23953 15023 23959 15049
rect 25321 15023 25327 15049
rect 25353 15023 25359 15049
rect 672 14909 39312 14926
rect 672 14883 4574 14909
rect 4600 14883 4636 14909
rect 4662 14883 4698 14909
rect 4724 14883 4760 14909
rect 4786 14883 4822 14909
rect 4848 14883 4884 14909
rect 4910 14883 4946 14909
rect 4972 14883 5008 14909
rect 5034 14883 9574 14909
rect 9600 14883 9636 14909
rect 9662 14883 9698 14909
rect 9724 14883 9760 14909
rect 9786 14883 9822 14909
rect 9848 14883 9884 14909
rect 9910 14883 9946 14909
rect 9972 14883 10008 14909
rect 10034 14883 14574 14909
rect 14600 14883 14636 14909
rect 14662 14883 14698 14909
rect 14724 14883 14760 14909
rect 14786 14883 14822 14909
rect 14848 14883 14884 14909
rect 14910 14883 14946 14909
rect 14972 14883 15008 14909
rect 15034 14883 19574 14909
rect 19600 14883 19636 14909
rect 19662 14883 19698 14909
rect 19724 14883 19760 14909
rect 19786 14883 19822 14909
rect 19848 14883 19884 14909
rect 19910 14883 19946 14909
rect 19972 14883 20008 14909
rect 20034 14883 24574 14909
rect 24600 14883 24636 14909
rect 24662 14883 24698 14909
rect 24724 14883 24760 14909
rect 24786 14883 24822 14909
rect 24848 14883 24884 14909
rect 24910 14883 24946 14909
rect 24972 14883 25008 14909
rect 25034 14883 29574 14909
rect 29600 14883 29636 14909
rect 29662 14883 29698 14909
rect 29724 14883 29760 14909
rect 29786 14883 29822 14909
rect 29848 14883 29884 14909
rect 29910 14883 29946 14909
rect 29972 14883 30008 14909
rect 30034 14883 34574 14909
rect 34600 14883 34636 14909
rect 34662 14883 34698 14909
rect 34724 14883 34760 14909
rect 34786 14883 34822 14909
rect 34848 14883 34884 14909
rect 34910 14883 34946 14909
rect 34972 14883 35008 14909
rect 35034 14883 39312 14909
rect 672 14866 39312 14883
rect 4489 14743 4495 14769
rect 4521 14743 4527 14769
rect 7009 14743 7015 14769
rect 7041 14743 7047 14769
rect 8465 14743 8471 14769
rect 8497 14743 8503 14769
rect 12441 14743 12447 14769
rect 12473 14743 12479 14769
rect 16361 14743 16367 14769
rect 16393 14743 16399 14769
rect 17929 14743 17935 14769
rect 17961 14743 17967 14769
rect 19441 14743 19447 14769
rect 19473 14743 19479 14769
rect 23417 14743 23423 14769
rect 23449 14743 23455 14769
rect 2361 14687 2367 14713
rect 2393 14687 2399 14713
rect 2473 14687 2479 14713
rect 2505 14687 2511 14713
rect 2753 14687 2759 14713
rect 2785 14687 2791 14713
rect 3313 14687 3319 14713
rect 3345 14687 3351 14713
rect 4489 14687 4495 14713
rect 4521 14687 4527 14713
rect 6113 14687 6119 14713
rect 6145 14687 6151 14713
rect 7009 14687 7015 14713
rect 7041 14687 7047 14713
rect 7569 14687 7575 14713
rect 7601 14687 7607 14713
rect 8465 14687 8471 14713
rect 8497 14687 8503 14713
rect 10033 14687 10039 14713
rect 10065 14687 10071 14713
rect 10369 14687 10375 14713
rect 10401 14687 10407 14713
rect 10481 14687 10487 14713
rect 10513 14687 10519 14713
rect 11265 14687 11271 14713
rect 11297 14687 11303 14713
rect 12441 14687 12447 14713
rect 12473 14687 12479 14713
rect 13729 14687 13735 14713
rect 13761 14687 13767 14713
rect 14289 14687 14295 14713
rect 14321 14687 14327 14713
rect 14457 14687 14463 14713
rect 14489 14687 14495 14713
rect 15185 14687 15191 14713
rect 15217 14687 15223 14713
rect 16361 14687 16367 14713
rect 16393 14687 16399 14713
rect 16809 14687 16815 14713
rect 16841 14687 16847 14713
rect 17929 14687 17935 14713
rect 17961 14687 17967 14713
rect 18265 14687 18271 14713
rect 18297 14687 18303 14713
rect 19441 14687 19447 14713
rect 19473 14687 19479 14713
rect 20785 14687 20791 14713
rect 20817 14687 20823 14713
rect 21233 14687 21239 14713
rect 21265 14687 21271 14713
rect 21457 14687 21463 14713
rect 21489 14687 21495 14713
rect 22521 14687 22527 14713
rect 22553 14687 22559 14713
rect 23417 14687 23423 14713
rect 23449 14687 23455 14713
rect 25041 14687 25047 14713
rect 25073 14687 25079 14713
rect 25321 14687 25327 14713
rect 25353 14687 25359 14713
rect 25433 14687 25439 14713
rect 25465 14687 25471 14713
rect 672 14517 39312 14534
rect 672 14491 2074 14517
rect 2100 14491 2136 14517
rect 2162 14491 2198 14517
rect 2224 14491 2260 14517
rect 2286 14491 2322 14517
rect 2348 14491 2384 14517
rect 2410 14491 2446 14517
rect 2472 14491 2508 14517
rect 2534 14491 7074 14517
rect 7100 14491 7136 14517
rect 7162 14491 7198 14517
rect 7224 14491 7260 14517
rect 7286 14491 7322 14517
rect 7348 14491 7384 14517
rect 7410 14491 7446 14517
rect 7472 14491 7508 14517
rect 7534 14491 12074 14517
rect 12100 14491 12136 14517
rect 12162 14491 12198 14517
rect 12224 14491 12260 14517
rect 12286 14491 12322 14517
rect 12348 14491 12384 14517
rect 12410 14491 12446 14517
rect 12472 14491 12508 14517
rect 12534 14491 17074 14517
rect 17100 14491 17136 14517
rect 17162 14491 17198 14517
rect 17224 14491 17260 14517
rect 17286 14491 17322 14517
rect 17348 14491 17384 14517
rect 17410 14491 17446 14517
rect 17472 14491 17508 14517
rect 17534 14491 22074 14517
rect 22100 14491 22136 14517
rect 22162 14491 22198 14517
rect 22224 14491 22260 14517
rect 22286 14491 22322 14517
rect 22348 14491 22384 14517
rect 22410 14491 22446 14517
rect 22472 14491 22508 14517
rect 22534 14491 27074 14517
rect 27100 14491 27136 14517
rect 27162 14491 27198 14517
rect 27224 14491 27260 14517
rect 27286 14491 27322 14517
rect 27348 14491 27384 14517
rect 27410 14491 27446 14517
rect 27472 14491 27508 14517
rect 27534 14491 32074 14517
rect 32100 14491 32136 14517
rect 32162 14491 32198 14517
rect 32224 14491 32260 14517
rect 32286 14491 32322 14517
rect 32348 14491 32384 14517
rect 32410 14491 32446 14517
rect 32472 14491 32508 14517
rect 32534 14491 37074 14517
rect 37100 14491 37136 14517
rect 37162 14491 37198 14517
rect 37224 14491 37260 14517
rect 37286 14491 37322 14517
rect 37348 14491 37384 14517
rect 37410 14491 37446 14517
rect 37472 14491 37508 14517
rect 37534 14491 39312 14517
rect 672 14474 39312 14491
rect 1745 14295 1751 14321
rect 1777 14295 1783 14321
rect 2473 14295 2479 14321
rect 2505 14295 2511 14321
rect 3817 14295 3823 14321
rect 3849 14295 3855 14321
rect 4377 14295 4383 14321
rect 4409 14295 4415 14321
rect 4489 14295 4495 14321
rect 4521 14295 4527 14321
rect 5553 14295 5559 14321
rect 5585 14295 5591 14321
rect 5833 14295 5839 14321
rect 5865 14295 5871 14321
rect 6449 14295 6455 14321
rect 6481 14295 6487 14321
rect 8073 14295 8079 14321
rect 8105 14295 8111 14321
rect 8969 14295 8975 14321
rect 9001 14295 9007 14321
rect 9473 14295 9479 14321
rect 9505 14295 9511 14321
rect 10369 14295 10375 14321
rect 10401 14295 10407 14321
rect 11769 14295 11775 14321
rect 11801 14295 11807 14321
rect 12609 14295 12615 14321
rect 12641 14295 12647 14321
rect 13281 14295 13287 14321
rect 13313 14295 13319 14321
rect 14401 14295 14407 14321
rect 14433 14295 14439 14321
rect 15073 14295 15079 14321
rect 15105 14295 15111 14321
rect 15969 14295 15975 14321
rect 16001 14295 16007 14321
rect 16249 14295 16255 14321
rect 16281 14295 16287 14321
rect 17425 14295 17431 14321
rect 17457 14295 17463 14321
rect 18825 14295 18831 14321
rect 18857 14295 18863 14321
rect 19329 14295 19335 14321
rect 19361 14295 19367 14321
rect 19441 14295 19447 14321
rect 19473 14295 19479 14321
rect 20505 14295 20511 14321
rect 20537 14295 20543 14321
rect 20673 14295 20679 14321
rect 20705 14295 20711 14321
rect 21009 14295 21015 14321
rect 21041 14295 21047 14321
rect 23025 14295 23031 14321
rect 23057 14295 23063 14321
rect 23921 14295 23927 14321
rect 23953 14295 23959 14321
rect 24481 14295 24487 14321
rect 24513 14295 24519 14321
rect 25377 14295 25383 14321
rect 25409 14295 25415 14321
rect 26721 14295 26727 14321
rect 26753 14295 26759 14321
rect 27673 14295 27679 14321
rect 27705 14295 27711 14321
rect 28457 14295 28463 14321
rect 28489 14295 28495 14321
rect 29353 14295 29359 14321
rect 29385 14295 29391 14321
rect 1521 14239 1527 14265
rect 1553 14239 1559 14265
rect 8969 14239 8975 14265
rect 9001 14239 9007 14265
rect 10369 14239 10375 14265
rect 10401 14239 10407 14265
rect 12721 14239 12727 14265
rect 12753 14239 12759 14265
rect 14401 14239 14407 14265
rect 14433 14239 14439 14265
rect 15969 14239 15975 14265
rect 16001 14239 16007 14265
rect 17425 14239 17431 14265
rect 17457 14239 17463 14265
rect 23921 14239 23927 14265
rect 23953 14239 23959 14265
rect 25377 14239 25383 14265
rect 25409 14239 25415 14265
rect 27673 14239 27679 14265
rect 27705 14239 27711 14265
rect 29353 14239 29359 14265
rect 29385 14239 29391 14265
rect 672 14125 39312 14142
rect 672 14099 4574 14125
rect 4600 14099 4636 14125
rect 4662 14099 4698 14125
rect 4724 14099 4760 14125
rect 4786 14099 4822 14125
rect 4848 14099 4884 14125
rect 4910 14099 4946 14125
rect 4972 14099 5008 14125
rect 5034 14099 9574 14125
rect 9600 14099 9636 14125
rect 9662 14099 9698 14125
rect 9724 14099 9760 14125
rect 9786 14099 9822 14125
rect 9848 14099 9884 14125
rect 9910 14099 9946 14125
rect 9972 14099 10008 14125
rect 10034 14099 14574 14125
rect 14600 14099 14636 14125
rect 14662 14099 14698 14125
rect 14724 14099 14760 14125
rect 14786 14099 14822 14125
rect 14848 14099 14884 14125
rect 14910 14099 14946 14125
rect 14972 14099 15008 14125
rect 15034 14099 19574 14125
rect 19600 14099 19636 14125
rect 19662 14099 19698 14125
rect 19724 14099 19760 14125
rect 19786 14099 19822 14125
rect 19848 14099 19884 14125
rect 19910 14099 19946 14125
rect 19972 14099 20008 14125
rect 20034 14099 24574 14125
rect 24600 14099 24636 14125
rect 24662 14099 24698 14125
rect 24724 14099 24760 14125
rect 24786 14099 24822 14125
rect 24848 14099 24884 14125
rect 24910 14099 24946 14125
rect 24972 14099 25008 14125
rect 25034 14099 29574 14125
rect 29600 14099 29636 14125
rect 29662 14099 29698 14125
rect 29724 14099 29760 14125
rect 29786 14099 29822 14125
rect 29848 14099 29884 14125
rect 29910 14099 29946 14125
rect 29972 14099 30008 14125
rect 30034 14099 34574 14125
rect 34600 14099 34636 14125
rect 34662 14099 34698 14125
rect 34724 14099 34760 14125
rect 34786 14099 34822 14125
rect 34848 14099 34884 14125
rect 34910 14099 34946 14125
rect 34972 14099 35008 14125
rect 35034 14099 39312 14125
rect 672 14082 39312 14099
rect 1969 13959 1975 13985
rect 2001 13959 2007 13985
rect 4489 13959 4495 13985
rect 4521 13959 4527 13985
rect 7009 13959 7015 13985
rect 7041 13959 7047 13985
rect 8465 13959 8471 13985
rect 8497 13959 8503 13985
rect 10761 13959 10767 13985
rect 10793 13959 10799 13985
rect 12441 13959 12447 13985
rect 12473 13959 12479 13985
rect 14905 13959 14911 13985
rect 14937 13959 14943 13985
rect 16361 13959 16367 13985
rect 16393 13959 16399 13985
rect 17929 13959 17935 13985
rect 17961 13959 17967 13985
rect 19441 13959 19447 13985
rect 19473 13959 19479 13985
rect 23417 13959 23423 13985
rect 23449 13959 23455 13985
rect 25937 13959 25943 13985
rect 25969 13959 25975 13985
rect 27393 13959 27399 13985
rect 27425 13959 27431 13985
rect 1969 13903 1975 13929
rect 2001 13903 2007 13929
rect 2753 13903 2759 13929
rect 2785 13903 2791 13929
rect 3313 13903 3319 13929
rect 3345 13903 3351 13929
rect 4489 13903 4495 13929
rect 4521 13903 4527 13929
rect 6113 13903 6119 13929
rect 6145 13903 6151 13929
rect 7009 13903 7015 13929
rect 7041 13903 7047 13929
rect 7569 13903 7575 13929
rect 7601 13903 7607 13929
rect 8465 13903 8471 13929
rect 8497 13903 8503 13929
rect 10089 13903 10095 13929
rect 10121 13903 10127 13929
rect 10761 13903 10767 13929
rect 10793 13903 10799 13929
rect 11265 13903 11271 13929
rect 11297 13903 11303 13929
rect 12441 13903 12447 13929
rect 12473 13903 12479 13929
rect 13729 13903 13735 13929
rect 13761 13903 13767 13929
rect 14905 13903 14911 13929
rect 14937 13903 14943 13929
rect 15185 13903 15191 13929
rect 15217 13903 15223 13929
rect 16361 13903 16367 13929
rect 16393 13903 16399 13929
rect 16809 13903 16815 13929
rect 16841 13903 16847 13929
rect 17929 13903 17935 13929
rect 17961 13903 17967 13929
rect 18265 13903 18271 13929
rect 18297 13903 18303 13929
rect 19441 13903 19447 13929
rect 19473 13903 19479 13929
rect 20953 13903 20959 13929
rect 20985 13903 20991 13929
rect 21233 13903 21239 13929
rect 21265 13903 21271 13929
rect 21457 13903 21463 13929
rect 21489 13903 21495 13929
rect 22521 13903 22527 13929
rect 22553 13903 22559 13929
rect 23417 13903 23423 13929
rect 23449 13903 23455 13929
rect 25041 13903 25047 13929
rect 25073 13903 25079 13929
rect 25937 13903 25943 13929
rect 25969 13903 25975 13929
rect 26217 13903 26223 13929
rect 26249 13903 26255 13929
rect 27393 13903 27399 13929
rect 27425 13903 27431 13929
rect 672 13733 39312 13750
rect 672 13707 2074 13733
rect 2100 13707 2136 13733
rect 2162 13707 2198 13733
rect 2224 13707 2260 13733
rect 2286 13707 2322 13733
rect 2348 13707 2384 13733
rect 2410 13707 2446 13733
rect 2472 13707 2508 13733
rect 2534 13707 7074 13733
rect 7100 13707 7136 13733
rect 7162 13707 7198 13733
rect 7224 13707 7260 13733
rect 7286 13707 7322 13733
rect 7348 13707 7384 13733
rect 7410 13707 7446 13733
rect 7472 13707 7508 13733
rect 7534 13707 12074 13733
rect 12100 13707 12136 13733
rect 12162 13707 12198 13733
rect 12224 13707 12260 13733
rect 12286 13707 12322 13733
rect 12348 13707 12384 13733
rect 12410 13707 12446 13733
rect 12472 13707 12508 13733
rect 12534 13707 17074 13733
rect 17100 13707 17136 13733
rect 17162 13707 17198 13733
rect 17224 13707 17260 13733
rect 17286 13707 17322 13733
rect 17348 13707 17384 13733
rect 17410 13707 17446 13733
rect 17472 13707 17508 13733
rect 17534 13707 22074 13733
rect 22100 13707 22136 13733
rect 22162 13707 22198 13733
rect 22224 13707 22260 13733
rect 22286 13707 22322 13733
rect 22348 13707 22384 13733
rect 22410 13707 22446 13733
rect 22472 13707 22508 13733
rect 22534 13707 27074 13733
rect 27100 13707 27136 13733
rect 27162 13707 27198 13733
rect 27224 13707 27260 13733
rect 27286 13707 27322 13733
rect 27348 13707 27384 13733
rect 27410 13707 27446 13733
rect 27472 13707 27508 13733
rect 27534 13707 32074 13733
rect 32100 13707 32136 13733
rect 32162 13707 32198 13733
rect 32224 13707 32260 13733
rect 32286 13707 32322 13733
rect 32348 13707 32384 13733
rect 32410 13707 32446 13733
rect 32472 13707 32508 13733
rect 32534 13707 37074 13733
rect 37100 13707 37136 13733
rect 37162 13707 37198 13733
rect 37224 13707 37260 13733
rect 37286 13707 37322 13733
rect 37348 13707 37384 13733
rect 37410 13707 37446 13733
rect 37472 13707 37508 13733
rect 37534 13707 39312 13733
rect 672 13690 39312 13707
rect 1801 13511 1807 13537
rect 1833 13511 1839 13537
rect 1969 13511 1975 13537
rect 2001 13511 2007 13537
rect 2473 13511 2479 13537
rect 2505 13511 2511 13537
rect 3817 13511 3823 13537
rect 3849 13511 3855 13537
rect 4377 13511 4383 13537
rect 4409 13511 4415 13537
rect 4489 13511 4495 13537
rect 4521 13511 4527 13537
rect 5497 13511 5503 13537
rect 5529 13511 5535 13537
rect 5833 13511 5839 13537
rect 5865 13511 5871 13537
rect 6449 13511 6455 13537
rect 6481 13511 6487 13537
rect 8073 13511 8079 13537
rect 8105 13511 8111 13537
rect 8353 13511 8359 13537
rect 8385 13511 8391 13537
rect 8465 13511 8471 13537
rect 8497 13511 8503 13537
rect 9473 13511 9479 13537
rect 9505 13511 9511 13537
rect 10425 13511 10431 13537
rect 10457 13511 10463 13537
rect 11769 13511 11775 13537
rect 11801 13511 11807 13537
rect 12945 13511 12951 13537
rect 12977 13511 12983 13537
rect 13281 13511 13287 13537
rect 13313 13511 13319 13537
rect 14121 13511 14127 13537
rect 14153 13511 14159 13537
rect 15465 13511 15471 13537
rect 15497 13511 15503 13537
rect 16249 13511 16255 13537
rect 16281 13511 16287 13537
rect 16809 13511 16815 13537
rect 16841 13511 16847 13537
rect 17929 13511 17935 13537
rect 17961 13511 17967 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 19329 13511 19335 13537
rect 19361 13511 19367 13537
rect 19441 13511 19447 13537
rect 19473 13511 19479 13537
rect 20505 13511 20511 13537
rect 20537 13511 20543 13537
rect 21009 13511 21015 13537
rect 21041 13511 21047 13537
rect 23025 13511 23031 13537
rect 23057 13511 23063 13537
rect 23921 13511 23927 13537
rect 23953 13511 23959 13537
rect 24481 13511 24487 13537
rect 24513 13511 24519 13537
rect 25377 13511 25383 13537
rect 25409 13511 25415 13537
rect 26721 13511 26727 13537
rect 26753 13511 26759 13537
rect 27673 13511 27679 13537
rect 27705 13511 27711 13537
rect 28457 13511 28463 13537
rect 28489 13511 28495 13537
rect 29353 13511 29359 13537
rect 29385 13511 29391 13537
rect 10425 13455 10431 13481
rect 10457 13455 10463 13481
rect 12945 13455 12951 13481
rect 12977 13455 12983 13481
rect 14401 13455 14407 13481
rect 14433 13455 14439 13481
rect 16249 13455 16255 13481
rect 16281 13455 16287 13481
rect 17929 13455 17935 13481
rect 17961 13455 17967 13481
rect 21177 13455 21183 13481
rect 21209 13455 21215 13481
rect 23921 13455 23927 13481
rect 23953 13455 23959 13481
rect 25377 13455 25383 13481
rect 25409 13455 25415 13481
rect 27673 13455 27679 13481
rect 27705 13455 27711 13481
rect 29353 13455 29359 13481
rect 29385 13455 29391 13481
rect 672 13341 39312 13358
rect 672 13315 4574 13341
rect 4600 13315 4636 13341
rect 4662 13315 4698 13341
rect 4724 13315 4760 13341
rect 4786 13315 4822 13341
rect 4848 13315 4884 13341
rect 4910 13315 4946 13341
rect 4972 13315 5008 13341
rect 5034 13315 9574 13341
rect 9600 13315 9636 13341
rect 9662 13315 9698 13341
rect 9724 13315 9760 13341
rect 9786 13315 9822 13341
rect 9848 13315 9884 13341
rect 9910 13315 9946 13341
rect 9972 13315 10008 13341
rect 10034 13315 14574 13341
rect 14600 13315 14636 13341
rect 14662 13315 14698 13341
rect 14724 13315 14760 13341
rect 14786 13315 14822 13341
rect 14848 13315 14884 13341
rect 14910 13315 14946 13341
rect 14972 13315 15008 13341
rect 15034 13315 19574 13341
rect 19600 13315 19636 13341
rect 19662 13315 19698 13341
rect 19724 13315 19760 13341
rect 19786 13315 19822 13341
rect 19848 13315 19884 13341
rect 19910 13315 19946 13341
rect 19972 13315 20008 13341
rect 20034 13315 24574 13341
rect 24600 13315 24636 13341
rect 24662 13315 24698 13341
rect 24724 13315 24760 13341
rect 24786 13315 24822 13341
rect 24848 13315 24884 13341
rect 24910 13315 24946 13341
rect 24972 13315 25008 13341
rect 25034 13315 29574 13341
rect 29600 13315 29636 13341
rect 29662 13315 29698 13341
rect 29724 13315 29760 13341
rect 29786 13315 29822 13341
rect 29848 13315 29884 13341
rect 29910 13315 29946 13341
rect 29972 13315 30008 13341
rect 30034 13315 34574 13341
rect 34600 13315 34636 13341
rect 34662 13315 34698 13341
rect 34724 13315 34760 13341
rect 34786 13315 34822 13341
rect 34848 13315 34884 13341
rect 34910 13315 34946 13341
rect 34972 13315 35008 13341
rect 35034 13315 39312 13341
rect 672 13298 39312 13315
rect 4489 13175 4495 13201
rect 4521 13175 4527 13201
rect 7009 13175 7015 13201
rect 7041 13175 7047 13201
rect 8353 13175 8359 13201
rect 8385 13175 8391 13201
rect 10761 13175 10767 13201
rect 10793 13175 10799 13201
rect 14345 13175 14351 13201
rect 14377 13175 14383 13201
rect 16025 13175 16031 13201
rect 16057 13175 16063 13201
rect 17985 13175 17991 13201
rect 18017 13175 18023 13201
rect 19441 13175 19447 13201
rect 19473 13175 19479 13201
rect 23417 13175 23423 13201
rect 23449 13175 23455 13201
rect 25937 13175 25943 13201
rect 25969 13175 25975 13201
rect 2361 13119 2367 13145
rect 2393 13119 2399 13145
rect 2585 13119 2591 13145
rect 2617 13119 2623 13145
rect 2753 13119 2759 13145
rect 2785 13119 2791 13145
rect 3593 13119 3599 13145
rect 3625 13119 3631 13145
rect 4489 13119 4495 13145
rect 4521 13119 4527 13145
rect 6113 13119 6119 13145
rect 6145 13119 6151 13145
rect 7009 13119 7015 13145
rect 7041 13119 7047 13145
rect 7569 13119 7575 13145
rect 7601 13119 7607 13145
rect 8353 13119 8359 13145
rect 8385 13119 8391 13145
rect 10089 13119 10095 13145
rect 10121 13119 10127 13145
rect 10761 13119 10767 13145
rect 10793 13119 10799 13145
rect 11265 13119 11271 13145
rect 11297 13119 11303 13145
rect 11825 13119 11831 13145
rect 11857 13119 11863 13145
rect 11993 13119 11999 13145
rect 12025 13119 12031 13145
rect 13393 13119 13399 13145
rect 13425 13119 13431 13145
rect 14177 13119 14183 13145
rect 14209 13119 14215 13145
rect 15129 13119 15135 13145
rect 15161 13119 15167 13145
rect 16025 13119 16031 13145
rect 16057 13119 16063 13145
rect 16977 13119 16983 13145
rect 17009 13119 17015 13145
rect 17985 13119 17991 13145
rect 18017 13119 18023 13145
rect 18545 13119 18551 13145
rect 18577 13119 18583 13145
rect 19441 13119 19447 13145
rect 19473 13119 19479 13145
rect 20953 13119 20959 13145
rect 20985 13119 20991 13145
rect 21233 13119 21239 13145
rect 21265 13119 21271 13145
rect 21457 13119 21463 13145
rect 21489 13119 21495 13145
rect 22521 13119 22527 13145
rect 22553 13119 22559 13145
rect 23417 13119 23423 13145
rect 23449 13119 23455 13145
rect 25041 13119 25047 13145
rect 25073 13119 25079 13145
rect 25937 13119 25943 13145
rect 25969 13119 25975 13145
rect 26497 13119 26503 13145
rect 26529 13119 26535 13145
rect 26777 13119 26783 13145
rect 26809 13119 26815 13145
rect 26889 13119 26895 13145
rect 26921 13119 26927 13145
rect 29017 13119 29023 13145
rect 29049 13119 29055 13145
rect 29297 13119 29303 13145
rect 29329 13119 29335 13145
rect 29409 13119 29415 13145
rect 29441 13119 29447 13145
rect 672 12949 39312 12966
rect 672 12923 2074 12949
rect 2100 12923 2136 12949
rect 2162 12923 2198 12949
rect 2224 12923 2260 12949
rect 2286 12923 2322 12949
rect 2348 12923 2384 12949
rect 2410 12923 2446 12949
rect 2472 12923 2508 12949
rect 2534 12923 7074 12949
rect 7100 12923 7136 12949
rect 7162 12923 7198 12949
rect 7224 12923 7260 12949
rect 7286 12923 7322 12949
rect 7348 12923 7384 12949
rect 7410 12923 7446 12949
rect 7472 12923 7508 12949
rect 7534 12923 12074 12949
rect 12100 12923 12136 12949
rect 12162 12923 12198 12949
rect 12224 12923 12260 12949
rect 12286 12923 12322 12949
rect 12348 12923 12384 12949
rect 12410 12923 12446 12949
rect 12472 12923 12508 12949
rect 12534 12923 17074 12949
rect 17100 12923 17136 12949
rect 17162 12923 17198 12949
rect 17224 12923 17260 12949
rect 17286 12923 17322 12949
rect 17348 12923 17384 12949
rect 17410 12923 17446 12949
rect 17472 12923 17508 12949
rect 17534 12923 22074 12949
rect 22100 12923 22136 12949
rect 22162 12923 22198 12949
rect 22224 12923 22260 12949
rect 22286 12923 22322 12949
rect 22348 12923 22384 12949
rect 22410 12923 22446 12949
rect 22472 12923 22508 12949
rect 22534 12923 27074 12949
rect 27100 12923 27136 12949
rect 27162 12923 27198 12949
rect 27224 12923 27260 12949
rect 27286 12923 27322 12949
rect 27348 12923 27384 12949
rect 27410 12923 27446 12949
rect 27472 12923 27508 12949
rect 27534 12923 32074 12949
rect 32100 12923 32136 12949
rect 32162 12923 32198 12949
rect 32224 12923 32260 12949
rect 32286 12923 32322 12949
rect 32348 12923 32384 12949
rect 32410 12923 32446 12949
rect 32472 12923 32508 12949
rect 32534 12923 37074 12949
rect 37100 12923 37136 12949
rect 37162 12923 37198 12949
rect 37224 12923 37260 12949
rect 37286 12923 37322 12949
rect 37348 12923 37384 12949
rect 37410 12923 37446 12949
rect 37472 12923 37508 12949
rect 37534 12923 39312 12949
rect 672 12906 39312 12923
rect 1801 12727 1807 12753
rect 1833 12727 1839 12753
rect 1969 12727 1975 12753
rect 2001 12727 2007 12753
rect 2473 12727 2479 12753
rect 2505 12727 2511 12753
rect 3817 12727 3823 12753
rect 3849 12727 3855 12753
rect 4993 12727 4999 12753
rect 5025 12727 5031 12753
rect 5553 12727 5559 12753
rect 5585 12727 5591 12753
rect 6449 12727 6455 12753
rect 6481 12727 6487 12753
rect 8073 12727 8079 12753
rect 8105 12727 8111 12753
rect 8353 12727 8359 12753
rect 8385 12727 8391 12753
rect 8465 12727 8471 12753
rect 8497 12727 8503 12753
rect 9473 12727 9479 12753
rect 9505 12727 9511 12753
rect 10425 12727 10431 12753
rect 10457 12727 10463 12753
rect 11769 12727 11775 12753
rect 11801 12727 11807 12753
rect 12217 12727 12223 12753
rect 12249 12727 12255 12753
rect 12441 12727 12447 12753
rect 12473 12727 12479 12753
rect 13225 12727 13231 12753
rect 13257 12727 13263 12753
rect 14177 12727 14183 12753
rect 14209 12727 14215 12753
rect 15745 12727 15751 12753
rect 15777 12727 15783 12753
rect 16641 12727 16647 12753
rect 16673 12727 16679 12753
rect 16921 12727 16927 12753
rect 16953 12727 16959 12753
rect 17873 12727 17879 12753
rect 17905 12727 17911 12753
rect 18769 12727 18775 12753
rect 18801 12727 18807 12753
rect 19945 12727 19951 12753
rect 19977 12727 19983 12753
rect 20505 12727 20511 12753
rect 20537 12727 20543 12753
rect 21177 12727 21183 12753
rect 21209 12727 21215 12753
rect 22745 12727 22751 12753
rect 22777 12727 22783 12753
rect 23305 12727 23311 12753
rect 23337 12727 23343 12753
rect 23417 12727 23423 12753
rect 23449 12727 23455 12753
rect 24369 12727 24375 12753
rect 24401 12727 24407 12753
rect 24649 12727 24655 12753
rect 24681 12727 24687 12753
rect 24873 12727 24879 12753
rect 24905 12727 24911 12753
rect 26721 12727 26727 12753
rect 26753 12727 26759 12753
rect 27169 12727 27175 12753
rect 27201 12727 27207 12753
rect 27393 12727 27399 12753
rect 27425 12727 27431 12753
rect 28457 12727 28463 12753
rect 28489 12727 28495 12753
rect 29353 12727 29359 12753
rect 29385 12727 29391 12753
rect 4993 12671 4999 12697
rect 5025 12671 5031 12697
rect 6449 12671 6455 12697
rect 6481 12671 6487 12697
rect 10425 12671 10431 12697
rect 10457 12671 10463 12697
rect 14177 12671 14183 12697
rect 14209 12671 14215 12697
rect 16641 12671 16647 12697
rect 16673 12671 16679 12697
rect 17873 12671 17879 12697
rect 17905 12671 17911 12697
rect 19945 12671 19951 12697
rect 19977 12671 19983 12697
rect 21177 12671 21183 12697
rect 21209 12671 21215 12697
rect 29353 12671 29359 12697
rect 29385 12671 29391 12697
rect 672 12557 39312 12574
rect 672 12531 4574 12557
rect 4600 12531 4636 12557
rect 4662 12531 4698 12557
rect 4724 12531 4760 12557
rect 4786 12531 4822 12557
rect 4848 12531 4884 12557
rect 4910 12531 4946 12557
rect 4972 12531 5008 12557
rect 5034 12531 9574 12557
rect 9600 12531 9636 12557
rect 9662 12531 9698 12557
rect 9724 12531 9760 12557
rect 9786 12531 9822 12557
rect 9848 12531 9884 12557
rect 9910 12531 9946 12557
rect 9972 12531 10008 12557
rect 10034 12531 14574 12557
rect 14600 12531 14636 12557
rect 14662 12531 14698 12557
rect 14724 12531 14760 12557
rect 14786 12531 14822 12557
rect 14848 12531 14884 12557
rect 14910 12531 14946 12557
rect 14972 12531 15008 12557
rect 15034 12531 19574 12557
rect 19600 12531 19636 12557
rect 19662 12531 19698 12557
rect 19724 12531 19760 12557
rect 19786 12531 19822 12557
rect 19848 12531 19884 12557
rect 19910 12531 19946 12557
rect 19972 12531 20008 12557
rect 20034 12531 24574 12557
rect 24600 12531 24636 12557
rect 24662 12531 24698 12557
rect 24724 12531 24760 12557
rect 24786 12531 24822 12557
rect 24848 12531 24884 12557
rect 24910 12531 24946 12557
rect 24972 12531 25008 12557
rect 25034 12531 29574 12557
rect 29600 12531 29636 12557
rect 29662 12531 29698 12557
rect 29724 12531 29760 12557
rect 29786 12531 29822 12557
rect 29848 12531 29884 12557
rect 29910 12531 29946 12557
rect 29972 12531 30008 12557
rect 30034 12531 34574 12557
rect 34600 12531 34636 12557
rect 34662 12531 34698 12557
rect 34724 12531 34760 12557
rect 34786 12531 34822 12557
rect 34848 12531 34884 12557
rect 34910 12531 34946 12557
rect 34972 12531 35008 12557
rect 35034 12531 39312 12557
rect 672 12514 39312 12531
rect 3033 12391 3039 12417
rect 3065 12391 3071 12417
rect 4489 12391 4495 12417
rect 4521 12391 4527 12417
rect 7009 12391 7015 12417
rect 7041 12391 7047 12417
rect 8353 12391 8359 12417
rect 8385 12391 8391 12417
rect 14961 12391 14967 12417
rect 14993 12391 14999 12417
rect 16417 12391 16423 12417
rect 16449 12391 16455 12417
rect 17873 12391 17879 12417
rect 17905 12391 17911 12417
rect 19441 12391 19447 12417
rect 19473 12391 19479 12417
rect 23417 12391 23423 12417
rect 23449 12391 23455 12417
rect 27169 12391 27175 12417
rect 27201 12391 27207 12417
rect 29689 12391 29695 12417
rect 29721 12391 29727 12417
rect 31145 12391 31151 12417
rect 31177 12391 31183 12417
rect 1913 12335 1919 12361
rect 1945 12335 1951 12361
rect 3033 12335 3039 12361
rect 3065 12335 3071 12361
rect 3593 12335 3599 12361
rect 3625 12335 3631 12361
rect 4489 12335 4495 12361
rect 4521 12335 4527 12361
rect 6113 12335 6119 12361
rect 6145 12335 6151 12361
rect 7009 12335 7015 12361
rect 7041 12335 7047 12361
rect 7569 12335 7575 12361
rect 7601 12335 7607 12361
rect 8353 12335 8359 12361
rect 8385 12335 8391 12361
rect 10089 12335 10095 12361
rect 10121 12335 10127 12361
rect 10369 12335 10375 12361
rect 10401 12335 10407 12361
rect 10481 12335 10487 12361
rect 10513 12335 10519 12361
rect 11265 12335 11271 12361
rect 11297 12335 11303 12361
rect 11825 12335 11831 12361
rect 11857 12335 11863 12361
rect 11993 12335 11999 12361
rect 12025 12335 12031 12361
rect 14065 12335 14071 12361
rect 14097 12335 14103 12361
rect 14961 12335 14967 12361
rect 14993 12335 14999 12361
rect 15521 12335 15527 12361
rect 15553 12335 15559 12361
rect 16417 12335 16423 12361
rect 16449 12335 16455 12361
rect 16921 12335 16927 12361
rect 16953 12335 16959 12361
rect 17873 12335 17879 12361
rect 17905 12335 17911 12361
rect 18545 12335 18551 12361
rect 18577 12335 18583 12361
rect 19441 12335 19447 12361
rect 19473 12335 19479 12361
rect 20953 12335 20959 12361
rect 20985 12335 20991 12361
rect 21233 12335 21239 12361
rect 21265 12335 21271 12361
rect 21457 12335 21463 12361
rect 21489 12335 21495 12361
rect 22521 12335 22527 12361
rect 22553 12335 22559 12361
rect 23417 12335 23423 12361
rect 23449 12335 23455 12361
rect 24761 12335 24767 12361
rect 24793 12335 24799 12361
rect 25209 12335 25215 12361
rect 25241 12335 25247 12361
rect 25433 12335 25439 12361
rect 25465 12335 25471 12361
rect 26497 12335 26503 12361
rect 26529 12335 26535 12361
rect 26889 12335 26895 12361
rect 26921 12335 26927 12361
rect 29017 12335 29023 12361
rect 29049 12335 29055 12361
rect 29465 12335 29471 12361
rect 29497 12335 29503 12361
rect 30473 12335 30479 12361
rect 30505 12335 30511 12361
rect 31089 12335 31095 12361
rect 31121 12335 31127 12361
rect 672 12165 39312 12182
rect 672 12139 2074 12165
rect 2100 12139 2136 12165
rect 2162 12139 2198 12165
rect 2224 12139 2260 12165
rect 2286 12139 2322 12165
rect 2348 12139 2384 12165
rect 2410 12139 2446 12165
rect 2472 12139 2508 12165
rect 2534 12139 7074 12165
rect 7100 12139 7136 12165
rect 7162 12139 7198 12165
rect 7224 12139 7260 12165
rect 7286 12139 7322 12165
rect 7348 12139 7384 12165
rect 7410 12139 7446 12165
rect 7472 12139 7508 12165
rect 7534 12139 12074 12165
rect 12100 12139 12136 12165
rect 12162 12139 12198 12165
rect 12224 12139 12260 12165
rect 12286 12139 12322 12165
rect 12348 12139 12384 12165
rect 12410 12139 12446 12165
rect 12472 12139 12508 12165
rect 12534 12139 17074 12165
rect 17100 12139 17136 12165
rect 17162 12139 17198 12165
rect 17224 12139 17260 12165
rect 17286 12139 17322 12165
rect 17348 12139 17384 12165
rect 17410 12139 17446 12165
rect 17472 12139 17508 12165
rect 17534 12139 22074 12165
rect 22100 12139 22136 12165
rect 22162 12139 22198 12165
rect 22224 12139 22260 12165
rect 22286 12139 22322 12165
rect 22348 12139 22384 12165
rect 22410 12139 22446 12165
rect 22472 12139 22508 12165
rect 22534 12139 27074 12165
rect 27100 12139 27136 12165
rect 27162 12139 27198 12165
rect 27224 12139 27260 12165
rect 27286 12139 27322 12165
rect 27348 12139 27384 12165
rect 27410 12139 27446 12165
rect 27472 12139 27508 12165
rect 27534 12139 32074 12165
rect 32100 12139 32136 12165
rect 32162 12139 32198 12165
rect 32224 12139 32260 12165
rect 32286 12139 32322 12165
rect 32348 12139 32384 12165
rect 32410 12139 32446 12165
rect 32472 12139 32508 12165
rect 32534 12139 37074 12165
rect 37100 12139 37136 12165
rect 37162 12139 37198 12165
rect 37224 12139 37260 12165
rect 37286 12139 37322 12165
rect 37348 12139 37384 12165
rect 37410 12139 37446 12165
rect 37472 12139 37508 12165
rect 37534 12139 39312 12165
rect 672 12122 39312 12139
rect 1577 11943 1583 11969
rect 1609 11943 1615 11969
rect 2473 11943 2479 11969
rect 2505 11943 2511 11969
rect 3817 11943 3823 11969
rect 3849 11943 3855 11969
rect 4993 11943 4999 11969
rect 5025 11943 5031 11969
rect 5553 11943 5559 11969
rect 5585 11943 5591 11969
rect 6449 11943 6455 11969
rect 6481 11943 6487 11969
rect 8073 11943 8079 11969
rect 8105 11943 8111 11969
rect 8969 11943 8975 11969
rect 9001 11943 9007 11969
rect 9529 11943 9535 11969
rect 9561 11943 9567 11969
rect 9697 11943 9703 11969
rect 9729 11943 9735 11969
rect 10369 11943 10375 11969
rect 10401 11943 10407 11969
rect 11769 11943 11775 11969
rect 11801 11943 11807 11969
rect 12217 11943 12223 11969
rect 12249 11943 12255 11969
rect 12441 11943 12447 11969
rect 12473 11943 12479 11969
rect 13225 11943 13231 11969
rect 13257 11943 13263 11969
rect 14401 11943 14407 11969
rect 14433 11943 14439 11969
rect 15857 11943 15863 11969
rect 15889 11943 15895 11969
rect 16753 11943 16759 11969
rect 16785 11943 16791 11969
rect 17033 11943 17039 11969
rect 17065 11943 17071 11969
rect 17873 11943 17879 11969
rect 17905 11943 17911 11969
rect 18769 11943 18775 11969
rect 18801 11943 18807 11969
rect 19945 11943 19951 11969
rect 19977 11943 19983 11969
rect 20505 11943 20511 11969
rect 20537 11943 20543 11969
rect 21177 11943 21183 11969
rect 21209 11943 21215 11969
rect 22801 11943 22807 11969
rect 22833 11943 22839 11969
rect 23921 11943 23927 11969
rect 23953 11943 23959 11969
rect 24369 11943 24375 11969
rect 24401 11943 24407 11969
rect 25153 11943 25159 11969
rect 25185 11943 25191 11969
rect 27001 11943 27007 11969
rect 27033 11943 27039 11969
rect 27561 11943 27567 11969
rect 27593 11943 27599 11969
rect 28457 11943 28463 11969
rect 28489 11943 28495 11969
rect 28961 11943 28967 11969
rect 28993 11943 28999 11969
rect 30977 11943 30983 11969
rect 31009 11943 31015 11969
rect 31145 11943 31151 11969
rect 31177 11943 31183 11969
rect 31369 11943 31375 11969
rect 31401 11943 31407 11969
rect 32153 11943 32159 11969
rect 32185 11943 32191 11969
rect 32825 11943 32831 11969
rect 32857 11943 32863 11969
rect 2473 11887 2479 11913
rect 2505 11887 2511 11913
rect 4993 11887 4999 11913
rect 5025 11887 5031 11913
rect 6449 11887 6455 11913
rect 6481 11887 6487 11913
rect 8969 11887 8975 11913
rect 9001 11887 9007 11913
rect 14401 11887 14407 11913
rect 14433 11887 14439 11913
rect 16753 11887 16759 11913
rect 16785 11887 16791 11913
rect 17985 11887 17991 11913
rect 18017 11887 18023 11913
rect 19945 11887 19951 11913
rect 19977 11887 19983 11913
rect 21177 11887 21183 11913
rect 21209 11887 21215 11913
rect 23921 11887 23927 11913
rect 23953 11887 23959 11913
rect 25153 11887 25159 11913
rect 25185 11887 25191 11913
rect 27673 11887 27679 11913
rect 27705 11887 27711 11913
rect 29129 11887 29135 11913
rect 29161 11887 29167 11913
rect 33105 11887 33111 11913
rect 33137 11887 33143 11913
rect 672 11773 39312 11790
rect 672 11747 4574 11773
rect 4600 11747 4636 11773
rect 4662 11747 4698 11773
rect 4724 11747 4760 11773
rect 4786 11747 4822 11773
rect 4848 11747 4884 11773
rect 4910 11747 4946 11773
rect 4972 11747 5008 11773
rect 5034 11747 9574 11773
rect 9600 11747 9636 11773
rect 9662 11747 9698 11773
rect 9724 11747 9760 11773
rect 9786 11747 9822 11773
rect 9848 11747 9884 11773
rect 9910 11747 9946 11773
rect 9972 11747 10008 11773
rect 10034 11747 14574 11773
rect 14600 11747 14636 11773
rect 14662 11747 14698 11773
rect 14724 11747 14760 11773
rect 14786 11747 14822 11773
rect 14848 11747 14884 11773
rect 14910 11747 14946 11773
rect 14972 11747 15008 11773
rect 15034 11747 19574 11773
rect 19600 11747 19636 11773
rect 19662 11747 19698 11773
rect 19724 11747 19760 11773
rect 19786 11747 19822 11773
rect 19848 11747 19884 11773
rect 19910 11747 19946 11773
rect 19972 11747 20008 11773
rect 20034 11747 24574 11773
rect 24600 11747 24636 11773
rect 24662 11747 24698 11773
rect 24724 11747 24760 11773
rect 24786 11747 24822 11773
rect 24848 11747 24884 11773
rect 24910 11747 24946 11773
rect 24972 11747 25008 11773
rect 25034 11747 29574 11773
rect 29600 11747 29636 11773
rect 29662 11747 29698 11773
rect 29724 11747 29760 11773
rect 29786 11747 29822 11773
rect 29848 11747 29884 11773
rect 29910 11747 29946 11773
rect 29972 11747 30008 11773
rect 30034 11747 34574 11773
rect 34600 11747 34636 11773
rect 34662 11747 34698 11773
rect 34724 11747 34760 11773
rect 34786 11747 34822 11773
rect 34848 11747 34884 11773
rect 34910 11747 34946 11773
rect 34972 11747 35008 11773
rect 35034 11747 39312 11773
rect 672 11730 39312 11747
rect 3033 11607 3039 11633
rect 3065 11607 3071 11633
rect 4489 11607 4495 11633
rect 4521 11607 4527 11633
rect 8465 11607 8471 11633
rect 8497 11607 8503 11633
rect 14961 11607 14967 11633
rect 14993 11607 14999 11633
rect 16193 11607 16199 11633
rect 16225 11607 16231 11633
rect 17985 11607 17991 11633
rect 18017 11607 18023 11633
rect 19329 11607 19335 11633
rect 19361 11607 19367 11633
rect 23305 11607 23311 11633
rect 23337 11607 23343 11633
rect 29913 11607 29919 11633
rect 29945 11607 29951 11633
rect 31369 11607 31375 11633
rect 31401 11607 31407 11633
rect 33889 11607 33895 11633
rect 33921 11607 33927 11633
rect 1913 11551 1919 11577
rect 1945 11551 1951 11577
rect 3033 11551 3039 11577
rect 3065 11551 3071 11577
rect 3593 11551 3599 11577
rect 3625 11551 3631 11577
rect 4489 11551 4495 11577
rect 4521 11551 4527 11577
rect 5833 11551 5839 11577
rect 5865 11551 5871 11577
rect 6393 11551 6399 11577
rect 6425 11551 6431 11577
rect 6505 11551 6511 11577
rect 6537 11551 6543 11577
rect 7569 11551 7575 11577
rect 7601 11551 7607 11577
rect 8465 11551 8471 11577
rect 8497 11551 8503 11577
rect 9809 11551 9815 11577
rect 9841 11551 9847 11577
rect 10369 11551 10375 11577
rect 10401 11551 10407 11577
rect 10481 11551 10487 11577
rect 10513 11551 10519 11577
rect 11321 11551 11327 11577
rect 11353 11551 11359 11577
rect 11825 11551 11831 11577
rect 11857 11551 11863 11577
rect 11993 11551 11999 11577
rect 12025 11551 12031 11577
rect 14065 11551 14071 11577
rect 14097 11551 14103 11577
rect 14961 11551 14967 11577
rect 14993 11551 14999 11577
rect 15465 11551 15471 11577
rect 15497 11551 15503 11577
rect 16193 11551 16199 11577
rect 16225 11551 16231 11577
rect 16977 11551 16983 11577
rect 17009 11551 17015 11577
rect 17985 11551 17991 11577
rect 18017 11551 18023 11577
rect 18545 11551 18551 11577
rect 18577 11551 18583 11577
rect 19329 11551 19335 11577
rect 19361 11551 19367 11577
rect 20953 11551 20959 11577
rect 20985 11551 20991 11577
rect 21233 11551 21239 11577
rect 21265 11551 21271 11577
rect 21457 11551 21463 11577
rect 21489 11551 21495 11577
rect 22521 11551 22527 11577
rect 22553 11551 22559 11577
rect 23305 11551 23311 11577
rect 23337 11551 23343 11577
rect 24761 11551 24767 11577
rect 24793 11551 24799 11577
rect 25321 11551 25327 11577
rect 25353 11551 25359 11577
rect 25433 11551 25439 11577
rect 25465 11551 25471 11577
rect 26721 11551 26727 11577
rect 26753 11551 26759 11577
rect 26945 11551 26951 11577
rect 26977 11551 26983 11577
rect 27393 11551 27399 11577
rect 27425 11551 27431 11577
rect 29017 11551 29023 11577
rect 29049 11551 29055 11577
rect 29913 11551 29919 11577
rect 29945 11551 29951 11577
rect 30473 11551 30479 11577
rect 30505 11551 30511 11577
rect 31369 11551 31375 11577
rect 31401 11551 31407 11577
rect 32769 11551 32775 11577
rect 32801 11551 32807 11577
rect 33889 11551 33895 11577
rect 33921 11551 33927 11577
rect 672 11381 39312 11398
rect 672 11355 2074 11381
rect 2100 11355 2136 11381
rect 2162 11355 2198 11381
rect 2224 11355 2260 11381
rect 2286 11355 2322 11381
rect 2348 11355 2384 11381
rect 2410 11355 2446 11381
rect 2472 11355 2508 11381
rect 2534 11355 7074 11381
rect 7100 11355 7136 11381
rect 7162 11355 7198 11381
rect 7224 11355 7260 11381
rect 7286 11355 7322 11381
rect 7348 11355 7384 11381
rect 7410 11355 7446 11381
rect 7472 11355 7508 11381
rect 7534 11355 12074 11381
rect 12100 11355 12136 11381
rect 12162 11355 12198 11381
rect 12224 11355 12260 11381
rect 12286 11355 12322 11381
rect 12348 11355 12384 11381
rect 12410 11355 12446 11381
rect 12472 11355 12508 11381
rect 12534 11355 17074 11381
rect 17100 11355 17136 11381
rect 17162 11355 17198 11381
rect 17224 11355 17260 11381
rect 17286 11355 17322 11381
rect 17348 11355 17384 11381
rect 17410 11355 17446 11381
rect 17472 11355 17508 11381
rect 17534 11355 22074 11381
rect 22100 11355 22136 11381
rect 22162 11355 22198 11381
rect 22224 11355 22260 11381
rect 22286 11355 22322 11381
rect 22348 11355 22384 11381
rect 22410 11355 22446 11381
rect 22472 11355 22508 11381
rect 22534 11355 27074 11381
rect 27100 11355 27136 11381
rect 27162 11355 27198 11381
rect 27224 11355 27260 11381
rect 27286 11355 27322 11381
rect 27348 11355 27384 11381
rect 27410 11355 27446 11381
rect 27472 11355 27508 11381
rect 27534 11355 32074 11381
rect 32100 11355 32136 11381
rect 32162 11355 32198 11381
rect 32224 11355 32260 11381
rect 32286 11355 32322 11381
rect 32348 11355 32384 11381
rect 32410 11355 32446 11381
rect 32472 11355 32508 11381
rect 32534 11355 37074 11381
rect 37100 11355 37136 11381
rect 37162 11355 37198 11381
rect 37224 11355 37260 11381
rect 37286 11355 37322 11381
rect 37348 11355 37384 11381
rect 37410 11355 37446 11381
rect 37472 11355 37508 11381
rect 37534 11355 39312 11381
rect 672 11338 39312 11355
rect 1577 11159 1583 11185
rect 1609 11159 1615 11185
rect 2473 11159 2479 11185
rect 2505 11159 2511 11185
rect 3817 11159 3823 11185
rect 3849 11159 3855 11185
rect 4993 11159 4999 11185
rect 5025 11159 5031 11185
rect 5553 11159 5559 11185
rect 5585 11159 5591 11185
rect 6393 11159 6399 11185
rect 6425 11159 6431 11185
rect 8073 11159 8079 11185
rect 8105 11159 8111 11185
rect 8969 11159 8975 11185
rect 9001 11159 9007 11185
rect 9473 11159 9479 11185
rect 9505 11159 9511 11185
rect 10369 11159 10375 11185
rect 10401 11159 10407 11185
rect 11769 11159 11775 11185
rect 11801 11159 11807 11185
rect 12945 11159 12951 11185
rect 12977 11159 12983 11185
rect 13505 11159 13511 11185
rect 13537 11159 13543 11185
rect 14401 11159 14407 11185
rect 14433 11159 14439 11185
rect 15689 11159 15695 11185
rect 15721 11159 15727 11185
rect 16193 11159 16199 11185
rect 16225 11159 16231 11185
rect 16305 11159 16311 11185
rect 16337 11159 16343 11185
rect 17089 11159 17095 11185
rect 17121 11159 17127 11185
rect 17985 11159 17991 11185
rect 18017 11159 18023 11185
rect 18769 11159 18775 11185
rect 18801 11159 18807 11185
rect 19329 11159 19335 11185
rect 19361 11159 19367 11185
rect 19497 11159 19503 11185
rect 19529 11159 19535 11185
rect 20505 11159 20511 11185
rect 20537 11159 20543 11185
rect 21009 11159 21015 11185
rect 21041 11159 21047 11185
rect 22745 11159 22751 11185
rect 22777 11159 22783 11185
rect 23305 11159 23311 11185
rect 23337 11159 23343 11185
rect 23417 11159 23423 11185
rect 23449 11159 23455 11185
rect 24369 11159 24375 11185
rect 24401 11159 24407 11185
rect 25153 11159 25159 11185
rect 25185 11159 25191 11185
rect 27225 11159 27231 11185
rect 27257 11159 27263 11185
rect 27449 11159 27455 11185
rect 27481 11159 27487 11185
rect 27841 11159 27847 11185
rect 27873 11159 27879 11185
rect 28457 11159 28463 11185
rect 28489 11159 28495 11185
rect 28625 11159 28631 11185
rect 28657 11159 28663 11185
rect 28849 11159 28855 11185
rect 28881 11159 28887 11185
rect 30697 11159 30703 11185
rect 30729 11159 30735 11185
rect 31257 11159 31263 11185
rect 31289 11159 31295 11185
rect 31369 11159 31375 11185
rect 31401 11159 31407 11185
rect 32433 11159 32439 11185
rect 32465 11159 32471 11185
rect 33105 11159 33111 11185
rect 33137 11159 33143 11185
rect 34953 11159 34959 11185
rect 34985 11159 34991 11185
rect 35233 11159 35239 11185
rect 35265 11159 35271 11185
rect 35849 11159 35855 11185
rect 35881 11159 35887 11185
rect 36185 11159 36191 11185
rect 36217 11159 36223 11185
rect 36689 11159 36695 11185
rect 36721 11159 36727 11185
rect 36801 11159 36807 11185
rect 36833 11159 36839 11185
rect 2473 11103 2479 11129
rect 2505 11103 2511 11129
rect 4993 11103 4999 11129
rect 5025 11103 5031 11129
rect 6393 11103 6399 11129
rect 6425 11103 6431 11129
rect 8969 11103 8975 11129
rect 9001 11103 9007 11129
rect 10369 11103 10375 11129
rect 10401 11103 10407 11129
rect 12945 11103 12951 11129
rect 12977 11103 12983 11129
rect 14401 11103 14407 11129
rect 14433 11103 14439 11129
rect 18041 11103 18047 11129
rect 18073 11103 18079 11129
rect 21177 11103 21183 11129
rect 21209 11103 21215 11129
rect 25153 11103 25159 11129
rect 25185 11103 25191 11129
rect 33105 11103 33111 11129
rect 33137 11103 33143 11129
rect 672 10989 39312 11006
rect 672 10963 4574 10989
rect 4600 10963 4636 10989
rect 4662 10963 4698 10989
rect 4724 10963 4760 10989
rect 4786 10963 4822 10989
rect 4848 10963 4884 10989
rect 4910 10963 4946 10989
rect 4972 10963 5008 10989
rect 5034 10963 9574 10989
rect 9600 10963 9636 10989
rect 9662 10963 9698 10989
rect 9724 10963 9760 10989
rect 9786 10963 9822 10989
rect 9848 10963 9884 10989
rect 9910 10963 9946 10989
rect 9972 10963 10008 10989
rect 10034 10963 14574 10989
rect 14600 10963 14636 10989
rect 14662 10963 14698 10989
rect 14724 10963 14760 10989
rect 14786 10963 14822 10989
rect 14848 10963 14884 10989
rect 14910 10963 14946 10989
rect 14972 10963 15008 10989
rect 15034 10963 19574 10989
rect 19600 10963 19636 10989
rect 19662 10963 19698 10989
rect 19724 10963 19760 10989
rect 19786 10963 19822 10989
rect 19848 10963 19884 10989
rect 19910 10963 19946 10989
rect 19972 10963 20008 10989
rect 20034 10963 24574 10989
rect 24600 10963 24636 10989
rect 24662 10963 24698 10989
rect 24724 10963 24760 10989
rect 24786 10963 24822 10989
rect 24848 10963 24884 10989
rect 24910 10963 24946 10989
rect 24972 10963 25008 10989
rect 25034 10963 29574 10989
rect 29600 10963 29636 10989
rect 29662 10963 29698 10989
rect 29724 10963 29760 10989
rect 29786 10963 29822 10989
rect 29848 10963 29884 10989
rect 29910 10963 29946 10989
rect 29972 10963 30008 10989
rect 30034 10963 34574 10989
rect 34600 10963 34636 10989
rect 34662 10963 34698 10989
rect 34724 10963 34760 10989
rect 34786 10963 34822 10989
rect 34848 10963 34884 10989
rect 34910 10963 34946 10989
rect 34972 10963 35008 10989
rect 35034 10963 39312 10989
rect 672 10946 39312 10963
rect 3033 10823 3039 10849
rect 3065 10823 3071 10849
rect 4489 10823 4495 10849
rect 4521 10823 4527 10849
rect 8297 10823 8303 10849
rect 8329 10823 8335 10849
rect 16193 10823 16199 10849
rect 16225 10823 16231 10849
rect 17985 10823 17991 10849
rect 18017 10823 18023 10849
rect 19441 10823 19447 10849
rect 19473 10823 19479 10849
rect 21737 10823 21743 10849
rect 21769 10823 21775 10849
rect 23361 10823 23367 10849
rect 23393 10823 23399 10849
rect 25937 10823 25943 10849
rect 25969 10823 25975 10849
rect 27281 10823 27287 10849
rect 27313 10823 27319 10849
rect 29913 10823 29919 10849
rect 29945 10823 29951 10849
rect 31145 10823 31151 10849
rect 31177 10823 31183 10849
rect 33889 10823 33895 10849
rect 33921 10823 33927 10849
rect 35345 10823 35351 10849
rect 35377 10823 35383 10849
rect 1913 10767 1919 10793
rect 1945 10767 1951 10793
rect 3033 10767 3039 10793
rect 3065 10767 3071 10793
rect 3593 10767 3599 10793
rect 3625 10767 3631 10793
rect 4489 10767 4495 10793
rect 4521 10767 4527 10793
rect 5833 10767 5839 10793
rect 5865 10767 5871 10793
rect 6393 10767 6399 10793
rect 6425 10767 6431 10793
rect 6505 10767 6511 10793
rect 6537 10767 6543 10793
rect 7569 10767 7575 10793
rect 7601 10767 7607 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 9809 10767 9815 10793
rect 9841 10767 9847 10793
rect 10369 10767 10375 10793
rect 10401 10767 10407 10793
rect 10481 10767 10487 10793
rect 10513 10767 10519 10793
rect 11321 10767 11327 10793
rect 11353 10767 11359 10793
rect 11825 10767 11831 10793
rect 11857 10767 11863 10793
rect 11993 10767 11999 10793
rect 12025 10767 12031 10793
rect 14065 10767 14071 10793
rect 14097 10767 14103 10793
rect 14345 10767 14351 10793
rect 14377 10767 14383 10793
rect 14457 10767 14463 10793
rect 14489 10767 14495 10793
rect 15465 10767 15471 10793
rect 15497 10767 15503 10793
rect 16137 10767 16143 10793
rect 16169 10767 16175 10793
rect 16977 10767 16983 10793
rect 17009 10767 17015 10793
rect 17985 10767 17991 10793
rect 18017 10767 18023 10793
rect 18545 10767 18551 10793
rect 18577 10767 18583 10793
rect 19441 10767 19447 10793
rect 19473 10767 19479 10793
rect 20785 10767 20791 10793
rect 20817 10767 20823 10793
rect 21737 10767 21743 10793
rect 21769 10767 21775 10793
rect 22521 10767 22527 10793
rect 22553 10767 22559 10793
rect 23361 10767 23367 10793
rect 23393 10767 23399 10793
rect 24761 10767 24767 10793
rect 24793 10767 24799 10793
rect 25937 10767 25943 10793
rect 25969 10767 25975 10793
rect 26217 10767 26223 10793
rect 26249 10767 26255 10793
rect 27281 10767 27287 10793
rect 27313 10767 27319 10793
rect 29017 10767 29023 10793
rect 29049 10767 29055 10793
rect 29913 10767 29919 10793
rect 29945 10767 29951 10793
rect 30249 10767 30255 10793
rect 30281 10767 30287 10793
rect 31089 10767 31095 10793
rect 31121 10767 31127 10793
rect 32993 10767 32999 10793
rect 33025 10767 33031 10793
rect 33889 10767 33895 10793
rect 33921 10767 33927 10793
rect 34225 10767 34231 10793
rect 34257 10767 34263 10793
rect 35345 10767 35351 10793
rect 35377 10767 35383 10793
rect 672 10597 39312 10614
rect 672 10571 2074 10597
rect 2100 10571 2136 10597
rect 2162 10571 2198 10597
rect 2224 10571 2260 10597
rect 2286 10571 2322 10597
rect 2348 10571 2384 10597
rect 2410 10571 2446 10597
rect 2472 10571 2508 10597
rect 2534 10571 7074 10597
rect 7100 10571 7136 10597
rect 7162 10571 7198 10597
rect 7224 10571 7260 10597
rect 7286 10571 7322 10597
rect 7348 10571 7384 10597
rect 7410 10571 7446 10597
rect 7472 10571 7508 10597
rect 7534 10571 12074 10597
rect 12100 10571 12136 10597
rect 12162 10571 12198 10597
rect 12224 10571 12260 10597
rect 12286 10571 12322 10597
rect 12348 10571 12384 10597
rect 12410 10571 12446 10597
rect 12472 10571 12508 10597
rect 12534 10571 17074 10597
rect 17100 10571 17136 10597
rect 17162 10571 17198 10597
rect 17224 10571 17260 10597
rect 17286 10571 17322 10597
rect 17348 10571 17384 10597
rect 17410 10571 17446 10597
rect 17472 10571 17508 10597
rect 17534 10571 22074 10597
rect 22100 10571 22136 10597
rect 22162 10571 22198 10597
rect 22224 10571 22260 10597
rect 22286 10571 22322 10597
rect 22348 10571 22384 10597
rect 22410 10571 22446 10597
rect 22472 10571 22508 10597
rect 22534 10571 27074 10597
rect 27100 10571 27136 10597
rect 27162 10571 27198 10597
rect 27224 10571 27260 10597
rect 27286 10571 27322 10597
rect 27348 10571 27384 10597
rect 27410 10571 27446 10597
rect 27472 10571 27508 10597
rect 27534 10571 32074 10597
rect 32100 10571 32136 10597
rect 32162 10571 32198 10597
rect 32224 10571 32260 10597
rect 32286 10571 32322 10597
rect 32348 10571 32384 10597
rect 32410 10571 32446 10597
rect 32472 10571 32508 10597
rect 32534 10571 37074 10597
rect 37100 10571 37136 10597
rect 37162 10571 37198 10597
rect 37224 10571 37260 10597
rect 37286 10571 37322 10597
rect 37348 10571 37384 10597
rect 37410 10571 37446 10597
rect 37472 10571 37508 10597
rect 37534 10571 39312 10597
rect 672 10554 39312 10571
rect 1577 10375 1583 10401
rect 1609 10375 1615 10401
rect 2473 10375 2479 10401
rect 2505 10375 2511 10401
rect 3817 10375 3823 10401
rect 3849 10375 3855 10401
rect 4993 10375 4999 10401
rect 5025 10375 5031 10401
rect 5553 10375 5559 10401
rect 5585 10375 5591 10401
rect 6449 10375 6455 10401
rect 6481 10375 6487 10401
rect 7793 10375 7799 10401
rect 7825 10375 7831 10401
rect 8297 10375 8303 10401
rect 8329 10375 8335 10401
rect 8465 10375 8471 10401
rect 8497 10375 8503 10401
rect 9473 10375 9479 10401
rect 9505 10375 9511 10401
rect 10369 10375 10375 10401
rect 10401 10375 10407 10401
rect 11881 10375 11887 10401
rect 11913 10375 11919 10401
rect 12945 10375 12951 10401
rect 12977 10375 12983 10401
rect 13505 10375 13511 10401
rect 13537 10375 13543 10401
rect 14401 10375 14407 10401
rect 14433 10375 14439 10401
rect 15689 10375 15695 10401
rect 15721 10375 15727 10401
rect 16137 10375 16143 10401
rect 16169 10375 16175 10401
rect 16361 10375 16367 10401
rect 16393 10375 16399 10401
rect 17145 10375 17151 10401
rect 17177 10375 17183 10401
rect 17985 10375 17991 10401
rect 18017 10375 18023 10401
rect 18769 10375 18775 10401
rect 18801 10375 18807 10401
rect 19945 10375 19951 10401
rect 19977 10375 19983 10401
rect 20225 10375 20231 10401
rect 20257 10375 20263 10401
rect 21401 10375 21407 10401
rect 21433 10375 21439 10401
rect 22745 10375 22751 10401
rect 22777 10375 22783 10401
rect 23697 10375 23703 10401
rect 23729 10375 23735 10401
rect 24481 10375 24487 10401
rect 24513 10375 24519 10401
rect 25377 10375 25383 10401
rect 25409 10375 25415 10401
rect 26721 10375 26727 10401
rect 26753 10375 26759 10401
rect 27561 10375 27567 10401
rect 27593 10375 27599 10401
rect 28177 10375 28183 10401
rect 28209 10375 28215 10401
rect 29129 10375 29135 10401
rect 29161 10375 29167 10401
rect 30697 10375 30703 10401
rect 30729 10375 30735 10401
rect 31649 10375 31655 10401
rect 31681 10375 31687 10401
rect 32153 10375 32159 10401
rect 32185 10375 32191 10401
rect 33105 10375 33111 10401
rect 33137 10375 33143 10401
rect 34673 10375 34679 10401
rect 34705 10375 34711 10401
rect 35625 10375 35631 10401
rect 35657 10375 35663 10401
rect 36129 10375 36135 10401
rect 36161 10375 36167 10401
rect 36689 10375 36695 10401
rect 36721 10375 36727 10401
rect 36857 10375 36863 10401
rect 36889 10375 36895 10401
rect 2473 10319 2479 10345
rect 2505 10319 2511 10345
rect 4993 10319 4999 10345
rect 5025 10319 5031 10345
rect 6449 10319 6455 10345
rect 6481 10319 6487 10345
rect 10369 10319 10375 10345
rect 10401 10319 10407 10345
rect 12945 10319 12951 10345
rect 12977 10319 12983 10345
rect 14401 10319 14407 10345
rect 14433 10319 14439 10345
rect 18097 10319 18103 10345
rect 18129 10319 18135 10345
rect 19945 10319 19951 10345
rect 19977 10319 19983 10345
rect 21401 10319 21407 10345
rect 21433 10319 21439 10345
rect 23697 10319 23703 10345
rect 23729 10319 23735 10345
rect 25377 10319 25383 10345
rect 25409 10319 25415 10345
rect 27673 10319 27679 10345
rect 27705 10319 27711 10345
rect 29129 10319 29135 10345
rect 29161 10319 29167 10345
rect 31649 10319 31655 10345
rect 31681 10319 31687 10345
rect 33105 10319 33111 10345
rect 33137 10319 33143 10345
rect 35625 10319 35631 10345
rect 35657 10319 35663 10345
rect 672 10205 39312 10222
rect 672 10179 4574 10205
rect 4600 10179 4636 10205
rect 4662 10179 4698 10205
rect 4724 10179 4760 10205
rect 4786 10179 4822 10205
rect 4848 10179 4884 10205
rect 4910 10179 4946 10205
rect 4972 10179 5008 10205
rect 5034 10179 9574 10205
rect 9600 10179 9636 10205
rect 9662 10179 9698 10205
rect 9724 10179 9760 10205
rect 9786 10179 9822 10205
rect 9848 10179 9884 10205
rect 9910 10179 9946 10205
rect 9972 10179 10008 10205
rect 10034 10179 14574 10205
rect 14600 10179 14636 10205
rect 14662 10179 14698 10205
rect 14724 10179 14760 10205
rect 14786 10179 14822 10205
rect 14848 10179 14884 10205
rect 14910 10179 14946 10205
rect 14972 10179 15008 10205
rect 15034 10179 19574 10205
rect 19600 10179 19636 10205
rect 19662 10179 19698 10205
rect 19724 10179 19760 10205
rect 19786 10179 19822 10205
rect 19848 10179 19884 10205
rect 19910 10179 19946 10205
rect 19972 10179 20008 10205
rect 20034 10179 24574 10205
rect 24600 10179 24636 10205
rect 24662 10179 24698 10205
rect 24724 10179 24760 10205
rect 24786 10179 24822 10205
rect 24848 10179 24884 10205
rect 24910 10179 24946 10205
rect 24972 10179 25008 10205
rect 25034 10179 29574 10205
rect 29600 10179 29636 10205
rect 29662 10179 29698 10205
rect 29724 10179 29760 10205
rect 29786 10179 29822 10205
rect 29848 10179 29884 10205
rect 29910 10179 29946 10205
rect 29972 10179 30008 10205
rect 30034 10179 34574 10205
rect 34600 10179 34636 10205
rect 34662 10179 34698 10205
rect 34724 10179 34760 10205
rect 34786 10179 34822 10205
rect 34848 10179 34884 10205
rect 34910 10179 34946 10205
rect 34972 10179 35008 10205
rect 35034 10179 39312 10205
rect 672 10162 39312 10179
rect 3033 10039 3039 10065
rect 3065 10039 3071 10065
rect 4489 10039 4495 10065
rect 4521 10039 4527 10065
rect 7009 10039 7015 10065
rect 7041 10039 7047 10065
rect 8353 10039 8359 10065
rect 8385 10039 8391 10065
rect 12441 10039 12447 10065
rect 12473 10039 12479 10065
rect 17985 10039 17991 10065
rect 18017 10039 18023 10065
rect 21737 10039 21743 10065
rect 21769 10039 21775 10065
rect 25937 10039 25943 10065
rect 25969 10039 25975 10065
rect 31257 10039 31263 10065
rect 31289 10039 31295 10065
rect 33833 10039 33839 10065
rect 33865 10039 33871 10065
rect 35345 10039 35351 10065
rect 35377 10039 35383 10065
rect 37641 10039 37647 10065
rect 37673 10039 37679 10065
rect 1913 9983 1919 10009
rect 1945 9983 1951 10009
rect 3033 9983 3039 10009
rect 3065 9983 3071 10009
rect 3593 9983 3599 10009
rect 3625 9983 3631 10009
rect 4489 9983 4495 10009
rect 4521 9983 4527 10009
rect 5833 9983 5839 10009
rect 5865 9983 5871 10009
rect 7009 9983 7015 10009
rect 7041 9983 7047 10009
rect 7569 9983 7575 10009
rect 7601 9983 7607 10009
rect 8353 9983 8359 10009
rect 8385 9983 8391 10009
rect 9809 9983 9815 10009
rect 9841 9983 9847 10009
rect 10369 9983 10375 10009
rect 10401 9983 10407 10009
rect 10481 9983 10487 10009
rect 10513 9983 10519 10009
rect 11265 9983 11271 10009
rect 11297 9983 11303 10009
rect 12441 9983 12447 10009
rect 12473 9983 12479 10009
rect 14065 9983 14071 10009
rect 14097 9983 14103 10009
rect 14345 9983 14351 10009
rect 14377 9983 14383 10009
rect 14457 9983 14463 10009
rect 14489 9983 14495 10009
rect 15465 9983 15471 10009
rect 15497 9983 15503 10009
rect 15801 9983 15807 10009
rect 15833 9983 15839 10009
rect 15913 9983 15919 10009
rect 15945 9983 15951 10009
rect 16977 9983 16983 10009
rect 17009 9983 17015 10009
rect 17985 9983 17991 10009
rect 18017 9983 18023 10009
rect 18545 9983 18551 10009
rect 18577 9983 18583 10009
rect 18713 9983 18719 10009
rect 18745 9983 18751 10009
rect 18937 9983 18943 10009
rect 18969 9983 18975 10009
rect 20785 9983 20791 10009
rect 20817 9983 20823 10009
rect 21737 9983 21743 10009
rect 21769 9983 21775 10009
rect 22521 9983 22527 10009
rect 22553 9983 22559 10009
rect 22689 9983 22695 10009
rect 22721 9983 22727 10009
rect 22913 9983 22919 10009
rect 22945 9983 22951 10009
rect 25041 9983 25047 10009
rect 25073 9983 25079 10009
rect 25937 9983 25943 10009
rect 25969 9983 25975 10009
rect 26721 9983 26727 10009
rect 26753 9983 26759 10009
rect 26945 9983 26951 10009
rect 26977 9983 26983 10009
rect 27393 9983 27399 10009
rect 27425 9983 27431 10009
rect 28737 9983 28743 10009
rect 28769 9983 28775 10009
rect 29297 9983 29303 10009
rect 29329 9983 29335 10009
rect 29409 9983 29415 10009
rect 29441 9983 29447 10009
rect 30417 9983 30423 10009
rect 30449 9983 30455 10009
rect 31089 9983 31095 10009
rect 31121 9983 31127 10009
rect 32769 9983 32775 10009
rect 32801 9983 32807 10009
rect 33833 9983 33839 10009
rect 33865 9983 33871 10009
rect 34449 9983 34455 10009
rect 34481 9983 34487 10009
rect 35345 9983 35351 10009
rect 35377 9983 35383 10009
rect 36689 9983 36695 10009
rect 36721 9983 36727 10009
rect 37641 9983 37647 10009
rect 37673 9983 37679 10009
rect 672 9813 39312 9830
rect 672 9787 2074 9813
rect 2100 9787 2136 9813
rect 2162 9787 2198 9813
rect 2224 9787 2260 9813
rect 2286 9787 2322 9813
rect 2348 9787 2384 9813
rect 2410 9787 2446 9813
rect 2472 9787 2508 9813
rect 2534 9787 7074 9813
rect 7100 9787 7136 9813
rect 7162 9787 7198 9813
rect 7224 9787 7260 9813
rect 7286 9787 7322 9813
rect 7348 9787 7384 9813
rect 7410 9787 7446 9813
rect 7472 9787 7508 9813
rect 7534 9787 12074 9813
rect 12100 9787 12136 9813
rect 12162 9787 12198 9813
rect 12224 9787 12260 9813
rect 12286 9787 12322 9813
rect 12348 9787 12384 9813
rect 12410 9787 12446 9813
rect 12472 9787 12508 9813
rect 12534 9787 17074 9813
rect 17100 9787 17136 9813
rect 17162 9787 17198 9813
rect 17224 9787 17260 9813
rect 17286 9787 17322 9813
rect 17348 9787 17384 9813
rect 17410 9787 17446 9813
rect 17472 9787 17508 9813
rect 17534 9787 22074 9813
rect 22100 9787 22136 9813
rect 22162 9787 22198 9813
rect 22224 9787 22260 9813
rect 22286 9787 22322 9813
rect 22348 9787 22384 9813
rect 22410 9787 22446 9813
rect 22472 9787 22508 9813
rect 22534 9787 27074 9813
rect 27100 9787 27136 9813
rect 27162 9787 27198 9813
rect 27224 9787 27260 9813
rect 27286 9787 27322 9813
rect 27348 9787 27384 9813
rect 27410 9787 27446 9813
rect 27472 9787 27508 9813
rect 27534 9787 32074 9813
rect 32100 9787 32136 9813
rect 32162 9787 32198 9813
rect 32224 9787 32260 9813
rect 32286 9787 32322 9813
rect 32348 9787 32384 9813
rect 32410 9787 32446 9813
rect 32472 9787 32508 9813
rect 32534 9787 37074 9813
rect 37100 9787 37136 9813
rect 37162 9787 37198 9813
rect 37224 9787 37260 9813
rect 37286 9787 37322 9813
rect 37348 9787 37384 9813
rect 37410 9787 37446 9813
rect 37472 9787 37508 9813
rect 37534 9787 39312 9813
rect 672 9770 39312 9787
rect 1577 9591 1583 9617
rect 1609 9591 1615 9617
rect 2473 9591 2479 9617
rect 2505 9591 2511 9617
rect 3929 9591 3935 9617
rect 3961 9591 3967 9617
rect 4993 9591 4999 9617
rect 5025 9591 5031 9617
rect 5553 9591 5559 9617
rect 5585 9591 5591 9617
rect 6449 9591 6455 9617
rect 6481 9591 6487 9617
rect 7793 9591 7799 9617
rect 7825 9591 7831 9617
rect 8353 9591 8359 9617
rect 8385 9591 8391 9617
rect 8465 9591 8471 9617
rect 8497 9591 8503 9617
rect 9473 9591 9479 9617
rect 9505 9591 9511 9617
rect 10425 9591 10431 9617
rect 10457 9591 10463 9617
rect 12049 9591 12055 9617
rect 12081 9591 12087 9617
rect 12945 9591 12951 9617
rect 12977 9591 12983 9617
rect 13505 9591 13511 9617
rect 13537 9591 13543 9617
rect 14401 9591 14407 9617
rect 14433 9591 14439 9617
rect 15521 9591 15527 9617
rect 15553 9591 15559 9617
rect 15969 9591 15975 9617
rect 16001 9591 16007 9617
rect 16193 9591 16199 9617
rect 16225 9591 16231 9617
rect 17089 9591 17095 9617
rect 17121 9591 17127 9617
rect 18265 9591 18271 9617
rect 18297 9591 18303 9617
rect 18769 9591 18775 9617
rect 18801 9591 18807 9617
rect 19217 9591 19223 9617
rect 19249 9591 19255 9617
rect 19441 9591 19447 9617
rect 19473 9591 19479 9617
rect 20225 9591 20231 9617
rect 20257 9591 20263 9617
rect 21289 9591 21295 9617
rect 21321 9591 21327 9617
rect 22745 9591 22751 9617
rect 22777 9591 22783 9617
rect 23305 9591 23311 9617
rect 23337 9591 23343 9617
rect 23417 9591 23423 9617
rect 23449 9591 23455 9617
rect 24369 9591 24375 9617
rect 24401 9591 24407 9617
rect 24649 9591 24655 9617
rect 24681 9591 24687 9617
rect 24873 9591 24879 9617
rect 24905 9591 24911 9617
rect 27225 9591 27231 9617
rect 27257 9591 27263 9617
rect 27449 9591 27455 9617
rect 27481 9591 27487 9617
rect 27897 9591 27903 9617
rect 27929 9591 27935 9617
rect 28457 9591 28463 9617
rect 28489 9591 28495 9617
rect 28737 9591 28743 9617
rect 28769 9591 28775 9617
rect 28961 9591 28967 9617
rect 28993 9591 28999 9617
rect 30977 9591 30983 9617
rect 31009 9591 31015 9617
rect 31145 9591 31151 9617
rect 31177 9591 31183 9617
rect 31369 9591 31375 9617
rect 31401 9591 31407 9617
rect 32433 9591 32439 9617
rect 32465 9591 32471 9617
rect 32825 9591 32831 9617
rect 32857 9591 32863 9617
rect 34953 9591 34959 9617
rect 34985 9591 34991 9617
rect 35849 9591 35855 9617
rect 35881 9591 35887 9617
rect 36129 9591 36135 9617
rect 36161 9591 36167 9617
rect 37305 9591 37311 9617
rect 37337 9591 37343 9617
rect 2473 9535 2479 9561
rect 2505 9535 2511 9561
rect 4993 9535 4999 9561
rect 5025 9535 5031 9561
rect 6449 9535 6455 9561
rect 6481 9535 6487 9561
rect 10425 9535 10431 9561
rect 10457 9535 10463 9561
rect 12945 9535 12951 9561
rect 12977 9535 12983 9561
rect 14401 9535 14407 9561
rect 14433 9535 14439 9561
rect 18265 9535 18271 9561
rect 18297 9535 18303 9561
rect 21289 9535 21295 9561
rect 21321 9535 21327 9561
rect 33105 9535 33111 9561
rect 33137 9535 33143 9561
rect 35849 9535 35855 9561
rect 35881 9535 35887 9561
rect 37305 9535 37311 9561
rect 37337 9535 37343 9561
rect 672 9421 39312 9438
rect 672 9395 4574 9421
rect 4600 9395 4636 9421
rect 4662 9395 4698 9421
rect 4724 9395 4760 9421
rect 4786 9395 4822 9421
rect 4848 9395 4884 9421
rect 4910 9395 4946 9421
rect 4972 9395 5008 9421
rect 5034 9395 9574 9421
rect 9600 9395 9636 9421
rect 9662 9395 9698 9421
rect 9724 9395 9760 9421
rect 9786 9395 9822 9421
rect 9848 9395 9884 9421
rect 9910 9395 9946 9421
rect 9972 9395 10008 9421
rect 10034 9395 14574 9421
rect 14600 9395 14636 9421
rect 14662 9395 14698 9421
rect 14724 9395 14760 9421
rect 14786 9395 14822 9421
rect 14848 9395 14884 9421
rect 14910 9395 14946 9421
rect 14972 9395 15008 9421
rect 15034 9395 19574 9421
rect 19600 9395 19636 9421
rect 19662 9395 19698 9421
rect 19724 9395 19760 9421
rect 19786 9395 19822 9421
rect 19848 9395 19884 9421
rect 19910 9395 19946 9421
rect 19972 9395 20008 9421
rect 20034 9395 24574 9421
rect 24600 9395 24636 9421
rect 24662 9395 24698 9421
rect 24724 9395 24760 9421
rect 24786 9395 24822 9421
rect 24848 9395 24884 9421
rect 24910 9395 24946 9421
rect 24972 9395 25008 9421
rect 25034 9395 29574 9421
rect 29600 9395 29636 9421
rect 29662 9395 29698 9421
rect 29724 9395 29760 9421
rect 29786 9395 29822 9421
rect 29848 9395 29884 9421
rect 29910 9395 29946 9421
rect 29972 9395 30008 9421
rect 30034 9395 34574 9421
rect 34600 9395 34636 9421
rect 34662 9395 34698 9421
rect 34724 9395 34760 9421
rect 34786 9395 34822 9421
rect 34848 9395 34884 9421
rect 34910 9395 34946 9421
rect 34972 9395 35008 9421
rect 35034 9395 39312 9421
rect 672 9378 39312 9395
rect 3033 9255 3039 9281
rect 3065 9255 3071 9281
rect 4265 9255 4271 9281
rect 4297 9255 4303 9281
rect 7009 9255 7015 9281
rect 7041 9255 7047 9281
rect 8353 9255 8359 9281
rect 8385 9255 8391 9281
rect 10873 9255 10879 9281
rect 10905 9255 10911 9281
rect 18265 9255 18271 9281
rect 18297 9255 18303 9281
rect 23417 9255 23423 9281
rect 23449 9255 23455 9281
rect 27393 9255 27399 9281
rect 27425 9255 27431 9281
rect 29689 9255 29695 9281
rect 29721 9255 29727 9281
rect 31369 9255 31375 9281
rect 31401 9255 31407 9281
rect 37641 9255 37647 9281
rect 37673 9255 37679 9281
rect 1913 9199 1919 9225
rect 1945 9199 1951 9225
rect 3033 9199 3039 9225
rect 3065 9199 3071 9225
rect 3593 9199 3599 9225
rect 3625 9199 3631 9225
rect 4265 9199 4271 9225
rect 4297 9199 4303 9225
rect 5833 9199 5839 9225
rect 5865 9199 5871 9225
rect 7009 9199 7015 9225
rect 7041 9199 7047 9225
rect 7569 9199 7575 9225
rect 7601 9199 7607 9225
rect 8353 9199 8359 9225
rect 8385 9199 8391 9225
rect 9809 9199 9815 9225
rect 9841 9199 9847 9225
rect 10873 9199 10879 9225
rect 10905 9199 10911 9225
rect 11545 9199 11551 9225
rect 11577 9199 11583 9225
rect 11769 9199 11775 9225
rect 11801 9199 11807 9225
rect 11937 9199 11943 9225
rect 11969 9199 11975 9225
rect 14065 9199 14071 9225
rect 14097 9199 14103 9225
rect 14345 9199 14351 9225
rect 14377 9199 14383 9225
rect 14457 9199 14463 9225
rect 14489 9199 14495 9225
rect 15241 9199 15247 9225
rect 15273 9199 15279 9225
rect 15801 9199 15807 9225
rect 15833 9199 15839 9225
rect 15913 9199 15919 9225
rect 15945 9199 15951 9225
rect 17201 9199 17207 9225
rect 17233 9199 17239 9225
rect 18265 9199 18271 9225
rect 18297 9199 18303 9225
rect 18769 9199 18775 9225
rect 18801 9199 18807 9225
rect 19217 9199 19223 9225
rect 19249 9199 19255 9225
rect 19329 9199 19335 9225
rect 19361 9199 19367 9225
rect 20785 9199 20791 9225
rect 20817 9199 20823 9225
rect 21289 9199 21295 9225
rect 21321 9199 21327 9225
rect 21457 9199 21463 9225
rect 21489 9199 21495 9225
rect 22521 9199 22527 9225
rect 22553 9199 22559 9225
rect 23417 9199 23423 9225
rect 23449 9199 23455 9225
rect 24761 9199 24767 9225
rect 24793 9199 24799 9225
rect 25209 9199 25215 9225
rect 25241 9199 25247 9225
rect 25433 9199 25439 9225
rect 25465 9199 25471 9225
rect 26497 9199 26503 9225
rect 26529 9199 26535 9225
rect 27393 9199 27399 9225
rect 27425 9199 27431 9225
rect 29017 9199 29023 9225
rect 29049 9199 29055 9225
rect 29409 9199 29415 9225
rect 29441 9199 29447 9225
rect 30417 9199 30423 9225
rect 30449 9199 30455 9225
rect 31369 9199 31375 9225
rect 31401 9199 31407 9225
rect 32937 9199 32943 9225
rect 32969 9199 32975 9225
rect 33161 9199 33167 9225
rect 33193 9199 33199 9225
rect 33385 9199 33391 9225
rect 33417 9199 33423 9225
rect 34169 9199 34175 9225
rect 34201 9199 34207 9225
rect 34617 9199 34623 9225
rect 34649 9199 34655 9225
rect 34841 9199 34847 9225
rect 34873 9199 34879 9225
rect 36689 9199 36695 9225
rect 36721 9199 36727 9225
rect 37585 9199 37591 9225
rect 37617 9199 37623 9225
rect 672 9029 39312 9046
rect 672 9003 2074 9029
rect 2100 9003 2136 9029
rect 2162 9003 2198 9029
rect 2224 9003 2260 9029
rect 2286 9003 2322 9029
rect 2348 9003 2384 9029
rect 2410 9003 2446 9029
rect 2472 9003 2508 9029
rect 2534 9003 7074 9029
rect 7100 9003 7136 9029
rect 7162 9003 7198 9029
rect 7224 9003 7260 9029
rect 7286 9003 7322 9029
rect 7348 9003 7384 9029
rect 7410 9003 7446 9029
rect 7472 9003 7508 9029
rect 7534 9003 12074 9029
rect 12100 9003 12136 9029
rect 12162 9003 12198 9029
rect 12224 9003 12260 9029
rect 12286 9003 12322 9029
rect 12348 9003 12384 9029
rect 12410 9003 12446 9029
rect 12472 9003 12508 9029
rect 12534 9003 17074 9029
rect 17100 9003 17136 9029
rect 17162 9003 17198 9029
rect 17224 9003 17260 9029
rect 17286 9003 17322 9029
rect 17348 9003 17384 9029
rect 17410 9003 17446 9029
rect 17472 9003 17508 9029
rect 17534 9003 22074 9029
rect 22100 9003 22136 9029
rect 22162 9003 22198 9029
rect 22224 9003 22260 9029
rect 22286 9003 22322 9029
rect 22348 9003 22384 9029
rect 22410 9003 22446 9029
rect 22472 9003 22508 9029
rect 22534 9003 27074 9029
rect 27100 9003 27136 9029
rect 27162 9003 27198 9029
rect 27224 9003 27260 9029
rect 27286 9003 27322 9029
rect 27348 9003 27384 9029
rect 27410 9003 27446 9029
rect 27472 9003 27508 9029
rect 27534 9003 32074 9029
rect 32100 9003 32136 9029
rect 32162 9003 32198 9029
rect 32224 9003 32260 9029
rect 32286 9003 32322 9029
rect 32348 9003 32384 9029
rect 32410 9003 32446 9029
rect 32472 9003 32508 9029
rect 32534 9003 37074 9029
rect 37100 9003 37136 9029
rect 37162 9003 37198 9029
rect 37224 9003 37260 9029
rect 37286 9003 37322 9029
rect 37348 9003 37384 9029
rect 37410 9003 37446 9029
rect 37472 9003 37508 9029
rect 37534 9003 39312 9029
rect 672 8986 39312 9003
rect 1577 8807 1583 8833
rect 1609 8807 1615 8833
rect 1745 8807 1751 8833
rect 1777 8807 1783 8833
rect 1969 8807 1975 8833
rect 2001 8807 2007 8833
rect 3929 8807 3935 8833
rect 3961 8807 3967 8833
rect 4265 8807 4271 8833
rect 4297 8807 4303 8833
rect 4489 8807 4495 8833
rect 4521 8807 4527 8833
rect 5553 8807 5559 8833
rect 5585 8807 5591 8833
rect 5945 8807 5951 8833
rect 5977 8807 5983 8833
rect 7793 8807 7799 8833
rect 7825 8807 7831 8833
rect 8353 8807 8359 8833
rect 8385 8807 8391 8833
rect 8465 8807 8471 8833
rect 8497 8807 8503 8833
rect 9249 8807 9255 8833
rect 9281 8807 9287 8833
rect 10257 8807 10263 8833
rect 10289 8807 10295 8833
rect 11993 8807 11999 8833
rect 12025 8807 12031 8833
rect 12217 8807 12223 8833
rect 12249 8807 12255 8833
rect 12441 8807 12447 8833
rect 12473 8807 12479 8833
rect 13505 8807 13511 8833
rect 13537 8807 13543 8833
rect 14401 8807 14407 8833
rect 14433 8807 14439 8833
rect 15465 8807 15471 8833
rect 15497 8807 15503 8833
rect 15913 8807 15919 8833
rect 15945 8807 15951 8833
rect 16137 8807 16143 8833
rect 16169 8807 16175 8833
rect 17201 8807 17207 8833
rect 17233 8807 17239 8833
rect 18265 8807 18271 8833
rect 18297 8807 18303 8833
rect 18769 8807 18775 8833
rect 18801 8807 18807 8833
rect 19329 8807 19335 8833
rect 19361 8807 19367 8833
rect 19497 8807 19503 8833
rect 19529 8807 19535 8833
rect 20225 8807 20231 8833
rect 20257 8807 20263 8833
rect 21289 8807 21295 8833
rect 21321 8807 21327 8833
rect 22745 8807 22751 8833
rect 22777 8807 22783 8833
rect 23305 8807 23311 8833
rect 23337 8807 23343 8833
rect 23417 8807 23423 8833
rect 23449 8807 23455 8833
rect 24369 8807 24375 8833
rect 24401 8807 24407 8833
rect 25209 8807 25215 8833
rect 25241 8807 25247 8833
rect 26721 8807 26727 8833
rect 26753 8807 26759 8833
rect 27281 8807 27287 8833
rect 27313 8807 27319 8833
rect 27505 8807 27511 8833
rect 27537 8807 27543 8833
rect 28457 8807 28463 8833
rect 28489 8807 28495 8833
rect 29353 8807 29359 8833
rect 29385 8807 29391 8833
rect 30977 8807 30983 8833
rect 31009 8807 31015 8833
rect 31873 8807 31879 8833
rect 31905 8807 31911 8833
rect 32153 8807 32159 8833
rect 32185 8807 32191 8833
rect 32713 8807 32719 8833
rect 32745 8807 32751 8833
rect 32825 8807 32831 8833
rect 32857 8807 32863 8833
rect 34953 8807 34959 8833
rect 34985 8807 34991 8833
rect 35849 8807 35855 8833
rect 35881 8807 35887 8833
rect 36353 8807 36359 8833
rect 36385 8807 36391 8833
rect 37305 8807 37311 8833
rect 37337 8807 37343 8833
rect 6225 8751 6231 8777
rect 6257 8751 6263 8777
rect 10257 8751 10263 8777
rect 10289 8751 10295 8777
rect 14401 8751 14407 8777
rect 14433 8751 14439 8777
rect 18265 8751 18271 8777
rect 18297 8751 18303 8777
rect 21289 8751 21295 8777
rect 21321 8751 21327 8777
rect 25153 8751 25159 8777
rect 25185 8751 25191 8777
rect 29353 8751 29359 8777
rect 29385 8751 29391 8777
rect 31873 8751 31879 8777
rect 31905 8751 31911 8777
rect 35849 8751 35855 8777
rect 35881 8751 35887 8777
rect 37305 8751 37311 8777
rect 37337 8751 37343 8777
rect 672 8637 39312 8654
rect 672 8611 4574 8637
rect 4600 8611 4636 8637
rect 4662 8611 4698 8637
rect 4724 8611 4760 8637
rect 4786 8611 4822 8637
rect 4848 8611 4884 8637
rect 4910 8611 4946 8637
rect 4972 8611 5008 8637
rect 5034 8611 9574 8637
rect 9600 8611 9636 8637
rect 9662 8611 9698 8637
rect 9724 8611 9760 8637
rect 9786 8611 9822 8637
rect 9848 8611 9884 8637
rect 9910 8611 9946 8637
rect 9972 8611 10008 8637
rect 10034 8611 14574 8637
rect 14600 8611 14636 8637
rect 14662 8611 14698 8637
rect 14724 8611 14760 8637
rect 14786 8611 14822 8637
rect 14848 8611 14884 8637
rect 14910 8611 14946 8637
rect 14972 8611 15008 8637
rect 15034 8611 19574 8637
rect 19600 8611 19636 8637
rect 19662 8611 19698 8637
rect 19724 8611 19760 8637
rect 19786 8611 19822 8637
rect 19848 8611 19884 8637
rect 19910 8611 19946 8637
rect 19972 8611 20008 8637
rect 20034 8611 24574 8637
rect 24600 8611 24636 8637
rect 24662 8611 24698 8637
rect 24724 8611 24760 8637
rect 24786 8611 24822 8637
rect 24848 8611 24884 8637
rect 24910 8611 24946 8637
rect 24972 8611 25008 8637
rect 25034 8611 29574 8637
rect 29600 8611 29636 8637
rect 29662 8611 29698 8637
rect 29724 8611 29760 8637
rect 29786 8611 29822 8637
rect 29848 8611 29884 8637
rect 29910 8611 29946 8637
rect 29972 8611 30008 8637
rect 30034 8611 34574 8637
rect 34600 8611 34636 8637
rect 34662 8611 34698 8637
rect 34724 8611 34760 8637
rect 34786 8611 34822 8637
rect 34848 8611 34884 8637
rect 34910 8611 34946 8637
rect 34972 8611 35008 8637
rect 35034 8611 39312 8637
rect 672 8594 39312 8611
rect 4265 8471 4271 8497
rect 4297 8471 4303 8497
rect 8353 8471 8359 8497
rect 8385 8471 8391 8497
rect 14961 8471 14967 8497
rect 14993 8471 14999 8497
rect 18265 8471 18271 8497
rect 18297 8471 18303 8497
rect 19497 8471 19503 8497
rect 19529 8471 19535 8497
rect 23417 8471 23423 8497
rect 23449 8471 23455 8497
rect 27169 8471 27175 8497
rect 27201 8471 27207 8497
rect 29913 8471 29919 8497
rect 29945 8471 29951 8497
rect 31145 8471 31151 8497
rect 31177 8471 31183 8497
rect 33889 8471 33895 8497
rect 33921 8471 33927 8497
rect 35121 8471 35127 8497
rect 35153 8471 35159 8497
rect 37641 8471 37647 8497
rect 37673 8471 37679 8497
rect 32047 8441 32073 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 2305 8415 2311 8441
rect 2337 8415 2343 8441
rect 2529 8415 2535 8441
rect 2561 8415 2567 8441
rect 3593 8415 3599 8441
rect 3625 8415 3631 8441
rect 4209 8415 4215 8441
rect 4241 8415 4247 8441
rect 5833 8415 5839 8441
rect 5865 8415 5871 8441
rect 6281 8415 6287 8441
rect 6313 8415 6319 8441
rect 6505 8415 6511 8441
rect 6537 8415 6543 8441
rect 7569 8415 7575 8441
rect 7601 8415 7607 8441
rect 8353 8415 8359 8441
rect 8385 8415 8391 8441
rect 9809 8415 9815 8441
rect 9841 8415 9847 8441
rect 10257 8415 10263 8441
rect 10289 8415 10295 8441
rect 10481 8415 10487 8441
rect 10513 8415 10519 8441
rect 11545 8415 11551 8441
rect 11577 8415 11583 8441
rect 11769 8415 11775 8441
rect 11801 8415 11807 8441
rect 11937 8415 11943 8441
rect 11969 8415 11975 8441
rect 14065 8415 14071 8441
rect 14097 8415 14103 8441
rect 14961 8415 14967 8441
rect 14993 8415 14999 8441
rect 15241 8415 15247 8441
rect 15273 8415 15279 8441
rect 15689 8415 15695 8441
rect 15721 8415 15727 8441
rect 15913 8415 15919 8441
rect 15945 8415 15951 8441
rect 17089 8415 17095 8441
rect 17121 8415 17127 8441
rect 18265 8415 18271 8441
rect 18297 8415 18303 8441
rect 18769 8415 18775 8441
rect 18801 8415 18807 8441
rect 19329 8415 19335 8441
rect 19361 8415 19367 8441
rect 20785 8415 20791 8441
rect 20817 8415 20823 8441
rect 21289 8415 21295 8441
rect 21321 8415 21327 8441
rect 21457 8415 21463 8441
rect 21489 8415 21495 8441
rect 22521 8415 22527 8441
rect 22553 8415 22559 8441
rect 23417 8415 23423 8441
rect 23449 8415 23455 8441
rect 24761 8415 24767 8441
rect 24793 8415 24799 8441
rect 25209 8415 25215 8441
rect 25241 8415 25247 8441
rect 25433 8415 25439 8441
rect 25465 8415 25471 8441
rect 26217 8415 26223 8441
rect 26249 8415 26255 8441
rect 26889 8415 26895 8441
rect 26921 8415 26927 8441
rect 29017 8415 29023 8441
rect 29049 8415 29055 8441
rect 29913 8415 29919 8441
rect 29945 8415 29951 8441
rect 30473 8415 30479 8441
rect 30505 8415 30511 8441
rect 31145 8415 31151 8441
rect 31177 8415 31183 8441
rect 32047 8409 32073 8415
rect 32215 8441 32241 8447
rect 32215 8409 32241 8415
rect 32327 8441 32353 8447
rect 32881 8415 32887 8441
rect 32913 8415 32919 8441
rect 33889 8415 33895 8441
rect 33921 8415 33927 8441
rect 34393 8415 34399 8441
rect 34425 8415 34431 8441
rect 35065 8415 35071 8441
rect 35097 8415 35103 8441
rect 36689 8415 36695 8441
rect 36721 8415 36727 8441
rect 37641 8415 37647 8441
rect 37673 8415 37679 8441
rect 32327 8409 32353 8415
rect 672 8245 39312 8262
rect 672 8219 2074 8245
rect 2100 8219 2136 8245
rect 2162 8219 2198 8245
rect 2224 8219 2260 8245
rect 2286 8219 2322 8245
rect 2348 8219 2384 8245
rect 2410 8219 2446 8245
rect 2472 8219 2508 8245
rect 2534 8219 7074 8245
rect 7100 8219 7136 8245
rect 7162 8219 7198 8245
rect 7224 8219 7260 8245
rect 7286 8219 7322 8245
rect 7348 8219 7384 8245
rect 7410 8219 7446 8245
rect 7472 8219 7508 8245
rect 7534 8219 12074 8245
rect 12100 8219 12136 8245
rect 12162 8219 12198 8245
rect 12224 8219 12260 8245
rect 12286 8219 12322 8245
rect 12348 8219 12384 8245
rect 12410 8219 12446 8245
rect 12472 8219 12508 8245
rect 12534 8219 17074 8245
rect 17100 8219 17136 8245
rect 17162 8219 17198 8245
rect 17224 8219 17260 8245
rect 17286 8219 17322 8245
rect 17348 8219 17384 8245
rect 17410 8219 17446 8245
rect 17472 8219 17508 8245
rect 17534 8219 22074 8245
rect 22100 8219 22136 8245
rect 22162 8219 22198 8245
rect 22224 8219 22260 8245
rect 22286 8219 22322 8245
rect 22348 8219 22384 8245
rect 22410 8219 22446 8245
rect 22472 8219 22508 8245
rect 22534 8219 27074 8245
rect 27100 8219 27136 8245
rect 27162 8219 27198 8245
rect 27224 8219 27260 8245
rect 27286 8219 27322 8245
rect 27348 8219 27384 8245
rect 27410 8219 27446 8245
rect 27472 8219 27508 8245
rect 27534 8219 32074 8245
rect 32100 8219 32136 8245
rect 32162 8219 32198 8245
rect 32224 8219 32260 8245
rect 32286 8219 32322 8245
rect 32348 8219 32384 8245
rect 32410 8219 32446 8245
rect 32472 8219 32508 8245
rect 32534 8219 37074 8245
rect 37100 8219 37136 8245
rect 37162 8219 37198 8245
rect 37224 8219 37260 8245
rect 37286 8219 37322 8245
rect 37348 8219 37384 8245
rect 37410 8219 37446 8245
rect 37472 8219 37508 8245
rect 37534 8219 39312 8245
rect 672 8202 39312 8219
rect 33727 8049 33753 8055
rect 1577 8023 1583 8049
rect 1609 8023 1615 8049
rect 1969 8023 1975 8049
rect 2001 8023 2007 8049
rect 3929 8023 3935 8049
rect 3961 8023 3967 8049
rect 4265 8023 4271 8049
rect 4297 8023 4303 8049
rect 4489 8023 4495 8049
rect 4521 8023 4527 8049
rect 5553 8023 5559 8049
rect 5585 8023 5591 8049
rect 6225 8023 6231 8049
rect 6257 8023 6263 8049
rect 7793 8023 7799 8049
rect 7825 8023 7831 8049
rect 8353 8023 8359 8049
rect 8385 8023 8391 8049
rect 8465 8023 8471 8049
rect 8497 8023 8503 8049
rect 9249 8023 9255 8049
rect 9281 8023 9287 8049
rect 10257 8023 10263 8049
rect 10289 8023 10295 8049
rect 12049 8023 12055 8049
rect 12081 8023 12087 8049
rect 12217 8023 12223 8049
rect 12249 8023 12255 8049
rect 12441 8023 12447 8049
rect 12473 8023 12479 8049
rect 13393 8023 13399 8049
rect 13425 8023 13431 8049
rect 14177 8023 14183 8049
rect 14209 8023 14215 8049
rect 15297 8023 15303 8049
rect 15329 8023 15335 8049
rect 16417 8023 16423 8049
rect 16449 8023 16455 8049
rect 16865 8023 16871 8049
rect 16897 8023 16903 8049
rect 17705 8023 17711 8049
rect 17737 8023 17743 8049
rect 18769 8023 18775 8049
rect 18801 8023 18807 8049
rect 19329 8023 19335 8049
rect 19361 8023 19367 8049
rect 19441 8023 19447 8049
rect 19473 8023 19479 8049
rect 20225 8023 20231 8049
rect 20257 8023 20263 8049
rect 21289 8023 21295 8049
rect 21321 8023 21327 8049
rect 22745 8023 22751 8049
rect 22777 8023 22783 8049
rect 23305 8023 23311 8049
rect 23337 8023 23343 8049
rect 23417 8023 23423 8049
rect 23449 8023 23455 8049
rect 24369 8023 24375 8049
rect 24401 8023 24407 8049
rect 24761 8023 24767 8049
rect 24793 8023 24799 8049
rect 24873 8023 24879 8049
rect 24905 8023 24911 8049
rect 26721 8023 26727 8049
rect 26753 8023 26759 8049
rect 27169 8023 27175 8049
rect 27201 8023 27207 8049
rect 27393 8023 27399 8049
rect 27425 8023 27431 8049
rect 28457 8023 28463 8049
rect 28489 8023 28495 8049
rect 29353 8023 29359 8049
rect 29385 8023 29391 8049
rect 30977 8023 30983 8049
rect 31009 8023 31015 8049
rect 31145 8023 31151 8049
rect 31177 8023 31183 8049
rect 31369 8023 31375 8049
rect 31401 8023 31407 8049
rect 32433 8023 32439 8049
rect 32465 8023 32471 8049
rect 33329 8023 33335 8049
rect 33361 8023 33367 8049
rect 34953 8023 34959 8049
rect 34985 8023 34991 8049
rect 35849 8023 35855 8049
rect 35881 8023 35887 8049
rect 36409 8023 36415 8049
rect 36441 8023 36447 8049
rect 37305 8023 37311 8049
rect 37337 8023 37343 8049
rect 33727 8017 33753 8023
rect 33615 7993 33641 7999
rect 2249 7967 2255 7993
rect 2281 7967 2287 7993
rect 6225 7967 6231 7993
rect 6257 7967 6263 7993
rect 10257 7967 10263 7993
rect 10289 7967 10295 7993
rect 14177 7967 14183 7993
rect 14209 7967 14215 7993
rect 16417 7967 16423 7993
rect 16449 7967 16455 7993
rect 17705 7967 17711 7993
rect 17737 7967 17743 7993
rect 21289 7967 21295 7993
rect 21321 7967 21327 7993
rect 29353 7967 29359 7993
rect 29385 7967 29391 7993
rect 33329 7967 33335 7993
rect 33361 7967 33367 7993
rect 33615 7961 33641 7967
rect 33895 7993 33921 7999
rect 35849 7967 35855 7993
rect 35881 7967 35887 7993
rect 37305 7967 37311 7993
rect 37337 7967 37343 7993
rect 33895 7961 33921 7967
rect 672 7853 39312 7870
rect 672 7827 4574 7853
rect 4600 7827 4636 7853
rect 4662 7827 4698 7853
rect 4724 7827 4760 7853
rect 4786 7827 4822 7853
rect 4848 7827 4884 7853
rect 4910 7827 4946 7853
rect 4972 7827 5008 7853
rect 5034 7827 9574 7853
rect 9600 7827 9636 7853
rect 9662 7827 9698 7853
rect 9724 7827 9760 7853
rect 9786 7827 9822 7853
rect 9848 7827 9884 7853
rect 9910 7827 9946 7853
rect 9972 7827 10008 7853
rect 10034 7827 14574 7853
rect 14600 7827 14636 7853
rect 14662 7827 14698 7853
rect 14724 7827 14760 7853
rect 14786 7827 14822 7853
rect 14848 7827 14884 7853
rect 14910 7827 14946 7853
rect 14972 7827 15008 7853
rect 15034 7827 19574 7853
rect 19600 7827 19636 7853
rect 19662 7827 19698 7853
rect 19724 7827 19760 7853
rect 19786 7827 19822 7853
rect 19848 7827 19884 7853
rect 19910 7827 19946 7853
rect 19972 7827 20008 7853
rect 20034 7827 24574 7853
rect 24600 7827 24636 7853
rect 24662 7827 24698 7853
rect 24724 7827 24760 7853
rect 24786 7827 24822 7853
rect 24848 7827 24884 7853
rect 24910 7827 24946 7853
rect 24972 7827 25008 7853
rect 25034 7827 29574 7853
rect 29600 7827 29636 7853
rect 29662 7827 29698 7853
rect 29724 7827 29760 7853
rect 29786 7827 29822 7853
rect 29848 7827 29884 7853
rect 29910 7827 29946 7853
rect 29972 7827 30008 7853
rect 30034 7827 34574 7853
rect 34600 7827 34636 7853
rect 34662 7827 34698 7853
rect 34724 7827 34760 7853
rect 34786 7827 34822 7853
rect 34848 7827 34884 7853
rect 34910 7827 34946 7853
rect 34972 7827 35008 7853
rect 35034 7827 39312 7853
rect 672 7810 39312 7827
rect 3033 7687 3039 7713
rect 3065 7687 3071 7713
rect 4265 7687 4271 7713
rect 4297 7687 4303 7713
rect 14961 7687 14967 7713
rect 14993 7687 14999 7713
rect 16417 7687 16423 7713
rect 16449 7687 16455 7713
rect 17761 7687 17767 7713
rect 17793 7687 17799 7713
rect 19329 7687 19335 7713
rect 19361 7687 19367 7713
rect 23417 7687 23423 7713
rect 23449 7687 23455 7713
rect 31369 7687 31375 7713
rect 31401 7687 31407 7713
rect 33833 7687 33839 7713
rect 33865 7687 33871 7713
rect 35233 7687 35239 7713
rect 35265 7687 35271 7713
rect 37641 7687 37647 7713
rect 37673 7687 37679 7713
rect 32103 7657 32129 7663
rect 1857 7631 1863 7657
rect 1889 7631 1895 7657
rect 3033 7631 3039 7657
rect 3065 7631 3071 7657
rect 3593 7631 3599 7657
rect 3625 7631 3631 7657
rect 4209 7631 4215 7657
rect 4241 7631 4247 7657
rect 5833 7631 5839 7657
rect 5865 7631 5871 7657
rect 6281 7631 6287 7657
rect 6313 7631 6319 7657
rect 6505 7631 6511 7657
rect 6537 7631 6543 7657
rect 7569 7631 7575 7657
rect 7601 7631 7607 7657
rect 7737 7631 7743 7657
rect 7769 7631 7775 7657
rect 7961 7631 7967 7657
rect 7993 7631 7999 7657
rect 9809 7631 9815 7657
rect 9841 7631 9847 7657
rect 10257 7631 10263 7657
rect 10289 7631 10295 7657
rect 10481 7631 10487 7657
rect 10513 7631 10519 7657
rect 11265 7631 11271 7657
rect 11297 7631 11303 7657
rect 11769 7631 11775 7657
rect 11801 7631 11807 7657
rect 11937 7631 11943 7657
rect 11969 7631 11975 7657
rect 14065 7631 14071 7657
rect 14097 7631 14103 7657
rect 14961 7631 14967 7657
rect 14993 7631 14999 7657
rect 15241 7631 15247 7657
rect 15273 7631 15279 7657
rect 16417 7631 16423 7657
rect 16449 7631 16455 7657
rect 16865 7631 16871 7657
rect 16897 7631 16903 7657
rect 17705 7631 17711 7657
rect 17737 7631 17743 7657
rect 18545 7631 18551 7657
rect 18577 7631 18583 7657
rect 19329 7631 19335 7657
rect 19361 7631 19367 7657
rect 20785 7631 20791 7657
rect 20817 7631 20823 7657
rect 21289 7631 21295 7657
rect 21321 7631 21327 7657
rect 21457 7631 21463 7657
rect 21489 7631 21495 7657
rect 22521 7631 22527 7657
rect 22553 7631 22559 7657
rect 23417 7631 23423 7657
rect 23449 7631 23455 7657
rect 24761 7631 24767 7657
rect 24793 7631 24799 7657
rect 25209 7631 25215 7657
rect 25241 7631 25247 7657
rect 25433 7631 25439 7657
rect 25465 7631 25471 7657
rect 26217 7631 26223 7657
rect 26249 7631 26255 7657
rect 26777 7631 26783 7657
rect 26809 7631 26815 7657
rect 26889 7631 26895 7657
rect 26921 7631 26927 7657
rect 29017 7631 29023 7657
rect 29049 7631 29055 7657
rect 29297 7631 29303 7657
rect 29329 7631 29335 7657
rect 29465 7631 29471 7657
rect 29497 7631 29503 7657
rect 30473 7631 30479 7657
rect 30505 7631 30511 7657
rect 31369 7631 31375 7657
rect 31401 7631 31407 7657
rect 32103 7625 32129 7631
rect 32159 7657 32185 7663
rect 32159 7625 32185 7631
rect 32327 7657 32353 7663
rect 32937 7631 32943 7657
rect 32969 7631 32975 7657
rect 33833 7631 33839 7657
rect 33865 7631 33871 7657
rect 34393 7631 34399 7657
rect 34425 7631 34431 7657
rect 35233 7631 35239 7657
rect 35265 7631 35271 7657
rect 36689 7631 36695 7657
rect 36721 7631 36727 7657
rect 37641 7631 37647 7657
rect 37673 7631 37679 7657
rect 32327 7625 32353 7631
rect 672 7461 39312 7478
rect 672 7435 2074 7461
rect 2100 7435 2136 7461
rect 2162 7435 2198 7461
rect 2224 7435 2260 7461
rect 2286 7435 2322 7461
rect 2348 7435 2384 7461
rect 2410 7435 2446 7461
rect 2472 7435 2508 7461
rect 2534 7435 7074 7461
rect 7100 7435 7136 7461
rect 7162 7435 7198 7461
rect 7224 7435 7260 7461
rect 7286 7435 7322 7461
rect 7348 7435 7384 7461
rect 7410 7435 7446 7461
rect 7472 7435 7508 7461
rect 7534 7435 12074 7461
rect 12100 7435 12136 7461
rect 12162 7435 12198 7461
rect 12224 7435 12260 7461
rect 12286 7435 12322 7461
rect 12348 7435 12384 7461
rect 12410 7435 12446 7461
rect 12472 7435 12508 7461
rect 12534 7435 17074 7461
rect 17100 7435 17136 7461
rect 17162 7435 17198 7461
rect 17224 7435 17260 7461
rect 17286 7435 17322 7461
rect 17348 7435 17384 7461
rect 17410 7435 17446 7461
rect 17472 7435 17508 7461
rect 17534 7435 22074 7461
rect 22100 7435 22136 7461
rect 22162 7435 22198 7461
rect 22224 7435 22260 7461
rect 22286 7435 22322 7461
rect 22348 7435 22384 7461
rect 22410 7435 22446 7461
rect 22472 7435 22508 7461
rect 22534 7435 27074 7461
rect 27100 7435 27136 7461
rect 27162 7435 27198 7461
rect 27224 7435 27260 7461
rect 27286 7435 27322 7461
rect 27348 7435 27384 7461
rect 27410 7435 27446 7461
rect 27472 7435 27508 7461
rect 27534 7435 32074 7461
rect 32100 7435 32136 7461
rect 32162 7435 32198 7461
rect 32224 7435 32260 7461
rect 32286 7435 32322 7461
rect 32348 7435 32384 7461
rect 32410 7435 32446 7461
rect 32472 7435 32508 7461
rect 32534 7435 37074 7461
rect 37100 7435 37136 7461
rect 37162 7435 37198 7461
rect 37224 7435 37260 7461
rect 37286 7435 37322 7461
rect 37348 7435 37384 7461
rect 37410 7435 37446 7461
rect 37472 7435 37508 7461
rect 37534 7435 39312 7461
rect 672 7418 39312 7435
rect 33671 7265 33697 7271
rect 1801 7239 1807 7265
rect 1833 7239 1839 7265
rect 2025 7239 2031 7265
rect 2057 7239 2063 7265
rect 2473 7239 2479 7265
rect 2505 7239 2511 7265
rect 4097 7239 4103 7265
rect 4129 7239 4135 7265
rect 4993 7239 4999 7265
rect 5025 7239 5031 7265
rect 5273 7239 5279 7265
rect 5305 7239 5311 7265
rect 6449 7239 6455 7265
rect 6481 7239 6487 7265
rect 8073 7239 8079 7265
rect 8105 7239 8111 7265
rect 8745 7239 8751 7265
rect 8777 7239 8783 7265
rect 9417 7239 9423 7265
rect 9449 7239 9455 7265
rect 10201 7239 10207 7265
rect 10233 7239 10239 7265
rect 11825 7239 11831 7265
rect 11857 7239 11863 7265
rect 12217 7239 12223 7265
rect 12249 7239 12255 7265
rect 12441 7239 12447 7265
rect 12473 7239 12479 7265
rect 13505 7239 13511 7265
rect 13537 7239 13543 7265
rect 14401 7239 14407 7265
rect 14433 7239 14439 7265
rect 15185 7239 15191 7265
rect 15217 7239 15223 7265
rect 15689 7239 15695 7265
rect 15721 7239 15727 7265
rect 15801 7239 15807 7265
rect 15833 7239 15839 7265
rect 16809 7239 16815 7265
rect 16841 7239 16847 7265
rect 17257 7239 17263 7265
rect 17289 7239 17295 7265
rect 17369 7239 17375 7265
rect 17401 7239 17407 7265
rect 18769 7239 18775 7265
rect 18801 7239 18807 7265
rect 19329 7239 19335 7265
rect 19361 7239 19367 7265
rect 19441 7239 19447 7265
rect 19473 7239 19479 7265
rect 20225 7239 20231 7265
rect 20257 7239 20263 7265
rect 21289 7239 21295 7265
rect 21321 7239 21327 7265
rect 22745 7239 22751 7265
rect 22777 7239 22783 7265
rect 23305 7239 23311 7265
rect 23337 7239 23343 7265
rect 23417 7239 23423 7265
rect 23449 7239 23455 7265
rect 24369 7239 24375 7265
rect 24401 7239 24407 7265
rect 25097 7239 25103 7265
rect 25129 7239 25135 7265
rect 26721 7239 26727 7265
rect 26753 7239 26759 7265
rect 27169 7239 27175 7265
rect 27201 7239 27207 7265
rect 27393 7239 27399 7265
rect 27425 7239 27431 7265
rect 28457 7239 28463 7265
rect 28489 7239 28495 7265
rect 29185 7239 29191 7265
rect 29217 7239 29223 7265
rect 30977 7239 30983 7265
rect 31009 7239 31015 7265
rect 31817 7239 31823 7265
rect 31849 7239 31855 7265
rect 32433 7239 32439 7265
rect 32465 7239 32471 7265
rect 33329 7239 33335 7265
rect 33361 7239 33367 7265
rect 33671 7233 33697 7239
rect 33727 7265 33753 7271
rect 34673 7239 34679 7265
rect 34705 7239 34711 7265
rect 35121 7239 35127 7265
rect 35153 7239 35159 7265
rect 35345 7239 35351 7265
rect 35377 7239 35383 7265
rect 36409 7239 36415 7265
rect 36441 7239 36447 7265
rect 37305 7239 37311 7265
rect 37337 7239 37343 7265
rect 33727 7233 33753 7239
rect 33895 7209 33921 7215
rect 4993 7183 4999 7209
rect 5025 7183 5031 7209
rect 6449 7183 6455 7209
rect 6481 7183 6487 7209
rect 8745 7183 8751 7209
rect 8777 7183 8783 7209
rect 10201 7183 10207 7209
rect 10233 7183 10239 7209
rect 14401 7183 14407 7209
rect 14433 7183 14439 7209
rect 21289 7183 21295 7209
rect 21321 7183 21327 7209
rect 25153 7183 25159 7209
rect 25185 7183 25191 7209
rect 29185 7183 29191 7209
rect 29217 7183 29223 7209
rect 31817 7183 31823 7209
rect 31849 7183 31855 7209
rect 33329 7183 33335 7209
rect 33361 7183 33367 7209
rect 37305 7183 37311 7209
rect 37337 7183 37343 7209
rect 33895 7177 33921 7183
rect 672 7069 39312 7086
rect 672 7043 4574 7069
rect 4600 7043 4636 7069
rect 4662 7043 4698 7069
rect 4724 7043 4760 7069
rect 4786 7043 4822 7069
rect 4848 7043 4884 7069
rect 4910 7043 4946 7069
rect 4972 7043 5008 7069
rect 5034 7043 9574 7069
rect 9600 7043 9636 7069
rect 9662 7043 9698 7069
rect 9724 7043 9760 7069
rect 9786 7043 9822 7069
rect 9848 7043 9884 7069
rect 9910 7043 9946 7069
rect 9972 7043 10008 7069
rect 10034 7043 14574 7069
rect 14600 7043 14636 7069
rect 14662 7043 14698 7069
rect 14724 7043 14760 7069
rect 14786 7043 14822 7069
rect 14848 7043 14884 7069
rect 14910 7043 14946 7069
rect 14972 7043 15008 7069
rect 15034 7043 19574 7069
rect 19600 7043 19636 7069
rect 19662 7043 19698 7069
rect 19724 7043 19760 7069
rect 19786 7043 19822 7069
rect 19848 7043 19884 7069
rect 19910 7043 19946 7069
rect 19972 7043 20008 7069
rect 20034 7043 24574 7069
rect 24600 7043 24636 7069
rect 24662 7043 24698 7069
rect 24724 7043 24760 7069
rect 24786 7043 24822 7069
rect 24848 7043 24884 7069
rect 24910 7043 24946 7069
rect 24972 7043 25008 7069
rect 25034 7043 29574 7069
rect 29600 7043 29636 7069
rect 29662 7043 29698 7069
rect 29724 7043 29760 7069
rect 29786 7043 29822 7069
rect 29848 7043 29884 7069
rect 29910 7043 29946 7069
rect 29972 7043 30008 7069
rect 30034 7043 34574 7069
rect 34600 7043 34636 7069
rect 34662 7043 34698 7069
rect 34724 7043 34760 7069
rect 34786 7043 34822 7069
rect 34848 7043 34884 7069
rect 34910 7043 34946 7069
rect 34972 7043 35008 7069
rect 35034 7043 39312 7069
rect 672 7026 39312 7043
rect 35631 6929 35657 6935
rect 4489 6903 4495 6929
rect 4521 6903 4527 6929
rect 7009 6903 7015 6929
rect 7041 6903 7047 6929
rect 8353 6903 8359 6929
rect 8385 6903 8391 6929
rect 16193 6903 16199 6929
rect 16225 6903 16231 6929
rect 19329 6903 19335 6929
rect 19361 6903 19367 6929
rect 23417 6903 23423 6929
rect 23449 6903 23455 6929
rect 33665 6903 33671 6929
rect 33697 6903 33703 6929
rect 35121 6903 35127 6929
rect 35153 6903 35159 6929
rect 35631 6897 35657 6903
rect 35743 6929 35769 6935
rect 35743 6897 35769 6903
rect 35911 6929 35937 6935
rect 37641 6903 37647 6929
rect 37673 6903 37679 6929
rect 35911 6897 35937 6903
rect 32047 6873 32073 6879
rect 2361 6847 2367 6873
rect 2393 6847 2399 6873
rect 2473 6847 2479 6873
rect 2505 6847 2511 6873
rect 3033 6847 3039 6873
rect 3065 6847 3071 6873
rect 3593 6847 3599 6873
rect 3625 6847 3631 6873
rect 4489 6847 4495 6873
rect 4521 6847 4527 6873
rect 6113 6847 6119 6873
rect 6145 6847 6151 6873
rect 7009 6847 7015 6873
rect 7041 6847 7047 6873
rect 7569 6847 7575 6873
rect 7601 6847 7607 6873
rect 8353 6847 8359 6873
rect 8385 6847 8391 6873
rect 10033 6847 10039 6873
rect 10065 6847 10071 6873
rect 10257 6847 10263 6873
rect 10289 6847 10295 6873
rect 10537 6847 10543 6873
rect 10569 6847 10575 6873
rect 11545 6847 11551 6873
rect 11577 6847 11583 6873
rect 11769 6847 11775 6873
rect 11801 6847 11807 6873
rect 11993 6847 11999 6873
rect 12025 6847 12031 6873
rect 13729 6847 13735 6873
rect 13761 6847 13767 6873
rect 14289 6847 14295 6873
rect 14321 6847 14327 6873
rect 14401 6847 14407 6873
rect 14433 6847 14439 6873
rect 15241 6847 15247 6873
rect 15273 6847 15279 6873
rect 16193 6847 16199 6873
rect 16225 6847 16231 6873
rect 16809 6847 16815 6873
rect 16841 6847 16847 6873
rect 17369 6847 17375 6873
rect 17401 6847 17407 6873
rect 17593 6847 17599 6873
rect 17625 6847 17631 6873
rect 18545 6847 18551 6873
rect 18577 6847 18583 6873
rect 19329 6847 19335 6873
rect 19361 6847 19367 6873
rect 20785 6847 20791 6873
rect 20817 6847 20823 6873
rect 21289 6847 21295 6873
rect 21321 6847 21327 6873
rect 21457 6847 21463 6873
rect 21489 6847 21495 6873
rect 22521 6847 22527 6873
rect 22553 6847 22559 6873
rect 23417 6847 23423 6873
rect 23449 6847 23455 6873
rect 24761 6847 24767 6873
rect 24793 6847 24799 6873
rect 25209 6847 25215 6873
rect 25241 6847 25247 6873
rect 25433 6847 25439 6873
rect 25465 6847 25471 6873
rect 26217 6847 26223 6873
rect 26249 6847 26255 6873
rect 26777 6847 26783 6873
rect 26809 6847 26815 6873
rect 26889 6847 26895 6873
rect 26921 6847 26927 6873
rect 28737 6847 28743 6873
rect 28769 6847 28775 6873
rect 29185 6847 29191 6873
rect 29217 6847 29223 6873
rect 29409 6847 29415 6873
rect 29441 6847 29447 6873
rect 30473 6847 30479 6873
rect 30505 6847 30511 6873
rect 30641 6847 30647 6873
rect 30673 6847 30679 6873
rect 31369 6847 31375 6873
rect 31401 6847 31407 6873
rect 32047 6841 32073 6847
rect 32159 6873 32185 6879
rect 32159 6841 32185 6847
rect 32327 6873 32353 6879
rect 32993 6847 32999 6873
rect 33025 6847 33031 6873
rect 33665 6847 33671 6873
rect 33697 6847 33703 6873
rect 34393 6847 34399 6873
rect 34425 6847 34431 6873
rect 35121 6847 35127 6873
rect 35153 6847 35159 6873
rect 36689 6847 36695 6873
rect 36721 6847 36727 6873
rect 37641 6847 37647 6873
rect 37673 6847 37679 6873
rect 32327 6841 32353 6847
rect 672 6677 39312 6694
rect 672 6651 2074 6677
rect 2100 6651 2136 6677
rect 2162 6651 2198 6677
rect 2224 6651 2260 6677
rect 2286 6651 2322 6677
rect 2348 6651 2384 6677
rect 2410 6651 2446 6677
rect 2472 6651 2508 6677
rect 2534 6651 7074 6677
rect 7100 6651 7136 6677
rect 7162 6651 7198 6677
rect 7224 6651 7260 6677
rect 7286 6651 7322 6677
rect 7348 6651 7384 6677
rect 7410 6651 7446 6677
rect 7472 6651 7508 6677
rect 7534 6651 12074 6677
rect 12100 6651 12136 6677
rect 12162 6651 12198 6677
rect 12224 6651 12260 6677
rect 12286 6651 12322 6677
rect 12348 6651 12384 6677
rect 12410 6651 12446 6677
rect 12472 6651 12508 6677
rect 12534 6651 17074 6677
rect 17100 6651 17136 6677
rect 17162 6651 17198 6677
rect 17224 6651 17260 6677
rect 17286 6651 17322 6677
rect 17348 6651 17384 6677
rect 17410 6651 17446 6677
rect 17472 6651 17508 6677
rect 17534 6651 22074 6677
rect 22100 6651 22136 6677
rect 22162 6651 22198 6677
rect 22224 6651 22260 6677
rect 22286 6651 22322 6677
rect 22348 6651 22384 6677
rect 22410 6651 22446 6677
rect 22472 6651 22508 6677
rect 22534 6651 27074 6677
rect 27100 6651 27136 6677
rect 27162 6651 27198 6677
rect 27224 6651 27260 6677
rect 27286 6651 27322 6677
rect 27348 6651 27384 6677
rect 27410 6651 27446 6677
rect 27472 6651 27508 6677
rect 27534 6651 32074 6677
rect 32100 6651 32136 6677
rect 32162 6651 32198 6677
rect 32224 6651 32260 6677
rect 32286 6651 32322 6677
rect 32348 6651 32384 6677
rect 32410 6651 32446 6677
rect 32472 6651 32508 6677
rect 32534 6651 37074 6677
rect 37100 6651 37136 6677
rect 37162 6651 37198 6677
rect 37224 6651 37260 6677
rect 37286 6651 37322 6677
rect 37348 6651 37384 6677
rect 37410 6651 37446 6677
rect 37472 6651 37508 6677
rect 37534 6651 39312 6677
rect 672 6634 39312 6651
rect 30199 6481 30225 6487
rect 1801 6455 1807 6481
rect 1833 6455 1839 6481
rect 1969 6455 1975 6481
rect 2001 6455 2007 6481
rect 2473 6455 2479 6481
rect 2505 6455 2511 6481
rect 4097 6455 4103 6481
rect 4129 6455 4135 6481
rect 4377 6455 4383 6481
rect 4409 6455 4415 6481
rect 4489 6455 4495 6481
rect 4521 6455 4527 6481
rect 5273 6455 5279 6481
rect 5305 6455 5311 6481
rect 6449 6455 6455 6481
rect 6481 6455 6487 6481
rect 8073 6455 8079 6481
rect 8105 6455 8111 6481
rect 8969 6455 8975 6481
rect 9001 6455 9007 6481
rect 9417 6455 9423 6481
rect 9449 6455 9455 6481
rect 10313 6455 10319 6481
rect 10345 6455 10351 6481
rect 11825 6455 11831 6481
rect 11857 6455 11863 6481
rect 12329 6455 12335 6481
rect 12361 6455 12367 6481
rect 12441 6455 12447 6481
rect 12473 6455 12479 6481
rect 13505 6455 13511 6481
rect 13537 6455 13543 6481
rect 14233 6455 14239 6481
rect 14265 6455 14271 6481
rect 16361 6455 16367 6481
rect 16393 6455 16399 6481
rect 17313 6455 17319 6481
rect 17345 6455 17351 6481
rect 18769 6455 18775 6481
rect 18801 6455 18807 6481
rect 19329 6455 19335 6481
rect 19361 6455 19367 6481
rect 19441 6455 19447 6481
rect 19473 6455 19479 6481
rect 20225 6455 20231 6481
rect 20257 6455 20263 6481
rect 21289 6455 21295 6481
rect 21321 6455 21327 6481
rect 22745 6455 22751 6481
rect 22777 6455 22783 6481
rect 23193 6455 23199 6481
rect 23225 6455 23231 6481
rect 23417 6455 23423 6481
rect 23449 6455 23455 6481
rect 24369 6455 24375 6481
rect 24401 6455 24407 6481
rect 25209 6455 25215 6481
rect 25241 6455 25247 6481
rect 26721 6455 26727 6481
rect 26753 6455 26759 6481
rect 27169 6455 27175 6481
rect 27201 6455 27207 6481
rect 27393 6455 27399 6481
rect 27425 6455 27431 6481
rect 28457 6455 28463 6481
rect 28489 6455 28495 6481
rect 28681 6455 28687 6481
rect 28713 6455 28719 6481
rect 28849 6455 28855 6481
rect 28881 6455 28887 6481
rect 30199 6449 30225 6455
rect 30311 6481 30337 6487
rect 30921 6455 30927 6481
rect 30953 6455 30959 6481
rect 31873 6455 31879 6481
rect 31905 6455 31911 6481
rect 32153 6455 32159 6481
rect 32185 6455 32191 6481
rect 33273 6455 33279 6481
rect 33305 6455 33311 6481
rect 34673 6455 34679 6481
rect 34705 6455 34711 6481
rect 35233 6455 35239 6481
rect 35265 6455 35271 6481
rect 35345 6455 35351 6481
rect 35377 6455 35383 6481
rect 36129 6455 36135 6481
rect 36161 6455 36167 6481
rect 37305 6455 37311 6481
rect 37337 6455 37343 6481
rect 30311 6449 30337 6455
rect 30031 6425 30057 6431
rect 33615 6425 33641 6431
rect 6449 6399 6455 6425
rect 6481 6399 6487 6425
rect 8969 6399 8975 6425
rect 9001 6399 9007 6425
rect 10313 6399 10319 6425
rect 10345 6399 10351 6425
rect 14233 6399 14239 6425
rect 14265 6399 14271 6425
rect 17313 6399 17319 6425
rect 17345 6399 17351 6425
rect 21289 6399 21295 6425
rect 21321 6399 21327 6425
rect 25209 6399 25215 6425
rect 25241 6399 25247 6425
rect 31873 6399 31879 6425
rect 31905 6399 31911 6425
rect 33273 6399 33279 6425
rect 33305 6399 33311 6425
rect 30031 6393 30057 6399
rect 33615 6393 33641 6399
rect 33727 6425 33753 6431
rect 33727 6393 33753 6399
rect 33895 6425 33921 6431
rect 37305 6399 37311 6425
rect 37337 6399 37343 6425
rect 33895 6393 33921 6399
rect 672 6285 39312 6302
rect 672 6259 4574 6285
rect 4600 6259 4636 6285
rect 4662 6259 4698 6285
rect 4724 6259 4760 6285
rect 4786 6259 4822 6285
rect 4848 6259 4884 6285
rect 4910 6259 4946 6285
rect 4972 6259 5008 6285
rect 5034 6259 9574 6285
rect 9600 6259 9636 6285
rect 9662 6259 9698 6285
rect 9724 6259 9760 6285
rect 9786 6259 9822 6285
rect 9848 6259 9884 6285
rect 9910 6259 9946 6285
rect 9972 6259 10008 6285
rect 10034 6259 14574 6285
rect 14600 6259 14636 6285
rect 14662 6259 14698 6285
rect 14724 6259 14760 6285
rect 14786 6259 14822 6285
rect 14848 6259 14884 6285
rect 14910 6259 14946 6285
rect 14972 6259 15008 6285
rect 15034 6259 19574 6285
rect 19600 6259 19636 6285
rect 19662 6259 19698 6285
rect 19724 6259 19760 6285
rect 19786 6259 19822 6285
rect 19848 6259 19884 6285
rect 19910 6259 19946 6285
rect 19972 6259 20008 6285
rect 20034 6259 24574 6285
rect 24600 6259 24636 6285
rect 24662 6259 24698 6285
rect 24724 6259 24760 6285
rect 24786 6259 24822 6285
rect 24848 6259 24884 6285
rect 24910 6259 24946 6285
rect 24972 6259 25008 6285
rect 25034 6259 29574 6285
rect 29600 6259 29636 6285
rect 29662 6259 29698 6285
rect 29724 6259 29760 6285
rect 29786 6259 29822 6285
rect 29848 6259 29884 6285
rect 29910 6259 29946 6285
rect 29972 6259 30008 6285
rect 30034 6259 34574 6285
rect 34600 6259 34636 6285
rect 34662 6259 34698 6285
rect 34724 6259 34760 6285
rect 34786 6259 34822 6285
rect 34848 6259 34884 6285
rect 34910 6259 34946 6285
rect 34972 6259 35008 6285
rect 35034 6259 39312 6285
rect 672 6242 39312 6259
rect 1969 6119 1975 6145
rect 2001 6119 2007 6145
rect 4489 6119 4495 6145
rect 4521 6119 4527 6145
rect 7009 6119 7015 6145
rect 7041 6119 7047 6145
rect 8465 6119 8471 6145
rect 8497 6119 8503 6145
rect 12441 6119 12447 6145
rect 12473 6119 12479 6145
rect 14849 6119 14855 6145
rect 14881 6119 14887 6145
rect 17761 6119 17767 6145
rect 17793 6119 17799 6145
rect 19441 6119 19447 6145
rect 19473 6119 19479 6145
rect 27169 6119 27175 6145
rect 27201 6119 27207 6145
rect 29913 6119 29919 6145
rect 29945 6119 29951 6145
rect 31369 6119 31375 6145
rect 31401 6119 31407 6145
rect 33777 6119 33783 6145
rect 33809 6119 33815 6145
rect 35121 6119 35127 6145
rect 35153 6119 35159 6145
rect 37641 6119 37647 6145
rect 37673 6119 37679 6145
rect 32047 6089 32073 6095
rect 1969 6063 1975 6089
rect 2001 6063 2007 6089
rect 3033 6063 3039 6089
rect 3065 6063 3071 6089
rect 3593 6063 3599 6089
rect 3625 6063 3631 6089
rect 4489 6063 4495 6089
rect 4521 6063 4527 6089
rect 6113 6063 6119 6089
rect 6145 6063 6151 6089
rect 7009 6063 7015 6089
rect 7041 6063 7047 6089
rect 7569 6063 7575 6089
rect 7601 6063 7607 6089
rect 8465 6063 8471 6089
rect 8497 6063 8503 6089
rect 10033 6063 10039 6089
rect 10065 6063 10071 6089
rect 10313 6063 10319 6089
rect 10345 6063 10351 6089
rect 10481 6063 10487 6089
rect 10513 6063 10519 6089
rect 11545 6063 11551 6089
rect 11577 6063 11583 6089
rect 12441 6063 12447 6089
rect 12473 6063 12479 6089
rect 13953 6063 13959 6089
rect 13985 6063 13991 6089
rect 14849 6063 14855 6089
rect 14881 6063 14887 6089
rect 15185 6063 15191 6089
rect 15217 6063 15223 6089
rect 15689 6063 15695 6089
rect 15721 6063 15727 6089
rect 15857 6063 15863 6089
rect 15889 6063 15895 6089
rect 16809 6063 16815 6089
rect 16841 6063 16847 6089
rect 17705 6063 17711 6089
rect 17737 6063 17743 6089
rect 18545 6063 18551 6089
rect 18577 6063 18583 6089
rect 19441 6063 19447 6089
rect 19473 6063 19479 6089
rect 20785 6063 20791 6089
rect 20817 6063 20823 6089
rect 21289 6063 21295 6089
rect 21321 6063 21327 6089
rect 21457 6063 21463 6089
rect 21489 6063 21495 6089
rect 22241 6063 22247 6089
rect 22273 6063 22279 6089
rect 22689 6063 22695 6089
rect 22721 6063 22727 6089
rect 22913 6063 22919 6089
rect 22945 6063 22951 6089
rect 24761 6063 24767 6089
rect 24793 6063 24799 6089
rect 25209 6063 25215 6089
rect 25241 6063 25247 6089
rect 25433 6063 25439 6089
rect 25465 6063 25471 6089
rect 26217 6063 26223 6089
rect 26249 6063 26255 6089
rect 26889 6063 26895 6089
rect 26921 6063 26927 6089
rect 28737 6063 28743 6089
rect 28769 6063 28775 6089
rect 29913 6063 29919 6089
rect 29945 6063 29951 6089
rect 30249 6063 30255 6089
rect 30281 6063 30287 6089
rect 31369 6063 31375 6089
rect 31401 6063 31407 6089
rect 32047 6057 32073 6063
rect 32159 6089 32185 6095
rect 32159 6057 32185 6063
rect 32327 6089 32353 6095
rect 35631 6089 35657 6095
rect 32713 6063 32719 6089
rect 32745 6063 32751 6089
rect 33609 6063 33615 6089
rect 33641 6063 33647 6089
rect 34393 6063 34399 6089
rect 34425 6063 34431 6089
rect 35121 6063 35127 6089
rect 35153 6063 35159 6089
rect 32327 6057 32353 6063
rect 35631 6057 35657 6063
rect 35743 6089 35769 6095
rect 35743 6057 35769 6063
rect 35911 6089 35937 6095
rect 36689 6063 36695 6089
rect 36721 6063 36727 6089
rect 37641 6063 37647 6089
rect 37673 6063 37679 6089
rect 35911 6057 35937 6063
rect 672 5893 39312 5910
rect 672 5867 2074 5893
rect 2100 5867 2136 5893
rect 2162 5867 2198 5893
rect 2224 5867 2260 5893
rect 2286 5867 2322 5893
rect 2348 5867 2384 5893
rect 2410 5867 2446 5893
rect 2472 5867 2508 5893
rect 2534 5867 7074 5893
rect 7100 5867 7136 5893
rect 7162 5867 7198 5893
rect 7224 5867 7260 5893
rect 7286 5867 7322 5893
rect 7348 5867 7384 5893
rect 7410 5867 7446 5893
rect 7472 5867 7508 5893
rect 7534 5867 12074 5893
rect 12100 5867 12136 5893
rect 12162 5867 12198 5893
rect 12224 5867 12260 5893
rect 12286 5867 12322 5893
rect 12348 5867 12384 5893
rect 12410 5867 12446 5893
rect 12472 5867 12508 5893
rect 12534 5867 17074 5893
rect 17100 5867 17136 5893
rect 17162 5867 17198 5893
rect 17224 5867 17260 5893
rect 17286 5867 17322 5893
rect 17348 5867 17384 5893
rect 17410 5867 17446 5893
rect 17472 5867 17508 5893
rect 17534 5867 22074 5893
rect 22100 5867 22136 5893
rect 22162 5867 22198 5893
rect 22224 5867 22260 5893
rect 22286 5867 22322 5893
rect 22348 5867 22384 5893
rect 22410 5867 22446 5893
rect 22472 5867 22508 5893
rect 22534 5867 27074 5893
rect 27100 5867 27136 5893
rect 27162 5867 27198 5893
rect 27224 5867 27260 5893
rect 27286 5867 27322 5893
rect 27348 5867 27384 5893
rect 27410 5867 27446 5893
rect 27472 5867 27508 5893
rect 27534 5867 32074 5893
rect 32100 5867 32136 5893
rect 32162 5867 32198 5893
rect 32224 5867 32260 5893
rect 32286 5867 32322 5893
rect 32348 5867 32384 5893
rect 32410 5867 32446 5893
rect 32472 5867 32508 5893
rect 32534 5867 37074 5893
rect 37100 5867 37136 5893
rect 37162 5867 37198 5893
rect 37224 5867 37260 5893
rect 37286 5867 37322 5893
rect 37348 5867 37384 5893
rect 37410 5867 37446 5893
rect 37472 5867 37508 5893
rect 37534 5867 39312 5893
rect 672 5850 39312 5867
rect 30087 5697 30113 5703
rect 33671 5697 33697 5703
rect 1801 5671 1807 5697
rect 1833 5671 1839 5697
rect 1969 5671 1975 5697
rect 2001 5671 2007 5697
rect 2473 5671 2479 5697
rect 2505 5671 2511 5697
rect 4097 5671 4103 5697
rect 4129 5671 4135 5697
rect 4993 5671 4999 5697
rect 5025 5671 5031 5697
rect 5273 5671 5279 5697
rect 5305 5671 5311 5697
rect 5833 5671 5839 5697
rect 5865 5671 5871 5697
rect 5945 5671 5951 5697
rect 5977 5671 5983 5697
rect 8073 5671 8079 5697
rect 8105 5671 8111 5697
rect 8969 5671 8975 5697
rect 9001 5671 9007 5697
rect 9417 5671 9423 5697
rect 9449 5671 9455 5697
rect 10257 5671 10263 5697
rect 10289 5671 10295 5697
rect 11993 5671 11999 5697
rect 12025 5671 12031 5697
rect 12945 5671 12951 5697
rect 12977 5671 12983 5697
rect 13337 5671 13343 5697
rect 13369 5671 13375 5697
rect 14401 5671 14407 5697
rect 14433 5671 14439 5697
rect 15185 5671 15191 5697
rect 15217 5671 15223 5697
rect 15857 5671 15863 5697
rect 15889 5671 15895 5697
rect 16809 5671 16815 5697
rect 16841 5671 16847 5697
rect 17705 5671 17711 5697
rect 17737 5671 17743 5697
rect 18769 5671 18775 5697
rect 18801 5671 18807 5697
rect 19945 5671 19951 5697
rect 19977 5671 19983 5697
rect 20225 5671 20231 5697
rect 20257 5671 20263 5697
rect 21289 5671 21295 5697
rect 21321 5671 21327 5697
rect 22745 5671 22751 5697
rect 22777 5671 22783 5697
rect 23193 5671 23199 5697
rect 23225 5671 23231 5697
rect 23417 5671 23423 5697
rect 23449 5671 23455 5697
rect 24369 5671 24375 5697
rect 24401 5671 24407 5697
rect 25153 5671 25159 5697
rect 25185 5671 25191 5697
rect 26721 5671 26727 5697
rect 26753 5671 26759 5697
rect 27561 5671 27567 5697
rect 27593 5671 27599 5697
rect 28233 5671 28239 5697
rect 28265 5671 28271 5697
rect 29129 5671 29135 5697
rect 29161 5671 29167 5697
rect 30697 5671 30703 5697
rect 30729 5671 30735 5697
rect 31873 5671 31879 5697
rect 31905 5671 31911 5697
rect 32153 5671 32159 5697
rect 32185 5671 32191 5697
rect 33329 5671 33335 5697
rect 33361 5671 33367 5697
rect 34953 5671 34959 5697
rect 34985 5671 34991 5697
rect 35121 5671 35127 5697
rect 35153 5671 35159 5697
rect 35345 5671 35351 5697
rect 35377 5671 35383 5697
rect 36129 5671 36135 5697
rect 36161 5671 36167 5697
rect 37137 5671 37143 5697
rect 37169 5671 37175 5697
rect 30087 5665 30113 5671
rect 33671 5665 33697 5671
rect 30143 5641 30169 5647
rect 4993 5615 4999 5641
rect 5025 5615 5031 5641
rect 8969 5615 8975 5641
rect 9001 5615 9007 5641
rect 10257 5615 10263 5641
rect 10289 5615 10295 5641
rect 12945 5615 12951 5641
rect 12977 5615 12983 5641
rect 14401 5615 14407 5641
rect 14433 5615 14439 5641
rect 16025 5615 16031 5641
rect 16057 5615 16063 5641
rect 17705 5615 17711 5641
rect 17737 5615 17743 5641
rect 19945 5615 19951 5641
rect 19977 5615 19983 5641
rect 21289 5615 21295 5641
rect 21321 5615 21327 5641
rect 25153 5615 25159 5641
rect 25185 5615 25191 5641
rect 27673 5615 27679 5641
rect 27705 5615 27711 5641
rect 29129 5615 29135 5641
rect 29161 5615 29167 5641
rect 30143 5609 30169 5615
rect 30311 5641 30337 5647
rect 33727 5641 33753 5647
rect 31873 5615 31879 5641
rect 31905 5615 31911 5641
rect 33329 5615 33335 5641
rect 33361 5615 33367 5641
rect 30311 5609 30337 5615
rect 33727 5609 33753 5615
rect 33895 5641 33921 5647
rect 37591 5641 37617 5647
rect 37137 5615 37143 5641
rect 37169 5615 37175 5641
rect 33895 5609 33921 5615
rect 37591 5609 37617 5615
rect 37703 5641 37729 5647
rect 37703 5609 37729 5615
rect 37871 5641 37897 5647
rect 37871 5609 37897 5615
rect 672 5501 39312 5518
rect 672 5475 4574 5501
rect 4600 5475 4636 5501
rect 4662 5475 4698 5501
rect 4724 5475 4760 5501
rect 4786 5475 4822 5501
rect 4848 5475 4884 5501
rect 4910 5475 4946 5501
rect 4972 5475 5008 5501
rect 5034 5475 9574 5501
rect 9600 5475 9636 5501
rect 9662 5475 9698 5501
rect 9724 5475 9760 5501
rect 9786 5475 9822 5501
rect 9848 5475 9884 5501
rect 9910 5475 9946 5501
rect 9972 5475 10008 5501
rect 10034 5475 14574 5501
rect 14600 5475 14636 5501
rect 14662 5475 14698 5501
rect 14724 5475 14760 5501
rect 14786 5475 14822 5501
rect 14848 5475 14884 5501
rect 14910 5475 14946 5501
rect 14972 5475 15008 5501
rect 15034 5475 19574 5501
rect 19600 5475 19636 5501
rect 19662 5475 19698 5501
rect 19724 5475 19760 5501
rect 19786 5475 19822 5501
rect 19848 5475 19884 5501
rect 19910 5475 19946 5501
rect 19972 5475 20008 5501
rect 20034 5475 24574 5501
rect 24600 5475 24636 5501
rect 24662 5475 24698 5501
rect 24724 5475 24760 5501
rect 24786 5475 24822 5501
rect 24848 5475 24884 5501
rect 24910 5475 24946 5501
rect 24972 5475 25008 5501
rect 25034 5475 29574 5501
rect 29600 5475 29636 5501
rect 29662 5475 29698 5501
rect 29724 5475 29760 5501
rect 29786 5475 29822 5501
rect 29848 5475 29884 5501
rect 29910 5475 29946 5501
rect 29972 5475 30008 5501
rect 30034 5475 34574 5501
rect 34600 5475 34636 5501
rect 34662 5475 34698 5501
rect 34724 5475 34760 5501
rect 34786 5475 34822 5501
rect 34848 5475 34884 5501
rect 34910 5475 34946 5501
rect 34972 5475 35008 5501
rect 35034 5475 39312 5501
rect 672 5458 39312 5475
rect 28071 5361 28097 5367
rect 1969 5335 1975 5361
rect 2001 5335 2007 5361
rect 4489 5335 4495 5361
rect 4521 5335 4527 5361
rect 6785 5335 6791 5361
rect 6817 5335 6823 5361
rect 8465 5335 8471 5361
rect 8497 5335 8503 5361
rect 12441 5335 12447 5361
rect 12473 5335 12479 5361
rect 14457 5335 14463 5361
rect 14489 5335 14495 5361
rect 15857 5335 15863 5361
rect 15889 5335 15895 5361
rect 17761 5335 17767 5361
rect 17793 5335 17799 5361
rect 19441 5335 19447 5361
rect 19473 5335 19479 5361
rect 23193 5335 23199 5361
rect 23225 5335 23231 5361
rect 29689 5335 29695 5361
rect 29721 5335 29727 5361
rect 31369 5335 31375 5361
rect 31401 5335 31407 5361
rect 33833 5335 33839 5361
rect 33865 5335 33871 5361
rect 35233 5335 35239 5361
rect 35265 5335 35271 5361
rect 28071 5329 28097 5335
rect 28183 5305 28209 5311
rect 1969 5279 1975 5305
rect 2001 5279 2007 5305
rect 3033 5279 3039 5305
rect 3065 5279 3071 5305
rect 3425 5279 3431 5305
rect 3457 5279 3463 5305
rect 4489 5279 4495 5305
rect 4521 5279 4527 5305
rect 6113 5279 6119 5305
rect 6145 5279 6151 5305
rect 6785 5279 6791 5305
rect 6817 5279 6823 5305
rect 7289 5279 7295 5305
rect 7321 5279 7327 5305
rect 8465 5279 8471 5305
rect 8497 5279 8503 5305
rect 10033 5279 10039 5305
rect 10065 5279 10071 5305
rect 10313 5279 10319 5305
rect 10345 5279 10351 5305
rect 10481 5279 10487 5305
rect 10513 5279 10519 5305
rect 11545 5279 11551 5305
rect 11577 5279 11583 5305
rect 12441 5279 12447 5305
rect 12473 5279 12479 5305
rect 13561 5279 13567 5305
rect 13593 5279 13599 5305
rect 14457 5279 14463 5305
rect 14489 5279 14495 5305
rect 15185 5279 15191 5305
rect 15217 5279 15223 5305
rect 15857 5279 15863 5305
rect 15889 5279 15895 5305
rect 16809 5279 16815 5305
rect 16841 5279 16847 5305
rect 17761 5279 17767 5305
rect 17793 5279 17799 5305
rect 18545 5279 18551 5305
rect 18577 5279 18583 5305
rect 19441 5279 19447 5305
rect 19473 5279 19479 5305
rect 20785 5279 20791 5305
rect 20817 5279 20823 5305
rect 21289 5279 21295 5305
rect 21321 5279 21327 5305
rect 21457 5279 21463 5305
rect 21489 5279 21495 5305
rect 22521 5279 22527 5305
rect 22553 5279 22559 5305
rect 23193 5279 23199 5305
rect 23225 5279 23231 5305
rect 24761 5279 24767 5305
rect 24793 5279 24799 5305
rect 25209 5279 25215 5305
rect 25241 5279 25247 5305
rect 25937 5279 25943 5305
rect 25969 5279 25975 5305
rect 26217 5279 26223 5305
rect 26249 5279 26255 5305
rect 26777 5279 26783 5305
rect 26809 5279 26815 5305
rect 26889 5279 26895 5305
rect 26921 5279 26927 5305
rect 28183 5273 28209 5279
rect 28407 5305 28433 5311
rect 32047 5305 32073 5311
rect 28737 5279 28743 5305
rect 28769 5279 28775 5305
rect 29465 5279 29471 5305
rect 29497 5279 29503 5305
rect 30361 5279 30367 5305
rect 30393 5279 30399 5305
rect 31369 5279 31375 5305
rect 31401 5279 31407 5305
rect 28407 5273 28433 5279
rect 32047 5273 32073 5279
rect 32159 5305 32185 5311
rect 32159 5273 32185 5279
rect 32327 5305 32353 5311
rect 35631 5305 35657 5311
rect 32769 5279 32775 5305
rect 32801 5279 32807 5305
rect 33833 5279 33839 5305
rect 33865 5279 33871 5305
rect 34169 5279 34175 5305
rect 34201 5279 34207 5305
rect 35233 5279 35239 5305
rect 35265 5279 35271 5305
rect 32327 5273 32353 5279
rect 35631 5273 35657 5279
rect 35743 5305 35769 5311
rect 35743 5273 35769 5279
rect 35911 5305 35937 5311
rect 38151 5305 38177 5311
rect 36689 5279 36695 5305
rect 36721 5279 36727 5305
rect 37137 5279 37143 5305
rect 37169 5279 37175 5305
rect 37361 5279 37367 5305
rect 37393 5279 37399 5305
rect 35911 5273 35937 5279
rect 38151 5273 38177 5279
rect 38263 5305 38289 5311
rect 38263 5273 38289 5279
rect 38431 5305 38457 5311
rect 38431 5273 38457 5279
rect 672 5109 39312 5126
rect 672 5083 2074 5109
rect 2100 5083 2136 5109
rect 2162 5083 2198 5109
rect 2224 5083 2260 5109
rect 2286 5083 2322 5109
rect 2348 5083 2384 5109
rect 2410 5083 2446 5109
rect 2472 5083 2508 5109
rect 2534 5083 7074 5109
rect 7100 5083 7136 5109
rect 7162 5083 7198 5109
rect 7224 5083 7260 5109
rect 7286 5083 7322 5109
rect 7348 5083 7384 5109
rect 7410 5083 7446 5109
rect 7472 5083 7508 5109
rect 7534 5083 12074 5109
rect 12100 5083 12136 5109
rect 12162 5083 12198 5109
rect 12224 5083 12260 5109
rect 12286 5083 12322 5109
rect 12348 5083 12384 5109
rect 12410 5083 12446 5109
rect 12472 5083 12508 5109
rect 12534 5083 17074 5109
rect 17100 5083 17136 5109
rect 17162 5083 17198 5109
rect 17224 5083 17260 5109
rect 17286 5083 17322 5109
rect 17348 5083 17384 5109
rect 17410 5083 17446 5109
rect 17472 5083 17508 5109
rect 17534 5083 22074 5109
rect 22100 5083 22136 5109
rect 22162 5083 22198 5109
rect 22224 5083 22260 5109
rect 22286 5083 22322 5109
rect 22348 5083 22384 5109
rect 22410 5083 22446 5109
rect 22472 5083 22508 5109
rect 22534 5083 27074 5109
rect 27100 5083 27136 5109
rect 27162 5083 27198 5109
rect 27224 5083 27260 5109
rect 27286 5083 27322 5109
rect 27348 5083 27384 5109
rect 27410 5083 27446 5109
rect 27472 5083 27508 5109
rect 27534 5083 32074 5109
rect 32100 5083 32136 5109
rect 32162 5083 32198 5109
rect 32224 5083 32260 5109
rect 32286 5083 32322 5109
rect 32348 5083 32384 5109
rect 32410 5083 32446 5109
rect 32472 5083 32508 5109
rect 32534 5083 37074 5109
rect 37100 5083 37136 5109
rect 37162 5083 37198 5109
rect 37224 5083 37260 5109
rect 37286 5083 37322 5109
rect 37348 5083 37384 5109
rect 37410 5083 37446 5109
rect 37472 5083 37508 5109
rect 37534 5083 39312 5109
rect 672 5066 39312 5083
rect 30087 4913 30113 4919
rect 1801 4887 1807 4913
rect 1833 4887 1839 4913
rect 1913 4887 1919 4913
rect 1945 4887 1951 4913
rect 2473 4887 2479 4913
rect 2505 4887 2511 4913
rect 4097 4887 4103 4913
rect 4129 4887 4135 4913
rect 4993 4887 4999 4913
rect 5025 4887 5031 4913
rect 5273 4887 5279 4913
rect 5305 4887 5311 4913
rect 6449 4887 6455 4913
rect 6481 4887 6487 4913
rect 8073 4887 8079 4913
rect 8105 4887 8111 4913
rect 8969 4887 8975 4913
rect 9001 4887 9007 4913
rect 9417 4887 9423 4913
rect 9449 4887 9455 4913
rect 10313 4887 10319 4913
rect 10345 4887 10351 4913
rect 11993 4887 11999 4913
rect 12025 4887 12031 4913
rect 12945 4887 12951 4913
rect 12977 4887 12983 4913
rect 13337 4887 13343 4913
rect 13369 4887 13375 4913
rect 14177 4887 14183 4913
rect 14209 4887 14215 4913
rect 15577 4887 15583 4913
rect 15609 4887 15615 4913
rect 15801 4887 15807 4913
rect 15833 4887 15839 4913
rect 16025 4887 16031 4913
rect 16057 4887 16063 4913
rect 16809 4887 16815 4913
rect 16841 4887 16847 4913
rect 17761 4887 17767 4913
rect 17793 4887 17799 4913
rect 18769 4887 18775 4913
rect 18801 4887 18807 4913
rect 19945 4887 19951 4913
rect 19977 4887 19983 4913
rect 20225 4887 20231 4913
rect 20257 4887 20263 4913
rect 21289 4887 21295 4913
rect 21321 4887 21327 4913
rect 22745 4887 22751 4913
rect 22777 4887 22783 4913
rect 23193 4887 23199 4913
rect 23225 4887 23231 4913
rect 23417 4887 23423 4913
rect 23449 4887 23455 4913
rect 24369 4887 24375 4913
rect 24401 4887 24407 4913
rect 25209 4887 25215 4913
rect 25241 4887 25247 4913
rect 26721 4887 26727 4913
rect 26753 4887 26759 4913
rect 27281 4887 27287 4913
rect 27313 4887 27319 4913
rect 27393 4887 27399 4913
rect 27425 4887 27431 4913
rect 28233 4887 28239 4913
rect 28265 4887 28271 4913
rect 29129 4887 29135 4913
rect 29161 4887 29167 4913
rect 30087 4881 30113 4887
rect 30199 4913 30225 4919
rect 30199 4881 30225 4887
rect 30311 4913 30337 4919
rect 33671 4913 33697 4919
rect 30697 4887 30703 4913
rect 30729 4887 30735 4913
rect 31873 4887 31879 4913
rect 31905 4887 31911 4913
rect 32153 4887 32159 4913
rect 32185 4887 32191 4913
rect 33329 4887 33335 4913
rect 33361 4887 33367 4913
rect 30311 4881 30337 4887
rect 33671 4881 33697 4887
rect 33783 4913 33809 4919
rect 33783 4881 33809 4887
rect 33895 4913 33921 4919
rect 37591 4913 37617 4919
rect 34673 4887 34679 4913
rect 34705 4887 34711 4913
rect 35849 4887 35855 4913
rect 35881 4887 35887 4913
rect 36129 4887 36135 4913
rect 36161 4887 36167 4913
rect 37305 4887 37311 4913
rect 37337 4887 37343 4913
rect 33895 4881 33921 4887
rect 37591 4881 37617 4887
rect 37759 4913 37785 4919
rect 37759 4881 37785 4887
rect 37871 4913 37897 4919
rect 37871 4881 37897 4887
rect 38655 4913 38681 4919
rect 38655 4881 38681 4887
rect 38767 4913 38793 4919
rect 38767 4881 38793 4887
rect 38879 4913 38905 4919
rect 38879 4881 38905 4887
rect 4993 4831 4999 4857
rect 5025 4831 5031 4857
rect 6449 4831 6455 4857
rect 6481 4831 6487 4857
rect 8969 4831 8975 4857
rect 9001 4831 9007 4857
rect 10313 4831 10319 4857
rect 10345 4831 10351 4857
rect 12945 4831 12951 4857
rect 12977 4831 12983 4857
rect 14177 4831 14183 4857
rect 14209 4831 14215 4857
rect 17761 4831 17767 4857
rect 17793 4831 17799 4857
rect 19945 4831 19951 4857
rect 19977 4831 19983 4857
rect 21289 4831 21295 4857
rect 21321 4831 21327 4857
rect 25209 4831 25215 4857
rect 25241 4831 25247 4857
rect 29129 4831 29135 4857
rect 29161 4831 29167 4857
rect 31873 4831 31879 4857
rect 31905 4831 31911 4857
rect 33329 4831 33335 4857
rect 33361 4831 33367 4857
rect 35849 4831 35855 4857
rect 35881 4831 35887 4857
rect 37305 4831 37311 4857
rect 37337 4831 37343 4857
rect 672 4717 39312 4734
rect 672 4691 4574 4717
rect 4600 4691 4636 4717
rect 4662 4691 4698 4717
rect 4724 4691 4760 4717
rect 4786 4691 4822 4717
rect 4848 4691 4884 4717
rect 4910 4691 4946 4717
rect 4972 4691 5008 4717
rect 5034 4691 9574 4717
rect 9600 4691 9636 4717
rect 9662 4691 9698 4717
rect 9724 4691 9760 4717
rect 9786 4691 9822 4717
rect 9848 4691 9884 4717
rect 9910 4691 9946 4717
rect 9972 4691 10008 4717
rect 10034 4691 14574 4717
rect 14600 4691 14636 4717
rect 14662 4691 14698 4717
rect 14724 4691 14760 4717
rect 14786 4691 14822 4717
rect 14848 4691 14884 4717
rect 14910 4691 14946 4717
rect 14972 4691 15008 4717
rect 15034 4691 19574 4717
rect 19600 4691 19636 4717
rect 19662 4691 19698 4717
rect 19724 4691 19760 4717
rect 19786 4691 19822 4717
rect 19848 4691 19884 4717
rect 19910 4691 19946 4717
rect 19972 4691 20008 4717
rect 20034 4691 24574 4717
rect 24600 4691 24636 4717
rect 24662 4691 24698 4717
rect 24724 4691 24760 4717
rect 24786 4691 24822 4717
rect 24848 4691 24884 4717
rect 24910 4691 24946 4717
rect 24972 4691 25008 4717
rect 25034 4691 29574 4717
rect 29600 4691 29636 4717
rect 29662 4691 29698 4717
rect 29724 4691 29760 4717
rect 29786 4691 29822 4717
rect 29848 4691 29884 4717
rect 29910 4691 29946 4717
rect 29972 4691 30008 4717
rect 30034 4691 34574 4717
rect 34600 4691 34636 4717
rect 34662 4691 34698 4717
rect 34724 4691 34760 4717
rect 34786 4691 34822 4717
rect 34848 4691 34884 4717
rect 34910 4691 34946 4717
rect 34972 4691 35008 4717
rect 35034 4691 39312 4717
rect 672 4674 39312 4691
rect 28183 4577 28209 4583
rect 35911 4577 35937 4583
rect 38151 4577 38177 4583
rect 1857 4551 1863 4577
rect 1889 4551 1895 4577
rect 4489 4551 4495 4577
rect 4521 4551 4527 4577
rect 6785 4551 6791 4577
rect 6817 4551 6823 4577
rect 8465 4551 8471 4577
rect 8497 4551 8503 4577
rect 12441 4551 12447 4577
rect 12473 4551 12479 4577
rect 17761 4551 17767 4577
rect 17793 4551 17799 4577
rect 19441 4551 19447 4577
rect 19473 4551 19479 4577
rect 21793 4551 21799 4577
rect 21825 4551 21831 4577
rect 27393 4551 27399 4577
rect 27425 4551 27431 4577
rect 31369 4551 31375 4577
rect 31401 4551 31407 4577
rect 33833 4551 33839 4577
rect 33865 4551 33871 4577
rect 37641 4551 37647 4577
rect 37673 4551 37679 4577
rect 28183 4545 28209 4551
rect 35911 4545 35937 4551
rect 38151 4545 38177 4551
rect 38263 4577 38289 4583
rect 38263 4545 38289 4551
rect 38431 4577 38457 4583
rect 38431 4545 38457 4551
rect 38711 4577 38737 4583
rect 38711 4545 38737 4551
rect 28127 4521 28153 4527
rect 1857 4495 1863 4521
rect 1889 4495 1895 4521
rect 3033 4495 3039 4521
rect 3065 4495 3071 4521
rect 3425 4495 3431 4521
rect 3457 4495 3463 4521
rect 4489 4495 4495 4521
rect 4521 4495 4527 4521
rect 6113 4495 6119 4521
rect 6145 4495 6151 4521
rect 6785 4495 6791 4521
rect 6817 4495 6823 4521
rect 7569 4495 7575 4521
rect 7601 4495 7607 4521
rect 8465 4495 8471 4521
rect 8497 4495 8503 4521
rect 10033 4495 10039 4521
rect 10065 4495 10071 4521
rect 10313 4495 10319 4521
rect 10345 4495 10351 4521
rect 10481 4495 10487 4521
rect 10513 4495 10519 4521
rect 11545 4495 11551 4521
rect 11577 4495 11583 4521
rect 12441 4495 12447 4521
rect 12473 4495 12479 4521
rect 13561 4495 13567 4521
rect 13593 4495 13599 4521
rect 14121 4495 14127 4521
rect 14153 4495 14159 4521
rect 14233 4495 14239 4521
rect 14265 4495 14271 4521
rect 15129 4495 15135 4521
rect 15161 4495 15167 4521
rect 15465 4495 15471 4521
rect 15497 4495 15503 4521
rect 15689 4495 15695 4521
rect 15721 4495 15727 4521
rect 16809 4495 16815 4521
rect 16841 4495 16847 4521
rect 17761 4495 17767 4521
rect 17793 4495 17799 4521
rect 18545 4495 18551 4521
rect 18577 4495 18583 4521
rect 19441 4495 19447 4521
rect 19473 4495 19479 4521
rect 20785 4495 20791 4521
rect 20817 4495 20823 4521
rect 21793 4495 21799 4521
rect 21825 4495 21831 4521
rect 22521 4495 22527 4521
rect 22553 4495 22559 4521
rect 22689 4495 22695 4521
rect 22721 4495 22727 4521
rect 22913 4495 22919 4521
rect 22945 4495 22951 4521
rect 24761 4495 24767 4521
rect 24793 4495 24799 4521
rect 25209 4495 25215 4521
rect 25241 4495 25247 4521
rect 25937 4495 25943 4521
rect 25969 4495 25975 4521
rect 26273 4495 26279 4521
rect 26305 4495 26311 4521
rect 27393 4495 27399 4521
rect 27425 4495 27431 4521
rect 28127 4489 28153 4495
rect 28351 4521 28377 4527
rect 32047 4521 32073 4527
rect 28737 4495 28743 4521
rect 28769 4495 28775 4521
rect 29185 4495 29191 4521
rect 29217 4495 29223 4521
rect 29409 4495 29415 4521
rect 29441 4495 29447 4521
rect 30361 4495 30367 4521
rect 30393 4495 30399 4521
rect 31369 4495 31375 4521
rect 31401 4495 31407 4521
rect 28351 4489 28377 4495
rect 32047 4489 32073 4495
rect 32215 4521 32241 4527
rect 32215 4489 32241 4495
rect 32383 4521 32409 4527
rect 35687 4521 35713 4527
rect 32769 4495 32775 4521
rect 32801 4495 32807 4521
rect 33833 4495 33839 4521
rect 33865 4495 33871 4521
rect 34169 4495 34175 4521
rect 34201 4495 34207 4521
rect 34617 4495 34623 4521
rect 34649 4495 34655 4521
rect 34841 4495 34847 4521
rect 34873 4495 34879 4521
rect 32383 4489 32409 4495
rect 35687 4489 35713 4495
rect 35799 4521 35825 4527
rect 38823 4521 38849 4527
rect 36689 4495 36695 4521
rect 36721 4495 36727 4521
rect 37641 4495 37647 4521
rect 37673 4495 37679 4521
rect 35799 4489 35825 4495
rect 38823 4489 38849 4495
rect 38935 4521 38961 4527
rect 38935 4489 38961 4495
rect 672 4325 39312 4342
rect 672 4299 2074 4325
rect 2100 4299 2136 4325
rect 2162 4299 2198 4325
rect 2224 4299 2260 4325
rect 2286 4299 2322 4325
rect 2348 4299 2384 4325
rect 2410 4299 2446 4325
rect 2472 4299 2508 4325
rect 2534 4299 7074 4325
rect 7100 4299 7136 4325
rect 7162 4299 7198 4325
rect 7224 4299 7260 4325
rect 7286 4299 7322 4325
rect 7348 4299 7384 4325
rect 7410 4299 7446 4325
rect 7472 4299 7508 4325
rect 7534 4299 12074 4325
rect 12100 4299 12136 4325
rect 12162 4299 12198 4325
rect 12224 4299 12260 4325
rect 12286 4299 12322 4325
rect 12348 4299 12384 4325
rect 12410 4299 12446 4325
rect 12472 4299 12508 4325
rect 12534 4299 17074 4325
rect 17100 4299 17136 4325
rect 17162 4299 17198 4325
rect 17224 4299 17260 4325
rect 17286 4299 17322 4325
rect 17348 4299 17384 4325
rect 17410 4299 17446 4325
rect 17472 4299 17508 4325
rect 17534 4299 22074 4325
rect 22100 4299 22136 4325
rect 22162 4299 22198 4325
rect 22224 4299 22260 4325
rect 22286 4299 22322 4325
rect 22348 4299 22384 4325
rect 22410 4299 22446 4325
rect 22472 4299 22508 4325
rect 22534 4299 27074 4325
rect 27100 4299 27136 4325
rect 27162 4299 27198 4325
rect 27224 4299 27260 4325
rect 27286 4299 27322 4325
rect 27348 4299 27384 4325
rect 27410 4299 27446 4325
rect 27472 4299 27508 4325
rect 27534 4299 32074 4325
rect 32100 4299 32136 4325
rect 32162 4299 32198 4325
rect 32224 4299 32260 4325
rect 32286 4299 32322 4325
rect 32348 4299 32384 4325
rect 32410 4299 32446 4325
rect 32472 4299 32508 4325
rect 32534 4299 37074 4325
rect 37100 4299 37136 4325
rect 37162 4299 37198 4325
rect 37224 4299 37260 4325
rect 37286 4299 37322 4325
rect 37348 4299 37384 4325
rect 37410 4299 37446 4325
rect 37472 4299 37508 4325
rect 37534 4299 39312 4325
rect 672 4282 39312 4299
rect 30199 4129 30225 4135
rect 1801 4103 1807 4129
rect 1833 4103 1839 4129
rect 1913 4103 1919 4129
rect 1945 4103 1951 4129
rect 2473 4103 2479 4129
rect 2505 4103 2511 4129
rect 4097 4103 4103 4129
rect 4129 4103 4135 4129
rect 4769 4103 4775 4129
rect 4801 4103 4807 4129
rect 5273 4103 5279 4129
rect 5305 4103 5311 4129
rect 6449 4103 6455 4129
rect 6481 4103 6487 4129
rect 8073 4103 8079 4129
rect 8105 4103 8111 4129
rect 8969 4103 8975 4129
rect 9001 4103 9007 4129
rect 9529 4103 9535 4129
rect 9561 4103 9567 4129
rect 10313 4103 10319 4129
rect 10345 4103 10351 4129
rect 11993 4103 11999 4129
rect 12025 4103 12031 4129
rect 12721 4103 12727 4129
rect 12753 4103 12759 4129
rect 13337 4103 13343 4129
rect 13369 4103 13375 4129
rect 14233 4103 14239 4129
rect 14265 4103 14271 4129
rect 15521 4103 15527 4129
rect 15553 4103 15559 4129
rect 15801 4103 15807 4129
rect 15833 4103 15839 4129
rect 16025 4103 16031 4129
rect 16057 4103 16063 4129
rect 16809 4103 16815 4129
rect 16841 4103 16847 4129
rect 17761 4103 17767 4129
rect 17793 4103 17799 4129
rect 18769 4103 18775 4129
rect 18801 4103 18807 4129
rect 19945 4103 19951 4129
rect 19977 4103 19983 4129
rect 20225 4103 20231 4129
rect 20257 4103 20263 4129
rect 21177 4103 21183 4129
rect 21209 4103 21215 4129
rect 22745 4103 22751 4129
rect 22777 4103 22783 4129
rect 23305 4103 23311 4129
rect 23337 4103 23343 4129
rect 23417 4103 23423 4129
rect 23449 4103 23455 4129
rect 24369 4103 24375 4129
rect 24401 4103 24407 4129
rect 24649 4103 24655 4129
rect 24681 4103 24687 4129
rect 24873 4103 24879 4129
rect 24905 4103 24911 4129
rect 26721 4103 26727 4129
rect 26753 4103 26759 4129
rect 27169 4103 27175 4129
rect 27201 4103 27207 4129
rect 27393 4103 27399 4129
rect 27425 4103 27431 4129
rect 28457 4103 28463 4129
rect 28489 4103 28495 4129
rect 29353 4103 29359 4129
rect 29385 4103 29391 4129
rect 30199 4097 30225 4103
rect 30311 4129 30337 4135
rect 33671 4129 33697 4135
rect 30697 4103 30703 4129
rect 30729 4103 30735 4129
rect 31873 4103 31879 4129
rect 31905 4103 31911 4129
rect 32153 4103 32159 4129
rect 32185 4103 32191 4129
rect 33329 4103 33335 4129
rect 33361 4103 33367 4129
rect 30311 4097 30337 4103
rect 33671 4097 33697 4103
rect 33783 4129 33809 4135
rect 33783 4097 33809 4103
rect 33951 4129 33977 4135
rect 37591 4129 37617 4135
rect 34673 4103 34679 4129
rect 34705 4103 34711 4129
rect 35177 4103 35183 4129
rect 35209 4103 35215 4129
rect 35345 4103 35351 4129
rect 35377 4103 35383 4129
rect 36129 4103 36135 4129
rect 36161 4103 36167 4129
rect 37081 4103 37087 4129
rect 37113 4103 37119 4129
rect 33951 4097 33977 4103
rect 37591 4097 37617 4103
rect 37703 4129 37729 4135
rect 37703 4097 37729 4103
rect 37871 4129 37897 4135
rect 37871 4097 37897 4103
rect 38655 4129 38681 4135
rect 38655 4097 38681 4103
rect 38767 4129 38793 4135
rect 38767 4097 38793 4103
rect 30031 4073 30057 4079
rect 38935 4073 38961 4079
rect 4769 4047 4775 4073
rect 4801 4047 4807 4073
rect 6449 4047 6455 4073
rect 6481 4047 6487 4073
rect 8969 4047 8975 4073
rect 9001 4047 9007 4073
rect 10313 4047 10319 4073
rect 10345 4047 10351 4073
rect 12721 4047 12727 4073
rect 12753 4047 12759 4073
rect 14233 4047 14239 4073
rect 14265 4047 14271 4073
rect 17761 4047 17767 4073
rect 17793 4047 17799 4073
rect 19945 4047 19951 4073
rect 19977 4047 19983 4073
rect 21177 4047 21183 4073
rect 21209 4047 21215 4073
rect 29353 4047 29359 4073
rect 29385 4047 29391 4073
rect 31873 4047 31879 4073
rect 31905 4047 31911 4073
rect 33329 4047 33335 4073
rect 33361 4047 33367 4073
rect 37081 4047 37087 4073
rect 37113 4047 37119 4073
rect 30031 4041 30057 4047
rect 38935 4041 38961 4047
rect 672 3933 39312 3950
rect 672 3907 4574 3933
rect 4600 3907 4636 3933
rect 4662 3907 4698 3933
rect 4724 3907 4760 3933
rect 4786 3907 4822 3933
rect 4848 3907 4884 3933
rect 4910 3907 4946 3933
rect 4972 3907 5008 3933
rect 5034 3907 9574 3933
rect 9600 3907 9636 3933
rect 9662 3907 9698 3933
rect 9724 3907 9760 3933
rect 9786 3907 9822 3933
rect 9848 3907 9884 3933
rect 9910 3907 9946 3933
rect 9972 3907 10008 3933
rect 10034 3907 14574 3933
rect 14600 3907 14636 3933
rect 14662 3907 14698 3933
rect 14724 3907 14760 3933
rect 14786 3907 14822 3933
rect 14848 3907 14884 3933
rect 14910 3907 14946 3933
rect 14972 3907 15008 3933
rect 15034 3907 19574 3933
rect 19600 3907 19636 3933
rect 19662 3907 19698 3933
rect 19724 3907 19760 3933
rect 19786 3907 19822 3933
rect 19848 3907 19884 3933
rect 19910 3907 19946 3933
rect 19972 3907 20008 3933
rect 20034 3907 24574 3933
rect 24600 3907 24636 3933
rect 24662 3907 24698 3933
rect 24724 3907 24760 3933
rect 24786 3907 24822 3933
rect 24848 3907 24884 3933
rect 24910 3907 24946 3933
rect 24972 3907 25008 3933
rect 25034 3907 29574 3933
rect 29600 3907 29636 3933
rect 29662 3907 29698 3933
rect 29724 3907 29760 3933
rect 29786 3907 29822 3933
rect 29848 3907 29884 3933
rect 29910 3907 29946 3933
rect 29972 3907 30008 3933
rect 30034 3907 34574 3933
rect 34600 3907 34636 3933
rect 34662 3907 34698 3933
rect 34724 3907 34760 3933
rect 34786 3907 34822 3933
rect 34848 3907 34884 3933
rect 34910 3907 34946 3933
rect 34972 3907 35008 3933
rect 35034 3907 39312 3933
rect 672 3890 39312 3907
rect 28351 3793 28377 3799
rect 35743 3793 35769 3799
rect 1913 3767 1919 3793
rect 1945 3767 1951 3793
rect 4489 3767 4495 3793
rect 4521 3767 4527 3793
rect 6953 3767 6959 3793
rect 6985 3767 6991 3793
rect 8353 3767 8359 3793
rect 8385 3767 8391 3793
rect 12441 3767 12447 3793
rect 12473 3767 12479 3793
rect 17761 3767 17767 3793
rect 17793 3767 17799 3793
rect 19441 3767 19447 3793
rect 19473 3767 19479 3793
rect 21737 3767 21743 3793
rect 21769 3767 21775 3793
rect 27169 3767 27175 3793
rect 27201 3767 27207 3793
rect 29913 3767 29919 3793
rect 29945 3767 29951 3793
rect 31313 3767 31319 3793
rect 31345 3767 31351 3793
rect 33889 3767 33895 3793
rect 33921 3767 33927 3793
rect 35121 3767 35127 3793
rect 35153 3767 35159 3793
rect 28351 3761 28377 3767
rect 35743 3761 35769 3767
rect 35911 3793 35937 3799
rect 38263 3793 38289 3799
rect 36913 3767 36919 3793
rect 36945 3767 36951 3793
rect 35911 3761 35937 3767
rect 38263 3761 38289 3767
rect 38431 3793 38457 3799
rect 38431 3761 38457 3767
rect 38711 3793 38737 3799
rect 38711 3761 38737 3767
rect 28071 3737 28097 3743
rect 1913 3711 1919 3737
rect 1945 3711 1951 3737
rect 3033 3711 3039 3737
rect 3065 3711 3071 3737
rect 3481 3711 3487 3737
rect 3513 3711 3519 3737
rect 4489 3711 4495 3737
rect 4521 3711 4527 3737
rect 5833 3711 5839 3737
rect 5865 3711 5871 3737
rect 6953 3711 6959 3737
rect 6985 3711 6991 3737
rect 7569 3711 7575 3737
rect 7601 3711 7607 3737
rect 8353 3711 8359 3737
rect 8385 3711 8391 3737
rect 10033 3711 10039 3737
rect 10065 3711 10071 3737
rect 10257 3711 10263 3737
rect 10289 3711 10295 3737
rect 10481 3711 10487 3737
rect 10513 3711 10519 3737
rect 11545 3711 11551 3737
rect 11577 3711 11583 3737
rect 12441 3711 12447 3737
rect 12473 3711 12479 3737
rect 13673 3711 13679 3737
rect 13705 3711 13711 3737
rect 14121 3711 14127 3737
rect 14153 3711 14159 3737
rect 14345 3711 14351 3737
rect 14377 3711 14383 3737
rect 15129 3711 15135 3737
rect 15161 3711 15167 3737
rect 15577 3711 15583 3737
rect 15609 3711 15615 3737
rect 15801 3711 15807 3737
rect 15833 3711 15839 3737
rect 16809 3711 16815 3737
rect 16841 3711 16847 3737
rect 17761 3711 17767 3737
rect 17793 3711 17799 3737
rect 18545 3711 18551 3737
rect 18577 3711 18583 3737
rect 19441 3711 19447 3737
rect 19473 3711 19479 3737
rect 20785 3711 20791 3737
rect 20817 3711 20823 3737
rect 21737 3711 21743 3737
rect 21769 3711 21775 3737
rect 22521 3711 22527 3737
rect 22553 3711 22559 3737
rect 22801 3711 22807 3737
rect 22833 3711 22839 3737
rect 22913 3711 22919 3737
rect 22945 3711 22951 3737
rect 24761 3711 24767 3737
rect 24793 3711 24799 3737
rect 25209 3711 25215 3737
rect 25241 3711 25247 3737
rect 25433 3711 25439 3737
rect 25465 3711 25471 3737
rect 26273 3711 26279 3737
rect 26305 3711 26311 3737
rect 26889 3711 26895 3737
rect 26921 3711 26927 3737
rect 28071 3705 28097 3711
rect 28239 3737 28265 3743
rect 32047 3737 32073 3743
rect 29017 3711 29023 3737
rect 29049 3711 29055 3737
rect 29913 3711 29919 3737
rect 29945 3711 29951 3737
rect 30361 3711 30367 3737
rect 30393 3711 30399 3737
rect 31313 3711 31319 3737
rect 31345 3711 31351 3737
rect 28239 3705 28265 3711
rect 32047 3705 32073 3711
rect 32215 3737 32241 3743
rect 32215 3705 32241 3711
rect 32383 3737 32409 3743
rect 35687 3737 35713 3743
rect 38151 3737 38177 3743
rect 32769 3711 32775 3737
rect 32801 3711 32807 3737
rect 33889 3711 33895 3737
rect 33921 3711 33927 3737
rect 34169 3711 34175 3737
rect 34201 3711 34207 3737
rect 35065 3711 35071 3737
rect 35097 3711 35103 3737
rect 36969 3711 36975 3737
rect 37001 3711 37007 3737
rect 37641 3711 37647 3737
rect 37673 3711 37679 3737
rect 32383 3705 32409 3711
rect 35687 3705 35713 3711
rect 38151 3705 38177 3711
rect 38823 3737 38849 3743
rect 38823 3705 38849 3711
rect 38991 3737 39017 3743
rect 38991 3705 39017 3711
rect 672 3541 39312 3558
rect 672 3515 2074 3541
rect 2100 3515 2136 3541
rect 2162 3515 2198 3541
rect 2224 3515 2260 3541
rect 2286 3515 2322 3541
rect 2348 3515 2384 3541
rect 2410 3515 2446 3541
rect 2472 3515 2508 3541
rect 2534 3515 7074 3541
rect 7100 3515 7136 3541
rect 7162 3515 7198 3541
rect 7224 3515 7260 3541
rect 7286 3515 7322 3541
rect 7348 3515 7384 3541
rect 7410 3515 7446 3541
rect 7472 3515 7508 3541
rect 7534 3515 12074 3541
rect 12100 3515 12136 3541
rect 12162 3515 12198 3541
rect 12224 3515 12260 3541
rect 12286 3515 12322 3541
rect 12348 3515 12384 3541
rect 12410 3515 12446 3541
rect 12472 3515 12508 3541
rect 12534 3515 17074 3541
rect 17100 3515 17136 3541
rect 17162 3515 17198 3541
rect 17224 3515 17260 3541
rect 17286 3515 17322 3541
rect 17348 3515 17384 3541
rect 17410 3515 17446 3541
rect 17472 3515 17508 3541
rect 17534 3515 22074 3541
rect 22100 3515 22136 3541
rect 22162 3515 22198 3541
rect 22224 3515 22260 3541
rect 22286 3515 22322 3541
rect 22348 3515 22384 3541
rect 22410 3515 22446 3541
rect 22472 3515 22508 3541
rect 22534 3515 27074 3541
rect 27100 3515 27136 3541
rect 27162 3515 27198 3541
rect 27224 3515 27260 3541
rect 27286 3515 27322 3541
rect 27348 3515 27384 3541
rect 27410 3515 27446 3541
rect 27472 3515 27508 3541
rect 27534 3515 32074 3541
rect 32100 3515 32136 3541
rect 32162 3515 32198 3541
rect 32224 3515 32260 3541
rect 32286 3515 32322 3541
rect 32348 3515 32384 3541
rect 32410 3515 32446 3541
rect 32472 3515 32508 3541
rect 32534 3515 37074 3541
rect 37100 3515 37136 3541
rect 37162 3515 37198 3541
rect 37224 3515 37260 3541
rect 37286 3515 37322 3541
rect 37348 3515 37384 3541
rect 37410 3515 37446 3541
rect 37472 3515 37508 3541
rect 37534 3515 39312 3541
rect 672 3498 39312 3515
rect 26055 3345 26081 3351
rect 1801 3319 1807 3345
rect 1833 3319 1839 3345
rect 1913 3319 1919 3345
rect 1945 3319 1951 3345
rect 2473 3319 2479 3345
rect 2505 3319 2511 3345
rect 3817 3319 3823 3345
rect 3849 3319 3855 3345
rect 4377 3319 4383 3345
rect 4409 3319 4415 3345
rect 4489 3319 4495 3345
rect 4521 3319 4527 3345
rect 5273 3319 5279 3345
rect 5305 3319 5311 3345
rect 6449 3319 6455 3345
rect 6481 3319 6487 3345
rect 8073 3319 8079 3345
rect 8105 3319 8111 3345
rect 8969 3319 8975 3345
rect 9001 3319 9007 3345
rect 9529 3319 9535 3345
rect 9561 3319 9567 3345
rect 10425 3319 10431 3345
rect 10457 3319 10463 3345
rect 12049 3319 12055 3345
rect 12081 3319 12087 3345
rect 12721 3319 12727 3345
rect 12753 3319 12759 3345
rect 13337 3319 13343 3345
rect 13369 3319 13375 3345
rect 13673 3319 13679 3345
rect 13705 3319 13711 3345
rect 13897 3319 13903 3345
rect 13929 3319 13935 3345
rect 15521 3319 15527 3345
rect 15553 3319 15559 3345
rect 15969 3319 15975 3345
rect 16001 3319 16007 3345
rect 16193 3319 16199 3345
rect 16225 3319 16231 3345
rect 16977 3319 16983 3345
rect 17009 3319 17015 3345
rect 17761 3319 17767 3345
rect 17793 3319 17799 3345
rect 18769 3319 18775 3345
rect 18801 3319 18807 3345
rect 19217 3319 19223 3345
rect 19249 3319 19255 3345
rect 19441 3319 19447 3345
rect 19473 3319 19479 3345
rect 20225 3319 20231 3345
rect 20257 3319 20263 3345
rect 21009 3319 21015 3345
rect 21041 3319 21047 3345
rect 22745 3319 22751 3345
rect 22777 3319 22783 3345
rect 23193 3319 23199 3345
rect 23225 3319 23231 3345
rect 23417 3319 23423 3345
rect 23449 3319 23455 3345
rect 24369 3319 24375 3345
rect 24401 3319 24407 3345
rect 25209 3319 25215 3345
rect 25241 3319 25247 3345
rect 26055 3313 26081 3319
rect 26167 3345 26193 3351
rect 26167 3313 26193 3319
rect 26335 3345 26361 3351
rect 30199 3345 30225 3351
rect 33671 3345 33697 3351
rect 26721 3319 26727 3345
rect 26753 3319 26759 3345
rect 27169 3319 27175 3345
rect 27201 3319 27207 3345
rect 27393 3319 27399 3345
rect 27425 3319 27431 3345
rect 28457 3319 28463 3345
rect 28489 3319 28495 3345
rect 29353 3319 29359 3345
rect 29385 3319 29391 3345
rect 30697 3319 30703 3345
rect 30729 3319 30735 3345
rect 31873 3319 31879 3345
rect 31905 3319 31911 3345
rect 32153 3319 32159 3345
rect 32185 3319 32191 3345
rect 33329 3319 33335 3345
rect 33361 3319 33367 3345
rect 26335 3313 26361 3319
rect 30199 3313 30225 3319
rect 33671 3313 33697 3319
rect 33783 3345 33809 3351
rect 33783 3313 33809 3319
rect 33951 3345 33977 3351
rect 37591 3345 37617 3351
rect 34673 3319 34679 3345
rect 34705 3319 34711 3345
rect 35177 3319 35183 3345
rect 35209 3319 35215 3345
rect 35737 3319 35743 3345
rect 35769 3319 35775 3345
rect 36129 3319 36135 3345
rect 36161 3319 36167 3345
rect 36689 3319 36695 3345
rect 36721 3319 36727 3345
rect 36857 3319 36863 3345
rect 36889 3319 36895 3345
rect 33951 3313 33977 3319
rect 37591 3313 37617 3319
rect 37927 3345 37953 3351
rect 37927 3313 37953 3319
rect 38655 3345 38681 3351
rect 38655 3313 38681 3319
rect 38767 3345 38793 3351
rect 38767 3313 38793 3319
rect 38879 3345 38905 3351
rect 38879 3313 38905 3319
rect 30031 3289 30057 3295
rect 6449 3263 6455 3289
rect 6481 3263 6487 3289
rect 8969 3263 8975 3289
rect 9001 3263 9007 3289
rect 10425 3263 10431 3289
rect 10457 3263 10463 3289
rect 12721 3263 12727 3289
rect 12753 3263 12759 3289
rect 17929 3263 17935 3289
rect 17961 3263 17967 3289
rect 21177 3263 21183 3289
rect 21209 3263 21215 3289
rect 25209 3263 25215 3289
rect 25241 3263 25247 3289
rect 29353 3263 29359 3289
rect 29385 3263 29391 3289
rect 30031 3257 30057 3263
rect 30311 3289 30337 3295
rect 37703 3289 37729 3295
rect 31873 3263 31879 3289
rect 31905 3263 31911 3289
rect 33329 3263 33335 3289
rect 33361 3263 33367 3289
rect 30311 3257 30337 3263
rect 37703 3257 37729 3263
rect 672 3149 39312 3166
rect 672 3123 4574 3149
rect 4600 3123 4636 3149
rect 4662 3123 4698 3149
rect 4724 3123 4760 3149
rect 4786 3123 4822 3149
rect 4848 3123 4884 3149
rect 4910 3123 4946 3149
rect 4972 3123 5008 3149
rect 5034 3123 9574 3149
rect 9600 3123 9636 3149
rect 9662 3123 9698 3149
rect 9724 3123 9760 3149
rect 9786 3123 9822 3149
rect 9848 3123 9884 3149
rect 9910 3123 9946 3149
rect 9972 3123 10008 3149
rect 10034 3123 14574 3149
rect 14600 3123 14636 3149
rect 14662 3123 14698 3149
rect 14724 3123 14760 3149
rect 14786 3123 14822 3149
rect 14848 3123 14884 3149
rect 14910 3123 14946 3149
rect 14972 3123 15008 3149
rect 15034 3123 19574 3149
rect 19600 3123 19636 3149
rect 19662 3123 19698 3149
rect 19724 3123 19760 3149
rect 19786 3123 19822 3149
rect 19848 3123 19884 3149
rect 19910 3123 19946 3149
rect 19972 3123 20008 3149
rect 20034 3123 24574 3149
rect 24600 3123 24636 3149
rect 24662 3123 24698 3149
rect 24724 3123 24760 3149
rect 24786 3123 24822 3149
rect 24848 3123 24884 3149
rect 24910 3123 24946 3149
rect 24972 3123 25008 3149
rect 25034 3123 29574 3149
rect 29600 3123 29636 3149
rect 29662 3123 29698 3149
rect 29724 3123 29760 3149
rect 29786 3123 29822 3149
rect 29848 3123 29884 3149
rect 29910 3123 29946 3149
rect 29972 3123 30008 3149
rect 30034 3123 34574 3149
rect 34600 3123 34636 3149
rect 34662 3123 34698 3149
rect 34724 3123 34760 3149
rect 34786 3123 34822 3149
rect 34848 3123 34884 3149
rect 34910 3123 34946 3149
rect 34972 3123 35008 3149
rect 35034 3123 39312 3149
rect 672 3106 39312 3123
rect 28351 3009 28377 3015
rect 32047 3009 32073 3015
rect 35743 3009 35769 3015
rect 1913 2983 1919 3009
rect 1945 2983 1951 3009
rect 4489 2983 4495 3009
rect 4521 2983 4527 3009
rect 7009 2983 7015 3009
rect 7041 2983 7047 3009
rect 8465 2983 8471 3009
rect 8497 2983 8503 3009
rect 10761 2983 10767 3009
rect 10793 2983 10799 3009
rect 12441 2983 12447 3009
rect 12473 2983 12479 3009
rect 14233 2983 14239 3009
rect 14265 2983 14271 3009
rect 17761 2983 17767 3009
rect 17793 2983 17799 3009
rect 19217 2983 19223 3009
rect 19249 2983 19255 3009
rect 21737 2983 21743 3009
rect 21769 2983 21775 3009
rect 23417 2983 23423 3009
rect 23449 2983 23455 3009
rect 31369 2983 31375 3009
rect 31401 2983 31407 3009
rect 33889 2983 33895 3009
rect 33921 2983 33927 3009
rect 35177 2983 35183 3009
rect 35209 2983 35215 3009
rect 28351 2977 28377 2983
rect 32047 2977 32073 2983
rect 35743 2977 35769 2983
rect 35911 3009 35937 3015
rect 35911 2977 35937 2983
rect 38151 3009 38177 3015
rect 38151 2977 38177 2983
rect 38263 3009 38289 3015
rect 38263 2977 38289 2983
rect 38431 3009 38457 3015
rect 38431 2977 38457 2983
rect 38711 3009 38737 3015
rect 38711 2977 38737 2983
rect 28015 2953 28041 2959
rect 1913 2927 1919 2953
rect 1945 2927 1951 2953
rect 3033 2927 3039 2953
rect 3065 2927 3071 2953
rect 3481 2927 3487 2953
rect 3513 2927 3519 2953
rect 4489 2927 4495 2953
rect 4521 2927 4527 2953
rect 5833 2927 5839 2953
rect 5865 2927 5871 2953
rect 7009 2927 7015 2953
rect 7041 2927 7047 2953
rect 7569 2927 7575 2953
rect 7601 2927 7607 2953
rect 8465 2927 8471 2953
rect 8497 2927 8503 2953
rect 10033 2927 10039 2953
rect 10065 2927 10071 2953
rect 10761 2927 10767 2953
rect 10793 2927 10799 2953
rect 11545 2927 11551 2953
rect 11577 2927 11583 2953
rect 12441 2927 12447 2953
rect 12473 2927 12479 2953
rect 13337 2927 13343 2953
rect 13369 2927 13375 2953
rect 14233 2927 14239 2953
rect 14265 2927 14271 2953
rect 15073 2927 15079 2953
rect 15105 2927 15111 2953
rect 15241 2927 15247 2953
rect 15273 2927 15279 2953
rect 15465 2927 15471 2953
rect 15497 2927 15503 2953
rect 16809 2927 16815 2953
rect 16841 2927 16847 2953
rect 17649 2927 17655 2953
rect 17681 2927 17687 2953
rect 18265 2927 18271 2953
rect 18297 2927 18303 2953
rect 19217 2927 19223 2953
rect 19249 2927 19255 2953
rect 20785 2927 20791 2953
rect 20817 2927 20823 2953
rect 21737 2927 21743 2953
rect 21769 2927 21775 2953
rect 22241 2927 22247 2953
rect 22273 2927 22279 2953
rect 23417 2927 23423 2953
rect 23449 2927 23455 2953
rect 24761 2927 24767 2953
rect 24793 2927 24799 2953
rect 25209 2927 25215 2953
rect 25241 2927 25247 2953
rect 25433 2927 25439 2953
rect 25465 2927 25471 2953
rect 26273 2927 26279 2953
rect 26305 2927 26311 2953
rect 26777 2927 26783 2953
rect 26809 2927 26815 2953
rect 26889 2927 26895 2953
rect 26921 2927 26927 2953
rect 28015 2921 28041 2927
rect 28183 2953 28209 2959
rect 32215 2953 32241 2959
rect 29017 2927 29023 2953
rect 29049 2927 29055 2953
rect 29297 2927 29303 2953
rect 29329 2927 29335 2953
rect 29465 2927 29471 2953
rect 29497 2927 29503 2953
rect 30361 2927 30367 2953
rect 30393 2927 30399 2953
rect 31369 2927 31375 2953
rect 31401 2927 31407 2953
rect 28183 2921 28209 2927
rect 32215 2921 32241 2927
rect 32383 2953 32409 2959
rect 35687 2953 35713 2959
rect 38823 2953 38849 2959
rect 32769 2927 32775 2953
rect 32801 2927 32807 2953
rect 33889 2927 33895 2953
rect 33921 2927 33927 2953
rect 34449 2927 34455 2953
rect 34481 2927 34487 2953
rect 35177 2927 35183 2953
rect 35209 2927 35215 2953
rect 36689 2927 36695 2953
rect 36721 2927 36727 2953
rect 37137 2927 37143 2953
rect 37169 2927 37175 2953
rect 37361 2927 37367 2953
rect 37393 2927 37399 2953
rect 32383 2921 32409 2927
rect 35687 2921 35713 2927
rect 38823 2921 38849 2927
rect 38935 2953 38961 2959
rect 38935 2921 38961 2927
rect 672 2757 39312 2774
rect 672 2731 2074 2757
rect 2100 2731 2136 2757
rect 2162 2731 2198 2757
rect 2224 2731 2260 2757
rect 2286 2731 2322 2757
rect 2348 2731 2384 2757
rect 2410 2731 2446 2757
rect 2472 2731 2508 2757
rect 2534 2731 7074 2757
rect 7100 2731 7136 2757
rect 7162 2731 7198 2757
rect 7224 2731 7260 2757
rect 7286 2731 7322 2757
rect 7348 2731 7384 2757
rect 7410 2731 7446 2757
rect 7472 2731 7508 2757
rect 7534 2731 12074 2757
rect 12100 2731 12136 2757
rect 12162 2731 12198 2757
rect 12224 2731 12260 2757
rect 12286 2731 12322 2757
rect 12348 2731 12384 2757
rect 12410 2731 12446 2757
rect 12472 2731 12508 2757
rect 12534 2731 17074 2757
rect 17100 2731 17136 2757
rect 17162 2731 17198 2757
rect 17224 2731 17260 2757
rect 17286 2731 17322 2757
rect 17348 2731 17384 2757
rect 17410 2731 17446 2757
rect 17472 2731 17508 2757
rect 17534 2731 22074 2757
rect 22100 2731 22136 2757
rect 22162 2731 22198 2757
rect 22224 2731 22260 2757
rect 22286 2731 22322 2757
rect 22348 2731 22384 2757
rect 22410 2731 22446 2757
rect 22472 2731 22508 2757
rect 22534 2731 27074 2757
rect 27100 2731 27136 2757
rect 27162 2731 27198 2757
rect 27224 2731 27260 2757
rect 27286 2731 27322 2757
rect 27348 2731 27384 2757
rect 27410 2731 27446 2757
rect 27472 2731 27508 2757
rect 27534 2731 32074 2757
rect 32100 2731 32136 2757
rect 32162 2731 32198 2757
rect 32224 2731 32260 2757
rect 32286 2731 32322 2757
rect 32348 2731 32384 2757
rect 32410 2731 32446 2757
rect 32472 2731 32508 2757
rect 32534 2731 37074 2757
rect 37100 2731 37136 2757
rect 37162 2731 37198 2757
rect 37224 2731 37260 2757
rect 37286 2731 37322 2757
rect 37348 2731 37384 2757
rect 37410 2731 37446 2757
rect 37472 2731 37508 2757
rect 37534 2731 39312 2757
rect 672 2714 39312 2731
rect 30031 2561 30057 2567
rect 1801 2535 1807 2561
rect 1833 2535 1839 2561
rect 2025 2535 2031 2561
rect 2057 2535 2063 2561
rect 2473 2535 2479 2561
rect 2505 2535 2511 2561
rect 3817 2535 3823 2561
rect 3849 2535 3855 2561
rect 4993 2535 4999 2561
rect 5025 2535 5031 2561
rect 5273 2535 5279 2561
rect 5305 2535 5311 2561
rect 6449 2535 6455 2561
rect 6481 2535 6487 2561
rect 7793 2535 7799 2561
rect 7825 2535 7831 2561
rect 8969 2535 8975 2561
rect 9001 2535 9007 2561
rect 9529 2535 9535 2561
rect 9561 2535 9567 2561
rect 10257 2535 10263 2561
rect 10289 2535 10295 2561
rect 11881 2535 11887 2561
rect 11913 2535 11919 2561
rect 12721 2535 12727 2561
rect 12753 2535 12759 2561
rect 13337 2535 13343 2561
rect 13369 2535 13375 2561
rect 14233 2535 14239 2561
rect 14265 2535 14271 2561
rect 15241 2535 15247 2561
rect 15273 2535 15279 2561
rect 15689 2535 15695 2561
rect 15721 2535 15727 2561
rect 15913 2535 15919 2561
rect 15945 2535 15951 2561
rect 16809 2535 16815 2561
rect 16841 2535 16847 2561
rect 17145 2535 17151 2561
rect 17177 2535 17183 2561
rect 17369 2535 17375 2561
rect 17401 2535 17407 2561
rect 20113 2535 20119 2561
rect 20145 2535 20151 2561
rect 20953 2535 20959 2561
rect 20985 2535 20991 2561
rect 22745 2535 22751 2561
rect 22777 2535 22783 2561
rect 23193 2535 23199 2561
rect 23225 2535 23231 2561
rect 23529 2535 23535 2561
rect 23561 2535 23567 2561
rect 24369 2535 24375 2561
rect 24401 2535 24407 2561
rect 24649 2535 24655 2561
rect 24681 2535 24687 2561
rect 24873 2535 24879 2561
rect 24905 2535 24911 2561
rect 26721 2535 26727 2561
rect 26753 2535 26759 2561
rect 27169 2535 27175 2561
rect 27201 2535 27207 2561
rect 27393 2535 27399 2561
rect 27425 2535 27431 2561
rect 28457 2535 28463 2561
rect 28489 2535 28495 2561
rect 29353 2535 29359 2561
rect 29385 2535 29391 2561
rect 30031 2529 30057 2535
rect 30199 2561 30225 2567
rect 33671 2561 33697 2567
rect 30697 2535 30703 2561
rect 30729 2535 30735 2561
rect 31257 2535 31263 2561
rect 31289 2535 31295 2561
rect 31369 2535 31375 2561
rect 31401 2535 31407 2561
rect 32433 2535 32439 2561
rect 32465 2535 32471 2561
rect 33329 2535 33335 2561
rect 33361 2535 33367 2561
rect 30199 2529 30225 2535
rect 33671 2529 33697 2535
rect 33783 2561 33809 2567
rect 33783 2529 33809 2535
rect 33895 2561 33921 2567
rect 37591 2561 37617 2567
rect 34673 2535 34679 2561
rect 34705 2535 34711 2561
rect 35177 2535 35183 2561
rect 35209 2535 35215 2561
rect 35345 2535 35351 2561
rect 35377 2535 35383 2561
rect 36129 2535 36135 2561
rect 36161 2535 36167 2561
rect 36689 2535 36695 2561
rect 36721 2535 36727 2561
rect 36857 2535 36863 2561
rect 36889 2535 36895 2561
rect 33895 2529 33921 2535
rect 37591 2529 37617 2535
rect 37703 2561 37729 2567
rect 37703 2529 37729 2535
rect 37871 2561 37897 2567
rect 37871 2529 37897 2535
rect 38767 2561 38793 2567
rect 38767 2529 38793 2535
rect 38879 2561 38905 2567
rect 38879 2529 38905 2535
rect 26055 2505 26081 2511
rect 4993 2479 4999 2505
rect 5025 2479 5031 2505
rect 6449 2479 6455 2505
rect 6481 2479 6487 2505
rect 8969 2479 8975 2505
rect 9001 2479 9007 2505
rect 10257 2479 10263 2505
rect 10289 2479 10295 2505
rect 12721 2479 12727 2505
rect 12753 2479 12759 2505
rect 14233 2479 14239 2505
rect 14265 2479 14271 2505
rect 20953 2479 20959 2505
rect 20985 2479 20991 2505
rect 26055 2473 26081 2479
rect 26223 2505 26249 2511
rect 26223 2473 26249 2479
rect 26335 2505 26361 2511
rect 30311 2505 30337 2511
rect 38655 2505 38681 2511
rect 29353 2479 29359 2505
rect 29385 2479 29391 2505
rect 33329 2479 33335 2505
rect 33361 2479 33367 2505
rect 26335 2473 26361 2479
rect 30311 2473 30337 2479
rect 38655 2473 38681 2479
rect 672 2365 39312 2382
rect 672 2339 4574 2365
rect 4600 2339 4636 2365
rect 4662 2339 4698 2365
rect 4724 2339 4760 2365
rect 4786 2339 4822 2365
rect 4848 2339 4884 2365
rect 4910 2339 4946 2365
rect 4972 2339 5008 2365
rect 5034 2339 9574 2365
rect 9600 2339 9636 2365
rect 9662 2339 9698 2365
rect 9724 2339 9760 2365
rect 9786 2339 9822 2365
rect 9848 2339 9884 2365
rect 9910 2339 9946 2365
rect 9972 2339 10008 2365
rect 10034 2339 14574 2365
rect 14600 2339 14636 2365
rect 14662 2339 14698 2365
rect 14724 2339 14760 2365
rect 14786 2339 14822 2365
rect 14848 2339 14884 2365
rect 14910 2339 14946 2365
rect 14972 2339 15008 2365
rect 15034 2339 19574 2365
rect 19600 2339 19636 2365
rect 19662 2339 19698 2365
rect 19724 2339 19760 2365
rect 19786 2339 19822 2365
rect 19848 2339 19884 2365
rect 19910 2339 19946 2365
rect 19972 2339 20008 2365
rect 20034 2339 24574 2365
rect 24600 2339 24636 2365
rect 24662 2339 24698 2365
rect 24724 2339 24760 2365
rect 24786 2339 24822 2365
rect 24848 2339 24884 2365
rect 24910 2339 24946 2365
rect 24972 2339 25008 2365
rect 25034 2339 29574 2365
rect 29600 2339 29636 2365
rect 29662 2339 29698 2365
rect 29724 2339 29760 2365
rect 29786 2339 29822 2365
rect 29848 2339 29884 2365
rect 29910 2339 29946 2365
rect 29972 2339 30008 2365
rect 30034 2339 34574 2365
rect 34600 2339 34636 2365
rect 34662 2339 34698 2365
rect 34724 2339 34760 2365
rect 34786 2339 34822 2365
rect 34848 2339 34884 2365
rect 34910 2339 34946 2365
rect 34972 2339 35008 2365
rect 35034 2339 39312 2365
rect 672 2322 39312 2339
rect 24095 2225 24121 2231
rect 4433 2199 4439 2225
rect 4465 2199 4471 2225
rect 8465 2199 8471 2225
rect 8497 2199 8503 2225
rect 10761 2199 10767 2225
rect 10793 2199 10799 2225
rect 12441 2199 12447 2225
rect 12473 2199 12479 2225
rect 17761 2199 17767 2225
rect 17793 2199 17799 2225
rect 19217 2199 19223 2225
rect 19249 2199 19255 2225
rect 21737 2199 21743 2225
rect 21769 2199 21775 2225
rect 23193 2199 23199 2225
rect 23225 2199 23231 2225
rect 24095 2193 24121 2199
rect 24375 2225 24401 2231
rect 24375 2193 24401 2199
rect 28071 2225 28097 2231
rect 28071 2193 28097 2199
rect 28239 2225 28265 2231
rect 31935 2225 31961 2231
rect 35911 2225 35937 2231
rect 31257 2199 31263 2225
rect 31289 2199 31295 2225
rect 35177 2199 35183 2225
rect 35209 2199 35215 2225
rect 28239 2193 28265 2199
rect 31935 2193 31961 2199
rect 35911 2193 35937 2199
rect 38711 2225 38737 2231
rect 38711 2193 38737 2199
rect 38879 2225 38905 2231
rect 38879 2193 38905 2199
rect 38991 2225 39017 2231
rect 38991 2193 39017 2199
rect 24207 2169 24233 2175
rect 28295 2169 28321 2175
rect 31655 2169 31681 2175
rect 2361 2143 2367 2169
rect 2393 2143 2399 2169
rect 2473 2143 2479 2169
rect 2505 2143 2511 2169
rect 3033 2143 3039 2169
rect 3065 2143 3071 2169
rect 3481 2143 3487 2169
rect 3513 2143 3519 2169
rect 4433 2143 4439 2169
rect 4465 2143 4471 2169
rect 5889 2143 5895 2169
rect 5921 2143 5927 2169
rect 6393 2143 6399 2169
rect 6425 2143 6431 2169
rect 6505 2143 6511 2169
rect 6537 2143 6543 2169
rect 7289 2143 7295 2169
rect 7321 2143 7327 2169
rect 8465 2143 8471 2169
rect 8497 2143 8503 2169
rect 10033 2143 10039 2169
rect 10065 2143 10071 2169
rect 10761 2143 10767 2169
rect 10793 2143 10799 2169
rect 11545 2143 11551 2169
rect 11577 2143 11583 2169
rect 12441 2143 12447 2169
rect 12473 2143 12479 2169
rect 13617 2143 13623 2169
rect 13649 2143 13655 2169
rect 14065 2143 14071 2169
rect 14097 2143 14103 2169
rect 14289 2143 14295 2169
rect 14321 2143 14327 2169
rect 15129 2143 15135 2169
rect 15161 2143 15167 2169
rect 15577 2143 15583 2169
rect 15609 2143 15615 2169
rect 15801 2143 15807 2169
rect 15833 2143 15839 2169
rect 16809 2143 16815 2169
rect 16841 2143 16847 2169
rect 17649 2143 17655 2169
rect 17681 2143 17687 2169
rect 18265 2143 18271 2169
rect 18297 2143 18303 2169
rect 19105 2143 19111 2169
rect 19137 2143 19143 2169
rect 20785 2143 20791 2169
rect 20817 2143 20823 2169
rect 21737 2143 21743 2169
rect 21769 2143 21775 2169
rect 22521 2143 22527 2169
rect 22553 2143 22559 2169
rect 23137 2143 23143 2169
rect 23169 2143 23175 2169
rect 24761 2143 24767 2169
rect 24793 2143 24799 2169
rect 25209 2143 25215 2169
rect 25241 2143 25247 2169
rect 25433 2143 25439 2169
rect 25465 2143 25471 2169
rect 26217 2143 26223 2169
rect 26249 2143 26255 2169
rect 26777 2143 26783 2169
rect 26809 2143 26815 2169
rect 26889 2143 26895 2169
rect 26921 2143 26927 2169
rect 29017 2143 29023 2169
rect 29049 2143 29055 2169
rect 29185 2143 29191 2169
rect 29217 2143 29223 2169
rect 29409 2143 29415 2169
rect 29441 2143 29447 2169
rect 30361 2143 30367 2169
rect 30393 2143 30399 2169
rect 31257 2143 31263 2169
rect 31289 2143 31295 2169
rect 24207 2137 24233 2143
rect 28295 2137 28321 2143
rect 31655 2137 31681 2143
rect 31823 2169 31849 2175
rect 35687 2169 35713 2175
rect 32713 2143 32719 2169
rect 32745 2143 32751 2169
rect 33273 2143 33279 2169
rect 33305 2143 33311 2169
rect 33441 2143 33447 2169
rect 33473 2143 33479 2169
rect 34393 2143 34399 2169
rect 34425 2143 34431 2169
rect 35177 2143 35183 2169
rect 35209 2143 35215 2169
rect 31823 2137 31849 2143
rect 35687 2137 35713 2143
rect 35799 2169 35825 2175
rect 38151 2169 38177 2175
rect 37193 2143 37199 2169
rect 37225 2143 37231 2169
rect 37305 2143 37311 2169
rect 37337 2143 37343 2169
rect 37585 2143 37591 2169
rect 37617 2143 37623 2169
rect 35799 2137 35825 2143
rect 38151 2137 38177 2143
rect 38319 2169 38345 2175
rect 38319 2137 38345 2143
rect 38487 2169 38513 2175
rect 38487 2137 38513 2143
rect 672 1973 39312 1990
rect 672 1947 2074 1973
rect 2100 1947 2136 1973
rect 2162 1947 2198 1973
rect 2224 1947 2260 1973
rect 2286 1947 2322 1973
rect 2348 1947 2384 1973
rect 2410 1947 2446 1973
rect 2472 1947 2508 1973
rect 2534 1947 7074 1973
rect 7100 1947 7136 1973
rect 7162 1947 7198 1973
rect 7224 1947 7260 1973
rect 7286 1947 7322 1973
rect 7348 1947 7384 1973
rect 7410 1947 7446 1973
rect 7472 1947 7508 1973
rect 7534 1947 12074 1973
rect 12100 1947 12136 1973
rect 12162 1947 12198 1973
rect 12224 1947 12260 1973
rect 12286 1947 12322 1973
rect 12348 1947 12384 1973
rect 12410 1947 12446 1973
rect 12472 1947 12508 1973
rect 12534 1947 17074 1973
rect 17100 1947 17136 1973
rect 17162 1947 17198 1973
rect 17224 1947 17260 1973
rect 17286 1947 17322 1973
rect 17348 1947 17384 1973
rect 17410 1947 17446 1973
rect 17472 1947 17508 1973
rect 17534 1947 22074 1973
rect 22100 1947 22136 1973
rect 22162 1947 22198 1973
rect 22224 1947 22260 1973
rect 22286 1947 22322 1973
rect 22348 1947 22384 1973
rect 22410 1947 22446 1973
rect 22472 1947 22508 1973
rect 22534 1947 27074 1973
rect 27100 1947 27136 1973
rect 27162 1947 27198 1973
rect 27224 1947 27260 1973
rect 27286 1947 27322 1973
rect 27348 1947 27384 1973
rect 27410 1947 27446 1973
rect 27472 1947 27508 1973
rect 27534 1947 32074 1973
rect 32100 1947 32136 1973
rect 32162 1947 32198 1973
rect 32224 1947 32260 1973
rect 32286 1947 32322 1973
rect 32348 1947 32384 1973
rect 32410 1947 32446 1973
rect 32472 1947 32508 1973
rect 32534 1947 37074 1973
rect 37100 1947 37136 1973
rect 37162 1947 37198 1973
rect 37224 1947 37260 1973
rect 37286 1947 37322 1973
rect 37348 1947 37384 1973
rect 37410 1947 37446 1973
rect 37472 1947 37508 1973
rect 37534 1947 39312 1973
rect 672 1930 39312 1947
rect 38151 1777 38177 1783
rect 1633 1751 1639 1777
rect 1665 1751 1671 1777
rect 2473 1751 2479 1777
rect 2505 1751 2511 1777
rect 3481 1751 3487 1777
rect 3513 1751 3519 1777
rect 4433 1751 4439 1777
rect 4465 1751 4471 1777
rect 5497 1751 5503 1777
rect 5529 1751 5535 1777
rect 6393 1751 6399 1777
rect 6425 1751 6431 1777
rect 7457 1751 7463 1777
rect 7489 1751 7495 1777
rect 8129 1751 8135 1777
rect 8161 1751 8167 1777
rect 9417 1751 9423 1777
rect 9449 1751 9455 1777
rect 10257 1751 10263 1777
rect 10289 1751 10295 1777
rect 11377 1751 11383 1777
rect 11409 1751 11415 1777
rect 11993 1751 11999 1777
rect 12025 1751 12031 1777
rect 13337 1751 13343 1777
rect 13369 1751 13375 1777
rect 13505 1751 13511 1777
rect 13537 1751 13543 1777
rect 13729 1751 13735 1777
rect 13761 1751 13767 1777
rect 15129 1751 15135 1777
rect 15161 1751 15167 1777
rect 15297 1751 15303 1777
rect 15329 1751 15335 1777
rect 15521 1751 15527 1777
rect 15553 1751 15559 1777
rect 16585 1751 16591 1777
rect 16617 1751 16623 1777
rect 17537 1751 17543 1777
rect 17569 1751 17575 1777
rect 18545 1751 18551 1777
rect 18577 1751 18583 1777
rect 19105 1751 19111 1777
rect 19137 1751 19143 1777
rect 19217 1751 19223 1777
rect 19249 1751 19255 1777
rect 21177 1751 21183 1777
rect 21209 1751 21215 1777
rect 21793 1751 21799 1777
rect 21825 1751 21831 1777
rect 22465 1751 22471 1777
rect 22497 1751 22503 1777
rect 22913 1751 22919 1777
rect 22945 1751 22951 1777
rect 23137 1751 23143 1777
rect 23169 1751 23175 1777
rect 24481 1751 24487 1777
rect 24513 1751 24519 1777
rect 25209 1751 25215 1777
rect 25241 1751 25247 1777
rect 26385 1751 26391 1777
rect 26417 1751 26423 1777
rect 26889 1751 26895 1777
rect 26921 1751 26927 1777
rect 27057 1751 27063 1777
rect 27089 1751 27095 1777
rect 28625 1751 28631 1777
rect 28657 1751 28663 1777
rect 28793 1751 28799 1777
rect 28825 1751 28831 1777
rect 29017 1751 29023 1777
rect 29049 1751 29055 1777
rect 30361 1751 30367 1777
rect 30393 1751 30399 1777
rect 31257 1751 31263 1777
rect 31289 1751 31295 1777
rect 32545 1751 32551 1777
rect 32577 1751 32583 1777
rect 33441 1751 33447 1777
rect 33473 1751 33479 1777
rect 34393 1751 34399 1777
rect 34425 1751 34431 1777
rect 35177 1751 35183 1777
rect 35209 1751 35215 1777
rect 36185 1751 36191 1777
rect 36217 1751 36223 1777
rect 37137 1751 37143 1777
rect 37169 1751 37175 1777
rect 38151 1745 38177 1751
rect 38263 1777 38289 1783
rect 38263 1745 38289 1751
rect 38431 1777 38457 1783
rect 38431 1745 38457 1751
rect 38655 1777 38681 1783
rect 38655 1745 38681 1751
rect 38823 1777 38849 1783
rect 38823 1745 38849 1751
rect 38935 1777 38961 1783
rect 38935 1745 38961 1751
rect 1521 1695 1527 1721
rect 1553 1695 1559 1721
rect 4433 1695 4439 1721
rect 4465 1695 4471 1721
rect 6393 1695 6399 1721
rect 6425 1695 6431 1721
rect 8129 1695 8135 1721
rect 8161 1695 8167 1721
rect 10257 1695 10263 1721
rect 10289 1695 10295 1721
rect 12049 1695 12055 1721
rect 12081 1695 12087 1721
rect 17537 1695 17543 1721
rect 17569 1695 17575 1721
rect 21849 1695 21855 1721
rect 21881 1695 21887 1721
rect 25377 1695 25383 1721
rect 25409 1695 25415 1721
rect 31257 1695 31263 1721
rect 31289 1695 31295 1721
rect 33441 1695 33447 1721
rect 33473 1695 33479 1721
rect 35177 1695 35183 1721
rect 35209 1695 35215 1721
rect 37137 1695 37143 1721
rect 37169 1695 37175 1721
rect 672 1581 39312 1598
rect 672 1555 4574 1581
rect 4600 1555 4636 1581
rect 4662 1555 4698 1581
rect 4724 1555 4760 1581
rect 4786 1555 4822 1581
rect 4848 1555 4884 1581
rect 4910 1555 4946 1581
rect 4972 1555 5008 1581
rect 5034 1555 9574 1581
rect 9600 1555 9636 1581
rect 9662 1555 9698 1581
rect 9724 1555 9760 1581
rect 9786 1555 9822 1581
rect 9848 1555 9884 1581
rect 9910 1555 9946 1581
rect 9972 1555 10008 1581
rect 10034 1555 14574 1581
rect 14600 1555 14636 1581
rect 14662 1555 14698 1581
rect 14724 1555 14760 1581
rect 14786 1555 14822 1581
rect 14848 1555 14884 1581
rect 14910 1555 14946 1581
rect 14972 1555 15008 1581
rect 15034 1555 19574 1581
rect 19600 1555 19636 1581
rect 19662 1555 19698 1581
rect 19724 1555 19760 1581
rect 19786 1555 19822 1581
rect 19848 1555 19884 1581
rect 19910 1555 19946 1581
rect 19972 1555 20008 1581
rect 20034 1555 24574 1581
rect 24600 1555 24636 1581
rect 24662 1555 24698 1581
rect 24724 1555 24760 1581
rect 24786 1555 24822 1581
rect 24848 1555 24884 1581
rect 24910 1555 24946 1581
rect 24972 1555 25008 1581
rect 25034 1555 29574 1581
rect 29600 1555 29636 1581
rect 29662 1555 29698 1581
rect 29724 1555 29760 1581
rect 29786 1555 29822 1581
rect 29848 1555 29884 1581
rect 29910 1555 29946 1581
rect 29972 1555 30008 1581
rect 30034 1555 34574 1581
rect 34600 1555 34636 1581
rect 34662 1555 34698 1581
rect 34724 1555 34760 1581
rect 34786 1555 34822 1581
rect 34848 1555 34884 1581
rect 34910 1555 34946 1581
rect 34972 1555 35008 1581
rect 35034 1555 39312 1581
rect 672 1538 39312 1555
<< via1 >>
rect 2074 18411 2100 18437
rect 2136 18411 2162 18437
rect 2198 18411 2224 18437
rect 2260 18411 2286 18437
rect 2322 18411 2348 18437
rect 2384 18411 2410 18437
rect 2446 18411 2472 18437
rect 2508 18411 2534 18437
rect 7074 18411 7100 18437
rect 7136 18411 7162 18437
rect 7198 18411 7224 18437
rect 7260 18411 7286 18437
rect 7322 18411 7348 18437
rect 7384 18411 7410 18437
rect 7446 18411 7472 18437
rect 7508 18411 7534 18437
rect 12074 18411 12100 18437
rect 12136 18411 12162 18437
rect 12198 18411 12224 18437
rect 12260 18411 12286 18437
rect 12322 18411 12348 18437
rect 12384 18411 12410 18437
rect 12446 18411 12472 18437
rect 12508 18411 12534 18437
rect 17074 18411 17100 18437
rect 17136 18411 17162 18437
rect 17198 18411 17224 18437
rect 17260 18411 17286 18437
rect 17322 18411 17348 18437
rect 17384 18411 17410 18437
rect 17446 18411 17472 18437
rect 17508 18411 17534 18437
rect 22074 18411 22100 18437
rect 22136 18411 22162 18437
rect 22198 18411 22224 18437
rect 22260 18411 22286 18437
rect 22322 18411 22348 18437
rect 22384 18411 22410 18437
rect 22446 18411 22472 18437
rect 22508 18411 22534 18437
rect 27074 18411 27100 18437
rect 27136 18411 27162 18437
rect 27198 18411 27224 18437
rect 27260 18411 27286 18437
rect 27322 18411 27348 18437
rect 27384 18411 27410 18437
rect 27446 18411 27472 18437
rect 27508 18411 27534 18437
rect 32074 18411 32100 18437
rect 32136 18411 32162 18437
rect 32198 18411 32224 18437
rect 32260 18411 32286 18437
rect 32322 18411 32348 18437
rect 32384 18411 32410 18437
rect 32446 18411 32472 18437
rect 32508 18411 32534 18437
rect 37074 18411 37100 18437
rect 37136 18411 37162 18437
rect 37198 18411 37224 18437
rect 37260 18411 37286 18437
rect 37322 18411 37348 18437
rect 37384 18411 37410 18437
rect 37446 18411 37472 18437
rect 37508 18411 37534 18437
rect 11103 18215 11129 18241
rect 11831 18215 11857 18241
rect 13343 18215 13369 18241
rect 14239 18215 14265 18241
rect 14631 18215 14657 18241
rect 15807 18215 15833 18241
rect 12055 18159 12081 18185
rect 14239 18159 14265 18185
rect 15807 18159 15833 18185
rect 4574 18019 4600 18045
rect 4636 18019 4662 18045
rect 4698 18019 4724 18045
rect 4760 18019 4786 18045
rect 4822 18019 4848 18045
rect 4884 18019 4910 18045
rect 4946 18019 4972 18045
rect 5008 18019 5034 18045
rect 9574 18019 9600 18045
rect 9636 18019 9662 18045
rect 9698 18019 9724 18045
rect 9760 18019 9786 18045
rect 9822 18019 9848 18045
rect 9884 18019 9910 18045
rect 9946 18019 9972 18045
rect 10008 18019 10034 18045
rect 14574 18019 14600 18045
rect 14636 18019 14662 18045
rect 14698 18019 14724 18045
rect 14760 18019 14786 18045
rect 14822 18019 14848 18045
rect 14884 18019 14910 18045
rect 14946 18019 14972 18045
rect 15008 18019 15034 18045
rect 19574 18019 19600 18045
rect 19636 18019 19662 18045
rect 19698 18019 19724 18045
rect 19760 18019 19786 18045
rect 19822 18019 19848 18045
rect 19884 18019 19910 18045
rect 19946 18019 19972 18045
rect 20008 18019 20034 18045
rect 24574 18019 24600 18045
rect 24636 18019 24662 18045
rect 24698 18019 24724 18045
rect 24760 18019 24786 18045
rect 24822 18019 24848 18045
rect 24884 18019 24910 18045
rect 24946 18019 24972 18045
rect 25008 18019 25034 18045
rect 29574 18019 29600 18045
rect 29636 18019 29662 18045
rect 29698 18019 29724 18045
rect 29760 18019 29786 18045
rect 29822 18019 29848 18045
rect 29884 18019 29910 18045
rect 29946 18019 29972 18045
rect 30008 18019 30034 18045
rect 34574 18019 34600 18045
rect 34636 18019 34662 18045
rect 34698 18019 34724 18045
rect 34760 18019 34786 18045
rect 34822 18019 34848 18045
rect 34884 18019 34910 18045
rect 34946 18019 34972 18045
rect 35008 18019 35034 18045
rect 14575 17879 14601 17905
rect 15919 17879 15945 17905
rect 9815 17823 9841 17849
rect 10263 17823 10289 17849
rect 10487 17823 10513 17849
rect 11271 17823 11297 17849
rect 11831 17823 11857 17849
rect 11943 17823 11969 17849
rect 13399 17823 13425 17849
rect 14575 17823 14601 17849
rect 15079 17823 15105 17849
rect 15919 17823 15945 17849
rect 2074 17627 2100 17653
rect 2136 17627 2162 17653
rect 2198 17627 2224 17653
rect 2260 17627 2286 17653
rect 2322 17627 2348 17653
rect 2384 17627 2410 17653
rect 2446 17627 2472 17653
rect 2508 17627 2534 17653
rect 7074 17627 7100 17653
rect 7136 17627 7162 17653
rect 7198 17627 7224 17653
rect 7260 17627 7286 17653
rect 7322 17627 7348 17653
rect 7384 17627 7410 17653
rect 7446 17627 7472 17653
rect 7508 17627 7534 17653
rect 12074 17627 12100 17653
rect 12136 17627 12162 17653
rect 12198 17627 12224 17653
rect 12260 17627 12286 17653
rect 12322 17627 12348 17653
rect 12384 17627 12410 17653
rect 12446 17627 12472 17653
rect 12508 17627 12534 17653
rect 17074 17627 17100 17653
rect 17136 17627 17162 17653
rect 17198 17627 17224 17653
rect 17260 17627 17286 17653
rect 17322 17627 17348 17653
rect 17384 17627 17410 17653
rect 17446 17627 17472 17653
rect 17508 17627 17534 17653
rect 22074 17627 22100 17653
rect 22136 17627 22162 17653
rect 22198 17627 22224 17653
rect 22260 17627 22286 17653
rect 22322 17627 22348 17653
rect 22384 17627 22410 17653
rect 22446 17627 22472 17653
rect 22508 17627 22534 17653
rect 27074 17627 27100 17653
rect 27136 17627 27162 17653
rect 27198 17627 27224 17653
rect 27260 17627 27286 17653
rect 27322 17627 27348 17653
rect 27384 17627 27410 17653
rect 27446 17627 27472 17653
rect 27508 17627 27534 17653
rect 32074 17627 32100 17653
rect 32136 17627 32162 17653
rect 32198 17627 32224 17653
rect 32260 17627 32286 17653
rect 32322 17627 32348 17653
rect 32384 17627 32410 17653
rect 32446 17627 32472 17653
rect 32508 17627 32534 17653
rect 37074 17627 37100 17653
rect 37136 17627 37162 17653
rect 37198 17627 37224 17653
rect 37260 17627 37286 17653
rect 37322 17627 37348 17653
rect 37384 17627 37410 17653
rect 37446 17627 37472 17653
rect 37508 17627 37534 17653
rect 9255 17431 9281 17457
rect 10375 17431 10401 17457
rect 11775 17431 11801 17457
rect 12223 17431 12249 17457
rect 12447 17431 12473 17457
rect 13287 17431 13313 17457
rect 14239 17431 14265 17457
rect 15079 17431 15105 17457
rect 15975 17431 16001 17457
rect 16255 17431 16281 17457
rect 16759 17431 16785 17457
rect 16927 17431 16953 17457
rect 10375 17375 10401 17401
rect 14239 17375 14265 17401
rect 15975 17375 16001 17401
rect 4574 17235 4600 17261
rect 4636 17235 4662 17261
rect 4698 17235 4724 17261
rect 4760 17235 4786 17261
rect 4822 17235 4848 17261
rect 4884 17235 4910 17261
rect 4946 17235 4972 17261
rect 5008 17235 5034 17261
rect 9574 17235 9600 17261
rect 9636 17235 9662 17261
rect 9698 17235 9724 17261
rect 9760 17235 9786 17261
rect 9822 17235 9848 17261
rect 9884 17235 9910 17261
rect 9946 17235 9972 17261
rect 10008 17235 10034 17261
rect 14574 17235 14600 17261
rect 14636 17235 14662 17261
rect 14698 17235 14724 17261
rect 14760 17235 14786 17261
rect 14822 17235 14848 17261
rect 14884 17235 14910 17261
rect 14946 17235 14972 17261
rect 15008 17235 15034 17261
rect 19574 17235 19600 17261
rect 19636 17235 19662 17261
rect 19698 17235 19724 17261
rect 19760 17235 19786 17261
rect 19822 17235 19848 17261
rect 19884 17235 19910 17261
rect 19946 17235 19972 17261
rect 20008 17235 20034 17261
rect 24574 17235 24600 17261
rect 24636 17235 24662 17261
rect 24698 17235 24724 17261
rect 24760 17235 24786 17261
rect 24822 17235 24848 17261
rect 24884 17235 24910 17261
rect 24946 17235 24972 17261
rect 25008 17235 25034 17261
rect 29574 17235 29600 17261
rect 29636 17235 29662 17261
rect 29698 17235 29724 17261
rect 29760 17235 29786 17261
rect 29822 17235 29848 17261
rect 29884 17235 29910 17261
rect 29946 17235 29972 17261
rect 30008 17235 30034 17261
rect 34574 17235 34600 17261
rect 34636 17235 34662 17261
rect 34698 17235 34724 17261
rect 34760 17235 34786 17261
rect 34822 17235 34848 17261
rect 34884 17235 34910 17261
rect 34946 17235 34972 17261
rect 35008 17235 35034 17261
rect 16143 17095 16169 17121
rect 17879 17095 17905 17121
rect 10095 17039 10121 17065
rect 10375 17039 10401 17065
rect 10487 17039 10513 17065
rect 11271 17039 11297 17065
rect 11831 17039 11857 17065
rect 11943 17039 11969 17065
rect 13735 17039 13761 17065
rect 14295 17039 14321 17065
rect 14463 17039 14489 17065
rect 15191 17039 15217 17065
rect 15975 17039 16001 17065
rect 16815 17039 16841 17065
rect 17879 17039 17905 17065
rect 2074 16843 2100 16869
rect 2136 16843 2162 16869
rect 2198 16843 2224 16869
rect 2260 16843 2286 16869
rect 2322 16843 2348 16869
rect 2384 16843 2410 16869
rect 2446 16843 2472 16869
rect 2508 16843 2534 16869
rect 7074 16843 7100 16869
rect 7136 16843 7162 16869
rect 7198 16843 7224 16869
rect 7260 16843 7286 16869
rect 7322 16843 7348 16869
rect 7384 16843 7410 16869
rect 7446 16843 7472 16869
rect 7508 16843 7534 16869
rect 12074 16843 12100 16869
rect 12136 16843 12162 16869
rect 12198 16843 12224 16869
rect 12260 16843 12286 16869
rect 12322 16843 12348 16869
rect 12384 16843 12410 16869
rect 12446 16843 12472 16869
rect 12508 16843 12534 16869
rect 17074 16843 17100 16869
rect 17136 16843 17162 16869
rect 17198 16843 17224 16869
rect 17260 16843 17286 16869
rect 17322 16843 17348 16869
rect 17384 16843 17410 16869
rect 17446 16843 17472 16869
rect 17508 16843 17534 16869
rect 22074 16843 22100 16869
rect 22136 16843 22162 16869
rect 22198 16843 22224 16869
rect 22260 16843 22286 16869
rect 22322 16843 22348 16869
rect 22384 16843 22410 16869
rect 22446 16843 22472 16869
rect 22508 16843 22534 16869
rect 27074 16843 27100 16869
rect 27136 16843 27162 16869
rect 27198 16843 27224 16869
rect 27260 16843 27286 16869
rect 27322 16843 27348 16869
rect 27384 16843 27410 16869
rect 27446 16843 27472 16869
rect 27508 16843 27534 16869
rect 32074 16843 32100 16869
rect 32136 16843 32162 16869
rect 32198 16843 32224 16869
rect 32260 16843 32286 16869
rect 32322 16843 32348 16869
rect 32384 16843 32410 16869
rect 32446 16843 32472 16869
rect 32508 16843 32534 16869
rect 37074 16843 37100 16869
rect 37136 16843 37162 16869
rect 37198 16843 37224 16869
rect 37260 16843 37286 16869
rect 37322 16843 37348 16869
rect 37384 16843 37410 16869
rect 37446 16843 37472 16869
rect 37508 16843 37534 16869
rect 7799 16647 7825 16673
rect 8975 16647 9001 16673
rect 9479 16647 9505 16673
rect 10431 16647 10457 16673
rect 11775 16647 11801 16673
rect 12223 16647 12249 16673
rect 12447 16647 12473 16673
rect 13287 16647 13313 16673
rect 14239 16647 14265 16673
rect 15079 16647 15105 16673
rect 15975 16647 16001 16673
rect 16255 16647 16281 16673
rect 16759 16647 16785 16673
rect 16927 16647 16953 16673
rect 8975 16591 9001 16617
rect 10431 16591 10457 16617
rect 14239 16591 14265 16617
rect 15975 16591 16001 16617
rect 4574 16451 4600 16477
rect 4636 16451 4662 16477
rect 4698 16451 4724 16477
rect 4760 16451 4786 16477
rect 4822 16451 4848 16477
rect 4884 16451 4910 16477
rect 4946 16451 4972 16477
rect 5008 16451 5034 16477
rect 9574 16451 9600 16477
rect 9636 16451 9662 16477
rect 9698 16451 9724 16477
rect 9760 16451 9786 16477
rect 9822 16451 9848 16477
rect 9884 16451 9910 16477
rect 9946 16451 9972 16477
rect 10008 16451 10034 16477
rect 14574 16451 14600 16477
rect 14636 16451 14662 16477
rect 14698 16451 14724 16477
rect 14760 16451 14786 16477
rect 14822 16451 14848 16477
rect 14884 16451 14910 16477
rect 14946 16451 14972 16477
rect 15008 16451 15034 16477
rect 19574 16451 19600 16477
rect 19636 16451 19662 16477
rect 19698 16451 19724 16477
rect 19760 16451 19786 16477
rect 19822 16451 19848 16477
rect 19884 16451 19910 16477
rect 19946 16451 19972 16477
rect 20008 16451 20034 16477
rect 24574 16451 24600 16477
rect 24636 16451 24662 16477
rect 24698 16451 24724 16477
rect 24760 16451 24786 16477
rect 24822 16451 24848 16477
rect 24884 16451 24910 16477
rect 24946 16451 24972 16477
rect 25008 16451 25034 16477
rect 29574 16451 29600 16477
rect 29636 16451 29662 16477
rect 29698 16451 29724 16477
rect 29760 16451 29786 16477
rect 29822 16451 29848 16477
rect 29884 16451 29910 16477
rect 29946 16451 29972 16477
rect 30008 16451 30034 16477
rect 34574 16451 34600 16477
rect 34636 16451 34662 16477
rect 34698 16451 34724 16477
rect 34760 16451 34786 16477
rect 34822 16451 34848 16477
rect 34884 16451 34910 16477
rect 34946 16451 34972 16477
rect 35008 16451 35034 16477
rect 10991 16311 11017 16337
rect 14631 16311 14657 16337
rect 16311 16311 16337 16337
rect 17879 16311 17905 16337
rect 10095 16255 10121 16281
rect 10991 16255 11017 16281
rect 11271 16255 11297 16281
rect 11831 16255 11857 16281
rect 11943 16255 11969 16281
rect 13735 16255 13761 16281
rect 14407 16255 14433 16281
rect 15135 16255 15161 16281
rect 16311 16255 16337 16281
rect 16815 16255 16841 16281
rect 17879 16255 17905 16281
rect 18271 16255 18297 16281
rect 18719 16255 18745 16281
rect 18943 16255 18969 16281
rect 2074 16059 2100 16085
rect 2136 16059 2162 16085
rect 2198 16059 2224 16085
rect 2260 16059 2286 16085
rect 2322 16059 2348 16085
rect 2384 16059 2410 16085
rect 2446 16059 2472 16085
rect 2508 16059 2534 16085
rect 7074 16059 7100 16085
rect 7136 16059 7162 16085
rect 7198 16059 7224 16085
rect 7260 16059 7286 16085
rect 7322 16059 7348 16085
rect 7384 16059 7410 16085
rect 7446 16059 7472 16085
rect 7508 16059 7534 16085
rect 12074 16059 12100 16085
rect 12136 16059 12162 16085
rect 12198 16059 12224 16085
rect 12260 16059 12286 16085
rect 12322 16059 12348 16085
rect 12384 16059 12410 16085
rect 12446 16059 12472 16085
rect 12508 16059 12534 16085
rect 17074 16059 17100 16085
rect 17136 16059 17162 16085
rect 17198 16059 17224 16085
rect 17260 16059 17286 16085
rect 17322 16059 17348 16085
rect 17384 16059 17410 16085
rect 17446 16059 17472 16085
rect 17508 16059 17534 16085
rect 22074 16059 22100 16085
rect 22136 16059 22162 16085
rect 22198 16059 22224 16085
rect 22260 16059 22286 16085
rect 22322 16059 22348 16085
rect 22384 16059 22410 16085
rect 22446 16059 22472 16085
rect 22508 16059 22534 16085
rect 27074 16059 27100 16085
rect 27136 16059 27162 16085
rect 27198 16059 27224 16085
rect 27260 16059 27286 16085
rect 27322 16059 27348 16085
rect 27384 16059 27410 16085
rect 27446 16059 27472 16085
rect 27508 16059 27534 16085
rect 32074 16059 32100 16085
rect 32136 16059 32162 16085
rect 32198 16059 32224 16085
rect 32260 16059 32286 16085
rect 32322 16059 32348 16085
rect 32384 16059 32410 16085
rect 32446 16059 32472 16085
rect 32508 16059 32534 16085
rect 37074 16059 37100 16085
rect 37136 16059 37162 16085
rect 37198 16059 37224 16085
rect 37260 16059 37286 16085
rect 37322 16059 37348 16085
rect 37384 16059 37410 16085
rect 37446 16059 37472 16085
rect 37508 16059 37534 16085
rect 8079 15863 8105 15889
rect 8975 15863 9001 15889
rect 9479 15863 9505 15889
rect 10431 15863 10457 15889
rect 11775 15863 11801 15889
rect 12223 15863 12249 15889
rect 12447 15863 12473 15889
rect 13287 15863 13313 15889
rect 14407 15863 14433 15889
rect 15079 15863 15105 15889
rect 15975 15863 16001 15889
rect 16255 15863 16281 15889
rect 16815 15863 16841 15889
rect 16927 15863 16953 15889
rect 18775 15863 18801 15889
rect 19223 15863 19249 15889
rect 19447 15863 19473 15889
rect 8975 15807 9001 15833
rect 10431 15807 10457 15833
rect 14407 15807 14433 15833
rect 15975 15807 16001 15833
rect 4574 15667 4600 15693
rect 4636 15667 4662 15693
rect 4698 15667 4724 15693
rect 4760 15667 4786 15693
rect 4822 15667 4848 15693
rect 4884 15667 4910 15693
rect 4946 15667 4972 15693
rect 5008 15667 5034 15693
rect 9574 15667 9600 15693
rect 9636 15667 9662 15693
rect 9698 15667 9724 15693
rect 9760 15667 9786 15693
rect 9822 15667 9848 15693
rect 9884 15667 9910 15693
rect 9946 15667 9972 15693
rect 10008 15667 10034 15693
rect 14574 15667 14600 15693
rect 14636 15667 14662 15693
rect 14698 15667 14724 15693
rect 14760 15667 14786 15693
rect 14822 15667 14848 15693
rect 14884 15667 14910 15693
rect 14946 15667 14972 15693
rect 15008 15667 15034 15693
rect 19574 15667 19600 15693
rect 19636 15667 19662 15693
rect 19698 15667 19724 15693
rect 19760 15667 19786 15693
rect 19822 15667 19848 15693
rect 19884 15667 19910 15693
rect 19946 15667 19972 15693
rect 20008 15667 20034 15693
rect 24574 15667 24600 15693
rect 24636 15667 24662 15693
rect 24698 15667 24724 15693
rect 24760 15667 24786 15693
rect 24822 15667 24848 15693
rect 24884 15667 24910 15693
rect 24946 15667 24972 15693
rect 25008 15667 25034 15693
rect 29574 15667 29600 15693
rect 29636 15667 29662 15693
rect 29698 15667 29724 15693
rect 29760 15667 29786 15693
rect 29822 15667 29848 15693
rect 29884 15667 29910 15693
rect 29946 15667 29972 15693
rect 30008 15667 30034 15693
rect 34574 15667 34600 15693
rect 34636 15667 34662 15693
rect 34698 15667 34724 15693
rect 34760 15667 34786 15693
rect 34822 15667 34848 15693
rect 34884 15667 34910 15693
rect 34946 15667 34972 15693
rect 35008 15667 35034 15693
rect 1863 15527 1889 15553
rect 4495 15527 4521 15553
rect 7015 15527 7041 15553
rect 8471 15527 8497 15553
rect 10991 15527 11017 15553
rect 16143 15527 16169 15553
rect 17879 15527 17905 15553
rect 23423 15527 23449 15553
rect 1863 15471 1889 15497
rect 2759 15471 2785 15497
rect 3319 15471 3345 15497
rect 4495 15471 4521 15497
rect 6119 15471 6145 15497
rect 7015 15471 7041 15497
rect 7575 15471 7601 15497
rect 8471 15471 8497 15497
rect 10039 15471 10065 15497
rect 10991 15471 11017 15497
rect 11271 15471 11297 15497
rect 11831 15471 11857 15497
rect 11943 15471 11969 15497
rect 13735 15471 13761 15497
rect 14295 15471 14321 15497
rect 14463 15471 14489 15497
rect 15191 15471 15217 15497
rect 15975 15471 16001 15497
rect 16815 15471 16841 15497
rect 17879 15471 17905 15497
rect 18271 15471 18297 15497
rect 18719 15471 18745 15497
rect 18943 15471 18969 15497
rect 20791 15471 20817 15497
rect 21239 15471 21265 15497
rect 21463 15471 21489 15497
rect 22527 15471 22553 15497
rect 23423 15471 23449 15497
rect 2074 15275 2100 15301
rect 2136 15275 2162 15301
rect 2198 15275 2224 15301
rect 2260 15275 2286 15301
rect 2322 15275 2348 15301
rect 2384 15275 2410 15301
rect 2446 15275 2472 15301
rect 2508 15275 2534 15301
rect 7074 15275 7100 15301
rect 7136 15275 7162 15301
rect 7198 15275 7224 15301
rect 7260 15275 7286 15301
rect 7322 15275 7348 15301
rect 7384 15275 7410 15301
rect 7446 15275 7472 15301
rect 7508 15275 7534 15301
rect 12074 15275 12100 15301
rect 12136 15275 12162 15301
rect 12198 15275 12224 15301
rect 12260 15275 12286 15301
rect 12322 15275 12348 15301
rect 12384 15275 12410 15301
rect 12446 15275 12472 15301
rect 12508 15275 12534 15301
rect 17074 15275 17100 15301
rect 17136 15275 17162 15301
rect 17198 15275 17224 15301
rect 17260 15275 17286 15301
rect 17322 15275 17348 15301
rect 17384 15275 17410 15301
rect 17446 15275 17472 15301
rect 17508 15275 17534 15301
rect 22074 15275 22100 15301
rect 22136 15275 22162 15301
rect 22198 15275 22224 15301
rect 22260 15275 22286 15301
rect 22322 15275 22348 15301
rect 22384 15275 22410 15301
rect 22446 15275 22472 15301
rect 22508 15275 22534 15301
rect 27074 15275 27100 15301
rect 27136 15275 27162 15301
rect 27198 15275 27224 15301
rect 27260 15275 27286 15301
rect 27322 15275 27348 15301
rect 27384 15275 27410 15301
rect 27446 15275 27472 15301
rect 27508 15275 27534 15301
rect 32074 15275 32100 15301
rect 32136 15275 32162 15301
rect 32198 15275 32224 15301
rect 32260 15275 32286 15301
rect 32322 15275 32348 15301
rect 32384 15275 32410 15301
rect 32446 15275 32472 15301
rect 32508 15275 32534 15301
rect 37074 15275 37100 15301
rect 37136 15275 37162 15301
rect 37198 15275 37224 15301
rect 37260 15275 37286 15301
rect 37322 15275 37348 15301
rect 37384 15275 37410 15301
rect 37446 15275 37472 15301
rect 37508 15275 37534 15301
rect 1527 15079 1553 15105
rect 2479 15079 2505 15105
rect 3823 15079 3849 15105
rect 4383 15079 4409 15105
rect 4495 15079 4521 15105
rect 5559 15079 5585 15105
rect 5839 15079 5865 15105
rect 6455 15079 6481 15105
rect 8079 15079 8105 15105
rect 8975 15079 9001 15105
rect 9479 15079 9505 15105
rect 10431 15079 10457 15105
rect 11775 15079 11801 15105
rect 12727 15079 12753 15105
rect 13287 15079 13313 15105
rect 14407 15079 14433 15105
rect 15079 15079 15105 15105
rect 15975 15079 16001 15105
rect 16255 15079 16281 15105
rect 16983 15079 17009 15105
rect 18831 15079 18857 15105
rect 19335 15079 19361 15105
rect 19447 15079 19473 15105
rect 20511 15079 20537 15105
rect 21015 15079 21041 15105
rect 23031 15079 23057 15105
rect 23927 15079 23953 15105
rect 24487 15079 24513 15105
rect 25327 15079 25353 15105
rect 1527 15023 1553 15049
rect 8975 15023 9001 15049
rect 10431 15023 10457 15049
rect 12727 15023 12753 15049
rect 14407 15023 14433 15049
rect 15975 15023 16001 15049
rect 17207 15023 17233 15049
rect 21183 15023 21209 15049
rect 23927 15023 23953 15049
rect 25327 15023 25353 15049
rect 4574 14883 4600 14909
rect 4636 14883 4662 14909
rect 4698 14883 4724 14909
rect 4760 14883 4786 14909
rect 4822 14883 4848 14909
rect 4884 14883 4910 14909
rect 4946 14883 4972 14909
rect 5008 14883 5034 14909
rect 9574 14883 9600 14909
rect 9636 14883 9662 14909
rect 9698 14883 9724 14909
rect 9760 14883 9786 14909
rect 9822 14883 9848 14909
rect 9884 14883 9910 14909
rect 9946 14883 9972 14909
rect 10008 14883 10034 14909
rect 14574 14883 14600 14909
rect 14636 14883 14662 14909
rect 14698 14883 14724 14909
rect 14760 14883 14786 14909
rect 14822 14883 14848 14909
rect 14884 14883 14910 14909
rect 14946 14883 14972 14909
rect 15008 14883 15034 14909
rect 19574 14883 19600 14909
rect 19636 14883 19662 14909
rect 19698 14883 19724 14909
rect 19760 14883 19786 14909
rect 19822 14883 19848 14909
rect 19884 14883 19910 14909
rect 19946 14883 19972 14909
rect 20008 14883 20034 14909
rect 24574 14883 24600 14909
rect 24636 14883 24662 14909
rect 24698 14883 24724 14909
rect 24760 14883 24786 14909
rect 24822 14883 24848 14909
rect 24884 14883 24910 14909
rect 24946 14883 24972 14909
rect 25008 14883 25034 14909
rect 29574 14883 29600 14909
rect 29636 14883 29662 14909
rect 29698 14883 29724 14909
rect 29760 14883 29786 14909
rect 29822 14883 29848 14909
rect 29884 14883 29910 14909
rect 29946 14883 29972 14909
rect 30008 14883 30034 14909
rect 34574 14883 34600 14909
rect 34636 14883 34662 14909
rect 34698 14883 34724 14909
rect 34760 14883 34786 14909
rect 34822 14883 34848 14909
rect 34884 14883 34910 14909
rect 34946 14883 34972 14909
rect 35008 14883 35034 14909
rect 4495 14743 4521 14769
rect 7015 14743 7041 14769
rect 8471 14743 8497 14769
rect 12447 14743 12473 14769
rect 16367 14743 16393 14769
rect 17935 14743 17961 14769
rect 19447 14743 19473 14769
rect 23423 14743 23449 14769
rect 2367 14687 2393 14713
rect 2479 14687 2505 14713
rect 2759 14687 2785 14713
rect 3319 14687 3345 14713
rect 4495 14687 4521 14713
rect 6119 14687 6145 14713
rect 7015 14687 7041 14713
rect 7575 14687 7601 14713
rect 8471 14687 8497 14713
rect 10039 14687 10065 14713
rect 10375 14687 10401 14713
rect 10487 14687 10513 14713
rect 11271 14687 11297 14713
rect 12447 14687 12473 14713
rect 13735 14687 13761 14713
rect 14295 14687 14321 14713
rect 14463 14687 14489 14713
rect 15191 14687 15217 14713
rect 16367 14687 16393 14713
rect 16815 14687 16841 14713
rect 17935 14687 17961 14713
rect 18271 14687 18297 14713
rect 19447 14687 19473 14713
rect 20791 14687 20817 14713
rect 21239 14687 21265 14713
rect 21463 14687 21489 14713
rect 22527 14687 22553 14713
rect 23423 14687 23449 14713
rect 25047 14687 25073 14713
rect 25327 14687 25353 14713
rect 25439 14687 25465 14713
rect 2074 14491 2100 14517
rect 2136 14491 2162 14517
rect 2198 14491 2224 14517
rect 2260 14491 2286 14517
rect 2322 14491 2348 14517
rect 2384 14491 2410 14517
rect 2446 14491 2472 14517
rect 2508 14491 2534 14517
rect 7074 14491 7100 14517
rect 7136 14491 7162 14517
rect 7198 14491 7224 14517
rect 7260 14491 7286 14517
rect 7322 14491 7348 14517
rect 7384 14491 7410 14517
rect 7446 14491 7472 14517
rect 7508 14491 7534 14517
rect 12074 14491 12100 14517
rect 12136 14491 12162 14517
rect 12198 14491 12224 14517
rect 12260 14491 12286 14517
rect 12322 14491 12348 14517
rect 12384 14491 12410 14517
rect 12446 14491 12472 14517
rect 12508 14491 12534 14517
rect 17074 14491 17100 14517
rect 17136 14491 17162 14517
rect 17198 14491 17224 14517
rect 17260 14491 17286 14517
rect 17322 14491 17348 14517
rect 17384 14491 17410 14517
rect 17446 14491 17472 14517
rect 17508 14491 17534 14517
rect 22074 14491 22100 14517
rect 22136 14491 22162 14517
rect 22198 14491 22224 14517
rect 22260 14491 22286 14517
rect 22322 14491 22348 14517
rect 22384 14491 22410 14517
rect 22446 14491 22472 14517
rect 22508 14491 22534 14517
rect 27074 14491 27100 14517
rect 27136 14491 27162 14517
rect 27198 14491 27224 14517
rect 27260 14491 27286 14517
rect 27322 14491 27348 14517
rect 27384 14491 27410 14517
rect 27446 14491 27472 14517
rect 27508 14491 27534 14517
rect 32074 14491 32100 14517
rect 32136 14491 32162 14517
rect 32198 14491 32224 14517
rect 32260 14491 32286 14517
rect 32322 14491 32348 14517
rect 32384 14491 32410 14517
rect 32446 14491 32472 14517
rect 32508 14491 32534 14517
rect 37074 14491 37100 14517
rect 37136 14491 37162 14517
rect 37198 14491 37224 14517
rect 37260 14491 37286 14517
rect 37322 14491 37348 14517
rect 37384 14491 37410 14517
rect 37446 14491 37472 14517
rect 37508 14491 37534 14517
rect 1751 14295 1777 14321
rect 2479 14295 2505 14321
rect 3823 14295 3849 14321
rect 4383 14295 4409 14321
rect 4495 14295 4521 14321
rect 5559 14295 5585 14321
rect 5839 14295 5865 14321
rect 6455 14295 6481 14321
rect 8079 14295 8105 14321
rect 8975 14295 9001 14321
rect 9479 14295 9505 14321
rect 10375 14295 10401 14321
rect 11775 14295 11801 14321
rect 12615 14295 12641 14321
rect 13287 14295 13313 14321
rect 14407 14295 14433 14321
rect 15079 14295 15105 14321
rect 15975 14295 16001 14321
rect 16255 14295 16281 14321
rect 17431 14295 17457 14321
rect 18831 14295 18857 14321
rect 19335 14295 19361 14321
rect 19447 14295 19473 14321
rect 20511 14295 20537 14321
rect 20679 14295 20705 14321
rect 21015 14295 21041 14321
rect 23031 14295 23057 14321
rect 23927 14295 23953 14321
rect 24487 14295 24513 14321
rect 25383 14295 25409 14321
rect 26727 14295 26753 14321
rect 27679 14295 27705 14321
rect 28463 14295 28489 14321
rect 29359 14295 29385 14321
rect 1527 14239 1553 14265
rect 8975 14239 9001 14265
rect 10375 14239 10401 14265
rect 12727 14239 12753 14265
rect 14407 14239 14433 14265
rect 15975 14239 16001 14265
rect 17431 14239 17457 14265
rect 23927 14239 23953 14265
rect 25383 14239 25409 14265
rect 27679 14239 27705 14265
rect 29359 14239 29385 14265
rect 4574 14099 4600 14125
rect 4636 14099 4662 14125
rect 4698 14099 4724 14125
rect 4760 14099 4786 14125
rect 4822 14099 4848 14125
rect 4884 14099 4910 14125
rect 4946 14099 4972 14125
rect 5008 14099 5034 14125
rect 9574 14099 9600 14125
rect 9636 14099 9662 14125
rect 9698 14099 9724 14125
rect 9760 14099 9786 14125
rect 9822 14099 9848 14125
rect 9884 14099 9910 14125
rect 9946 14099 9972 14125
rect 10008 14099 10034 14125
rect 14574 14099 14600 14125
rect 14636 14099 14662 14125
rect 14698 14099 14724 14125
rect 14760 14099 14786 14125
rect 14822 14099 14848 14125
rect 14884 14099 14910 14125
rect 14946 14099 14972 14125
rect 15008 14099 15034 14125
rect 19574 14099 19600 14125
rect 19636 14099 19662 14125
rect 19698 14099 19724 14125
rect 19760 14099 19786 14125
rect 19822 14099 19848 14125
rect 19884 14099 19910 14125
rect 19946 14099 19972 14125
rect 20008 14099 20034 14125
rect 24574 14099 24600 14125
rect 24636 14099 24662 14125
rect 24698 14099 24724 14125
rect 24760 14099 24786 14125
rect 24822 14099 24848 14125
rect 24884 14099 24910 14125
rect 24946 14099 24972 14125
rect 25008 14099 25034 14125
rect 29574 14099 29600 14125
rect 29636 14099 29662 14125
rect 29698 14099 29724 14125
rect 29760 14099 29786 14125
rect 29822 14099 29848 14125
rect 29884 14099 29910 14125
rect 29946 14099 29972 14125
rect 30008 14099 30034 14125
rect 34574 14099 34600 14125
rect 34636 14099 34662 14125
rect 34698 14099 34724 14125
rect 34760 14099 34786 14125
rect 34822 14099 34848 14125
rect 34884 14099 34910 14125
rect 34946 14099 34972 14125
rect 35008 14099 35034 14125
rect 1975 13959 2001 13985
rect 4495 13959 4521 13985
rect 7015 13959 7041 13985
rect 8471 13959 8497 13985
rect 10767 13959 10793 13985
rect 12447 13959 12473 13985
rect 14911 13959 14937 13985
rect 16367 13959 16393 13985
rect 17935 13959 17961 13985
rect 19447 13959 19473 13985
rect 23423 13959 23449 13985
rect 25943 13959 25969 13985
rect 27399 13959 27425 13985
rect 1975 13903 2001 13929
rect 2759 13903 2785 13929
rect 3319 13903 3345 13929
rect 4495 13903 4521 13929
rect 6119 13903 6145 13929
rect 7015 13903 7041 13929
rect 7575 13903 7601 13929
rect 8471 13903 8497 13929
rect 10095 13903 10121 13929
rect 10767 13903 10793 13929
rect 11271 13903 11297 13929
rect 12447 13903 12473 13929
rect 13735 13903 13761 13929
rect 14911 13903 14937 13929
rect 15191 13903 15217 13929
rect 16367 13903 16393 13929
rect 16815 13903 16841 13929
rect 17935 13903 17961 13929
rect 18271 13903 18297 13929
rect 19447 13903 19473 13929
rect 20959 13903 20985 13929
rect 21239 13903 21265 13929
rect 21463 13903 21489 13929
rect 22527 13903 22553 13929
rect 23423 13903 23449 13929
rect 25047 13903 25073 13929
rect 25943 13903 25969 13929
rect 26223 13903 26249 13929
rect 27399 13903 27425 13929
rect 2074 13707 2100 13733
rect 2136 13707 2162 13733
rect 2198 13707 2224 13733
rect 2260 13707 2286 13733
rect 2322 13707 2348 13733
rect 2384 13707 2410 13733
rect 2446 13707 2472 13733
rect 2508 13707 2534 13733
rect 7074 13707 7100 13733
rect 7136 13707 7162 13733
rect 7198 13707 7224 13733
rect 7260 13707 7286 13733
rect 7322 13707 7348 13733
rect 7384 13707 7410 13733
rect 7446 13707 7472 13733
rect 7508 13707 7534 13733
rect 12074 13707 12100 13733
rect 12136 13707 12162 13733
rect 12198 13707 12224 13733
rect 12260 13707 12286 13733
rect 12322 13707 12348 13733
rect 12384 13707 12410 13733
rect 12446 13707 12472 13733
rect 12508 13707 12534 13733
rect 17074 13707 17100 13733
rect 17136 13707 17162 13733
rect 17198 13707 17224 13733
rect 17260 13707 17286 13733
rect 17322 13707 17348 13733
rect 17384 13707 17410 13733
rect 17446 13707 17472 13733
rect 17508 13707 17534 13733
rect 22074 13707 22100 13733
rect 22136 13707 22162 13733
rect 22198 13707 22224 13733
rect 22260 13707 22286 13733
rect 22322 13707 22348 13733
rect 22384 13707 22410 13733
rect 22446 13707 22472 13733
rect 22508 13707 22534 13733
rect 27074 13707 27100 13733
rect 27136 13707 27162 13733
rect 27198 13707 27224 13733
rect 27260 13707 27286 13733
rect 27322 13707 27348 13733
rect 27384 13707 27410 13733
rect 27446 13707 27472 13733
rect 27508 13707 27534 13733
rect 32074 13707 32100 13733
rect 32136 13707 32162 13733
rect 32198 13707 32224 13733
rect 32260 13707 32286 13733
rect 32322 13707 32348 13733
rect 32384 13707 32410 13733
rect 32446 13707 32472 13733
rect 32508 13707 32534 13733
rect 37074 13707 37100 13733
rect 37136 13707 37162 13733
rect 37198 13707 37224 13733
rect 37260 13707 37286 13733
rect 37322 13707 37348 13733
rect 37384 13707 37410 13733
rect 37446 13707 37472 13733
rect 37508 13707 37534 13733
rect 1807 13511 1833 13537
rect 1975 13511 2001 13537
rect 2479 13511 2505 13537
rect 3823 13511 3849 13537
rect 4383 13511 4409 13537
rect 4495 13511 4521 13537
rect 5503 13511 5529 13537
rect 5839 13511 5865 13537
rect 6455 13511 6481 13537
rect 8079 13511 8105 13537
rect 8359 13511 8385 13537
rect 8471 13511 8497 13537
rect 9479 13511 9505 13537
rect 10431 13511 10457 13537
rect 11775 13511 11801 13537
rect 12951 13511 12977 13537
rect 13287 13511 13313 13537
rect 14127 13511 14153 13537
rect 15471 13511 15497 13537
rect 16255 13511 16281 13537
rect 16815 13511 16841 13537
rect 17935 13511 17961 13537
rect 18831 13511 18857 13537
rect 19335 13511 19361 13537
rect 19447 13511 19473 13537
rect 20511 13511 20537 13537
rect 21015 13511 21041 13537
rect 23031 13511 23057 13537
rect 23927 13511 23953 13537
rect 24487 13511 24513 13537
rect 25383 13511 25409 13537
rect 26727 13511 26753 13537
rect 27679 13511 27705 13537
rect 28463 13511 28489 13537
rect 29359 13511 29385 13537
rect 10431 13455 10457 13481
rect 12951 13455 12977 13481
rect 14407 13455 14433 13481
rect 16255 13455 16281 13481
rect 17935 13455 17961 13481
rect 21183 13455 21209 13481
rect 23927 13455 23953 13481
rect 25383 13455 25409 13481
rect 27679 13455 27705 13481
rect 29359 13455 29385 13481
rect 4574 13315 4600 13341
rect 4636 13315 4662 13341
rect 4698 13315 4724 13341
rect 4760 13315 4786 13341
rect 4822 13315 4848 13341
rect 4884 13315 4910 13341
rect 4946 13315 4972 13341
rect 5008 13315 5034 13341
rect 9574 13315 9600 13341
rect 9636 13315 9662 13341
rect 9698 13315 9724 13341
rect 9760 13315 9786 13341
rect 9822 13315 9848 13341
rect 9884 13315 9910 13341
rect 9946 13315 9972 13341
rect 10008 13315 10034 13341
rect 14574 13315 14600 13341
rect 14636 13315 14662 13341
rect 14698 13315 14724 13341
rect 14760 13315 14786 13341
rect 14822 13315 14848 13341
rect 14884 13315 14910 13341
rect 14946 13315 14972 13341
rect 15008 13315 15034 13341
rect 19574 13315 19600 13341
rect 19636 13315 19662 13341
rect 19698 13315 19724 13341
rect 19760 13315 19786 13341
rect 19822 13315 19848 13341
rect 19884 13315 19910 13341
rect 19946 13315 19972 13341
rect 20008 13315 20034 13341
rect 24574 13315 24600 13341
rect 24636 13315 24662 13341
rect 24698 13315 24724 13341
rect 24760 13315 24786 13341
rect 24822 13315 24848 13341
rect 24884 13315 24910 13341
rect 24946 13315 24972 13341
rect 25008 13315 25034 13341
rect 29574 13315 29600 13341
rect 29636 13315 29662 13341
rect 29698 13315 29724 13341
rect 29760 13315 29786 13341
rect 29822 13315 29848 13341
rect 29884 13315 29910 13341
rect 29946 13315 29972 13341
rect 30008 13315 30034 13341
rect 34574 13315 34600 13341
rect 34636 13315 34662 13341
rect 34698 13315 34724 13341
rect 34760 13315 34786 13341
rect 34822 13315 34848 13341
rect 34884 13315 34910 13341
rect 34946 13315 34972 13341
rect 35008 13315 35034 13341
rect 4495 13175 4521 13201
rect 7015 13175 7041 13201
rect 8359 13175 8385 13201
rect 10767 13175 10793 13201
rect 14351 13175 14377 13201
rect 16031 13175 16057 13201
rect 17991 13175 18017 13201
rect 19447 13175 19473 13201
rect 23423 13175 23449 13201
rect 25943 13175 25969 13201
rect 2367 13119 2393 13145
rect 2591 13119 2617 13145
rect 2759 13119 2785 13145
rect 3599 13119 3625 13145
rect 4495 13119 4521 13145
rect 6119 13119 6145 13145
rect 7015 13119 7041 13145
rect 7575 13119 7601 13145
rect 8359 13119 8385 13145
rect 10095 13119 10121 13145
rect 10767 13119 10793 13145
rect 11271 13119 11297 13145
rect 11831 13119 11857 13145
rect 11999 13119 12025 13145
rect 13399 13119 13425 13145
rect 14183 13119 14209 13145
rect 15135 13119 15161 13145
rect 16031 13119 16057 13145
rect 16983 13119 17009 13145
rect 17991 13119 18017 13145
rect 18551 13119 18577 13145
rect 19447 13119 19473 13145
rect 20959 13119 20985 13145
rect 21239 13119 21265 13145
rect 21463 13119 21489 13145
rect 22527 13119 22553 13145
rect 23423 13119 23449 13145
rect 25047 13119 25073 13145
rect 25943 13119 25969 13145
rect 26503 13119 26529 13145
rect 26783 13119 26809 13145
rect 26895 13119 26921 13145
rect 29023 13119 29049 13145
rect 29303 13119 29329 13145
rect 29415 13119 29441 13145
rect 2074 12923 2100 12949
rect 2136 12923 2162 12949
rect 2198 12923 2224 12949
rect 2260 12923 2286 12949
rect 2322 12923 2348 12949
rect 2384 12923 2410 12949
rect 2446 12923 2472 12949
rect 2508 12923 2534 12949
rect 7074 12923 7100 12949
rect 7136 12923 7162 12949
rect 7198 12923 7224 12949
rect 7260 12923 7286 12949
rect 7322 12923 7348 12949
rect 7384 12923 7410 12949
rect 7446 12923 7472 12949
rect 7508 12923 7534 12949
rect 12074 12923 12100 12949
rect 12136 12923 12162 12949
rect 12198 12923 12224 12949
rect 12260 12923 12286 12949
rect 12322 12923 12348 12949
rect 12384 12923 12410 12949
rect 12446 12923 12472 12949
rect 12508 12923 12534 12949
rect 17074 12923 17100 12949
rect 17136 12923 17162 12949
rect 17198 12923 17224 12949
rect 17260 12923 17286 12949
rect 17322 12923 17348 12949
rect 17384 12923 17410 12949
rect 17446 12923 17472 12949
rect 17508 12923 17534 12949
rect 22074 12923 22100 12949
rect 22136 12923 22162 12949
rect 22198 12923 22224 12949
rect 22260 12923 22286 12949
rect 22322 12923 22348 12949
rect 22384 12923 22410 12949
rect 22446 12923 22472 12949
rect 22508 12923 22534 12949
rect 27074 12923 27100 12949
rect 27136 12923 27162 12949
rect 27198 12923 27224 12949
rect 27260 12923 27286 12949
rect 27322 12923 27348 12949
rect 27384 12923 27410 12949
rect 27446 12923 27472 12949
rect 27508 12923 27534 12949
rect 32074 12923 32100 12949
rect 32136 12923 32162 12949
rect 32198 12923 32224 12949
rect 32260 12923 32286 12949
rect 32322 12923 32348 12949
rect 32384 12923 32410 12949
rect 32446 12923 32472 12949
rect 32508 12923 32534 12949
rect 37074 12923 37100 12949
rect 37136 12923 37162 12949
rect 37198 12923 37224 12949
rect 37260 12923 37286 12949
rect 37322 12923 37348 12949
rect 37384 12923 37410 12949
rect 37446 12923 37472 12949
rect 37508 12923 37534 12949
rect 1807 12727 1833 12753
rect 1975 12727 2001 12753
rect 2479 12727 2505 12753
rect 3823 12727 3849 12753
rect 4999 12727 5025 12753
rect 5559 12727 5585 12753
rect 6455 12727 6481 12753
rect 8079 12727 8105 12753
rect 8359 12727 8385 12753
rect 8471 12727 8497 12753
rect 9479 12727 9505 12753
rect 10431 12727 10457 12753
rect 11775 12727 11801 12753
rect 12223 12727 12249 12753
rect 12447 12727 12473 12753
rect 13231 12727 13257 12753
rect 14183 12727 14209 12753
rect 15751 12727 15777 12753
rect 16647 12727 16673 12753
rect 16927 12727 16953 12753
rect 17879 12727 17905 12753
rect 18775 12727 18801 12753
rect 19951 12727 19977 12753
rect 20511 12727 20537 12753
rect 21183 12727 21209 12753
rect 22751 12727 22777 12753
rect 23311 12727 23337 12753
rect 23423 12727 23449 12753
rect 24375 12727 24401 12753
rect 24655 12727 24681 12753
rect 24879 12727 24905 12753
rect 26727 12727 26753 12753
rect 27175 12727 27201 12753
rect 27399 12727 27425 12753
rect 28463 12727 28489 12753
rect 29359 12727 29385 12753
rect 4999 12671 5025 12697
rect 6455 12671 6481 12697
rect 10431 12671 10457 12697
rect 14183 12671 14209 12697
rect 16647 12671 16673 12697
rect 17879 12671 17905 12697
rect 19951 12671 19977 12697
rect 21183 12671 21209 12697
rect 29359 12671 29385 12697
rect 4574 12531 4600 12557
rect 4636 12531 4662 12557
rect 4698 12531 4724 12557
rect 4760 12531 4786 12557
rect 4822 12531 4848 12557
rect 4884 12531 4910 12557
rect 4946 12531 4972 12557
rect 5008 12531 5034 12557
rect 9574 12531 9600 12557
rect 9636 12531 9662 12557
rect 9698 12531 9724 12557
rect 9760 12531 9786 12557
rect 9822 12531 9848 12557
rect 9884 12531 9910 12557
rect 9946 12531 9972 12557
rect 10008 12531 10034 12557
rect 14574 12531 14600 12557
rect 14636 12531 14662 12557
rect 14698 12531 14724 12557
rect 14760 12531 14786 12557
rect 14822 12531 14848 12557
rect 14884 12531 14910 12557
rect 14946 12531 14972 12557
rect 15008 12531 15034 12557
rect 19574 12531 19600 12557
rect 19636 12531 19662 12557
rect 19698 12531 19724 12557
rect 19760 12531 19786 12557
rect 19822 12531 19848 12557
rect 19884 12531 19910 12557
rect 19946 12531 19972 12557
rect 20008 12531 20034 12557
rect 24574 12531 24600 12557
rect 24636 12531 24662 12557
rect 24698 12531 24724 12557
rect 24760 12531 24786 12557
rect 24822 12531 24848 12557
rect 24884 12531 24910 12557
rect 24946 12531 24972 12557
rect 25008 12531 25034 12557
rect 29574 12531 29600 12557
rect 29636 12531 29662 12557
rect 29698 12531 29724 12557
rect 29760 12531 29786 12557
rect 29822 12531 29848 12557
rect 29884 12531 29910 12557
rect 29946 12531 29972 12557
rect 30008 12531 30034 12557
rect 34574 12531 34600 12557
rect 34636 12531 34662 12557
rect 34698 12531 34724 12557
rect 34760 12531 34786 12557
rect 34822 12531 34848 12557
rect 34884 12531 34910 12557
rect 34946 12531 34972 12557
rect 35008 12531 35034 12557
rect 3039 12391 3065 12417
rect 4495 12391 4521 12417
rect 7015 12391 7041 12417
rect 8359 12391 8385 12417
rect 14967 12391 14993 12417
rect 16423 12391 16449 12417
rect 17879 12391 17905 12417
rect 19447 12391 19473 12417
rect 23423 12391 23449 12417
rect 27175 12391 27201 12417
rect 29695 12391 29721 12417
rect 31151 12391 31177 12417
rect 1919 12335 1945 12361
rect 3039 12335 3065 12361
rect 3599 12335 3625 12361
rect 4495 12335 4521 12361
rect 6119 12335 6145 12361
rect 7015 12335 7041 12361
rect 7575 12335 7601 12361
rect 8359 12335 8385 12361
rect 10095 12335 10121 12361
rect 10375 12335 10401 12361
rect 10487 12335 10513 12361
rect 11271 12335 11297 12361
rect 11831 12335 11857 12361
rect 11999 12335 12025 12361
rect 14071 12335 14097 12361
rect 14967 12335 14993 12361
rect 15527 12335 15553 12361
rect 16423 12335 16449 12361
rect 16927 12335 16953 12361
rect 17879 12335 17905 12361
rect 18551 12335 18577 12361
rect 19447 12335 19473 12361
rect 20959 12335 20985 12361
rect 21239 12335 21265 12361
rect 21463 12335 21489 12361
rect 22527 12335 22553 12361
rect 23423 12335 23449 12361
rect 24767 12335 24793 12361
rect 25215 12335 25241 12361
rect 25439 12335 25465 12361
rect 26503 12335 26529 12361
rect 26895 12335 26921 12361
rect 29023 12335 29049 12361
rect 29471 12335 29497 12361
rect 30479 12335 30505 12361
rect 31095 12335 31121 12361
rect 2074 12139 2100 12165
rect 2136 12139 2162 12165
rect 2198 12139 2224 12165
rect 2260 12139 2286 12165
rect 2322 12139 2348 12165
rect 2384 12139 2410 12165
rect 2446 12139 2472 12165
rect 2508 12139 2534 12165
rect 7074 12139 7100 12165
rect 7136 12139 7162 12165
rect 7198 12139 7224 12165
rect 7260 12139 7286 12165
rect 7322 12139 7348 12165
rect 7384 12139 7410 12165
rect 7446 12139 7472 12165
rect 7508 12139 7534 12165
rect 12074 12139 12100 12165
rect 12136 12139 12162 12165
rect 12198 12139 12224 12165
rect 12260 12139 12286 12165
rect 12322 12139 12348 12165
rect 12384 12139 12410 12165
rect 12446 12139 12472 12165
rect 12508 12139 12534 12165
rect 17074 12139 17100 12165
rect 17136 12139 17162 12165
rect 17198 12139 17224 12165
rect 17260 12139 17286 12165
rect 17322 12139 17348 12165
rect 17384 12139 17410 12165
rect 17446 12139 17472 12165
rect 17508 12139 17534 12165
rect 22074 12139 22100 12165
rect 22136 12139 22162 12165
rect 22198 12139 22224 12165
rect 22260 12139 22286 12165
rect 22322 12139 22348 12165
rect 22384 12139 22410 12165
rect 22446 12139 22472 12165
rect 22508 12139 22534 12165
rect 27074 12139 27100 12165
rect 27136 12139 27162 12165
rect 27198 12139 27224 12165
rect 27260 12139 27286 12165
rect 27322 12139 27348 12165
rect 27384 12139 27410 12165
rect 27446 12139 27472 12165
rect 27508 12139 27534 12165
rect 32074 12139 32100 12165
rect 32136 12139 32162 12165
rect 32198 12139 32224 12165
rect 32260 12139 32286 12165
rect 32322 12139 32348 12165
rect 32384 12139 32410 12165
rect 32446 12139 32472 12165
rect 32508 12139 32534 12165
rect 37074 12139 37100 12165
rect 37136 12139 37162 12165
rect 37198 12139 37224 12165
rect 37260 12139 37286 12165
rect 37322 12139 37348 12165
rect 37384 12139 37410 12165
rect 37446 12139 37472 12165
rect 37508 12139 37534 12165
rect 1583 11943 1609 11969
rect 2479 11943 2505 11969
rect 3823 11943 3849 11969
rect 4999 11943 5025 11969
rect 5559 11943 5585 11969
rect 6455 11943 6481 11969
rect 8079 11943 8105 11969
rect 8975 11943 9001 11969
rect 9535 11943 9561 11969
rect 9703 11943 9729 11969
rect 10375 11943 10401 11969
rect 11775 11943 11801 11969
rect 12223 11943 12249 11969
rect 12447 11943 12473 11969
rect 13231 11943 13257 11969
rect 14407 11943 14433 11969
rect 15863 11943 15889 11969
rect 16759 11943 16785 11969
rect 17039 11943 17065 11969
rect 17879 11943 17905 11969
rect 18775 11943 18801 11969
rect 19951 11943 19977 11969
rect 20511 11943 20537 11969
rect 21183 11943 21209 11969
rect 22807 11943 22833 11969
rect 23927 11943 23953 11969
rect 24375 11943 24401 11969
rect 25159 11943 25185 11969
rect 27007 11943 27033 11969
rect 27567 11943 27593 11969
rect 28463 11943 28489 11969
rect 28967 11943 28993 11969
rect 30983 11943 31009 11969
rect 31151 11943 31177 11969
rect 31375 11943 31401 11969
rect 32159 11943 32185 11969
rect 32831 11943 32857 11969
rect 2479 11887 2505 11913
rect 4999 11887 5025 11913
rect 6455 11887 6481 11913
rect 8975 11887 9001 11913
rect 14407 11887 14433 11913
rect 16759 11887 16785 11913
rect 17991 11887 18017 11913
rect 19951 11887 19977 11913
rect 21183 11887 21209 11913
rect 23927 11887 23953 11913
rect 25159 11887 25185 11913
rect 27679 11887 27705 11913
rect 29135 11887 29161 11913
rect 33111 11887 33137 11913
rect 4574 11747 4600 11773
rect 4636 11747 4662 11773
rect 4698 11747 4724 11773
rect 4760 11747 4786 11773
rect 4822 11747 4848 11773
rect 4884 11747 4910 11773
rect 4946 11747 4972 11773
rect 5008 11747 5034 11773
rect 9574 11747 9600 11773
rect 9636 11747 9662 11773
rect 9698 11747 9724 11773
rect 9760 11747 9786 11773
rect 9822 11747 9848 11773
rect 9884 11747 9910 11773
rect 9946 11747 9972 11773
rect 10008 11747 10034 11773
rect 14574 11747 14600 11773
rect 14636 11747 14662 11773
rect 14698 11747 14724 11773
rect 14760 11747 14786 11773
rect 14822 11747 14848 11773
rect 14884 11747 14910 11773
rect 14946 11747 14972 11773
rect 15008 11747 15034 11773
rect 19574 11747 19600 11773
rect 19636 11747 19662 11773
rect 19698 11747 19724 11773
rect 19760 11747 19786 11773
rect 19822 11747 19848 11773
rect 19884 11747 19910 11773
rect 19946 11747 19972 11773
rect 20008 11747 20034 11773
rect 24574 11747 24600 11773
rect 24636 11747 24662 11773
rect 24698 11747 24724 11773
rect 24760 11747 24786 11773
rect 24822 11747 24848 11773
rect 24884 11747 24910 11773
rect 24946 11747 24972 11773
rect 25008 11747 25034 11773
rect 29574 11747 29600 11773
rect 29636 11747 29662 11773
rect 29698 11747 29724 11773
rect 29760 11747 29786 11773
rect 29822 11747 29848 11773
rect 29884 11747 29910 11773
rect 29946 11747 29972 11773
rect 30008 11747 30034 11773
rect 34574 11747 34600 11773
rect 34636 11747 34662 11773
rect 34698 11747 34724 11773
rect 34760 11747 34786 11773
rect 34822 11747 34848 11773
rect 34884 11747 34910 11773
rect 34946 11747 34972 11773
rect 35008 11747 35034 11773
rect 3039 11607 3065 11633
rect 4495 11607 4521 11633
rect 8471 11607 8497 11633
rect 14967 11607 14993 11633
rect 16199 11607 16225 11633
rect 17991 11607 18017 11633
rect 19335 11607 19361 11633
rect 23311 11607 23337 11633
rect 29919 11607 29945 11633
rect 31375 11607 31401 11633
rect 33895 11607 33921 11633
rect 1919 11551 1945 11577
rect 3039 11551 3065 11577
rect 3599 11551 3625 11577
rect 4495 11551 4521 11577
rect 5839 11551 5865 11577
rect 6399 11551 6425 11577
rect 6511 11551 6537 11577
rect 7575 11551 7601 11577
rect 8471 11551 8497 11577
rect 9815 11551 9841 11577
rect 10375 11551 10401 11577
rect 10487 11551 10513 11577
rect 11327 11551 11353 11577
rect 11831 11551 11857 11577
rect 11999 11551 12025 11577
rect 14071 11551 14097 11577
rect 14967 11551 14993 11577
rect 15471 11551 15497 11577
rect 16199 11551 16225 11577
rect 16983 11551 17009 11577
rect 17991 11551 18017 11577
rect 18551 11551 18577 11577
rect 19335 11551 19361 11577
rect 20959 11551 20985 11577
rect 21239 11551 21265 11577
rect 21463 11551 21489 11577
rect 22527 11551 22553 11577
rect 23311 11551 23337 11577
rect 24767 11551 24793 11577
rect 25327 11551 25353 11577
rect 25439 11551 25465 11577
rect 26727 11551 26753 11577
rect 26951 11551 26977 11577
rect 27399 11551 27425 11577
rect 29023 11551 29049 11577
rect 29919 11551 29945 11577
rect 30479 11551 30505 11577
rect 31375 11551 31401 11577
rect 32775 11551 32801 11577
rect 33895 11551 33921 11577
rect 2074 11355 2100 11381
rect 2136 11355 2162 11381
rect 2198 11355 2224 11381
rect 2260 11355 2286 11381
rect 2322 11355 2348 11381
rect 2384 11355 2410 11381
rect 2446 11355 2472 11381
rect 2508 11355 2534 11381
rect 7074 11355 7100 11381
rect 7136 11355 7162 11381
rect 7198 11355 7224 11381
rect 7260 11355 7286 11381
rect 7322 11355 7348 11381
rect 7384 11355 7410 11381
rect 7446 11355 7472 11381
rect 7508 11355 7534 11381
rect 12074 11355 12100 11381
rect 12136 11355 12162 11381
rect 12198 11355 12224 11381
rect 12260 11355 12286 11381
rect 12322 11355 12348 11381
rect 12384 11355 12410 11381
rect 12446 11355 12472 11381
rect 12508 11355 12534 11381
rect 17074 11355 17100 11381
rect 17136 11355 17162 11381
rect 17198 11355 17224 11381
rect 17260 11355 17286 11381
rect 17322 11355 17348 11381
rect 17384 11355 17410 11381
rect 17446 11355 17472 11381
rect 17508 11355 17534 11381
rect 22074 11355 22100 11381
rect 22136 11355 22162 11381
rect 22198 11355 22224 11381
rect 22260 11355 22286 11381
rect 22322 11355 22348 11381
rect 22384 11355 22410 11381
rect 22446 11355 22472 11381
rect 22508 11355 22534 11381
rect 27074 11355 27100 11381
rect 27136 11355 27162 11381
rect 27198 11355 27224 11381
rect 27260 11355 27286 11381
rect 27322 11355 27348 11381
rect 27384 11355 27410 11381
rect 27446 11355 27472 11381
rect 27508 11355 27534 11381
rect 32074 11355 32100 11381
rect 32136 11355 32162 11381
rect 32198 11355 32224 11381
rect 32260 11355 32286 11381
rect 32322 11355 32348 11381
rect 32384 11355 32410 11381
rect 32446 11355 32472 11381
rect 32508 11355 32534 11381
rect 37074 11355 37100 11381
rect 37136 11355 37162 11381
rect 37198 11355 37224 11381
rect 37260 11355 37286 11381
rect 37322 11355 37348 11381
rect 37384 11355 37410 11381
rect 37446 11355 37472 11381
rect 37508 11355 37534 11381
rect 1583 11159 1609 11185
rect 2479 11159 2505 11185
rect 3823 11159 3849 11185
rect 4999 11159 5025 11185
rect 5559 11159 5585 11185
rect 6399 11159 6425 11185
rect 8079 11159 8105 11185
rect 8975 11159 9001 11185
rect 9479 11159 9505 11185
rect 10375 11159 10401 11185
rect 11775 11159 11801 11185
rect 12951 11159 12977 11185
rect 13511 11159 13537 11185
rect 14407 11159 14433 11185
rect 15695 11159 15721 11185
rect 16199 11159 16225 11185
rect 16311 11159 16337 11185
rect 17095 11159 17121 11185
rect 17991 11159 18017 11185
rect 18775 11159 18801 11185
rect 19335 11159 19361 11185
rect 19503 11159 19529 11185
rect 20511 11159 20537 11185
rect 21015 11159 21041 11185
rect 22751 11159 22777 11185
rect 23311 11159 23337 11185
rect 23423 11159 23449 11185
rect 24375 11159 24401 11185
rect 25159 11159 25185 11185
rect 27231 11159 27257 11185
rect 27455 11159 27481 11185
rect 27847 11159 27873 11185
rect 28463 11159 28489 11185
rect 28631 11159 28657 11185
rect 28855 11159 28881 11185
rect 30703 11159 30729 11185
rect 31263 11159 31289 11185
rect 31375 11159 31401 11185
rect 32439 11159 32465 11185
rect 33111 11159 33137 11185
rect 34959 11159 34985 11185
rect 35239 11159 35265 11185
rect 35855 11159 35881 11185
rect 36191 11159 36217 11185
rect 36695 11159 36721 11185
rect 36807 11159 36833 11185
rect 2479 11103 2505 11129
rect 4999 11103 5025 11129
rect 6399 11103 6425 11129
rect 8975 11103 9001 11129
rect 10375 11103 10401 11129
rect 12951 11103 12977 11129
rect 14407 11103 14433 11129
rect 18047 11103 18073 11129
rect 21183 11103 21209 11129
rect 25159 11103 25185 11129
rect 33111 11103 33137 11129
rect 4574 10963 4600 10989
rect 4636 10963 4662 10989
rect 4698 10963 4724 10989
rect 4760 10963 4786 10989
rect 4822 10963 4848 10989
rect 4884 10963 4910 10989
rect 4946 10963 4972 10989
rect 5008 10963 5034 10989
rect 9574 10963 9600 10989
rect 9636 10963 9662 10989
rect 9698 10963 9724 10989
rect 9760 10963 9786 10989
rect 9822 10963 9848 10989
rect 9884 10963 9910 10989
rect 9946 10963 9972 10989
rect 10008 10963 10034 10989
rect 14574 10963 14600 10989
rect 14636 10963 14662 10989
rect 14698 10963 14724 10989
rect 14760 10963 14786 10989
rect 14822 10963 14848 10989
rect 14884 10963 14910 10989
rect 14946 10963 14972 10989
rect 15008 10963 15034 10989
rect 19574 10963 19600 10989
rect 19636 10963 19662 10989
rect 19698 10963 19724 10989
rect 19760 10963 19786 10989
rect 19822 10963 19848 10989
rect 19884 10963 19910 10989
rect 19946 10963 19972 10989
rect 20008 10963 20034 10989
rect 24574 10963 24600 10989
rect 24636 10963 24662 10989
rect 24698 10963 24724 10989
rect 24760 10963 24786 10989
rect 24822 10963 24848 10989
rect 24884 10963 24910 10989
rect 24946 10963 24972 10989
rect 25008 10963 25034 10989
rect 29574 10963 29600 10989
rect 29636 10963 29662 10989
rect 29698 10963 29724 10989
rect 29760 10963 29786 10989
rect 29822 10963 29848 10989
rect 29884 10963 29910 10989
rect 29946 10963 29972 10989
rect 30008 10963 30034 10989
rect 34574 10963 34600 10989
rect 34636 10963 34662 10989
rect 34698 10963 34724 10989
rect 34760 10963 34786 10989
rect 34822 10963 34848 10989
rect 34884 10963 34910 10989
rect 34946 10963 34972 10989
rect 35008 10963 35034 10989
rect 3039 10823 3065 10849
rect 4495 10823 4521 10849
rect 8303 10823 8329 10849
rect 16199 10823 16225 10849
rect 17991 10823 18017 10849
rect 19447 10823 19473 10849
rect 21743 10823 21769 10849
rect 23367 10823 23393 10849
rect 25943 10823 25969 10849
rect 27287 10823 27313 10849
rect 29919 10823 29945 10849
rect 31151 10823 31177 10849
rect 33895 10823 33921 10849
rect 35351 10823 35377 10849
rect 1919 10767 1945 10793
rect 3039 10767 3065 10793
rect 3599 10767 3625 10793
rect 4495 10767 4521 10793
rect 5839 10767 5865 10793
rect 6399 10767 6425 10793
rect 6511 10767 6537 10793
rect 7575 10767 7601 10793
rect 8303 10767 8329 10793
rect 9815 10767 9841 10793
rect 10375 10767 10401 10793
rect 10487 10767 10513 10793
rect 11327 10767 11353 10793
rect 11831 10767 11857 10793
rect 11999 10767 12025 10793
rect 14071 10767 14097 10793
rect 14351 10767 14377 10793
rect 14463 10767 14489 10793
rect 15471 10767 15497 10793
rect 16143 10767 16169 10793
rect 16983 10767 17009 10793
rect 17991 10767 18017 10793
rect 18551 10767 18577 10793
rect 19447 10767 19473 10793
rect 20791 10767 20817 10793
rect 21743 10767 21769 10793
rect 22527 10767 22553 10793
rect 23367 10767 23393 10793
rect 24767 10767 24793 10793
rect 25943 10767 25969 10793
rect 26223 10767 26249 10793
rect 27287 10767 27313 10793
rect 29023 10767 29049 10793
rect 29919 10767 29945 10793
rect 30255 10767 30281 10793
rect 31095 10767 31121 10793
rect 32999 10767 33025 10793
rect 33895 10767 33921 10793
rect 34231 10767 34257 10793
rect 35351 10767 35377 10793
rect 2074 10571 2100 10597
rect 2136 10571 2162 10597
rect 2198 10571 2224 10597
rect 2260 10571 2286 10597
rect 2322 10571 2348 10597
rect 2384 10571 2410 10597
rect 2446 10571 2472 10597
rect 2508 10571 2534 10597
rect 7074 10571 7100 10597
rect 7136 10571 7162 10597
rect 7198 10571 7224 10597
rect 7260 10571 7286 10597
rect 7322 10571 7348 10597
rect 7384 10571 7410 10597
rect 7446 10571 7472 10597
rect 7508 10571 7534 10597
rect 12074 10571 12100 10597
rect 12136 10571 12162 10597
rect 12198 10571 12224 10597
rect 12260 10571 12286 10597
rect 12322 10571 12348 10597
rect 12384 10571 12410 10597
rect 12446 10571 12472 10597
rect 12508 10571 12534 10597
rect 17074 10571 17100 10597
rect 17136 10571 17162 10597
rect 17198 10571 17224 10597
rect 17260 10571 17286 10597
rect 17322 10571 17348 10597
rect 17384 10571 17410 10597
rect 17446 10571 17472 10597
rect 17508 10571 17534 10597
rect 22074 10571 22100 10597
rect 22136 10571 22162 10597
rect 22198 10571 22224 10597
rect 22260 10571 22286 10597
rect 22322 10571 22348 10597
rect 22384 10571 22410 10597
rect 22446 10571 22472 10597
rect 22508 10571 22534 10597
rect 27074 10571 27100 10597
rect 27136 10571 27162 10597
rect 27198 10571 27224 10597
rect 27260 10571 27286 10597
rect 27322 10571 27348 10597
rect 27384 10571 27410 10597
rect 27446 10571 27472 10597
rect 27508 10571 27534 10597
rect 32074 10571 32100 10597
rect 32136 10571 32162 10597
rect 32198 10571 32224 10597
rect 32260 10571 32286 10597
rect 32322 10571 32348 10597
rect 32384 10571 32410 10597
rect 32446 10571 32472 10597
rect 32508 10571 32534 10597
rect 37074 10571 37100 10597
rect 37136 10571 37162 10597
rect 37198 10571 37224 10597
rect 37260 10571 37286 10597
rect 37322 10571 37348 10597
rect 37384 10571 37410 10597
rect 37446 10571 37472 10597
rect 37508 10571 37534 10597
rect 1583 10375 1609 10401
rect 2479 10375 2505 10401
rect 3823 10375 3849 10401
rect 4999 10375 5025 10401
rect 5559 10375 5585 10401
rect 6455 10375 6481 10401
rect 7799 10375 7825 10401
rect 8303 10375 8329 10401
rect 8471 10375 8497 10401
rect 9479 10375 9505 10401
rect 10375 10375 10401 10401
rect 11887 10375 11913 10401
rect 12951 10375 12977 10401
rect 13511 10375 13537 10401
rect 14407 10375 14433 10401
rect 15695 10375 15721 10401
rect 16143 10375 16169 10401
rect 16367 10375 16393 10401
rect 17151 10375 17177 10401
rect 17991 10375 18017 10401
rect 18775 10375 18801 10401
rect 19951 10375 19977 10401
rect 20231 10375 20257 10401
rect 21407 10375 21433 10401
rect 22751 10375 22777 10401
rect 23703 10375 23729 10401
rect 24487 10375 24513 10401
rect 25383 10375 25409 10401
rect 26727 10375 26753 10401
rect 27567 10375 27593 10401
rect 28183 10375 28209 10401
rect 29135 10375 29161 10401
rect 30703 10375 30729 10401
rect 31655 10375 31681 10401
rect 32159 10375 32185 10401
rect 33111 10375 33137 10401
rect 34679 10375 34705 10401
rect 35631 10375 35657 10401
rect 36135 10375 36161 10401
rect 36695 10375 36721 10401
rect 36863 10375 36889 10401
rect 2479 10319 2505 10345
rect 4999 10319 5025 10345
rect 6455 10319 6481 10345
rect 10375 10319 10401 10345
rect 12951 10319 12977 10345
rect 14407 10319 14433 10345
rect 18103 10319 18129 10345
rect 19951 10319 19977 10345
rect 21407 10319 21433 10345
rect 23703 10319 23729 10345
rect 25383 10319 25409 10345
rect 27679 10319 27705 10345
rect 29135 10319 29161 10345
rect 31655 10319 31681 10345
rect 33111 10319 33137 10345
rect 35631 10319 35657 10345
rect 4574 10179 4600 10205
rect 4636 10179 4662 10205
rect 4698 10179 4724 10205
rect 4760 10179 4786 10205
rect 4822 10179 4848 10205
rect 4884 10179 4910 10205
rect 4946 10179 4972 10205
rect 5008 10179 5034 10205
rect 9574 10179 9600 10205
rect 9636 10179 9662 10205
rect 9698 10179 9724 10205
rect 9760 10179 9786 10205
rect 9822 10179 9848 10205
rect 9884 10179 9910 10205
rect 9946 10179 9972 10205
rect 10008 10179 10034 10205
rect 14574 10179 14600 10205
rect 14636 10179 14662 10205
rect 14698 10179 14724 10205
rect 14760 10179 14786 10205
rect 14822 10179 14848 10205
rect 14884 10179 14910 10205
rect 14946 10179 14972 10205
rect 15008 10179 15034 10205
rect 19574 10179 19600 10205
rect 19636 10179 19662 10205
rect 19698 10179 19724 10205
rect 19760 10179 19786 10205
rect 19822 10179 19848 10205
rect 19884 10179 19910 10205
rect 19946 10179 19972 10205
rect 20008 10179 20034 10205
rect 24574 10179 24600 10205
rect 24636 10179 24662 10205
rect 24698 10179 24724 10205
rect 24760 10179 24786 10205
rect 24822 10179 24848 10205
rect 24884 10179 24910 10205
rect 24946 10179 24972 10205
rect 25008 10179 25034 10205
rect 29574 10179 29600 10205
rect 29636 10179 29662 10205
rect 29698 10179 29724 10205
rect 29760 10179 29786 10205
rect 29822 10179 29848 10205
rect 29884 10179 29910 10205
rect 29946 10179 29972 10205
rect 30008 10179 30034 10205
rect 34574 10179 34600 10205
rect 34636 10179 34662 10205
rect 34698 10179 34724 10205
rect 34760 10179 34786 10205
rect 34822 10179 34848 10205
rect 34884 10179 34910 10205
rect 34946 10179 34972 10205
rect 35008 10179 35034 10205
rect 3039 10039 3065 10065
rect 4495 10039 4521 10065
rect 7015 10039 7041 10065
rect 8359 10039 8385 10065
rect 12447 10039 12473 10065
rect 17991 10039 18017 10065
rect 21743 10039 21769 10065
rect 25943 10039 25969 10065
rect 31263 10039 31289 10065
rect 33839 10039 33865 10065
rect 35351 10039 35377 10065
rect 37647 10039 37673 10065
rect 1919 9983 1945 10009
rect 3039 9983 3065 10009
rect 3599 9983 3625 10009
rect 4495 9983 4521 10009
rect 5839 9983 5865 10009
rect 7015 9983 7041 10009
rect 7575 9983 7601 10009
rect 8359 9983 8385 10009
rect 9815 9983 9841 10009
rect 10375 9983 10401 10009
rect 10487 9983 10513 10009
rect 11271 9983 11297 10009
rect 12447 9983 12473 10009
rect 14071 9983 14097 10009
rect 14351 9983 14377 10009
rect 14463 9983 14489 10009
rect 15471 9983 15497 10009
rect 15807 9983 15833 10009
rect 15919 9983 15945 10009
rect 16983 9983 17009 10009
rect 17991 9983 18017 10009
rect 18551 9983 18577 10009
rect 18719 9983 18745 10009
rect 18943 9983 18969 10009
rect 20791 9983 20817 10009
rect 21743 9983 21769 10009
rect 22527 9983 22553 10009
rect 22695 9983 22721 10009
rect 22919 9983 22945 10009
rect 25047 9983 25073 10009
rect 25943 9983 25969 10009
rect 26727 9983 26753 10009
rect 26951 9983 26977 10009
rect 27399 9983 27425 10009
rect 28743 9983 28769 10009
rect 29303 9983 29329 10009
rect 29415 9983 29441 10009
rect 30423 9983 30449 10009
rect 31095 9983 31121 10009
rect 32775 9983 32801 10009
rect 33839 9983 33865 10009
rect 34455 9983 34481 10009
rect 35351 9983 35377 10009
rect 36695 9983 36721 10009
rect 37647 9983 37673 10009
rect 2074 9787 2100 9813
rect 2136 9787 2162 9813
rect 2198 9787 2224 9813
rect 2260 9787 2286 9813
rect 2322 9787 2348 9813
rect 2384 9787 2410 9813
rect 2446 9787 2472 9813
rect 2508 9787 2534 9813
rect 7074 9787 7100 9813
rect 7136 9787 7162 9813
rect 7198 9787 7224 9813
rect 7260 9787 7286 9813
rect 7322 9787 7348 9813
rect 7384 9787 7410 9813
rect 7446 9787 7472 9813
rect 7508 9787 7534 9813
rect 12074 9787 12100 9813
rect 12136 9787 12162 9813
rect 12198 9787 12224 9813
rect 12260 9787 12286 9813
rect 12322 9787 12348 9813
rect 12384 9787 12410 9813
rect 12446 9787 12472 9813
rect 12508 9787 12534 9813
rect 17074 9787 17100 9813
rect 17136 9787 17162 9813
rect 17198 9787 17224 9813
rect 17260 9787 17286 9813
rect 17322 9787 17348 9813
rect 17384 9787 17410 9813
rect 17446 9787 17472 9813
rect 17508 9787 17534 9813
rect 22074 9787 22100 9813
rect 22136 9787 22162 9813
rect 22198 9787 22224 9813
rect 22260 9787 22286 9813
rect 22322 9787 22348 9813
rect 22384 9787 22410 9813
rect 22446 9787 22472 9813
rect 22508 9787 22534 9813
rect 27074 9787 27100 9813
rect 27136 9787 27162 9813
rect 27198 9787 27224 9813
rect 27260 9787 27286 9813
rect 27322 9787 27348 9813
rect 27384 9787 27410 9813
rect 27446 9787 27472 9813
rect 27508 9787 27534 9813
rect 32074 9787 32100 9813
rect 32136 9787 32162 9813
rect 32198 9787 32224 9813
rect 32260 9787 32286 9813
rect 32322 9787 32348 9813
rect 32384 9787 32410 9813
rect 32446 9787 32472 9813
rect 32508 9787 32534 9813
rect 37074 9787 37100 9813
rect 37136 9787 37162 9813
rect 37198 9787 37224 9813
rect 37260 9787 37286 9813
rect 37322 9787 37348 9813
rect 37384 9787 37410 9813
rect 37446 9787 37472 9813
rect 37508 9787 37534 9813
rect 1583 9591 1609 9617
rect 2479 9591 2505 9617
rect 3935 9591 3961 9617
rect 4999 9591 5025 9617
rect 5559 9591 5585 9617
rect 6455 9591 6481 9617
rect 7799 9591 7825 9617
rect 8359 9591 8385 9617
rect 8471 9591 8497 9617
rect 9479 9591 9505 9617
rect 10431 9591 10457 9617
rect 12055 9591 12081 9617
rect 12951 9591 12977 9617
rect 13511 9591 13537 9617
rect 14407 9591 14433 9617
rect 15527 9591 15553 9617
rect 15975 9591 16001 9617
rect 16199 9591 16225 9617
rect 17095 9591 17121 9617
rect 18271 9591 18297 9617
rect 18775 9591 18801 9617
rect 19223 9591 19249 9617
rect 19447 9591 19473 9617
rect 20231 9591 20257 9617
rect 21295 9591 21321 9617
rect 22751 9591 22777 9617
rect 23311 9591 23337 9617
rect 23423 9591 23449 9617
rect 24375 9591 24401 9617
rect 24655 9591 24681 9617
rect 24879 9591 24905 9617
rect 27231 9591 27257 9617
rect 27455 9591 27481 9617
rect 27903 9591 27929 9617
rect 28463 9591 28489 9617
rect 28743 9591 28769 9617
rect 28967 9591 28993 9617
rect 30983 9591 31009 9617
rect 31151 9591 31177 9617
rect 31375 9591 31401 9617
rect 32439 9591 32465 9617
rect 32831 9591 32857 9617
rect 34959 9591 34985 9617
rect 35855 9591 35881 9617
rect 36135 9591 36161 9617
rect 37311 9591 37337 9617
rect 2479 9535 2505 9561
rect 4999 9535 5025 9561
rect 6455 9535 6481 9561
rect 10431 9535 10457 9561
rect 12951 9535 12977 9561
rect 14407 9535 14433 9561
rect 18271 9535 18297 9561
rect 21295 9535 21321 9561
rect 33111 9535 33137 9561
rect 35855 9535 35881 9561
rect 37311 9535 37337 9561
rect 4574 9395 4600 9421
rect 4636 9395 4662 9421
rect 4698 9395 4724 9421
rect 4760 9395 4786 9421
rect 4822 9395 4848 9421
rect 4884 9395 4910 9421
rect 4946 9395 4972 9421
rect 5008 9395 5034 9421
rect 9574 9395 9600 9421
rect 9636 9395 9662 9421
rect 9698 9395 9724 9421
rect 9760 9395 9786 9421
rect 9822 9395 9848 9421
rect 9884 9395 9910 9421
rect 9946 9395 9972 9421
rect 10008 9395 10034 9421
rect 14574 9395 14600 9421
rect 14636 9395 14662 9421
rect 14698 9395 14724 9421
rect 14760 9395 14786 9421
rect 14822 9395 14848 9421
rect 14884 9395 14910 9421
rect 14946 9395 14972 9421
rect 15008 9395 15034 9421
rect 19574 9395 19600 9421
rect 19636 9395 19662 9421
rect 19698 9395 19724 9421
rect 19760 9395 19786 9421
rect 19822 9395 19848 9421
rect 19884 9395 19910 9421
rect 19946 9395 19972 9421
rect 20008 9395 20034 9421
rect 24574 9395 24600 9421
rect 24636 9395 24662 9421
rect 24698 9395 24724 9421
rect 24760 9395 24786 9421
rect 24822 9395 24848 9421
rect 24884 9395 24910 9421
rect 24946 9395 24972 9421
rect 25008 9395 25034 9421
rect 29574 9395 29600 9421
rect 29636 9395 29662 9421
rect 29698 9395 29724 9421
rect 29760 9395 29786 9421
rect 29822 9395 29848 9421
rect 29884 9395 29910 9421
rect 29946 9395 29972 9421
rect 30008 9395 30034 9421
rect 34574 9395 34600 9421
rect 34636 9395 34662 9421
rect 34698 9395 34724 9421
rect 34760 9395 34786 9421
rect 34822 9395 34848 9421
rect 34884 9395 34910 9421
rect 34946 9395 34972 9421
rect 35008 9395 35034 9421
rect 3039 9255 3065 9281
rect 4271 9255 4297 9281
rect 7015 9255 7041 9281
rect 8359 9255 8385 9281
rect 10879 9255 10905 9281
rect 18271 9255 18297 9281
rect 23423 9255 23449 9281
rect 27399 9255 27425 9281
rect 29695 9255 29721 9281
rect 31375 9255 31401 9281
rect 37647 9255 37673 9281
rect 1919 9199 1945 9225
rect 3039 9199 3065 9225
rect 3599 9199 3625 9225
rect 4271 9199 4297 9225
rect 5839 9199 5865 9225
rect 7015 9199 7041 9225
rect 7575 9199 7601 9225
rect 8359 9199 8385 9225
rect 9815 9199 9841 9225
rect 10879 9199 10905 9225
rect 11551 9199 11577 9225
rect 11775 9199 11801 9225
rect 11943 9199 11969 9225
rect 14071 9199 14097 9225
rect 14351 9199 14377 9225
rect 14463 9199 14489 9225
rect 15247 9199 15273 9225
rect 15807 9199 15833 9225
rect 15919 9199 15945 9225
rect 17207 9199 17233 9225
rect 18271 9199 18297 9225
rect 18775 9199 18801 9225
rect 19223 9199 19249 9225
rect 19335 9199 19361 9225
rect 20791 9199 20817 9225
rect 21295 9199 21321 9225
rect 21463 9199 21489 9225
rect 22527 9199 22553 9225
rect 23423 9199 23449 9225
rect 24767 9199 24793 9225
rect 25215 9199 25241 9225
rect 25439 9199 25465 9225
rect 26503 9199 26529 9225
rect 27399 9199 27425 9225
rect 29023 9199 29049 9225
rect 29415 9199 29441 9225
rect 30423 9199 30449 9225
rect 31375 9199 31401 9225
rect 32943 9199 32969 9225
rect 33167 9199 33193 9225
rect 33391 9199 33417 9225
rect 34175 9199 34201 9225
rect 34623 9199 34649 9225
rect 34847 9199 34873 9225
rect 36695 9199 36721 9225
rect 37591 9199 37617 9225
rect 2074 9003 2100 9029
rect 2136 9003 2162 9029
rect 2198 9003 2224 9029
rect 2260 9003 2286 9029
rect 2322 9003 2348 9029
rect 2384 9003 2410 9029
rect 2446 9003 2472 9029
rect 2508 9003 2534 9029
rect 7074 9003 7100 9029
rect 7136 9003 7162 9029
rect 7198 9003 7224 9029
rect 7260 9003 7286 9029
rect 7322 9003 7348 9029
rect 7384 9003 7410 9029
rect 7446 9003 7472 9029
rect 7508 9003 7534 9029
rect 12074 9003 12100 9029
rect 12136 9003 12162 9029
rect 12198 9003 12224 9029
rect 12260 9003 12286 9029
rect 12322 9003 12348 9029
rect 12384 9003 12410 9029
rect 12446 9003 12472 9029
rect 12508 9003 12534 9029
rect 17074 9003 17100 9029
rect 17136 9003 17162 9029
rect 17198 9003 17224 9029
rect 17260 9003 17286 9029
rect 17322 9003 17348 9029
rect 17384 9003 17410 9029
rect 17446 9003 17472 9029
rect 17508 9003 17534 9029
rect 22074 9003 22100 9029
rect 22136 9003 22162 9029
rect 22198 9003 22224 9029
rect 22260 9003 22286 9029
rect 22322 9003 22348 9029
rect 22384 9003 22410 9029
rect 22446 9003 22472 9029
rect 22508 9003 22534 9029
rect 27074 9003 27100 9029
rect 27136 9003 27162 9029
rect 27198 9003 27224 9029
rect 27260 9003 27286 9029
rect 27322 9003 27348 9029
rect 27384 9003 27410 9029
rect 27446 9003 27472 9029
rect 27508 9003 27534 9029
rect 32074 9003 32100 9029
rect 32136 9003 32162 9029
rect 32198 9003 32224 9029
rect 32260 9003 32286 9029
rect 32322 9003 32348 9029
rect 32384 9003 32410 9029
rect 32446 9003 32472 9029
rect 32508 9003 32534 9029
rect 37074 9003 37100 9029
rect 37136 9003 37162 9029
rect 37198 9003 37224 9029
rect 37260 9003 37286 9029
rect 37322 9003 37348 9029
rect 37384 9003 37410 9029
rect 37446 9003 37472 9029
rect 37508 9003 37534 9029
rect 1583 8807 1609 8833
rect 1751 8807 1777 8833
rect 1975 8807 2001 8833
rect 3935 8807 3961 8833
rect 4271 8807 4297 8833
rect 4495 8807 4521 8833
rect 5559 8807 5585 8833
rect 5951 8807 5977 8833
rect 7799 8807 7825 8833
rect 8359 8807 8385 8833
rect 8471 8807 8497 8833
rect 9255 8807 9281 8833
rect 10263 8807 10289 8833
rect 11999 8807 12025 8833
rect 12223 8807 12249 8833
rect 12447 8807 12473 8833
rect 13511 8807 13537 8833
rect 14407 8807 14433 8833
rect 15471 8807 15497 8833
rect 15919 8807 15945 8833
rect 16143 8807 16169 8833
rect 17207 8807 17233 8833
rect 18271 8807 18297 8833
rect 18775 8807 18801 8833
rect 19335 8807 19361 8833
rect 19503 8807 19529 8833
rect 20231 8807 20257 8833
rect 21295 8807 21321 8833
rect 22751 8807 22777 8833
rect 23311 8807 23337 8833
rect 23423 8807 23449 8833
rect 24375 8807 24401 8833
rect 25215 8807 25241 8833
rect 26727 8807 26753 8833
rect 27287 8807 27313 8833
rect 27511 8807 27537 8833
rect 28463 8807 28489 8833
rect 29359 8807 29385 8833
rect 30983 8807 31009 8833
rect 31879 8807 31905 8833
rect 32159 8807 32185 8833
rect 32719 8807 32745 8833
rect 32831 8807 32857 8833
rect 34959 8807 34985 8833
rect 35855 8807 35881 8833
rect 36359 8807 36385 8833
rect 37311 8807 37337 8833
rect 6231 8751 6257 8777
rect 10263 8751 10289 8777
rect 14407 8751 14433 8777
rect 18271 8751 18297 8777
rect 21295 8751 21321 8777
rect 25159 8751 25185 8777
rect 29359 8751 29385 8777
rect 31879 8751 31905 8777
rect 35855 8751 35881 8777
rect 37311 8751 37337 8777
rect 4574 8611 4600 8637
rect 4636 8611 4662 8637
rect 4698 8611 4724 8637
rect 4760 8611 4786 8637
rect 4822 8611 4848 8637
rect 4884 8611 4910 8637
rect 4946 8611 4972 8637
rect 5008 8611 5034 8637
rect 9574 8611 9600 8637
rect 9636 8611 9662 8637
rect 9698 8611 9724 8637
rect 9760 8611 9786 8637
rect 9822 8611 9848 8637
rect 9884 8611 9910 8637
rect 9946 8611 9972 8637
rect 10008 8611 10034 8637
rect 14574 8611 14600 8637
rect 14636 8611 14662 8637
rect 14698 8611 14724 8637
rect 14760 8611 14786 8637
rect 14822 8611 14848 8637
rect 14884 8611 14910 8637
rect 14946 8611 14972 8637
rect 15008 8611 15034 8637
rect 19574 8611 19600 8637
rect 19636 8611 19662 8637
rect 19698 8611 19724 8637
rect 19760 8611 19786 8637
rect 19822 8611 19848 8637
rect 19884 8611 19910 8637
rect 19946 8611 19972 8637
rect 20008 8611 20034 8637
rect 24574 8611 24600 8637
rect 24636 8611 24662 8637
rect 24698 8611 24724 8637
rect 24760 8611 24786 8637
rect 24822 8611 24848 8637
rect 24884 8611 24910 8637
rect 24946 8611 24972 8637
rect 25008 8611 25034 8637
rect 29574 8611 29600 8637
rect 29636 8611 29662 8637
rect 29698 8611 29724 8637
rect 29760 8611 29786 8637
rect 29822 8611 29848 8637
rect 29884 8611 29910 8637
rect 29946 8611 29972 8637
rect 30008 8611 30034 8637
rect 34574 8611 34600 8637
rect 34636 8611 34662 8637
rect 34698 8611 34724 8637
rect 34760 8611 34786 8637
rect 34822 8611 34848 8637
rect 34884 8611 34910 8637
rect 34946 8611 34972 8637
rect 35008 8611 35034 8637
rect 4271 8471 4297 8497
rect 8359 8471 8385 8497
rect 14967 8471 14993 8497
rect 18271 8471 18297 8497
rect 19503 8471 19529 8497
rect 23423 8471 23449 8497
rect 27175 8471 27201 8497
rect 29919 8471 29945 8497
rect 31151 8471 31177 8497
rect 33895 8471 33921 8497
rect 35127 8471 35153 8497
rect 37647 8471 37673 8497
rect 2143 8415 2169 8441
rect 2311 8415 2337 8441
rect 2535 8415 2561 8441
rect 3599 8415 3625 8441
rect 4215 8415 4241 8441
rect 5839 8415 5865 8441
rect 6287 8415 6313 8441
rect 6511 8415 6537 8441
rect 7575 8415 7601 8441
rect 8359 8415 8385 8441
rect 9815 8415 9841 8441
rect 10263 8415 10289 8441
rect 10487 8415 10513 8441
rect 11551 8415 11577 8441
rect 11775 8415 11801 8441
rect 11943 8415 11969 8441
rect 14071 8415 14097 8441
rect 14967 8415 14993 8441
rect 15247 8415 15273 8441
rect 15695 8415 15721 8441
rect 15919 8415 15945 8441
rect 17095 8415 17121 8441
rect 18271 8415 18297 8441
rect 18775 8415 18801 8441
rect 19335 8415 19361 8441
rect 20791 8415 20817 8441
rect 21295 8415 21321 8441
rect 21463 8415 21489 8441
rect 22527 8415 22553 8441
rect 23423 8415 23449 8441
rect 24767 8415 24793 8441
rect 25215 8415 25241 8441
rect 25439 8415 25465 8441
rect 26223 8415 26249 8441
rect 26895 8415 26921 8441
rect 29023 8415 29049 8441
rect 29919 8415 29945 8441
rect 30479 8415 30505 8441
rect 31151 8415 31177 8441
rect 32047 8415 32073 8441
rect 32215 8415 32241 8441
rect 32327 8415 32353 8441
rect 32887 8415 32913 8441
rect 33895 8415 33921 8441
rect 34399 8415 34425 8441
rect 35071 8415 35097 8441
rect 36695 8415 36721 8441
rect 37647 8415 37673 8441
rect 2074 8219 2100 8245
rect 2136 8219 2162 8245
rect 2198 8219 2224 8245
rect 2260 8219 2286 8245
rect 2322 8219 2348 8245
rect 2384 8219 2410 8245
rect 2446 8219 2472 8245
rect 2508 8219 2534 8245
rect 7074 8219 7100 8245
rect 7136 8219 7162 8245
rect 7198 8219 7224 8245
rect 7260 8219 7286 8245
rect 7322 8219 7348 8245
rect 7384 8219 7410 8245
rect 7446 8219 7472 8245
rect 7508 8219 7534 8245
rect 12074 8219 12100 8245
rect 12136 8219 12162 8245
rect 12198 8219 12224 8245
rect 12260 8219 12286 8245
rect 12322 8219 12348 8245
rect 12384 8219 12410 8245
rect 12446 8219 12472 8245
rect 12508 8219 12534 8245
rect 17074 8219 17100 8245
rect 17136 8219 17162 8245
rect 17198 8219 17224 8245
rect 17260 8219 17286 8245
rect 17322 8219 17348 8245
rect 17384 8219 17410 8245
rect 17446 8219 17472 8245
rect 17508 8219 17534 8245
rect 22074 8219 22100 8245
rect 22136 8219 22162 8245
rect 22198 8219 22224 8245
rect 22260 8219 22286 8245
rect 22322 8219 22348 8245
rect 22384 8219 22410 8245
rect 22446 8219 22472 8245
rect 22508 8219 22534 8245
rect 27074 8219 27100 8245
rect 27136 8219 27162 8245
rect 27198 8219 27224 8245
rect 27260 8219 27286 8245
rect 27322 8219 27348 8245
rect 27384 8219 27410 8245
rect 27446 8219 27472 8245
rect 27508 8219 27534 8245
rect 32074 8219 32100 8245
rect 32136 8219 32162 8245
rect 32198 8219 32224 8245
rect 32260 8219 32286 8245
rect 32322 8219 32348 8245
rect 32384 8219 32410 8245
rect 32446 8219 32472 8245
rect 32508 8219 32534 8245
rect 37074 8219 37100 8245
rect 37136 8219 37162 8245
rect 37198 8219 37224 8245
rect 37260 8219 37286 8245
rect 37322 8219 37348 8245
rect 37384 8219 37410 8245
rect 37446 8219 37472 8245
rect 37508 8219 37534 8245
rect 1583 8023 1609 8049
rect 1975 8023 2001 8049
rect 3935 8023 3961 8049
rect 4271 8023 4297 8049
rect 4495 8023 4521 8049
rect 5559 8023 5585 8049
rect 6231 8023 6257 8049
rect 7799 8023 7825 8049
rect 8359 8023 8385 8049
rect 8471 8023 8497 8049
rect 9255 8023 9281 8049
rect 10263 8023 10289 8049
rect 12055 8023 12081 8049
rect 12223 8023 12249 8049
rect 12447 8023 12473 8049
rect 13399 8023 13425 8049
rect 14183 8023 14209 8049
rect 15303 8023 15329 8049
rect 16423 8023 16449 8049
rect 16871 8023 16897 8049
rect 17711 8023 17737 8049
rect 18775 8023 18801 8049
rect 19335 8023 19361 8049
rect 19447 8023 19473 8049
rect 20231 8023 20257 8049
rect 21295 8023 21321 8049
rect 22751 8023 22777 8049
rect 23311 8023 23337 8049
rect 23423 8023 23449 8049
rect 24375 8023 24401 8049
rect 24767 8023 24793 8049
rect 24879 8023 24905 8049
rect 26727 8023 26753 8049
rect 27175 8023 27201 8049
rect 27399 8023 27425 8049
rect 28463 8023 28489 8049
rect 29359 8023 29385 8049
rect 30983 8023 31009 8049
rect 31151 8023 31177 8049
rect 31375 8023 31401 8049
rect 32439 8023 32465 8049
rect 33335 8023 33361 8049
rect 33727 8023 33753 8049
rect 34959 8023 34985 8049
rect 35855 8023 35881 8049
rect 36415 8023 36441 8049
rect 37311 8023 37337 8049
rect 2255 7967 2281 7993
rect 6231 7967 6257 7993
rect 10263 7967 10289 7993
rect 14183 7967 14209 7993
rect 16423 7967 16449 7993
rect 17711 7967 17737 7993
rect 21295 7967 21321 7993
rect 29359 7967 29385 7993
rect 33335 7967 33361 7993
rect 33615 7967 33641 7993
rect 33895 7967 33921 7993
rect 35855 7967 35881 7993
rect 37311 7967 37337 7993
rect 4574 7827 4600 7853
rect 4636 7827 4662 7853
rect 4698 7827 4724 7853
rect 4760 7827 4786 7853
rect 4822 7827 4848 7853
rect 4884 7827 4910 7853
rect 4946 7827 4972 7853
rect 5008 7827 5034 7853
rect 9574 7827 9600 7853
rect 9636 7827 9662 7853
rect 9698 7827 9724 7853
rect 9760 7827 9786 7853
rect 9822 7827 9848 7853
rect 9884 7827 9910 7853
rect 9946 7827 9972 7853
rect 10008 7827 10034 7853
rect 14574 7827 14600 7853
rect 14636 7827 14662 7853
rect 14698 7827 14724 7853
rect 14760 7827 14786 7853
rect 14822 7827 14848 7853
rect 14884 7827 14910 7853
rect 14946 7827 14972 7853
rect 15008 7827 15034 7853
rect 19574 7827 19600 7853
rect 19636 7827 19662 7853
rect 19698 7827 19724 7853
rect 19760 7827 19786 7853
rect 19822 7827 19848 7853
rect 19884 7827 19910 7853
rect 19946 7827 19972 7853
rect 20008 7827 20034 7853
rect 24574 7827 24600 7853
rect 24636 7827 24662 7853
rect 24698 7827 24724 7853
rect 24760 7827 24786 7853
rect 24822 7827 24848 7853
rect 24884 7827 24910 7853
rect 24946 7827 24972 7853
rect 25008 7827 25034 7853
rect 29574 7827 29600 7853
rect 29636 7827 29662 7853
rect 29698 7827 29724 7853
rect 29760 7827 29786 7853
rect 29822 7827 29848 7853
rect 29884 7827 29910 7853
rect 29946 7827 29972 7853
rect 30008 7827 30034 7853
rect 34574 7827 34600 7853
rect 34636 7827 34662 7853
rect 34698 7827 34724 7853
rect 34760 7827 34786 7853
rect 34822 7827 34848 7853
rect 34884 7827 34910 7853
rect 34946 7827 34972 7853
rect 35008 7827 35034 7853
rect 3039 7687 3065 7713
rect 4271 7687 4297 7713
rect 14967 7687 14993 7713
rect 16423 7687 16449 7713
rect 17767 7687 17793 7713
rect 19335 7687 19361 7713
rect 23423 7687 23449 7713
rect 31375 7687 31401 7713
rect 33839 7687 33865 7713
rect 35239 7687 35265 7713
rect 37647 7687 37673 7713
rect 1863 7631 1889 7657
rect 3039 7631 3065 7657
rect 3599 7631 3625 7657
rect 4215 7631 4241 7657
rect 5839 7631 5865 7657
rect 6287 7631 6313 7657
rect 6511 7631 6537 7657
rect 7575 7631 7601 7657
rect 7743 7631 7769 7657
rect 7967 7631 7993 7657
rect 9815 7631 9841 7657
rect 10263 7631 10289 7657
rect 10487 7631 10513 7657
rect 11271 7631 11297 7657
rect 11775 7631 11801 7657
rect 11943 7631 11969 7657
rect 14071 7631 14097 7657
rect 14967 7631 14993 7657
rect 15247 7631 15273 7657
rect 16423 7631 16449 7657
rect 16871 7631 16897 7657
rect 17711 7631 17737 7657
rect 18551 7631 18577 7657
rect 19335 7631 19361 7657
rect 20791 7631 20817 7657
rect 21295 7631 21321 7657
rect 21463 7631 21489 7657
rect 22527 7631 22553 7657
rect 23423 7631 23449 7657
rect 24767 7631 24793 7657
rect 25215 7631 25241 7657
rect 25439 7631 25465 7657
rect 26223 7631 26249 7657
rect 26783 7631 26809 7657
rect 26895 7631 26921 7657
rect 29023 7631 29049 7657
rect 29303 7631 29329 7657
rect 29471 7631 29497 7657
rect 30479 7631 30505 7657
rect 31375 7631 31401 7657
rect 32103 7631 32129 7657
rect 32159 7631 32185 7657
rect 32327 7631 32353 7657
rect 32943 7631 32969 7657
rect 33839 7631 33865 7657
rect 34399 7631 34425 7657
rect 35239 7631 35265 7657
rect 36695 7631 36721 7657
rect 37647 7631 37673 7657
rect 2074 7435 2100 7461
rect 2136 7435 2162 7461
rect 2198 7435 2224 7461
rect 2260 7435 2286 7461
rect 2322 7435 2348 7461
rect 2384 7435 2410 7461
rect 2446 7435 2472 7461
rect 2508 7435 2534 7461
rect 7074 7435 7100 7461
rect 7136 7435 7162 7461
rect 7198 7435 7224 7461
rect 7260 7435 7286 7461
rect 7322 7435 7348 7461
rect 7384 7435 7410 7461
rect 7446 7435 7472 7461
rect 7508 7435 7534 7461
rect 12074 7435 12100 7461
rect 12136 7435 12162 7461
rect 12198 7435 12224 7461
rect 12260 7435 12286 7461
rect 12322 7435 12348 7461
rect 12384 7435 12410 7461
rect 12446 7435 12472 7461
rect 12508 7435 12534 7461
rect 17074 7435 17100 7461
rect 17136 7435 17162 7461
rect 17198 7435 17224 7461
rect 17260 7435 17286 7461
rect 17322 7435 17348 7461
rect 17384 7435 17410 7461
rect 17446 7435 17472 7461
rect 17508 7435 17534 7461
rect 22074 7435 22100 7461
rect 22136 7435 22162 7461
rect 22198 7435 22224 7461
rect 22260 7435 22286 7461
rect 22322 7435 22348 7461
rect 22384 7435 22410 7461
rect 22446 7435 22472 7461
rect 22508 7435 22534 7461
rect 27074 7435 27100 7461
rect 27136 7435 27162 7461
rect 27198 7435 27224 7461
rect 27260 7435 27286 7461
rect 27322 7435 27348 7461
rect 27384 7435 27410 7461
rect 27446 7435 27472 7461
rect 27508 7435 27534 7461
rect 32074 7435 32100 7461
rect 32136 7435 32162 7461
rect 32198 7435 32224 7461
rect 32260 7435 32286 7461
rect 32322 7435 32348 7461
rect 32384 7435 32410 7461
rect 32446 7435 32472 7461
rect 32508 7435 32534 7461
rect 37074 7435 37100 7461
rect 37136 7435 37162 7461
rect 37198 7435 37224 7461
rect 37260 7435 37286 7461
rect 37322 7435 37348 7461
rect 37384 7435 37410 7461
rect 37446 7435 37472 7461
rect 37508 7435 37534 7461
rect 1807 7239 1833 7265
rect 2031 7239 2057 7265
rect 2479 7239 2505 7265
rect 4103 7239 4129 7265
rect 4999 7239 5025 7265
rect 5279 7239 5305 7265
rect 6455 7239 6481 7265
rect 8079 7239 8105 7265
rect 8751 7239 8777 7265
rect 9423 7239 9449 7265
rect 10207 7239 10233 7265
rect 11831 7239 11857 7265
rect 12223 7239 12249 7265
rect 12447 7239 12473 7265
rect 13511 7239 13537 7265
rect 14407 7239 14433 7265
rect 15191 7239 15217 7265
rect 15695 7239 15721 7265
rect 15807 7239 15833 7265
rect 16815 7239 16841 7265
rect 17263 7239 17289 7265
rect 17375 7239 17401 7265
rect 18775 7239 18801 7265
rect 19335 7239 19361 7265
rect 19447 7239 19473 7265
rect 20231 7239 20257 7265
rect 21295 7239 21321 7265
rect 22751 7239 22777 7265
rect 23311 7239 23337 7265
rect 23423 7239 23449 7265
rect 24375 7239 24401 7265
rect 25103 7239 25129 7265
rect 26727 7239 26753 7265
rect 27175 7239 27201 7265
rect 27399 7239 27425 7265
rect 28463 7239 28489 7265
rect 29191 7239 29217 7265
rect 30983 7239 31009 7265
rect 31823 7239 31849 7265
rect 32439 7239 32465 7265
rect 33335 7239 33361 7265
rect 33671 7239 33697 7265
rect 33727 7239 33753 7265
rect 34679 7239 34705 7265
rect 35127 7239 35153 7265
rect 35351 7239 35377 7265
rect 36415 7239 36441 7265
rect 37311 7239 37337 7265
rect 4999 7183 5025 7209
rect 6455 7183 6481 7209
rect 8751 7183 8777 7209
rect 10207 7183 10233 7209
rect 14407 7183 14433 7209
rect 21295 7183 21321 7209
rect 25159 7183 25185 7209
rect 29191 7183 29217 7209
rect 31823 7183 31849 7209
rect 33335 7183 33361 7209
rect 33895 7183 33921 7209
rect 37311 7183 37337 7209
rect 4574 7043 4600 7069
rect 4636 7043 4662 7069
rect 4698 7043 4724 7069
rect 4760 7043 4786 7069
rect 4822 7043 4848 7069
rect 4884 7043 4910 7069
rect 4946 7043 4972 7069
rect 5008 7043 5034 7069
rect 9574 7043 9600 7069
rect 9636 7043 9662 7069
rect 9698 7043 9724 7069
rect 9760 7043 9786 7069
rect 9822 7043 9848 7069
rect 9884 7043 9910 7069
rect 9946 7043 9972 7069
rect 10008 7043 10034 7069
rect 14574 7043 14600 7069
rect 14636 7043 14662 7069
rect 14698 7043 14724 7069
rect 14760 7043 14786 7069
rect 14822 7043 14848 7069
rect 14884 7043 14910 7069
rect 14946 7043 14972 7069
rect 15008 7043 15034 7069
rect 19574 7043 19600 7069
rect 19636 7043 19662 7069
rect 19698 7043 19724 7069
rect 19760 7043 19786 7069
rect 19822 7043 19848 7069
rect 19884 7043 19910 7069
rect 19946 7043 19972 7069
rect 20008 7043 20034 7069
rect 24574 7043 24600 7069
rect 24636 7043 24662 7069
rect 24698 7043 24724 7069
rect 24760 7043 24786 7069
rect 24822 7043 24848 7069
rect 24884 7043 24910 7069
rect 24946 7043 24972 7069
rect 25008 7043 25034 7069
rect 29574 7043 29600 7069
rect 29636 7043 29662 7069
rect 29698 7043 29724 7069
rect 29760 7043 29786 7069
rect 29822 7043 29848 7069
rect 29884 7043 29910 7069
rect 29946 7043 29972 7069
rect 30008 7043 30034 7069
rect 34574 7043 34600 7069
rect 34636 7043 34662 7069
rect 34698 7043 34724 7069
rect 34760 7043 34786 7069
rect 34822 7043 34848 7069
rect 34884 7043 34910 7069
rect 34946 7043 34972 7069
rect 35008 7043 35034 7069
rect 4495 6903 4521 6929
rect 7015 6903 7041 6929
rect 8359 6903 8385 6929
rect 16199 6903 16225 6929
rect 19335 6903 19361 6929
rect 23423 6903 23449 6929
rect 33671 6903 33697 6929
rect 35127 6903 35153 6929
rect 35631 6903 35657 6929
rect 35743 6903 35769 6929
rect 35911 6903 35937 6929
rect 37647 6903 37673 6929
rect 2367 6847 2393 6873
rect 2479 6847 2505 6873
rect 3039 6847 3065 6873
rect 3599 6847 3625 6873
rect 4495 6847 4521 6873
rect 6119 6847 6145 6873
rect 7015 6847 7041 6873
rect 7575 6847 7601 6873
rect 8359 6847 8385 6873
rect 10039 6847 10065 6873
rect 10263 6847 10289 6873
rect 10543 6847 10569 6873
rect 11551 6847 11577 6873
rect 11775 6847 11801 6873
rect 11999 6847 12025 6873
rect 13735 6847 13761 6873
rect 14295 6847 14321 6873
rect 14407 6847 14433 6873
rect 15247 6847 15273 6873
rect 16199 6847 16225 6873
rect 16815 6847 16841 6873
rect 17375 6847 17401 6873
rect 17599 6847 17625 6873
rect 18551 6847 18577 6873
rect 19335 6847 19361 6873
rect 20791 6847 20817 6873
rect 21295 6847 21321 6873
rect 21463 6847 21489 6873
rect 22527 6847 22553 6873
rect 23423 6847 23449 6873
rect 24767 6847 24793 6873
rect 25215 6847 25241 6873
rect 25439 6847 25465 6873
rect 26223 6847 26249 6873
rect 26783 6847 26809 6873
rect 26895 6847 26921 6873
rect 28743 6847 28769 6873
rect 29191 6847 29217 6873
rect 29415 6847 29441 6873
rect 30479 6847 30505 6873
rect 30647 6847 30673 6873
rect 31375 6847 31401 6873
rect 32047 6847 32073 6873
rect 32159 6847 32185 6873
rect 32327 6847 32353 6873
rect 32999 6847 33025 6873
rect 33671 6847 33697 6873
rect 34399 6847 34425 6873
rect 35127 6847 35153 6873
rect 36695 6847 36721 6873
rect 37647 6847 37673 6873
rect 2074 6651 2100 6677
rect 2136 6651 2162 6677
rect 2198 6651 2224 6677
rect 2260 6651 2286 6677
rect 2322 6651 2348 6677
rect 2384 6651 2410 6677
rect 2446 6651 2472 6677
rect 2508 6651 2534 6677
rect 7074 6651 7100 6677
rect 7136 6651 7162 6677
rect 7198 6651 7224 6677
rect 7260 6651 7286 6677
rect 7322 6651 7348 6677
rect 7384 6651 7410 6677
rect 7446 6651 7472 6677
rect 7508 6651 7534 6677
rect 12074 6651 12100 6677
rect 12136 6651 12162 6677
rect 12198 6651 12224 6677
rect 12260 6651 12286 6677
rect 12322 6651 12348 6677
rect 12384 6651 12410 6677
rect 12446 6651 12472 6677
rect 12508 6651 12534 6677
rect 17074 6651 17100 6677
rect 17136 6651 17162 6677
rect 17198 6651 17224 6677
rect 17260 6651 17286 6677
rect 17322 6651 17348 6677
rect 17384 6651 17410 6677
rect 17446 6651 17472 6677
rect 17508 6651 17534 6677
rect 22074 6651 22100 6677
rect 22136 6651 22162 6677
rect 22198 6651 22224 6677
rect 22260 6651 22286 6677
rect 22322 6651 22348 6677
rect 22384 6651 22410 6677
rect 22446 6651 22472 6677
rect 22508 6651 22534 6677
rect 27074 6651 27100 6677
rect 27136 6651 27162 6677
rect 27198 6651 27224 6677
rect 27260 6651 27286 6677
rect 27322 6651 27348 6677
rect 27384 6651 27410 6677
rect 27446 6651 27472 6677
rect 27508 6651 27534 6677
rect 32074 6651 32100 6677
rect 32136 6651 32162 6677
rect 32198 6651 32224 6677
rect 32260 6651 32286 6677
rect 32322 6651 32348 6677
rect 32384 6651 32410 6677
rect 32446 6651 32472 6677
rect 32508 6651 32534 6677
rect 37074 6651 37100 6677
rect 37136 6651 37162 6677
rect 37198 6651 37224 6677
rect 37260 6651 37286 6677
rect 37322 6651 37348 6677
rect 37384 6651 37410 6677
rect 37446 6651 37472 6677
rect 37508 6651 37534 6677
rect 1807 6455 1833 6481
rect 1975 6455 2001 6481
rect 2479 6455 2505 6481
rect 4103 6455 4129 6481
rect 4383 6455 4409 6481
rect 4495 6455 4521 6481
rect 5279 6455 5305 6481
rect 6455 6455 6481 6481
rect 8079 6455 8105 6481
rect 8975 6455 9001 6481
rect 9423 6455 9449 6481
rect 10319 6455 10345 6481
rect 11831 6455 11857 6481
rect 12335 6455 12361 6481
rect 12447 6455 12473 6481
rect 13511 6455 13537 6481
rect 14239 6455 14265 6481
rect 16367 6455 16393 6481
rect 17319 6455 17345 6481
rect 18775 6455 18801 6481
rect 19335 6455 19361 6481
rect 19447 6455 19473 6481
rect 20231 6455 20257 6481
rect 21295 6455 21321 6481
rect 22751 6455 22777 6481
rect 23199 6455 23225 6481
rect 23423 6455 23449 6481
rect 24375 6455 24401 6481
rect 25215 6455 25241 6481
rect 26727 6455 26753 6481
rect 27175 6455 27201 6481
rect 27399 6455 27425 6481
rect 28463 6455 28489 6481
rect 28687 6455 28713 6481
rect 28855 6455 28881 6481
rect 30199 6455 30225 6481
rect 30311 6455 30337 6481
rect 30927 6455 30953 6481
rect 31879 6455 31905 6481
rect 32159 6455 32185 6481
rect 33279 6455 33305 6481
rect 34679 6455 34705 6481
rect 35239 6455 35265 6481
rect 35351 6455 35377 6481
rect 36135 6455 36161 6481
rect 37311 6455 37337 6481
rect 6455 6399 6481 6425
rect 8975 6399 9001 6425
rect 10319 6399 10345 6425
rect 14239 6399 14265 6425
rect 17319 6399 17345 6425
rect 21295 6399 21321 6425
rect 25215 6399 25241 6425
rect 30031 6399 30057 6425
rect 31879 6399 31905 6425
rect 33279 6399 33305 6425
rect 33615 6399 33641 6425
rect 33727 6399 33753 6425
rect 33895 6399 33921 6425
rect 37311 6399 37337 6425
rect 4574 6259 4600 6285
rect 4636 6259 4662 6285
rect 4698 6259 4724 6285
rect 4760 6259 4786 6285
rect 4822 6259 4848 6285
rect 4884 6259 4910 6285
rect 4946 6259 4972 6285
rect 5008 6259 5034 6285
rect 9574 6259 9600 6285
rect 9636 6259 9662 6285
rect 9698 6259 9724 6285
rect 9760 6259 9786 6285
rect 9822 6259 9848 6285
rect 9884 6259 9910 6285
rect 9946 6259 9972 6285
rect 10008 6259 10034 6285
rect 14574 6259 14600 6285
rect 14636 6259 14662 6285
rect 14698 6259 14724 6285
rect 14760 6259 14786 6285
rect 14822 6259 14848 6285
rect 14884 6259 14910 6285
rect 14946 6259 14972 6285
rect 15008 6259 15034 6285
rect 19574 6259 19600 6285
rect 19636 6259 19662 6285
rect 19698 6259 19724 6285
rect 19760 6259 19786 6285
rect 19822 6259 19848 6285
rect 19884 6259 19910 6285
rect 19946 6259 19972 6285
rect 20008 6259 20034 6285
rect 24574 6259 24600 6285
rect 24636 6259 24662 6285
rect 24698 6259 24724 6285
rect 24760 6259 24786 6285
rect 24822 6259 24848 6285
rect 24884 6259 24910 6285
rect 24946 6259 24972 6285
rect 25008 6259 25034 6285
rect 29574 6259 29600 6285
rect 29636 6259 29662 6285
rect 29698 6259 29724 6285
rect 29760 6259 29786 6285
rect 29822 6259 29848 6285
rect 29884 6259 29910 6285
rect 29946 6259 29972 6285
rect 30008 6259 30034 6285
rect 34574 6259 34600 6285
rect 34636 6259 34662 6285
rect 34698 6259 34724 6285
rect 34760 6259 34786 6285
rect 34822 6259 34848 6285
rect 34884 6259 34910 6285
rect 34946 6259 34972 6285
rect 35008 6259 35034 6285
rect 1975 6119 2001 6145
rect 4495 6119 4521 6145
rect 7015 6119 7041 6145
rect 8471 6119 8497 6145
rect 12447 6119 12473 6145
rect 14855 6119 14881 6145
rect 17767 6119 17793 6145
rect 19447 6119 19473 6145
rect 27175 6119 27201 6145
rect 29919 6119 29945 6145
rect 31375 6119 31401 6145
rect 33783 6119 33809 6145
rect 35127 6119 35153 6145
rect 37647 6119 37673 6145
rect 1975 6063 2001 6089
rect 3039 6063 3065 6089
rect 3599 6063 3625 6089
rect 4495 6063 4521 6089
rect 6119 6063 6145 6089
rect 7015 6063 7041 6089
rect 7575 6063 7601 6089
rect 8471 6063 8497 6089
rect 10039 6063 10065 6089
rect 10319 6063 10345 6089
rect 10487 6063 10513 6089
rect 11551 6063 11577 6089
rect 12447 6063 12473 6089
rect 13959 6063 13985 6089
rect 14855 6063 14881 6089
rect 15191 6063 15217 6089
rect 15695 6063 15721 6089
rect 15863 6063 15889 6089
rect 16815 6063 16841 6089
rect 17711 6063 17737 6089
rect 18551 6063 18577 6089
rect 19447 6063 19473 6089
rect 20791 6063 20817 6089
rect 21295 6063 21321 6089
rect 21463 6063 21489 6089
rect 22247 6063 22273 6089
rect 22695 6063 22721 6089
rect 22919 6063 22945 6089
rect 24767 6063 24793 6089
rect 25215 6063 25241 6089
rect 25439 6063 25465 6089
rect 26223 6063 26249 6089
rect 26895 6063 26921 6089
rect 28743 6063 28769 6089
rect 29919 6063 29945 6089
rect 30255 6063 30281 6089
rect 31375 6063 31401 6089
rect 32047 6063 32073 6089
rect 32159 6063 32185 6089
rect 32327 6063 32353 6089
rect 32719 6063 32745 6089
rect 33615 6063 33641 6089
rect 34399 6063 34425 6089
rect 35127 6063 35153 6089
rect 35631 6063 35657 6089
rect 35743 6063 35769 6089
rect 35911 6063 35937 6089
rect 36695 6063 36721 6089
rect 37647 6063 37673 6089
rect 2074 5867 2100 5893
rect 2136 5867 2162 5893
rect 2198 5867 2224 5893
rect 2260 5867 2286 5893
rect 2322 5867 2348 5893
rect 2384 5867 2410 5893
rect 2446 5867 2472 5893
rect 2508 5867 2534 5893
rect 7074 5867 7100 5893
rect 7136 5867 7162 5893
rect 7198 5867 7224 5893
rect 7260 5867 7286 5893
rect 7322 5867 7348 5893
rect 7384 5867 7410 5893
rect 7446 5867 7472 5893
rect 7508 5867 7534 5893
rect 12074 5867 12100 5893
rect 12136 5867 12162 5893
rect 12198 5867 12224 5893
rect 12260 5867 12286 5893
rect 12322 5867 12348 5893
rect 12384 5867 12410 5893
rect 12446 5867 12472 5893
rect 12508 5867 12534 5893
rect 17074 5867 17100 5893
rect 17136 5867 17162 5893
rect 17198 5867 17224 5893
rect 17260 5867 17286 5893
rect 17322 5867 17348 5893
rect 17384 5867 17410 5893
rect 17446 5867 17472 5893
rect 17508 5867 17534 5893
rect 22074 5867 22100 5893
rect 22136 5867 22162 5893
rect 22198 5867 22224 5893
rect 22260 5867 22286 5893
rect 22322 5867 22348 5893
rect 22384 5867 22410 5893
rect 22446 5867 22472 5893
rect 22508 5867 22534 5893
rect 27074 5867 27100 5893
rect 27136 5867 27162 5893
rect 27198 5867 27224 5893
rect 27260 5867 27286 5893
rect 27322 5867 27348 5893
rect 27384 5867 27410 5893
rect 27446 5867 27472 5893
rect 27508 5867 27534 5893
rect 32074 5867 32100 5893
rect 32136 5867 32162 5893
rect 32198 5867 32224 5893
rect 32260 5867 32286 5893
rect 32322 5867 32348 5893
rect 32384 5867 32410 5893
rect 32446 5867 32472 5893
rect 32508 5867 32534 5893
rect 37074 5867 37100 5893
rect 37136 5867 37162 5893
rect 37198 5867 37224 5893
rect 37260 5867 37286 5893
rect 37322 5867 37348 5893
rect 37384 5867 37410 5893
rect 37446 5867 37472 5893
rect 37508 5867 37534 5893
rect 1807 5671 1833 5697
rect 1975 5671 2001 5697
rect 2479 5671 2505 5697
rect 4103 5671 4129 5697
rect 4999 5671 5025 5697
rect 5279 5671 5305 5697
rect 5839 5671 5865 5697
rect 5951 5671 5977 5697
rect 8079 5671 8105 5697
rect 8975 5671 9001 5697
rect 9423 5671 9449 5697
rect 10263 5671 10289 5697
rect 11999 5671 12025 5697
rect 12951 5671 12977 5697
rect 13343 5671 13369 5697
rect 14407 5671 14433 5697
rect 15191 5671 15217 5697
rect 15863 5671 15889 5697
rect 16815 5671 16841 5697
rect 17711 5671 17737 5697
rect 18775 5671 18801 5697
rect 19951 5671 19977 5697
rect 20231 5671 20257 5697
rect 21295 5671 21321 5697
rect 22751 5671 22777 5697
rect 23199 5671 23225 5697
rect 23423 5671 23449 5697
rect 24375 5671 24401 5697
rect 25159 5671 25185 5697
rect 26727 5671 26753 5697
rect 27567 5671 27593 5697
rect 28239 5671 28265 5697
rect 29135 5671 29161 5697
rect 30087 5671 30113 5697
rect 30703 5671 30729 5697
rect 31879 5671 31905 5697
rect 32159 5671 32185 5697
rect 33335 5671 33361 5697
rect 33671 5671 33697 5697
rect 34959 5671 34985 5697
rect 35127 5671 35153 5697
rect 35351 5671 35377 5697
rect 36135 5671 36161 5697
rect 37143 5671 37169 5697
rect 4999 5615 5025 5641
rect 8975 5615 9001 5641
rect 10263 5615 10289 5641
rect 12951 5615 12977 5641
rect 14407 5615 14433 5641
rect 16031 5615 16057 5641
rect 17711 5615 17737 5641
rect 19951 5615 19977 5641
rect 21295 5615 21321 5641
rect 25159 5615 25185 5641
rect 27679 5615 27705 5641
rect 29135 5615 29161 5641
rect 30143 5615 30169 5641
rect 30311 5615 30337 5641
rect 31879 5615 31905 5641
rect 33335 5615 33361 5641
rect 33727 5615 33753 5641
rect 33895 5615 33921 5641
rect 37143 5615 37169 5641
rect 37591 5615 37617 5641
rect 37703 5615 37729 5641
rect 37871 5615 37897 5641
rect 4574 5475 4600 5501
rect 4636 5475 4662 5501
rect 4698 5475 4724 5501
rect 4760 5475 4786 5501
rect 4822 5475 4848 5501
rect 4884 5475 4910 5501
rect 4946 5475 4972 5501
rect 5008 5475 5034 5501
rect 9574 5475 9600 5501
rect 9636 5475 9662 5501
rect 9698 5475 9724 5501
rect 9760 5475 9786 5501
rect 9822 5475 9848 5501
rect 9884 5475 9910 5501
rect 9946 5475 9972 5501
rect 10008 5475 10034 5501
rect 14574 5475 14600 5501
rect 14636 5475 14662 5501
rect 14698 5475 14724 5501
rect 14760 5475 14786 5501
rect 14822 5475 14848 5501
rect 14884 5475 14910 5501
rect 14946 5475 14972 5501
rect 15008 5475 15034 5501
rect 19574 5475 19600 5501
rect 19636 5475 19662 5501
rect 19698 5475 19724 5501
rect 19760 5475 19786 5501
rect 19822 5475 19848 5501
rect 19884 5475 19910 5501
rect 19946 5475 19972 5501
rect 20008 5475 20034 5501
rect 24574 5475 24600 5501
rect 24636 5475 24662 5501
rect 24698 5475 24724 5501
rect 24760 5475 24786 5501
rect 24822 5475 24848 5501
rect 24884 5475 24910 5501
rect 24946 5475 24972 5501
rect 25008 5475 25034 5501
rect 29574 5475 29600 5501
rect 29636 5475 29662 5501
rect 29698 5475 29724 5501
rect 29760 5475 29786 5501
rect 29822 5475 29848 5501
rect 29884 5475 29910 5501
rect 29946 5475 29972 5501
rect 30008 5475 30034 5501
rect 34574 5475 34600 5501
rect 34636 5475 34662 5501
rect 34698 5475 34724 5501
rect 34760 5475 34786 5501
rect 34822 5475 34848 5501
rect 34884 5475 34910 5501
rect 34946 5475 34972 5501
rect 35008 5475 35034 5501
rect 1975 5335 2001 5361
rect 4495 5335 4521 5361
rect 6791 5335 6817 5361
rect 8471 5335 8497 5361
rect 12447 5335 12473 5361
rect 14463 5335 14489 5361
rect 15863 5335 15889 5361
rect 17767 5335 17793 5361
rect 19447 5335 19473 5361
rect 23199 5335 23225 5361
rect 28071 5335 28097 5361
rect 29695 5335 29721 5361
rect 31375 5335 31401 5361
rect 33839 5335 33865 5361
rect 35239 5335 35265 5361
rect 1975 5279 2001 5305
rect 3039 5279 3065 5305
rect 3431 5279 3457 5305
rect 4495 5279 4521 5305
rect 6119 5279 6145 5305
rect 6791 5279 6817 5305
rect 7295 5279 7321 5305
rect 8471 5279 8497 5305
rect 10039 5279 10065 5305
rect 10319 5279 10345 5305
rect 10487 5279 10513 5305
rect 11551 5279 11577 5305
rect 12447 5279 12473 5305
rect 13567 5279 13593 5305
rect 14463 5279 14489 5305
rect 15191 5279 15217 5305
rect 15863 5279 15889 5305
rect 16815 5279 16841 5305
rect 17767 5279 17793 5305
rect 18551 5279 18577 5305
rect 19447 5279 19473 5305
rect 20791 5279 20817 5305
rect 21295 5279 21321 5305
rect 21463 5279 21489 5305
rect 22527 5279 22553 5305
rect 23199 5279 23225 5305
rect 24767 5279 24793 5305
rect 25215 5279 25241 5305
rect 25943 5279 25969 5305
rect 26223 5279 26249 5305
rect 26783 5279 26809 5305
rect 26895 5279 26921 5305
rect 28183 5279 28209 5305
rect 28407 5279 28433 5305
rect 28743 5279 28769 5305
rect 29471 5279 29497 5305
rect 30367 5279 30393 5305
rect 31375 5279 31401 5305
rect 32047 5279 32073 5305
rect 32159 5279 32185 5305
rect 32327 5279 32353 5305
rect 32775 5279 32801 5305
rect 33839 5279 33865 5305
rect 34175 5279 34201 5305
rect 35239 5279 35265 5305
rect 35631 5279 35657 5305
rect 35743 5279 35769 5305
rect 35911 5279 35937 5305
rect 36695 5279 36721 5305
rect 37143 5279 37169 5305
rect 37367 5279 37393 5305
rect 38151 5279 38177 5305
rect 38263 5279 38289 5305
rect 38431 5279 38457 5305
rect 2074 5083 2100 5109
rect 2136 5083 2162 5109
rect 2198 5083 2224 5109
rect 2260 5083 2286 5109
rect 2322 5083 2348 5109
rect 2384 5083 2410 5109
rect 2446 5083 2472 5109
rect 2508 5083 2534 5109
rect 7074 5083 7100 5109
rect 7136 5083 7162 5109
rect 7198 5083 7224 5109
rect 7260 5083 7286 5109
rect 7322 5083 7348 5109
rect 7384 5083 7410 5109
rect 7446 5083 7472 5109
rect 7508 5083 7534 5109
rect 12074 5083 12100 5109
rect 12136 5083 12162 5109
rect 12198 5083 12224 5109
rect 12260 5083 12286 5109
rect 12322 5083 12348 5109
rect 12384 5083 12410 5109
rect 12446 5083 12472 5109
rect 12508 5083 12534 5109
rect 17074 5083 17100 5109
rect 17136 5083 17162 5109
rect 17198 5083 17224 5109
rect 17260 5083 17286 5109
rect 17322 5083 17348 5109
rect 17384 5083 17410 5109
rect 17446 5083 17472 5109
rect 17508 5083 17534 5109
rect 22074 5083 22100 5109
rect 22136 5083 22162 5109
rect 22198 5083 22224 5109
rect 22260 5083 22286 5109
rect 22322 5083 22348 5109
rect 22384 5083 22410 5109
rect 22446 5083 22472 5109
rect 22508 5083 22534 5109
rect 27074 5083 27100 5109
rect 27136 5083 27162 5109
rect 27198 5083 27224 5109
rect 27260 5083 27286 5109
rect 27322 5083 27348 5109
rect 27384 5083 27410 5109
rect 27446 5083 27472 5109
rect 27508 5083 27534 5109
rect 32074 5083 32100 5109
rect 32136 5083 32162 5109
rect 32198 5083 32224 5109
rect 32260 5083 32286 5109
rect 32322 5083 32348 5109
rect 32384 5083 32410 5109
rect 32446 5083 32472 5109
rect 32508 5083 32534 5109
rect 37074 5083 37100 5109
rect 37136 5083 37162 5109
rect 37198 5083 37224 5109
rect 37260 5083 37286 5109
rect 37322 5083 37348 5109
rect 37384 5083 37410 5109
rect 37446 5083 37472 5109
rect 37508 5083 37534 5109
rect 1807 4887 1833 4913
rect 1919 4887 1945 4913
rect 2479 4887 2505 4913
rect 4103 4887 4129 4913
rect 4999 4887 5025 4913
rect 5279 4887 5305 4913
rect 6455 4887 6481 4913
rect 8079 4887 8105 4913
rect 8975 4887 9001 4913
rect 9423 4887 9449 4913
rect 10319 4887 10345 4913
rect 11999 4887 12025 4913
rect 12951 4887 12977 4913
rect 13343 4887 13369 4913
rect 14183 4887 14209 4913
rect 15583 4887 15609 4913
rect 15807 4887 15833 4913
rect 16031 4887 16057 4913
rect 16815 4887 16841 4913
rect 17767 4887 17793 4913
rect 18775 4887 18801 4913
rect 19951 4887 19977 4913
rect 20231 4887 20257 4913
rect 21295 4887 21321 4913
rect 22751 4887 22777 4913
rect 23199 4887 23225 4913
rect 23423 4887 23449 4913
rect 24375 4887 24401 4913
rect 25215 4887 25241 4913
rect 26727 4887 26753 4913
rect 27287 4887 27313 4913
rect 27399 4887 27425 4913
rect 28239 4887 28265 4913
rect 29135 4887 29161 4913
rect 30087 4887 30113 4913
rect 30199 4887 30225 4913
rect 30311 4887 30337 4913
rect 30703 4887 30729 4913
rect 31879 4887 31905 4913
rect 32159 4887 32185 4913
rect 33335 4887 33361 4913
rect 33671 4887 33697 4913
rect 33783 4887 33809 4913
rect 33895 4887 33921 4913
rect 34679 4887 34705 4913
rect 35855 4887 35881 4913
rect 36135 4887 36161 4913
rect 37311 4887 37337 4913
rect 37591 4887 37617 4913
rect 37759 4887 37785 4913
rect 37871 4887 37897 4913
rect 38655 4887 38681 4913
rect 38767 4887 38793 4913
rect 38879 4887 38905 4913
rect 4999 4831 5025 4857
rect 6455 4831 6481 4857
rect 8975 4831 9001 4857
rect 10319 4831 10345 4857
rect 12951 4831 12977 4857
rect 14183 4831 14209 4857
rect 17767 4831 17793 4857
rect 19951 4831 19977 4857
rect 21295 4831 21321 4857
rect 25215 4831 25241 4857
rect 29135 4831 29161 4857
rect 31879 4831 31905 4857
rect 33335 4831 33361 4857
rect 35855 4831 35881 4857
rect 37311 4831 37337 4857
rect 4574 4691 4600 4717
rect 4636 4691 4662 4717
rect 4698 4691 4724 4717
rect 4760 4691 4786 4717
rect 4822 4691 4848 4717
rect 4884 4691 4910 4717
rect 4946 4691 4972 4717
rect 5008 4691 5034 4717
rect 9574 4691 9600 4717
rect 9636 4691 9662 4717
rect 9698 4691 9724 4717
rect 9760 4691 9786 4717
rect 9822 4691 9848 4717
rect 9884 4691 9910 4717
rect 9946 4691 9972 4717
rect 10008 4691 10034 4717
rect 14574 4691 14600 4717
rect 14636 4691 14662 4717
rect 14698 4691 14724 4717
rect 14760 4691 14786 4717
rect 14822 4691 14848 4717
rect 14884 4691 14910 4717
rect 14946 4691 14972 4717
rect 15008 4691 15034 4717
rect 19574 4691 19600 4717
rect 19636 4691 19662 4717
rect 19698 4691 19724 4717
rect 19760 4691 19786 4717
rect 19822 4691 19848 4717
rect 19884 4691 19910 4717
rect 19946 4691 19972 4717
rect 20008 4691 20034 4717
rect 24574 4691 24600 4717
rect 24636 4691 24662 4717
rect 24698 4691 24724 4717
rect 24760 4691 24786 4717
rect 24822 4691 24848 4717
rect 24884 4691 24910 4717
rect 24946 4691 24972 4717
rect 25008 4691 25034 4717
rect 29574 4691 29600 4717
rect 29636 4691 29662 4717
rect 29698 4691 29724 4717
rect 29760 4691 29786 4717
rect 29822 4691 29848 4717
rect 29884 4691 29910 4717
rect 29946 4691 29972 4717
rect 30008 4691 30034 4717
rect 34574 4691 34600 4717
rect 34636 4691 34662 4717
rect 34698 4691 34724 4717
rect 34760 4691 34786 4717
rect 34822 4691 34848 4717
rect 34884 4691 34910 4717
rect 34946 4691 34972 4717
rect 35008 4691 35034 4717
rect 1863 4551 1889 4577
rect 4495 4551 4521 4577
rect 6791 4551 6817 4577
rect 8471 4551 8497 4577
rect 12447 4551 12473 4577
rect 17767 4551 17793 4577
rect 19447 4551 19473 4577
rect 21799 4551 21825 4577
rect 27399 4551 27425 4577
rect 28183 4551 28209 4577
rect 31375 4551 31401 4577
rect 33839 4551 33865 4577
rect 35911 4551 35937 4577
rect 37647 4551 37673 4577
rect 38151 4551 38177 4577
rect 38263 4551 38289 4577
rect 38431 4551 38457 4577
rect 38711 4551 38737 4577
rect 1863 4495 1889 4521
rect 3039 4495 3065 4521
rect 3431 4495 3457 4521
rect 4495 4495 4521 4521
rect 6119 4495 6145 4521
rect 6791 4495 6817 4521
rect 7575 4495 7601 4521
rect 8471 4495 8497 4521
rect 10039 4495 10065 4521
rect 10319 4495 10345 4521
rect 10487 4495 10513 4521
rect 11551 4495 11577 4521
rect 12447 4495 12473 4521
rect 13567 4495 13593 4521
rect 14127 4495 14153 4521
rect 14239 4495 14265 4521
rect 15135 4495 15161 4521
rect 15471 4495 15497 4521
rect 15695 4495 15721 4521
rect 16815 4495 16841 4521
rect 17767 4495 17793 4521
rect 18551 4495 18577 4521
rect 19447 4495 19473 4521
rect 20791 4495 20817 4521
rect 21799 4495 21825 4521
rect 22527 4495 22553 4521
rect 22695 4495 22721 4521
rect 22919 4495 22945 4521
rect 24767 4495 24793 4521
rect 25215 4495 25241 4521
rect 25943 4495 25969 4521
rect 26279 4495 26305 4521
rect 27399 4495 27425 4521
rect 28127 4495 28153 4521
rect 28351 4495 28377 4521
rect 28743 4495 28769 4521
rect 29191 4495 29217 4521
rect 29415 4495 29441 4521
rect 30367 4495 30393 4521
rect 31375 4495 31401 4521
rect 32047 4495 32073 4521
rect 32215 4495 32241 4521
rect 32383 4495 32409 4521
rect 32775 4495 32801 4521
rect 33839 4495 33865 4521
rect 34175 4495 34201 4521
rect 34623 4495 34649 4521
rect 34847 4495 34873 4521
rect 35687 4495 35713 4521
rect 35799 4495 35825 4521
rect 36695 4495 36721 4521
rect 37647 4495 37673 4521
rect 38823 4495 38849 4521
rect 38935 4495 38961 4521
rect 2074 4299 2100 4325
rect 2136 4299 2162 4325
rect 2198 4299 2224 4325
rect 2260 4299 2286 4325
rect 2322 4299 2348 4325
rect 2384 4299 2410 4325
rect 2446 4299 2472 4325
rect 2508 4299 2534 4325
rect 7074 4299 7100 4325
rect 7136 4299 7162 4325
rect 7198 4299 7224 4325
rect 7260 4299 7286 4325
rect 7322 4299 7348 4325
rect 7384 4299 7410 4325
rect 7446 4299 7472 4325
rect 7508 4299 7534 4325
rect 12074 4299 12100 4325
rect 12136 4299 12162 4325
rect 12198 4299 12224 4325
rect 12260 4299 12286 4325
rect 12322 4299 12348 4325
rect 12384 4299 12410 4325
rect 12446 4299 12472 4325
rect 12508 4299 12534 4325
rect 17074 4299 17100 4325
rect 17136 4299 17162 4325
rect 17198 4299 17224 4325
rect 17260 4299 17286 4325
rect 17322 4299 17348 4325
rect 17384 4299 17410 4325
rect 17446 4299 17472 4325
rect 17508 4299 17534 4325
rect 22074 4299 22100 4325
rect 22136 4299 22162 4325
rect 22198 4299 22224 4325
rect 22260 4299 22286 4325
rect 22322 4299 22348 4325
rect 22384 4299 22410 4325
rect 22446 4299 22472 4325
rect 22508 4299 22534 4325
rect 27074 4299 27100 4325
rect 27136 4299 27162 4325
rect 27198 4299 27224 4325
rect 27260 4299 27286 4325
rect 27322 4299 27348 4325
rect 27384 4299 27410 4325
rect 27446 4299 27472 4325
rect 27508 4299 27534 4325
rect 32074 4299 32100 4325
rect 32136 4299 32162 4325
rect 32198 4299 32224 4325
rect 32260 4299 32286 4325
rect 32322 4299 32348 4325
rect 32384 4299 32410 4325
rect 32446 4299 32472 4325
rect 32508 4299 32534 4325
rect 37074 4299 37100 4325
rect 37136 4299 37162 4325
rect 37198 4299 37224 4325
rect 37260 4299 37286 4325
rect 37322 4299 37348 4325
rect 37384 4299 37410 4325
rect 37446 4299 37472 4325
rect 37508 4299 37534 4325
rect 1807 4103 1833 4129
rect 1919 4103 1945 4129
rect 2479 4103 2505 4129
rect 4103 4103 4129 4129
rect 4775 4103 4801 4129
rect 5279 4103 5305 4129
rect 6455 4103 6481 4129
rect 8079 4103 8105 4129
rect 8975 4103 9001 4129
rect 9535 4103 9561 4129
rect 10319 4103 10345 4129
rect 11999 4103 12025 4129
rect 12727 4103 12753 4129
rect 13343 4103 13369 4129
rect 14239 4103 14265 4129
rect 15527 4103 15553 4129
rect 15807 4103 15833 4129
rect 16031 4103 16057 4129
rect 16815 4103 16841 4129
rect 17767 4103 17793 4129
rect 18775 4103 18801 4129
rect 19951 4103 19977 4129
rect 20231 4103 20257 4129
rect 21183 4103 21209 4129
rect 22751 4103 22777 4129
rect 23311 4103 23337 4129
rect 23423 4103 23449 4129
rect 24375 4103 24401 4129
rect 24655 4103 24681 4129
rect 24879 4103 24905 4129
rect 26727 4103 26753 4129
rect 27175 4103 27201 4129
rect 27399 4103 27425 4129
rect 28463 4103 28489 4129
rect 29359 4103 29385 4129
rect 30199 4103 30225 4129
rect 30311 4103 30337 4129
rect 30703 4103 30729 4129
rect 31879 4103 31905 4129
rect 32159 4103 32185 4129
rect 33335 4103 33361 4129
rect 33671 4103 33697 4129
rect 33783 4103 33809 4129
rect 33951 4103 33977 4129
rect 34679 4103 34705 4129
rect 35183 4103 35209 4129
rect 35351 4103 35377 4129
rect 36135 4103 36161 4129
rect 37087 4103 37113 4129
rect 37591 4103 37617 4129
rect 37703 4103 37729 4129
rect 37871 4103 37897 4129
rect 38655 4103 38681 4129
rect 38767 4103 38793 4129
rect 4775 4047 4801 4073
rect 6455 4047 6481 4073
rect 8975 4047 9001 4073
rect 10319 4047 10345 4073
rect 12727 4047 12753 4073
rect 14239 4047 14265 4073
rect 17767 4047 17793 4073
rect 19951 4047 19977 4073
rect 21183 4047 21209 4073
rect 29359 4047 29385 4073
rect 30031 4047 30057 4073
rect 31879 4047 31905 4073
rect 33335 4047 33361 4073
rect 37087 4047 37113 4073
rect 38935 4047 38961 4073
rect 4574 3907 4600 3933
rect 4636 3907 4662 3933
rect 4698 3907 4724 3933
rect 4760 3907 4786 3933
rect 4822 3907 4848 3933
rect 4884 3907 4910 3933
rect 4946 3907 4972 3933
rect 5008 3907 5034 3933
rect 9574 3907 9600 3933
rect 9636 3907 9662 3933
rect 9698 3907 9724 3933
rect 9760 3907 9786 3933
rect 9822 3907 9848 3933
rect 9884 3907 9910 3933
rect 9946 3907 9972 3933
rect 10008 3907 10034 3933
rect 14574 3907 14600 3933
rect 14636 3907 14662 3933
rect 14698 3907 14724 3933
rect 14760 3907 14786 3933
rect 14822 3907 14848 3933
rect 14884 3907 14910 3933
rect 14946 3907 14972 3933
rect 15008 3907 15034 3933
rect 19574 3907 19600 3933
rect 19636 3907 19662 3933
rect 19698 3907 19724 3933
rect 19760 3907 19786 3933
rect 19822 3907 19848 3933
rect 19884 3907 19910 3933
rect 19946 3907 19972 3933
rect 20008 3907 20034 3933
rect 24574 3907 24600 3933
rect 24636 3907 24662 3933
rect 24698 3907 24724 3933
rect 24760 3907 24786 3933
rect 24822 3907 24848 3933
rect 24884 3907 24910 3933
rect 24946 3907 24972 3933
rect 25008 3907 25034 3933
rect 29574 3907 29600 3933
rect 29636 3907 29662 3933
rect 29698 3907 29724 3933
rect 29760 3907 29786 3933
rect 29822 3907 29848 3933
rect 29884 3907 29910 3933
rect 29946 3907 29972 3933
rect 30008 3907 30034 3933
rect 34574 3907 34600 3933
rect 34636 3907 34662 3933
rect 34698 3907 34724 3933
rect 34760 3907 34786 3933
rect 34822 3907 34848 3933
rect 34884 3907 34910 3933
rect 34946 3907 34972 3933
rect 35008 3907 35034 3933
rect 1919 3767 1945 3793
rect 4495 3767 4521 3793
rect 6959 3767 6985 3793
rect 8359 3767 8385 3793
rect 12447 3767 12473 3793
rect 17767 3767 17793 3793
rect 19447 3767 19473 3793
rect 21743 3767 21769 3793
rect 27175 3767 27201 3793
rect 28351 3767 28377 3793
rect 29919 3767 29945 3793
rect 31319 3767 31345 3793
rect 33895 3767 33921 3793
rect 35127 3767 35153 3793
rect 35743 3767 35769 3793
rect 35911 3767 35937 3793
rect 36919 3767 36945 3793
rect 38263 3767 38289 3793
rect 38431 3767 38457 3793
rect 38711 3767 38737 3793
rect 1919 3711 1945 3737
rect 3039 3711 3065 3737
rect 3487 3711 3513 3737
rect 4495 3711 4521 3737
rect 5839 3711 5865 3737
rect 6959 3711 6985 3737
rect 7575 3711 7601 3737
rect 8359 3711 8385 3737
rect 10039 3711 10065 3737
rect 10263 3711 10289 3737
rect 10487 3711 10513 3737
rect 11551 3711 11577 3737
rect 12447 3711 12473 3737
rect 13679 3711 13705 3737
rect 14127 3711 14153 3737
rect 14351 3711 14377 3737
rect 15135 3711 15161 3737
rect 15583 3711 15609 3737
rect 15807 3711 15833 3737
rect 16815 3711 16841 3737
rect 17767 3711 17793 3737
rect 18551 3711 18577 3737
rect 19447 3711 19473 3737
rect 20791 3711 20817 3737
rect 21743 3711 21769 3737
rect 22527 3711 22553 3737
rect 22807 3711 22833 3737
rect 22919 3711 22945 3737
rect 24767 3711 24793 3737
rect 25215 3711 25241 3737
rect 25439 3711 25465 3737
rect 26279 3711 26305 3737
rect 26895 3711 26921 3737
rect 28071 3711 28097 3737
rect 28239 3711 28265 3737
rect 29023 3711 29049 3737
rect 29919 3711 29945 3737
rect 30367 3711 30393 3737
rect 31319 3711 31345 3737
rect 32047 3711 32073 3737
rect 32215 3711 32241 3737
rect 32383 3711 32409 3737
rect 32775 3711 32801 3737
rect 33895 3711 33921 3737
rect 34175 3711 34201 3737
rect 35071 3711 35097 3737
rect 35687 3711 35713 3737
rect 36975 3711 37001 3737
rect 37647 3711 37673 3737
rect 38151 3711 38177 3737
rect 38823 3711 38849 3737
rect 38991 3711 39017 3737
rect 2074 3515 2100 3541
rect 2136 3515 2162 3541
rect 2198 3515 2224 3541
rect 2260 3515 2286 3541
rect 2322 3515 2348 3541
rect 2384 3515 2410 3541
rect 2446 3515 2472 3541
rect 2508 3515 2534 3541
rect 7074 3515 7100 3541
rect 7136 3515 7162 3541
rect 7198 3515 7224 3541
rect 7260 3515 7286 3541
rect 7322 3515 7348 3541
rect 7384 3515 7410 3541
rect 7446 3515 7472 3541
rect 7508 3515 7534 3541
rect 12074 3515 12100 3541
rect 12136 3515 12162 3541
rect 12198 3515 12224 3541
rect 12260 3515 12286 3541
rect 12322 3515 12348 3541
rect 12384 3515 12410 3541
rect 12446 3515 12472 3541
rect 12508 3515 12534 3541
rect 17074 3515 17100 3541
rect 17136 3515 17162 3541
rect 17198 3515 17224 3541
rect 17260 3515 17286 3541
rect 17322 3515 17348 3541
rect 17384 3515 17410 3541
rect 17446 3515 17472 3541
rect 17508 3515 17534 3541
rect 22074 3515 22100 3541
rect 22136 3515 22162 3541
rect 22198 3515 22224 3541
rect 22260 3515 22286 3541
rect 22322 3515 22348 3541
rect 22384 3515 22410 3541
rect 22446 3515 22472 3541
rect 22508 3515 22534 3541
rect 27074 3515 27100 3541
rect 27136 3515 27162 3541
rect 27198 3515 27224 3541
rect 27260 3515 27286 3541
rect 27322 3515 27348 3541
rect 27384 3515 27410 3541
rect 27446 3515 27472 3541
rect 27508 3515 27534 3541
rect 32074 3515 32100 3541
rect 32136 3515 32162 3541
rect 32198 3515 32224 3541
rect 32260 3515 32286 3541
rect 32322 3515 32348 3541
rect 32384 3515 32410 3541
rect 32446 3515 32472 3541
rect 32508 3515 32534 3541
rect 37074 3515 37100 3541
rect 37136 3515 37162 3541
rect 37198 3515 37224 3541
rect 37260 3515 37286 3541
rect 37322 3515 37348 3541
rect 37384 3515 37410 3541
rect 37446 3515 37472 3541
rect 37508 3515 37534 3541
rect 1807 3319 1833 3345
rect 1919 3319 1945 3345
rect 2479 3319 2505 3345
rect 3823 3319 3849 3345
rect 4383 3319 4409 3345
rect 4495 3319 4521 3345
rect 5279 3319 5305 3345
rect 6455 3319 6481 3345
rect 8079 3319 8105 3345
rect 8975 3319 9001 3345
rect 9535 3319 9561 3345
rect 10431 3319 10457 3345
rect 12055 3319 12081 3345
rect 12727 3319 12753 3345
rect 13343 3319 13369 3345
rect 13679 3319 13705 3345
rect 13903 3319 13929 3345
rect 15527 3319 15553 3345
rect 15975 3319 16001 3345
rect 16199 3319 16225 3345
rect 16983 3319 17009 3345
rect 17767 3319 17793 3345
rect 18775 3319 18801 3345
rect 19223 3319 19249 3345
rect 19447 3319 19473 3345
rect 20231 3319 20257 3345
rect 21015 3319 21041 3345
rect 22751 3319 22777 3345
rect 23199 3319 23225 3345
rect 23423 3319 23449 3345
rect 24375 3319 24401 3345
rect 25215 3319 25241 3345
rect 26055 3319 26081 3345
rect 26167 3319 26193 3345
rect 26335 3319 26361 3345
rect 26727 3319 26753 3345
rect 27175 3319 27201 3345
rect 27399 3319 27425 3345
rect 28463 3319 28489 3345
rect 29359 3319 29385 3345
rect 30199 3319 30225 3345
rect 30703 3319 30729 3345
rect 31879 3319 31905 3345
rect 32159 3319 32185 3345
rect 33335 3319 33361 3345
rect 33671 3319 33697 3345
rect 33783 3319 33809 3345
rect 33951 3319 33977 3345
rect 34679 3319 34705 3345
rect 35183 3319 35209 3345
rect 35743 3319 35769 3345
rect 36135 3319 36161 3345
rect 36695 3319 36721 3345
rect 36863 3319 36889 3345
rect 37591 3319 37617 3345
rect 37927 3319 37953 3345
rect 38655 3319 38681 3345
rect 38767 3319 38793 3345
rect 38879 3319 38905 3345
rect 6455 3263 6481 3289
rect 8975 3263 9001 3289
rect 10431 3263 10457 3289
rect 12727 3263 12753 3289
rect 17935 3263 17961 3289
rect 21183 3263 21209 3289
rect 25215 3263 25241 3289
rect 29359 3263 29385 3289
rect 30031 3263 30057 3289
rect 30311 3263 30337 3289
rect 31879 3263 31905 3289
rect 33335 3263 33361 3289
rect 37703 3263 37729 3289
rect 4574 3123 4600 3149
rect 4636 3123 4662 3149
rect 4698 3123 4724 3149
rect 4760 3123 4786 3149
rect 4822 3123 4848 3149
rect 4884 3123 4910 3149
rect 4946 3123 4972 3149
rect 5008 3123 5034 3149
rect 9574 3123 9600 3149
rect 9636 3123 9662 3149
rect 9698 3123 9724 3149
rect 9760 3123 9786 3149
rect 9822 3123 9848 3149
rect 9884 3123 9910 3149
rect 9946 3123 9972 3149
rect 10008 3123 10034 3149
rect 14574 3123 14600 3149
rect 14636 3123 14662 3149
rect 14698 3123 14724 3149
rect 14760 3123 14786 3149
rect 14822 3123 14848 3149
rect 14884 3123 14910 3149
rect 14946 3123 14972 3149
rect 15008 3123 15034 3149
rect 19574 3123 19600 3149
rect 19636 3123 19662 3149
rect 19698 3123 19724 3149
rect 19760 3123 19786 3149
rect 19822 3123 19848 3149
rect 19884 3123 19910 3149
rect 19946 3123 19972 3149
rect 20008 3123 20034 3149
rect 24574 3123 24600 3149
rect 24636 3123 24662 3149
rect 24698 3123 24724 3149
rect 24760 3123 24786 3149
rect 24822 3123 24848 3149
rect 24884 3123 24910 3149
rect 24946 3123 24972 3149
rect 25008 3123 25034 3149
rect 29574 3123 29600 3149
rect 29636 3123 29662 3149
rect 29698 3123 29724 3149
rect 29760 3123 29786 3149
rect 29822 3123 29848 3149
rect 29884 3123 29910 3149
rect 29946 3123 29972 3149
rect 30008 3123 30034 3149
rect 34574 3123 34600 3149
rect 34636 3123 34662 3149
rect 34698 3123 34724 3149
rect 34760 3123 34786 3149
rect 34822 3123 34848 3149
rect 34884 3123 34910 3149
rect 34946 3123 34972 3149
rect 35008 3123 35034 3149
rect 1919 2983 1945 3009
rect 4495 2983 4521 3009
rect 7015 2983 7041 3009
rect 8471 2983 8497 3009
rect 10767 2983 10793 3009
rect 12447 2983 12473 3009
rect 14239 2983 14265 3009
rect 17767 2983 17793 3009
rect 19223 2983 19249 3009
rect 21743 2983 21769 3009
rect 23423 2983 23449 3009
rect 28351 2983 28377 3009
rect 31375 2983 31401 3009
rect 32047 2983 32073 3009
rect 33895 2983 33921 3009
rect 35183 2983 35209 3009
rect 35743 2983 35769 3009
rect 35911 2983 35937 3009
rect 38151 2983 38177 3009
rect 38263 2983 38289 3009
rect 38431 2983 38457 3009
rect 38711 2983 38737 3009
rect 1919 2927 1945 2953
rect 3039 2927 3065 2953
rect 3487 2927 3513 2953
rect 4495 2927 4521 2953
rect 5839 2927 5865 2953
rect 7015 2927 7041 2953
rect 7575 2927 7601 2953
rect 8471 2927 8497 2953
rect 10039 2927 10065 2953
rect 10767 2927 10793 2953
rect 11551 2927 11577 2953
rect 12447 2927 12473 2953
rect 13343 2927 13369 2953
rect 14239 2927 14265 2953
rect 15079 2927 15105 2953
rect 15247 2927 15273 2953
rect 15471 2927 15497 2953
rect 16815 2927 16841 2953
rect 17655 2927 17681 2953
rect 18271 2927 18297 2953
rect 19223 2927 19249 2953
rect 20791 2927 20817 2953
rect 21743 2927 21769 2953
rect 22247 2927 22273 2953
rect 23423 2927 23449 2953
rect 24767 2927 24793 2953
rect 25215 2927 25241 2953
rect 25439 2927 25465 2953
rect 26279 2927 26305 2953
rect 26783 2927 26809 2953
rect 26895 2927 26921 2953
rect 28015 2927 28041 2953
rect 28183 2927 28209 2953
rect 29023 2927 29049 2953
rect 29303 2927 29329 2953
rect 29471 2927 29497 2953
rect 30367 2927 30393 2953
rect 31375 2927 31401 2953
rect 32215 2927 32241 2953
rect 32383 2927 32409 2953
rect 32775 2927 32801 2953
rect 33895 2927 33921 2953
rect 34455 2927 34481 2953
rect 35183 2927 35209 2953
rect 35687 2927 35713 2953
rect 36695 2927 36721 2953
rect 37143 2927 37169 2953
rect 37367 2927 37393 2953
rect 38823 2927 38849 2953
rect 38935 2927 38961 2953
rect 2074 2731 2100 2757
rect 2136 2731 2162 2757
rect 2198 2731 2224 2757
rect 2260 2731 2286 2757
rect 2322 2731 2348 2757
rect 2384 2731 2410 2757
rect 2446 2731 2472 2757
rect 2508 2731 2534 2757
rect 7074 2731 7100 2757
rect 7136 2731 7162 2757
rect 7198 2731 7224 2757
rect 7260 2731 7286 2757
rect 7322 2731 7348 2757
rect 7384 2731 7410 2757
rect 7446 2731 7472 2757
rect 7508 2731 7534 2757
rect 12074 2731 12100 2757
rect 12136 2731 12162 2757
rect 12198 2731 12224 2757
rect 12260 2731 12286 2757
rect 12322 2731 12348 2757
rect 12384 2731 12410 2757
rect 12446 2731 12472 2757
rect 12508 2731 12534 2757
rect 17074 2731 17100 2757
rect 17136 2731 17162 2757
rect 17198 2731 17224 2757
rect 17260 2731 17286 2757
rect 17322 2731 17348 2757
rect 17384 2731 17410 2757
rect 17446 2731 17472 2757
rect 17508 2731 17534 2757
rect 22074 2731 22100 2757
rect 22136 2731 22162 2757
rect 22198 2731 22224 2757
rect 22260 2731 22286 2757
rect 22322 2731 22348 2757
rect 22384 2731 22410 2757
rect 22446 2731 22472 2757
rect 22508 2731 22534 2757
rect 27074 2731 27100 2757
rect 27136 2731 27162 2757
rect 27198 2731 27224 2757
rect 27260 2731 27286 2757
rect 27322 2731 27348 2757
rect 27384 2731 27410 2757
rect 27446 2731 27472 2757
rect 27508 2731 27534 2757
rect 32074 2731 32100 2757
rect 32136 2731 32162 2757
rect 32198 2731 32224 2757
rect 32260 2731 32286 2757
rect 32322 2731 32348 2757
rect 32384 2731 32410 2757
rect 32446 2731 32472 2757
rect 32508 2731 32534 2757
rect 37074 2731 37100 2757
rect 37136 2731 37162 2757
rect 37198 2731 37224 2757
rect 37260 2731 37286 2757
rect 37322 2731 37348 2757
rect 37384 2731 37410 2757
rect 37446 2731 37472 2757
rect 37508 2731 37534 2757
rect 1807 2535 1833 2561
rect 2031 2535 2057 2561
rect 2479 2535 2505 2561
rect 3823 2535 3849 2561
rect 4999 2535 5025 2561
rect 5279 2535 5305 2561
rect 6455 2535 6481 2561
rect 7799 2535 7825 2561
rect 8975 2535 9001 2561
rect 9535 2535 9561 2561
rect 10263 2535 10289 2561
rect 11887 2535 11913 2561
rect 12727 2535 12753 2561
rect 13343 2535 13369 2561
rect 14239 2535 14265 2561
rect 15247 2535 15273 2561
rect 15695 2535 15721 2561
rect 15919 2535 15945 2561
rect 16815 2535 16841 2561
rect 17151 2535 17177 2561
rect 17375 2535 17401 2561
rect 20119 2535 20145 2561
rect 20959 2535 20985 2561
rect 22751 2535 22777 2561
rect 23199 2535 23225 2561
rect 23535 2535 23561 2561
rect 24375 2535 24401 2561
rect 24655 2535 24681 2561
rect 24879 2535 24905 2561
rect 26727 2535 26753 2561
rect 27175 2535 27201 2561
rect 27399 2535 27425 2561
rect 28463 2535 28489 2561
rect 29359 2535 29385 2561
rect 30031 2535 30057 2561
rect 30199 2535 30225 2561
rect 30703 2535 30729 2561
rect 31263 2535 31289 2561
rect 31375 2535 31401 2561
rect 32439 2535 32465 2561
rect 33335 2535 33361 2561
rect 33671 2535 33697 2561
rect 33783 2535 33809 2561
rect 33895 2535 33921 2561
rect 34679 2535 34705 2561
rect 35183 2535 35209 2561
rect 35351 2535 35377 2561
rect 36135 2535 36161 2561
rect 36695 2535 36721 2561
rect 36863 2535 36889 2561
rect 37591 2535 37617 2561
rect 37703 2535 37729 2561
rect 37871 2535 37897 2561
rect 38767 2535 38793 2561
rect 38879 2535 38905 2561
rect 4999 2479 5025 2505
rect 6455 2479 6481 2505
rect 8975 2479 9001 2505
rect 10263 2479 10289 2505
rect 12727 2479 12753 2505
rect 14239 2479 14265 2505
rect 20959 2479 20985 2505
rect 26055 2479 26081 2505
rect 26223 2479 26249 2505
rect 26335 2479 26361 2505
rect 29359 2479 29385 2505
rect 30311 2479 30337 2505
rect 33335 2479 33361 2505
rect 38655 2479 38681 2505
rect 4574 2339 4600 2365
rect 4636 2339 4662 2365
rect 4698 2339 4724 2365
rect 4760 2339 4786 2365
rect 4822 2339 4848 2365
rect 4884 2339 4910 2365
rect 4946 2339 4972 2365
rect 5008 2339 5034 2365
rect 9574 2339 9600 2365
rect 9636 2339 9662 2365
rect 9698 2339 9724 2365
rect 9760 2339 9786 2365
rect 9822 2339 9848 2365
rect 9884 2339 9910 2365
rect 9946 2339 9972 2365
rect 10008 2339 10034 2365
rect 14574 2339 14600 2365
rect 14636 2339 14662 2365
rect 14698 2339 14724 2365
rect 14760 2339 14786 2365
rect 14822 2339 14848 2365
rect 14884 2339 14910 2365
rect 14946 2339 14972 2365
rect 15008 2339 15034 2365
rect 19574 2339 19600 2365
rect 19636 2339 19662 2365
rect 19698 2339 19724 2365
rect 19760 2339 19786 2365
rect 19822 2339 19848 2365
rect 19884 2339 19910 2365
rect 19946 2339 19972 2365
rect 20008 2339 20034 2365
rect 24574 2339 24600 2365
rect 24636 2339 24662 2365
rect 24698 2339 24724 2365
rect 24760 2339 24786 2365
rect 24822 2339 24848 2365
rect 24884 2339 24910 2365
rect 24946 2339 24972 2365
rect 25008 2339 25034 2365
rect 29574 2339 29600 2365
rect 29636 2339 29662 2365
rect 29698 2339 29724 2365
rect 29760 2339 29786 2365
rect 29822 2339 29848 2365
rect 29884 2339 29910 2365
rect 29946 2339 29972 2365
rect 30008 2339 30034 2365
rect 34574 2339 34600 2365
rect 34636 2339 34662 2365
rect 34698 2339 34724 2365
rect 34760 2339 34786 2365
rect 34822 2339 34848 2365
rect 34884 2339 34910 2365
rect 34946 2339 34972 2365
rect 35008 2339 35034 2365
rect 4439 2199 4465 2225
rect 8471 2199 8497 2225
rect 10767 2199 10793 2225
rect 12447 2199 12473 2225
rect 17767 2199 17793 2225
rect 19223 2199 19249 2225
rect 21743 2199 21769 2225
rect 23199 2199 23225 2225
rect 24095 2199 24121 2225
rect 24375 2199 24401 2225
rect 28071 2199 28097 2225
rect 28239 2199 28265 2225
rect 31263 2199 31289 2225
rect 31935 2199 31961 2225
rect 35183 2199 35209 2225
rect 35911 2199 35937 2225
rect 38711 2199 38737 2225
rect 38879 2199 38905 2225
rect 38991 2199 39017 2225
rect 2367 2143 2393 2169
rect 2479 2143 2505 2169
rect 3039 2143 3065 2169
rect 3487 2143 3513 2169
rect 4439 2143 4465 2169
rect 5895 2143 5921 2169
rect 6399 2143 6425 2169
rect 6511 2143 6537 2169
rect 7295 2143 7321 2169
rect 8471 2143 8497 2169
rect 10039 2143 10065 2169
rect 10767 2143 10793 2169
rect 11551 2143 11577 2169
rect 12447 2143 12473 2169
rect 13623 2143 13649 2169
rect 14071 2143 14097 2169
rect 14295 2143 14321 2169
rect 15135 2143 15161 2169
rect 15583 2143 15609 2169
rect 15807 2143 15833 2169
rect 16815 2143 16841 2169
rect 17655 2143 17681 2169
rect 18271 2143 18297 2169
rect 19111 2143 19137 2169
rect 20791 2143 20817 2169
rect 21743 2143 21769 2169
rect 22527 2143 22553 2169
rect 23143 2143 23169 2169
rect 24207 2143 24233 2169
rect 24767 2143 24793 2169
rect 25215 2143 25241 2169
rect 25439 2143 25465 2169
rect 26223 2143 26249 2169
rect 26783 2143 26809 2169
rect 26895 2143 26921 2169
rect 28295 2143 28321 2169
rect 29023 2143 29049 2169
rect 29191 2143 29217 2169
rect 29415 2143 29441 2169
rect 30367 2143 30393 2169
rect 31263 2143 31289 2169
rect 31655 2143 31681 2169
rect 31823 2143 31849 2169
rect 32719 2143 32745 2169
rect 33279 2143 33305 2169
rect 33447 2143 33473 2169
rect 34399 2143 34425 2169
rect 35183 2143 35209 2169
rect 35687 2143 35713 2169
rect 35799 2143 35825 2169
rect 37199 2143 37225 2169
rect 37311 2143 37337 2169
rect 37591 2143 37617 2169
rect 38151 2143 38177 2169
rect 38319 2143 38345 2169
rect 38487 2143 38513 2169
rect 2074 1947 2100 1973
rect 2136 1947 2162 1973
rect 2198 1947 2224 1973
rect 2260 1947 2286 1973
rect 2322 1947 2348 1973
rect 2384 1947 2410 1973
rect 2446 1947 2472 1973
rect 2508 1947 2534 1973
rect 7074 1947 7100 1973
rect 7136 1947 7162 1973
rect 7198 1947 7224 1973
rect 7260 1947 7286 1973
rect 7322 1947 7348 1973
rect 7384 1947 7410 1973
rect 7446 1947 7472 1973
rect 7508 1947 7534 1973
rect 12074 1947 12100 1973
rect 12136 1947 12162 1973
rect 12198 1947 12224 1973
rect 12260 1947 12286 1973
rect 12322 1947 12348 1973
rect 12384 1947 12410 1973
rect 12446 1947 12472 1973
rect 12508 1947 12534 1973
rect 17074 1947 17100 1973
rect 17136 1947 17162 1973
rect 17198 1947 17224 1973
rect 17260 1947 17286 1973
rect 17322 1947 17348 1973
rect 17384 1947 17410 1973
rect 17446 1947 17472 1973
rect 17508 1947 17534 1973
rect 22074 1947 22100 1973
rect 22136 1947 22162 1973
rect 22198 1947 22224 1973
rect 22260 1947 22286 1973
rect 22322 1947 22348 1973
rect 22384 1947 22410 1973
rect 22446 1947 22472 1973
rect 22508 1947 22534 1973
rect 27074 1947 27100 1973
rect 27136 1947 27162 1973
rect 27198 1947 27224 1973
rect 27260 1947 27286 1973
rect 27322 1947 27348 1973
rect 27384 1947 27410 1973
rect 27446 1947 27472 1973
rect 27508 1947 27534 1973
rect 32074 1947 32100 1973
rect 32136 1947 32162 1973
rect 32198 1947 32224 1973
rect 32260 1947 32286 1973
rect 32322 1947 32348 1973
rect 32384 1947 32410 1973
rect 32446 1947 32472 1973
rect 32508 1947 32534 1973
rect 37074 1947 37100 1973
rect 37136 1947 37162 1973
rect 37198 1947 37224 1973
rect 37260 1947 37286 1973
rect 37322 1947 37348 1973
rect 37384 1947 37410 1973
rect 37446 1947 37472 1973
rect 37508 1947 37534 1973
rect 1639 1751 1665 1777
rect 2479 1751 2505 1777
rect 3487 1751 3513 1777
rect 4439 1751 4465 1777
rect 5503 1751 5529 1777
rect 6399 1751 6425 1777
rect 7463 1751 7489 1777
rect 8135 1751 8161 1777
rect 9423 1751 9449 1777
rect 10263 1751 10289 1777
rect 11383 1751 11409 1777
rect 11999 1751 12025 1777
rect 13343 1751 13369 1777
rect 13511 1751 13537 1777
rect 13735 1751 13761 1777
rect 15135 1751 15161 1777
rect 15303 1751 15329 1777
rect 15527 1751 15553 1777
rect 16591 1751 16617 1777
rect 17543 1751 17569 1777
rect 18551 1751 18577 1777
rect 19111 1751 19137 1777
rect 19223 1751 19249 1777
rect 21183 1751 21209 1777
rect 21799 1751 21825 1777
rect 22471 1751 22497 1777
rect 22919 1751 22945 1777
rect 23143 1751 23169 1777
rect 24487 1751 24513 1777
rect 25215 1751 25241 1777
rect 26391 1751 26417 1777
rect 26895 1751 26921 1777
rect 27063 1751 27089 1777
rect 28631 1751 28657 1777
rect 28799 1751 28825 1777
rect 29023 1751 29049 1777
rect 30367 1751 30393 1777
rect 31263 1751 31289 1777
rect 32551 1751 32577 1777
rect 33447 1751 33473 1777
rect 34399 1751 34425 1777
rect 35183 1751 35209 1777
rect 36191 1751 36217 1777
rect 37143 1751 37169 1777
rect 38151 1751 38177 1777
rect 38263 1751 38289 1777
rect 38431 1751 38457 1777
rect 38655 1751 38681 1777
rect 38823 1751 38849 1777
rect 38935 1751 38961 1777
rect 1527 1695 1553 1721
rect 4439 1695 4465 1721
rect 6399 1695 6425 1721
rect 8135 1695 8161 1721
rect 10263 1695 10289 1721
rect 12055 1695 12081 1721
rect 17543 1695 17569 1721
rect 21855 1695 21881 1721
rect 25383 1695 25409 1721
rect 31263 1695 31289 1721
rect 33447 1695 33473 1721
rect 35183 1695 35209 1721
rect 37143 1695 37169 1721
rect 4574 1555 4600 1581
rect 4636 1555 4662 1581
rect 4698 1555 4724 1581
rect 4760 1555 4786 1581
rect 4822 1555 4848 1581
rect 4884 1555 4910 1581
rect 4946 1555 4972 1581
rect 5008 1555 5034 1581
rect 9574 1555 9600 1581
rect 9636 1555 9662 1581
rect 9698 1555 9724 1581
rect 9760 1555 9786 1581
rect 9822 1555 9848 1581
rect 9884 1555 9910 1581
rect 9946 1555 9972 1581
rect 10008 1555 10034 1581
rect 14574 1555 14600 1581
rect 14636 1555 14662 1581
rect 14698 1555 14724 1581
rect 14760 1555 14786 1581
rect 14822 1555 14848 1581
rect 14884 1555 14910 1581
rect 14946 1555 14972 1581
rect 15008 1555 15034 1581
rect 19574 1555 19600 1581
rect 19636 1555 19662 1581
rect 19698 1555 19724 1581
rect 19760 1555 19786 1581
rect 19822 1555 19848 1581
rect 19884 1555 19910 1581
rect 19946 1555 19972 1581
rect 20008 1555 20034 1581
rect 24574 1555 24600 1581
rect 24636 1555 24662 1581
rect 24698 1555 24724 1581
rect 24760 1555 24786 1581
rect 24822 1555 24848 1581
rect 24884 1555 24910 1581
rect 24946 1555 24972 1581
rect 25008 1555 25034 1581
rect 29574 1555 29600 1581
rect 29636 1555 29662 1581
rect 29698 1555 29724 1581
rect 29760 1555 29786 1581
rect 29822 1555 29848 1581
rect 29884 1555 29910 1581
rect 29946 1555 29972 1581
rect 30008 1555 30034 1581
rect 34574 1555 34600 1581
rect 34636 1555 34662 1581
rect 34698 1555 34724 1581
rect 34760 1555 34786 1581
rect 34822 1555 34848 1581
rect 34884 1555 34910 1581
rect 34946 1555 34972 1581
rect 35008 1555 35034 1581
<< metal2 >>
rect 2520 19600 2576 20000
rect 6790 19614 7378 19642
rect 2534 18522 2562 19600
rect 2534 18494 2674 18522
rect 2073 18438 2535 18443
rect 2073 18437 2082 18438
rect 2073 18411 2074 18437
rect 2073 18410 2082 18411
rect 2110 18410 2134 18438
rect 2162 18410 2186 18438
rect 2214 18437 2238 18438
rect 2266 18437 2290 18438
rect 2224 18411 2238 18437
rect 2286 18411 2290 18437
rect 2214 18410 2238 18411
rect 2266 18410 2290 18411
rect 2318 18437 2342 18438
rect 2370 18437 2394 18438
rect 2318 18411 2322 18437
rect 2370 18411 2384 18437
rect 2318 18410 2342 18411
rect 2370 18410 2394 18411
rect 2422 18410 2446 18438
rect 2474 18410 2498 18438
rect 2526 18437 2535 18438
rect 2534 18411 2535 18437
rect 2526 18410 2535 18411
rect 2073 18405 2535 18410
rect 2073 17654 2535 17659
rect 2073 17653 2082 17654
rect 2073 17627 2074 17653
rect 2073 17626 2082 17627
rect 2110 17626 2134 17654
rect 2162 17626 2186 17654
rect 2214 17653 2238 17654
rect 2266 17653 2290 17654
rect 2224 17627 2238 17653
rect 2286 17627 2290 17653
rect 2214 17626 2238 17627
rect 2266 17626 2290 17627
rect 2318 17653 2342 17654
rect 2370 17653 2394 17654
rect 2318 17627 2322 17653
rect 2370 17627 2384 17653
rect 2318 17626 2342 17627
rect 2370 17626 2394 17627
rect 2422 17626 2446 17654
rect 2474 17626 2498 17654
rect 2526 17653 2535 17654
rect 2534 17627 2535 17653
rect 2526 17626 2535 17627
rect 2073 17621 2535 17626
rect 2073 16870 2535 16875
rect 2073 16869 2082 16870
rect 2073 16843 2074 16869
rect 2073 16842 2082 16843
rect 2110 16842 2134 16870
rect 2162 16842 2186 16870
rect 2214 16869 2238 16870
rect 2266 16869 2290 16870
rect 2224 16843 2238 16869
rect 2286 16843 2290 16869
rect 2214 16842 2238 16843
rect 2266 16842 2290 16843
rect 2318 16869 2342 16870
rect 2370 16869 2394 16870
rect 2318 16843 2322 16869
rect 2370 16843 2384 16869
rect 2318 16842 2342 16843
rect 2370 16842 2394 16843
rect 2422 16842 2446 16870
rect 2474 16842 2498 16870
rect 2526 16869 2535 16870
rect 2534 16843 2535 16869
rect 2526 16842 2535 16843
rect 2073 16837 2535 16842
rect 2073 16086 2535 16091
rect 2073 16085 2082 16086
rect 2073 16059 2074 16085
rect 2073 16058 2082 16059
rect 2110 16058 2134 16086
rect 2162 16058 2186 16086
rect 2214 16085 2238 16086
rect 2266 16085 2290 16086
rect 2224 16059 2238 16085
rect 2286 16059 2290 16085
rect 2214 16058 2238 16059
rect 2266 16058 2290 16059
rect 2318 16085 2342 16086
rect 2370 16085 2394 16086
rect 2318 16059 2322 16085
rect 2370 16059 2384 16085
rect 2318 16058 2342 16059
rect 2370 16058 2394 16059
rect 2422 16058 2446 16086
rect 2474 16058 2498 16086
rect 2526 16085 2535 16086
rect 2534 16059 2535 16085
rect 2526 16058 2535 16059
rect 2073 16053 2535 16058
rect 1862 15553 1890 15559
rect 1862 15527 1863 15553
rect 1889 15527 1890 15553
rect 1862 15497 1890 15527
rect 1862 15471 1863 15497
rect 1889 15471 1890 15497
rect 1526 15106 1554 15111
rect 1862 15106 1890 15471
rect 2073 15302 2535 15307
rect 2073 15301 2082 15302
rect 2073 15275 2074 15301
rect 2073 15274 2082 15275
rect 2110 15274 2134 15302
rect 2162 15274 2186 15302
rect 2214 15301 2238 15302
rect 2266 15301 2290 15302
rect 2224 15275 2238 15301
rect 2286 15275 2290 15301
rect 2214 15274 2238 15275
rect 2266 15274 2290 15275
rect 2318 15301 2342 15302
rect 2370 15301 2394 15302
rect 2318 15275 2322 15301
rect 2370 15275 2384 15301
rect 2318 15274 2342 15275
rect 2370 15274 2394 15275
rect 2422 15274 2446 15302
rect 2474 15274 2498 15302
rect 2526 15301 2535 15302
rect 2534 15275 2535 15301
rect 2526 15274 2535 15275
rect 2073 15269 2535 15274
rect 1526 15105 1890 15106
rect 1526 15079 1527 15105
rect 1553 15079 1890 15105
rect 1526 15078 1890 15079
rect 2478 15106 2506 15111
rect 2478 15105 2618 15106
rect 2478 15079 2479 15105
rect 2505 15079 2618 15105
rect 2478 15078 2618 15079
rect 1526 15049 1554 15078
rect 2478 15073 2506 15078
rect 1526 15023 1527 15049
rect 1553 15023 1554 15049
rect 1526 14266 1554 15023
rect 1974 14714 2002 14719
rect 1750 14321 1778 14327
rect 1750 14295 1751 14321
rect 1777 14295 1778 14321
rect 1750 14266 1778 14295
rect 1526 14265 1778 14266
rect 1526 14239 1527 14265
rect 1553 14239 1778 14265
rect 1526 14238 1778 14239
rect 1526 14233 1554 14238
rect 1582 11969 1610 11975
rect 1582 11943 1583 11969
rect 1609 11943 1610 11969
rect 1582 11185 1610 11943
rect 1582 11159 1583 11185
rect 1609 11159 1610 11185
rect 1582 10401 1610 11159
rect 1582 10375 1583 10401
rect 1609 10375 1610 10401
rect 1582 9617 1610 10375
rect 1582 9591 1583 9617
rect 1609 9591 1610 9617
rect 1582 9226 1610 9591
rect 1582 8833 1610 9198
rect 1582 8807 1583 8833
rect 1609 8807 1610 8833
rect 1582 8050 1610 8807
rect 1750 8834 1778 14238
rect 1974 13985 2002 14686
rect 2366 14714 2394 14719
rect 2478 14714 2506 14719
rect 2366 14713 2478 14714
rect 2366 14687 2367 14713
rect 2393 14687 2478 14713
rect 2366 14686 2478 14687
rect 2366 14681 2394 14686
rect 2478 14667 2506 14686
rect 2073 14518 2535 14523
rect 2073 14517 2082 14518
rect 2073 14491 2074 14517
rect 2073 14490 2082 14491
rect 2110 14490 2134 14518
rect 2162 14490 2186 14518
rect 2214 14517 2238 14518
rect 2266 14517 2290 14518
rect 2224 14491 2238 14517
rect 2286 14491 2290 14517
rect 2214 14490 2238 14491
rect 2266 14490 2290 14491
rect 2318 14517 2342 14518
rect 2370 14517 2394 14518
rect 2318 14491 2322 14517
rect 2370 14491 2384 14517
rect 2318 14490 2342 14491
rect 2370 14490 2394 14491
rect 2422 14490 2446 14518
rect 2474 14490 2498 14518
rect 2526 14517 2535 14518
rect 2534 14491 2535 14517
rect 2526 14490 2535 14491
rect 2073 14485 2535 14490
rect 2478 14322 2506 14327
rect 2590 14322 2618 15078
rect 2646 14714 2674 18494
rect 4573 18046 5035 18051
rect 4573 18045 4582 18046
rect 4573 18019 4574 18045
rect 4573 18018 4582 18019
rect 4610 18018 4634 18046
rect 4662 18018 4686 18046
rect 4714 18045 4738 18046
rect 4766 18045 4790 18046
rect 4724 18019 4738 18045
rect 4786 18019 4790 18045
rect 4714 18018 4738 18019
rect 4766 18018 4790 18019
rect 4818 18045 4842 18046
rect 4870 18045 4894 18046
rect 4818 18019 4822 18045
rect 4870 18019 4884 18045
rect 4818 18018 4842 18019
rect 4870 18018 4894 18019
rect 4922 18018 4946 18046
rect 4974 18018 4998 18046
rect 5026 18045 5035 18046
rect 5034 18019 5035 18045
rect 5026 18018 5035 18019
rect 4573 18013 5035 18018
rect 4573 17262 5035 17267
rect 4573 17261 4582 17262
rect 4573 17235 4574 17261
rect 4573 17234 4582 17235
rect 4610 17234 4634 17262
rect 4662 17234 4686 17262
rect 4714 17261 4738 17262
rect 4766 17261 4790 17262
rect 4724 17235 4738 17261
rect 4786 17235 4790 17261
rect 4714 17234 4738 17235
rect 4766 17234 4790 17235
rect 4818 17261 4842 17262
rect 4870 17261 4894 17262
rect 4818 17235 4822 17261
rect 4870 17235 4884 17261
rect 4818 17234 4842 17235
rect 4870 17234 4894 17235
rect 4922 17234 4946 17262
rect 4974 17234 4998 17262
rect 5026 17261 5035 17262
rect 5034 17235 5035 17261
rect 5026 17234 5035 17235
rect 4573 17229 5035 17234
rect 4573 16478 5035 16483
rect 4573 16477 4582 16478
rect 4573 16451 4574 16477
rect 4573 16450 4582 16451
rect 4610 16450 4634 16478
rect 4662 16450 4686 16478
rect 4714 16477 4738 16478
rect 4766 16477 4790 16478
rect 4724 16451 4738 16477
rect 4786 16451 4790 16477
rect 4714 16450 4738 16451
rect 4766 16450 4790 16451
rect 4818 16477 4842 16478
rect 4870 16477 4894 16478
rect 4818 16451 4822 16477
rect 4870 16451 4884 16477
rect 4818 16450 4842 16451
rect 4870 16450 4894 16451
rect 4922 16450 4946 16478
rect 4974 16450 4998 16478
rect 5026 16477 5035 16478
rect 5034 16451 5035 16477
rect 5026 16450 5035 16451
rect 4573 16445 5035 16450
rect 4573 15694 5035 15699
rect 4573 15693 4582 15694
rect 4573 15667 4574 15693
rect 4573 15666 4582 15667
rect 4610 15666 4634 15694
rect 4662 15666 4686 15694
rect 4714 15693 4738 15694
rect 4766 15693 4790 15694
rect 4724 15667 4738 15693
rect 4786 15667 4790 15693
rect 4714 15666 4738 15667
rect 4766 15666 4790 15667
rect 4818 15693 4842 15694
rect 4870 15693 4894 15694
rect 4818 15667 4822 15693
rect 4870 15667 4884 15693
rect 4818 15666 4842 15667
rect 4870 15666 4894 15667
rect 4922 15666 4946 15694
rect 4974 15666 4998 15694
rect 5026 15693 5035 15694
rect 5034 15667 5035 15693
rect 5026 15666 5035 15667
rect 4573 15661 5035 15666
rect 4494 15553 4522 15559
rect 4494 15527 4495 15553
rect 4521 15527 4522 15553
rect 2646 14681 2674 14686
rect 2758 15497 2786 15503
rect 2758 15471 2759 15497
rect 2785 15471 2786 15497
rect 2758 14713 2786 15471
rect 2758 14687 2759 14713
rect 2785 14687 2786 14713
rect 2478 14321 2618 14322
rect 2478 14295 2479 14321
rect 2505 14295 2618 14321
rect 2478 14294 2618 14295
rect 2478 14289 2506 14294
rect 1974 13959 1975 13985
rect 2001 13959 2002 13985
rect 1974 13929 2002 13959
rect 1974 13903 1975 13929
rect 2001 13903 2002 13929
rect 1806 13537 1834 13543
rect 1806 13511 1807 13537
rect 1833 13511 1834 13537
rect 1806 13454 1834 13511
rect 1974 13537 2002 13903
rect 2073 13734 2535 13739
rect 2073 13733 2082 13734
rect 2073 13707 2074 13733
rect 2073 13706 2082 13707
rect 2110 13706 2134 13734
rect 2162 13706 2186 13734
rect 2214 13733 2238 13734
rect 2266 13733 2290 13734
rect 2224 13707 2238 13733
rect 2286 13707 2290 13733
rect 2214 13706 2238 13707
rect 2266 13706 2290 13707
rect 2318 13733 2342 13734
rect 2370 13733 2394 13734
rect 2318 13707 2322 13733
rect 2370 13707 2384 13733
rect 2318 13706 2342 13707
rect 2370 13706 2394 13707
rect 2422 13706 2446 13734
rect 2474 13706 2498 13734
rect 2526 13733 2535 13734
rect 2534 13707 2535 13733
rect 2526 13706 2535 13707
rect 2073 13701 2535 13706
rect 1974 13511 1975 13537
rect 2001 13511 2002 13537
rect 1974 13454 2002 13511
rect 2478 13538 2506 13543
rect 2590 13538 2618 14294
rect 2478 13537 2618 13538
rect 2478 13511 2479 13537
rect 2505 13511 2618 13537
rect 2478 13510 2618 13511
rect 2478 13505 2506 13510
rect 1806 13426 2002 13454
rect 2590 13454 2618 13510
rect 2758 14322 2786 14687
rect 2758 13929 2786 14294
rect 2758 13903 2759 13929
rect 2785 13903 2786 13929
rect 2758 13454 2786 13903
rect 3318 15497 3346 15503
rect 3318 15471 3319 15497
rect 3345 15471 3346 15497
rect 3318 14713 3346 15471
rect 4494 15497 4522 15527
rect 4494 15471 4495 15497
rect 4521 15471 4522 15497
rect 3318 14687 3319 14713
rect 3345 14687 3346 14713
rect 3318 14322 3346 14687
rect 3318 13929 3346 14294
rect 3822 15106 3850 15111
rect 3822 14322 3850 15078
rect 4382 15106 4410 15111
rect 4494 15106 4522 15471
rect 6118 15497 6146 15503
rect 6118 15471 6119 15497
rect 6145 15471 6146 15497
rect 4382 15105 4522 15106
rect 4382 15079 4383 15105
rect 4409 15079 4495 15105
rect 4521 15079 4522 15105
rect 4382 15078 4522 15079
rect 4382 15073 4410 15078
rect 4494 14769 4522 15078
rect 5558 15106 5586 15111
rect 5558 15059 5586 15078
rect 5838 15106 5866 15111
rect 6118 15106 6146 15471
rect 5838 15105 5922 15106
rect 5838 15079 5839 15105
rect 5865 15079 5922 15105
rect 5838 15078 5922 15079
rect 5838 15073 5866 15078
rect 4573 14910 5035 14915
rect 4573 14909 4582 14910
rect 4573 14883 4574 14909
rect 4573 14882 4582 14883
rect 4610 14882 4634 14910
rect 4662 14882 4686 14910
rect 4714 14909 4738 14910
rect 4766 14909 4790 14910
rect 4724 14883 4738 14909
rect 4786 14883 4790 14909
rect 4714 14882 4738 14883
rect 4766 14882 4790 14883
rect 4818 14909 4842 14910
rect 4870 14909 4894 14910
rect 4818 14883 4822 14909
rect 4870 14883 4884 14909
rect 4818 14882 4842 14883
rect 4870 14882 4894 14883
rect 4922 14882 4946 14910
rect 4974 14882 4998 14910
rect 5026 14909 5035 14910
rect 5034 14883 5035 14909
rect 5026 14882 5035 14883
rect 4573 14877 5035 14882
rect 4494 14743 4495 14769
rect 4521 14743 4522 14769
rect 4494 14713 4522 14743
rect 4494 14687 4495 14713
rect 4521 14687 4522 14713
rect 3822 14275 3850 14294
rect 4382 14322 4410 14327
rect 4494 14322 4522 14687
rect 4382 14321 4522 14322
rect 4382 14295 4383 14321
rect 4409 14295 4495 14321
rect 4521 14295 4522 14321
rect 4382 14294 4522 14295
rect 4382 14289 4410 14294
rect 3318 13903 3319 13929
rect 3345 13903 3346 13929
rect 3318 13897 3346 13903
rect 4494 13985 4522 14294
rect 5558 14714 5586 14719
rect 5558 14321 5586 14686
rect 5558 14295 5559 14321
rect 5585 14295 5586 14321
rect 4573 14126 5035 14131
rect 4573 14125 4582 14126
rect 4573 14099 4574 14125
rect 4573 14098 4582 14099
rect 4610 14098 4634 14126
rect 4662 14098 4686 14126
rect 4714 14125 4738 14126
rect 4766 14125 4790 14126
rect 4724 14099 4738 14125
rect 4786 14099 4790 14125
rect 4714 14098 4738 14099
rect 4766 14098 4790 14099
rect 4818 14125 4842 14126
rect 4870 14125 4894 14126
rect 4818 14099 4822 14125
rect 4870 14099 4884 14125
rect 4818 14098 4842 14099
rect 4870 14098 4894 14099
rect 4922 14098 4946 14126
rect 4974 14098 4998 14126
rect 5026 14125 5035 14126
rect 5034 14099 5035 14125
rect 5026 14098 5035 14099
rect 4573 14093 5035 14098
rect 4494 13959 4495 13985
rect 4521 13959 4522 13985
rect 4494 13929 4522 13959
rect 4494 13903 4495 13929
rect 4521 13903 4522 13929
rect 2590 13426 2786 13454
rect 1974 13146 2002 13426
rect 1806 12754 1834 12759
rect 1974 12754 2002 13118
rect 2366 13146 2394 13151
rect 2590 13146 2618 13151
rect 2394 13145 2618 13146
rect 2394 13119 2591 13145
rect 2617 13119 2618 13145
rect 2394 13118 2618 13119
rect 2366 13080 2394 13118
rect 2073 12950 2535 12955
rect 2073 12949 2082 12950
rect 2073 12923 2074 12949
rect 2073 12922 2082 12923
rect 2110 12922 2134 12950
rect 2162 12922 2186 12950
rect 2214 12949 2238 12950
rect 2266 12949 2290 12950
rect 2224 12923 2238 12949
rect 2286 12923 2290 12949
rect 2214 12922 2238 12923
rect 2266 12922 2290 12923
rect 2318 12949 2342 12950
rect 2370 12949 2394 12950
rect 2318 12923 2322 12949
rect 2370 12923 2384 12949
rect 2318 12922 2342 12923
rect 2370 12922 2394 12923
rect 2422 12922 2446 12950
rect 2474 12922 2498 12950
rect 2526 12949 2535 12950
rect 2534 12923 2535 12949
rect 2526 12922 2535 12923
rect 2073 12917 2535 12922
rect 2590 12922 2618 13118
rect 2758 13145 2786 13426
rect 3822 13537 3850 13543
rect 3822 13511 3823 13537
rect 3849 13511 3850 13537
rect 2758 13119 2759 13145
rect 2785 13119 2786 13145
rect 2590 12894 2730 12922
rect 1806 12753 2002 12754
rect 1806 12727 1807 12753
rect 1833 12727 1975 12753
rect 2001 12727 2002 12753
rect 1806 12726 2002 12727
rect 1806 12721 1834 12726
rect 1974 12721 2002 12726
rect 2478 12754 2506 12759
rect 2478 12707 2506 12726
rect 1750 8768 1778 8806
rect 1918 12361 1946 12367
rect 1918 12335 1919 12361
rect 1945 12335 1946 12361
rect 1918 11577 1946 12335
rect 2073 12166 2535 12171
rect 2073 12165 2082 12166
rect 2073 12139 2074 12165
rect 2073 12138 2082 12139
rect 2110 12138 2134 12166
rect 2162 12138 2186 12166
rect 2214 12165 2238 12166
rect 2266 12165 2290 12166
rect 2224 12139 2238 12165
rect 2286 12139 2290 12165
rect 2214 12138 2238 12139
rect 2266 12138 2290 12139
rect 2318 12165 2342 12166
rect 2370 12165 2394 12166
rect 2318 12139 2322 12165
rect 2370 12139 2384 12165
rect 2318 12138 2342 12139
rect 2370 12138 2394 12139
rect 2422 12138 2446 12166
rect 2474 12138 2498 12166
rect 2526 12165 2535 12166
rect 2534 12139 2535 12165
rect 2526 12138 2535 12139
rect 2073 12133 2535 12138
rect 2478 11970 2506 11975
rect 2702 11970 2730 12894
rect 2758 12754 2786 13119
rect 2758 12721 2786 12726
rect 3598 13146 3626 13151
rect 3822 13146 3850 13511
rect 4382 13538 4410 13543
rect 4494 13538 4522 13903
rect 4382 13537 4522 13538
rect 4382 13511 4383 13537
rect 4409 13511 4495 13537
rect 4521 13511 4522 13537
rect 4382 13510 4522 13511
rect 4382 13505 4410 13510
rect 3598 13145 3850 13146
rect 3598 13119 3599 13145
rect 3625 13119 3850 13145
rect 3598 13118 3850 13119
rect 3038 12417 3066 12423
rect 3038 12391 3039 12417
rect 3065 12391 3066 12417
rect 3038 12361 3066 12391
rect 3038 12335 3039 12361
rect 3065 12335 3066 12361
rect 3038 11970 3066 12335
rect 2478 11969 3066 11970
rect 2478 11943 2479 11969
rect 2505 11943 3066 11969
rect 2478 11942 3066 11943
rect 2478 11913 2506 11942
rect 2478 11887 2479 11913
rect 2505 11887 2506 11913
rect 2478 11881 2506 11887
rect 1918 11551 1919 11577
rect 1945 11551 1946 11577
rect 1918 10793 1946 11551
rect 2073 11382 2535 11387
rect 2073 11381 2082 11382
rect 2073 11355 2074 11381
rect 2073 11354 2082 11355
rect 2110 11354 2134 11382
rect 2162 11354 2186 11382
rect 2214 11381 2238 11382
rect 2266 11381 2290 11382
rect 2224 11355 2238 11381
rect 2286 11355 2290 11381
rect 2214 11354 2238 11355
rect 2266 11354 2290 11355
rect 2318 11381 2342 11382
rect 2370 11381 2394 11382
rect 2318 11355 2322 11381
rect 2370 11355 2384 11381
rect 2318 11354 2342 11355
rect 2370 11354 2394 11355
rect 2422 11354 2446 11382
rect 2474 11354 2498 11382
rect 2526 11381 2535 11382
rect 2534 11355 2535 11381
rect 2526 11354 2535 11355
rect 2073 11349 2535 11354
rect 2590 11242 2618 11942
rect 2478 11214 2618 11242
rect 3038 11633 3066 11942
rect 3038 11607 3039 11633
rect 3065 11607 3066 11633
rect 3038 11577 3066 11607
rect 3038 11551 3039 11577
rect 3065 11551 3066 11577
rect 2478 11185 2506 11214
rect 2478 11159 2479 11185
rect 2505 11159 2506 11185
rect 2478 11129 2506 11159
rect 2478 11103 2479 11129
rect 2505 11103 2506 11129
rect 2478 11097 2506 11103
rect 1918 10767 1919 10793
rect 1945 10767 1946 10793
rect 1918 10009 1946 10767
rect 3038 10849 3066 11551
rect 3038 10823 3039 10849
rect 3065 10823 3066 10849
rect 3038 10793 3066 10823
rect 3038 10767 3039 10793
rect 3065 10767 3066 10793
rect 2073 10598 2535 10603
rect 2073 10597 2082 10598
rect 2073 10571 2074 10597
rect 2073 10570 2082 10571
rect 2110 10570 2134 10598
rect 2162 10570 2186 10598
rect 2214 10597 2238 10598
rect 2266 10597 2290 10598
rect 2224 10571 2238 10597
rect 2286 10571 2290 10597
rect 2214 10570 2238 10571
rect 2266 10570 2290 10571
rect 2318 10597 2342 10598
rect 2370 10597 2394 10598
rect 2318 10571 2322 10597
rect 2370 10571 2384 10597
rect 2318 10570 2342 10571
rect 2370 10570 2394 10571
rect 2422 10570 2446 10598
rect 2474 10570 2498 10598
rect 2526 10597 2535 10598
rect 2534 10571 2535 10597
rect 2526 10570 2535 10571
rect 2073 10565 2535 10570
rect 2478 10401 2506 10407
rect 2478 10375 2479 10401
rect 2505 10375 2506 10401
rect 2478 10345 2506 10375
rect 2478 10319 2479 10345
rect 2505 10319 2506 10345
rect 2478 10290 2506 10319
rect 2478 10262 2618 10290
rect 1918 9983 1919 10009
rect 1945 9983 1946 10009
rect 1918 9226 1946 9983
rect 2073 9814 2535 9819
rect 2073 9813 2082 9814
rect 2073 9787 2074 9813
rect 2073 9786 2082 9787
rect 2110 9786 2134 9814
rect 2162 9786 2186 9814
rect 2214 9813 2238 9814
rect 2266 9813 2290 9814
rect 2224 9787 2238 9813
rect 2286 9787 2290 9813
rect 2214 9786 2238 9787
rect 2266 9786 2290 9787
rect 2318 9813 2342 9814
rect 2370 9813 2394 9814
rect 2318 9787 2322 9813
rect 2370 9787 2384 9813
rect 2318 9786 2342 9787
rect 2370 9786 2394 9787
rect 2422 9786 2446 9814
rect 2474 9786 2498 9814
rect 2526 9813 2535 9814
rect 2534 9787 2535 9813
rect 2526 9786 2535 9787
rect 2073 9781 2535 9786
rect 1918 8442 1946 9198
rect 2478 9618 2506 9623
rect 2590 9618 2618 10262
rect 2478 9617 2618 9618
rect 2478 9591 2479 9617
rect 2505 9591 2618 9617
rect 2478 9590 2618 9591
rect 3038 10065 3066 10767
rect 3038 10039 3039 10065
rect 3065 10039 3066 10065
rect 3038 10009 3066 10039
rect 3038 9983 3039 10009
rect 3065 9983 3066 10009
rect 2478 9561 2506 9590
rect 2478 9535 2479 9561
rect 2505 9535 2506 9561
rect 2478 9226 2506 9535
rect 2478 9193 2506 9198
rect 3038 9281 3066 9983
rect 3038 9255 3039 9281
rect 3065 9255 3066 9281
rect 3038 9226 3066 9255
rect 2073 9030 2535 9035
rect 2073 9029 2082 9030
rect 2073 9003 2074 9029
rect 2073 9002 2082 9003
rect 2110 9002 2134 9030
rect 2162 9002 2186 9030
rect 2214 9029 2238 9030
rect 2266 9029 2290 9030
rect 2224 9003 2238 9029
rect 2286 9003 2290 9029
rect 2214 9002 2238 9003
rect 2266 9002 2290 9003
rect 2318 9029 2342 9030
rect 2370 9029 2394 9030
rect 2318 9003 2322 9029
rect 2370 9003 2384 9029
rect 2318 9002 2342 9003
rect 2370 9002 2394 9003
rect 2422 9002 2446 9030
rect 2474 9002 2498 9030
rect 2526 9029 2535 9030
rect 2534 9003 2535 9029
rect 2526 9002 2535 9003
rect 2073 8997 2535 9002
rect 1918 8409 1946 8414
rect 1974 8834 2002 8839
rect 1582 8049 1890 8050
rect 1582 8023 1583 8049
rect 1609 8023 1890 8049
rect 1582 8022 1890 8023
rect 1582 8017 1610 8022
rect 1022 7994 1050 7999
rect 1022 400 1050 7966
rect 1862 7657 1890 8022
rect 1862 7631 1863 7657
rect 1889 7631 1890 7657
rect 1862 7625 1890 7631
rect 1974 8049 2002 8806
rect 2310 8834 2338 8839
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 2310 8442 2338 8806
rect 2534 8498 2562 8503
rect 2534 8442 2562 8470
rect 2310 8441 2562 8442
rect 2310 8415 2311 8441
rect 2337 8415 2535 8441
rect 2561 8415 2562 8441
rect 2310 8414 2562 8415
rect 2310 8409 2338 8414
rect 2534 8409 2562 8414
rect 2073 8246 2535 8251
rect 2073 8245 2082 8246
rect 2073 8219 2074 8245
rect 2073 8218 2082 8219
rect 2110 8218 2134 8246
rect 2162 8218 2186 8246
rect 2214 8245 2238 8246
rect 2266 8245 2290 8246
rect 2224 8219 2238 8245
rect 2286 8219 2290 8245
rect 2214 8218 2238 8219
rect 2266 8218 2290 8219
rect 2318 8245 2342 8246
rect 2370 8245 2394 8246
rect 2318 8219 2322 8245
rect 2370 8219 2384 8245
rect 2318 8218 2342 8219
rect 2370 8218 2394 8219
rect 2422 8218 2446 8246
rect 2474 8218 2498 8246
rect 2526 8245 2535 8246
rect 2534 8219 2535 8245
rect 2526 8218 2535 8219
rect 2073 8213 2535 8218
rect 1974 8023 1975 8049
rect 2001 8023 2002 8049
rect 1974 7994 2002 8023
rect 2926 8106 2954 8111
rect 2254 7994 2282 7999
rect 1974 7993 2282 7994
rect 1974 7967 2255 7993
rect 2281 7967 2282 7993
rect 1974 7966 2282 7967
rect 1806 7266 1834 7271
rect 1806 7219 1834 7238
rect 1806 6482 1834 6487
rect 1974 6482 2002 7966
rect 2254 7961 2282 7966
rect 2590 7658 2618 7663
rect 2073 7462 2535 7467
rect 2073 7461 2082 7462
rect 2073 7435 2074 7461
rect 2073 7434 2082 7435
rect 2110 7434 2134 7462
rect 2162 7434 2186 7462
rect 2214 7461 2238 7462
rect 2266 7461 2290 7462
rect 2224 7435 2238 7461
rect 2286 7435 2290 7461
rect 2214 7434 2238 7435
rect 2266 7434 2290 7435
rect 2318 7461 2342 7462
rect 2370 7461 2394 7462
rect 2318 7435 2322 7461
rect 2370 7435 2384 7461
rect 2318 7434 2342 7435
rect 2370 7434 2394 7435
rect 2422 7434 2446 7462
rect 2474 7434 2498 7462
rect 2526 7461 2535 7462
rect 2534 7435 2535 7461
rect 2526 7434 2535 7435
rect 2073 7429 2535 7434
rect 2590 7378 2618 7630
rect 2366 7350 2618 7378
rect 2030 7266 2058 7271
rect 2030 7219 2058 7238
rect 2366 7266 2394 7350
rect 2366 6874 2394 7238
rect 2478 7266 2506 7271
rect 2478 7265 2618 7266
rect 2478 7239 2479 7265
rect 2505 7239 2618 7265
rect 2478 7238 2618 7239
rect 2478 7233 2506 7238
rect 2478 6874 2506 6879
rect 2366 6873 2506 6874
rect 2366 6847 2367 6873
rect 2393 6847 2479 6873
rect 2505 6847 2506 6873
rect 2366 6846 2506 6847
rect 2366 6841 2394 6846
rect 2478 6841 2506 6846
rect 2073 6678 2535 6683
rect 2073 6677 2082 6678
rect 2073 6651 2074 6677
rect 2073 6650 2082 6651
rect 2110 6650 2134 6678
rect 2162 6650 2186 6678
rect 2214 6677 2238 6678
rect 2266 6677 2290 6678
rect 2224 6651 2238 6677
rect 2286 6651 2290 6677
rect 2214 6650 2238 6651
rect 2266 6650 2290 6651
rect 2318 6677 2342 6678
rect 2370 6677 2394 6678
rect 2318 6651 2322 6677
rect 2370 6651 2384 6677
rect 2318 6650 2342 6651
rect 2370 6650 2394 6651
rect 2422 6650 2446 6678
rect 2474 6650 2498 6678
rect 2526 6677 2535 6678
rect 2534 6651 2535 6677
rect 2526 6650 2535 6651
rect 2073 6645 2535 6650
rect 1806 6481 2002 6482
rect 1806 6455 1807 6481
rect 1833 6455 1975 6481
rect 2001 6455 2002 6481
rect 1806 6454 2002 6455
rect 1806 6449 1834 6454
rect 1974 6145 2002 6454
rect 1974 6119 1975 6145
rect 2001 6119 2002 6145
rect 1974 6089 2002 6119
rect 1974 6063 1975 6089
rect 2001 6063 2002 6089
rect 1806 5698 1834 5703
rect 1974 5698 2002 6063
rect 2478 6482 2506 6487
rect 2590 6482 2618 7238
rect 2478 6481 2618 6482
rect 2478 6455 2479 6481
rect 2505 6455 2618 6481
rect 2478 6454 2618 6455
rect 2478 6090 2506 6454
rect 2590 6090 2618 6095
rect 2478 6062 2590 6090
rect 2073 5894 2535 5899
rect 2073 5893 2082 5894
rect 2073 5867 2074 5893
rect 2073 5866 2082 5867
rect 2110 5866 2134 5894
rect 2162 5866 2186 5894
rect 2214 5893 2238 5894
rect 2266 5893 2290 5894
rect 2224 5867 2238 5893
rect 2286 5867 2290 5893
rect 2214 5866 2238 5867
rect 2266 5866 2290 5867
rect 2318 5893 2342 5894
rect 2370 5893 2394 5894
rect 2318 5867 2322 5893
rect 2370 5867 2384 5893
rect 2318 5866 2342 5867
rect 2370 5866 2394 5867
rect 2422 5866 2446 5894
rect 2474 5866 2498 5894
rect 2526 5893 2535 5894
rect 2534 5867 2535 5893
rect 2526 5866 2535 5867
rect 2073 5861 2535 5866
rect 1806 5697 2002 5698
rect 1806 5671 1807 5697
rect 1833 5671 1975 5697
rect 2001 5671 2002 5697
rect 1806 5670 2002 5671
rect 1806 5665 1834 5670
rect 1974 5361 2002 5670
rect 2478 5698 2506 5703
rect 2590 5698 2618 6062
rect 2478 5697 2618 5698
rect 2478 5671 2479 5697
rect 2505 5671 2618 5697
rect 2478 5670 2618 5671
rect 2478 5665 2506 5670
rect 1974 5335 1975 5361
rect 2001 5335 2002 5361
rect 1974 5305 2002 5335
rect 1974 5279 1975 5305
rect 2001 5279 2002 5305
rect 1974 5273 2002 5279
rect 2073 5110 2535 5115
rect 2073 5109 2082 5110
rect 2073 5083 2074 5109
rect 2073 5082 2082 5083
rect 2110 5082 2134 5110
rect 2162 5082 2186 5110
rect 2214 5109 2238 5110
rect 2266 5109 2290 5110
rect 2224 5083 2238 5109
rect 2286 5083 2290 5109
rect 2214 5082 2238 5083
rect 2266 5082 2290 5083
rect 2318 5109 2342 5110
rect 2370 5109 2394 5110
rect 2318 5083 2322 5109
rect 2370 5083 2384 5109
rect 2318 5082 2342 5083
rect 2370 5082 2394 5083
rect 2422 5082 2446 5110
rect 2474 5082 2498 5110
rect 2526 5109 2535 5110
rect 2534 5083 2535 5109
rect 2526 5082 2535 5083
rect 2073 5077 2535 5082
rect 1806 4914 1834 4919
rect 1918 4914 1946 4919
rect 1806 4913 1946 4914
rect 1806 4887 1807 4913
rect 1833 4887 1919 4913
rect 1945 4887 1946 4913
rect 1806 4886 1946 4887
rect 1806 4881 1834 4886
rect 1862 4577 1890 4886
rect 1918 4881 1946 4886
rect 2478 4914 2506 4919
rect 2478 4913 2618 4914
rect 2478 4887 2479 4913
rect 2505 4887 2618 4913
rect 2478 4886 2618 4887
rect 2478 4881 2506 4886
rect 1862 4551 1863 4577
rect 1889 4551 1890 4577
rect 1862 4521 1890 4551
rect 1862 4495 1863 4521
rect 1889 4495 1890 4521
rect 1862 4214 1890 4495
rect 2073 4326 2535 4331
rect 2073 4325 2082 4326
rect 2073 4299 2074 4325
rect 2073 4298 2082 4299
rect 2110 4298 2134 4326
rect 2162 4298 2186 4326
rect 2214 4325 2238 4326
rect 2266 4325 2290 4326
rect 2224 4299 2238 4325
rect 2286 4299 2290 4325
rect 2214 4298 2238 4299
rect 2266 4298 2290 4299
rect 2318 4325 2342 4326
rect 2370 4325 2394 4326
rect 2318 4299 2322 4325
rect 2370 4299 2384 4325
rect 2318 4298 2342 4299
rect 2370 4298 2394 4299
rect 2422 4298 2446 4326
rect 2474 4298 2498 4326
rect 2526 4325 2535 4326
rect 2534 4299 2535 4325
rect 2526 4298 2535 4299
rect 2073 4293 2535 4298
rect 1862 4186 2002 4214
rect 1806 4130 1834 4135
rect 1918 4130 1946 4135
rect 1974 4130 2002 4186
rect 2590 4186 2618 4886
rect 1806 4129 2002 4130
rect 1806 4103 1807 4129
rect 1833 4103 1919 4129
rect 1945 4103 2002 4129
rect 1806 4102 2002 4103
rect 2478 4130 2506 4135
rect 2590 4130 2618 4158
rect 2478 4129 2618 4130
rect 2478 4103 2479 4129
rect 2505 4103 2618 4129
rect 2478 4102 2618 4103
rect 1806 4097 1834 4102
rect 1918 3793 1946 4102
rect 2478 4097 2506 4102
rect 1918 3767 1919 3793
rect 1945 3767 1946 3793
rect 1918 3737 1946 3767
rect 1918 3711 1919 3737
rect 1945 3711 1946 3737
rect 1806 3346 1834 3351
rect 1918 3346 1946 3711
rect 2073 3542 2535 3547
rect 2073 3541 2082 3542
rect 2073 3515 2074 3541
rect 2073 3514 2082 3515
rect 2110 3514 2134 3542
rect 2162 3514 2186 3542
rect 2214 3541 2238 3542
rect 2266 3541 2290 3542
rect 2224 3515 2238 3541
rect 2286 3515 2290 3541
rect 2214 3514 2238 3515
rect 2266 3514 2290 3515
rect 2318 3541 2342 3542
rect 2370 3541 2394 3542
rect 2318 3515 2322 3541
rect 2370 3515 2384 3541
rect 2318 3514 2342 3515
rect 2370 3514 2394 3515
rect 2422 3514 2446 3542
rect 2474 3514 2498 3542
rect 2526 3541 2535 3542
rect 2534 3515 2535 3541
rect 2526 3514 2535 3515
rect 2073 3509 2535 3514
rect 1806 3345 1946 3346
rect 1806 3319 1807 3345
rect 1833 3319 1919 3345
rect 1945 3319 1946 3345
rect 1806 3318 1946 3319
rect 1806 3313 1834 3318
rect 1918 3009 1946 3318
rect 2478 3346 2506 3351
rect 2478 3299 2506 3318
rect 1918 2983 1919 3009
rect 1945 2983 1946 3009
rect 1918 2953 1946 2983
rect 1918 2927 1919 2953
rect 1945 2927 1946 2953
rect 1806 2562 1834 2567
rect 1918 2562 1946 2927
rect 2073 2758 2535 2763
rect 2073 2757 2082 2758
rect 2073 2731 2074 2757
rect 2073 2730 2082 2731
rect 2110 2730 2134 2758
rect 2162 2730 2186 2758
rect 2214 2757 2238 2758
rect 2266 2757 2290 2758
rect 2224 2731 2238 2757
rect 2286 2731 2290 2757
rect 2214 2730 2238 2731
rect 2266 2730 2290 2731
rect 2318 2757 2342 2758
rect 2370 2757 2394 2758
rect 2318 2731 2322 2757
rect 2370 2731 2384 2757
rect 2318 2730 2342 2731
rect 2370 2730 2394 2731
rect 2422 2730 2446 2758
rect 2474 2730 2498 2758
rect 2526 2757 2535 2758
rect 2534 2731 2535 2757
rect 2526 2730 2535 2731
rect 2073 2725 2535 2730
rect 2030 2562 2058 2567
rect 1806 2561 2058 2562
rect 1806 2535 1807 2561
rect 1833 2535 2031 2561
rect 2057 2535 2058 2561
rect 1806 2534 2058 2535
rect 1806 2529 1834 2534
rect 1638 2506 1666 2511
rect 1638 1777 1666 2478
rect 2030 2226 2058 2534
rect 2478 2562 2506 2567
rect 2478 2515 2506 2534
rect 2030 2193 2058 2198
rect 2478 2226 2506 2231
rect 2366 2170 2394 2175
rect 2478 2170 2506 2198
rect 2366 2169 2506 2170
rect 2366 2143 2367 2169
rect 2393 2143 2479 2169
rect 2505 2143 2506 2169
rect 2366 2142 2506 2143
rect 2366 2137 2394 2142
rect 2478 2137 2506 2142
rect 2073 1974 2535 1979
rect 2073 1973 2082 1974
rect 2073 1947 2074 1973
rect 2073 1946 2082 1947
rect 2110 1946 2134 1974
rect 2162 1946 2186 1974
rect 2214 1973 2238 1974
rect 2266 1973 2290 1974
rect 2224 1947 2238 1973
rect 2286 1947 2290 1973
rect 2214 1946 2238 1947
rect 2266 1946 2290 1947
rect 2318 1973 2342 1974
rect 2370 1973 2394 1974
rect 2318 1947 2322 1973
rect 2370 1947 2384 1973
rect 2318 1946 2342 1947
rect 2370 1946 2394 1947
rect 2422 1946 2446 1974
rect 2474 1946 2498 1974
rect 2526 1973 2535 1974
rect 2534 1947 2535 1973
rect 2526 1946 2535 1947
rect 2073 1941 2535 1946
rect 1638 1751 1639 1777
rect 1665 1751 1666 1777
rect 1526 1722 1554 1727
rect 1638 1722 1666 1751
rect 2478 1778 2506 1783
rect 2478 1777 2562 1778
rect 2478 1751 2479 1777
rect 2505 1751 2562 1777
rect 2478 1750 2562 1751
rect 2478 1745 2506 1750
rect 1526 1721 1666 1722
rect 1526 1695 1527 1721
rect 1553 1695 1666 1721
rect 1526 1694 1666 1695
rect 1526 1689 1554 1694
rect 2478 1666 2506 1671
rect 2478 400 2506 1638
rect 2534 1498 2562 1750
rect 2926 1722 2954 8078
rect 3038 7713 3066 9198
rect 3038 7687 3039 7713
rect 3065 7687 3066 7713
rect 3038 7658 3066 7687
rect 3038 7592 3066 7630
rect 3598 12361 3626 13118
rect 3598 12335 3599 12361
rect 3625 12335 3626 12361
rect 3598 11577 3626 12335
rect 3598 11551 3599 11577
rect 3625 11551 3626 11577
rect 3598 10793 3626 11551
rect 3598 10767 3599 10793
rect 3625 10767 3626 10793
rect 3598 10009 3626 10767
rect 3822 12753 3850 13118
rect 3822 12727 3823 12753
rect 3849 12727 3850 12753
rect 3822 11969 3850 12727
rect 3822 11943 3823 11969
rect 3849 11943 3850 11969
rect 3822 11185 3850 11943
rect 3822 11159 3823 11185
rect 3849 11159 3850 11185
rect 3822 10401 3850 11159
rect 3822 10375 3823 10401
rect 3849 10375 3850 10401
rect 3822 10369 3850 10375
rect 4494 13201 4522 13510
rect 5502 13537 5530 13543
rect 5502 13511 5503 13537
rect 5529 13511 5530 13537
rect 4573 13342 5035 13347
rect 4573 13341 4582 13342
rect 4573 13315 4574 13341
rect 4573 13314 4582 13315
rect 4610 13314 4634 13342
rect 4662 13314 4686 13342
rect 4714 13341 4738 13342
rect 4766 13341 4790 13342
rect 4724 13315 4738 13341
rect 4786 13315 4790 13341
rect 4714 13314 4738 13315
rect 4766 13314 4790 13315
rect 4818 13341 4842 13342
rect 4870 13341 4894 13342
rect 4818 13315 4822 13341
rect 4870 13315 4884 13341
rect 4818 13314 4842 13315
rect 4870 13314 4894 13315
rect 4922 13314 4946 13342
rect 4974 13314 4998 13342
rect 5026 13341 5035 13342
rect 5034 13315 5035 13341
rect 5026 13314 5035 13315
rect 4573 13309 5035 13314
rect 4494 13175 4495 13201
rect 4521 13175 4522 13201
rect 4494 13145 4522 13175
rect 4494 13119 4495 13145
rect 4521 13119 4522 13145
rect 4494 12417 4522 13119
rect 4998 12753 5026 12759
rect 4998 12727 4999 12753
rect 5025 12727 5026 12753
rect 4998 12697 5026 12727
rect 5502 12754 5530 13511
rect 5558 13454 5586 14295
rect 5838 14322 5866 14327
rect 5894 14322 5922 15078
rect 6118 14826 6146 15078
rect 6118 14793 6146 14798
rect 6454 15105 6482 15111
rect 6454 15079 6455 15105
rect 6481 15079 6482 15105
rect 6118 14714 6146 14719
rect 6118 14667 6146 14686
rect 5838 14321 5922 14322
rect 5838 14295 5839 14321
rect 5865 14295 5922 14321
rect 5838 14294 5922 14295
rect 5838 14289 5866 14294
rect 5838 13538 5866 13543
rect 5894 13538 5922 14294
rect 6454 14321 6482 15079
rect 6454 14295 6455 14321
rect 6481 14295 6482 14321
rect 5838 13537 5894 13538
rect 5838 13511 5839 13537
rect 5865 13511 5894 13537
rect 5838 13510 5894 13511
rect 5838 13505 5866 13510
rect 5894 13505 5922 13510
rect 6118 13929 6146 13935
rect 6118 13903 6119 13929
rect 6145 13903 6146 13929
rect 5558 13426 5642 13454
rect 5558 12754 5586 12759
rect 5502 12726 5558 12754
rect 5558 12707 5586 12726
rect 4998 12671 4999 12697
rect 5025 12671 5026 12697
rect 4998 12642 5026 12671
rect 4998 12614 5138 12642
rect 4573 12558 5035 12563
rect 4573 12557 4582 12558
rect 4573 12531 4574 12557
rect 4573 12530 4582 12531
rect 4610 12530 4634 12558
rect 4662 12530 4686 12558
rect 4714 12557 4738 12558
rect 4766 12557 4790 12558
rect 4724 12531 4738 12557
rect 4786 12531 4790 12557
rect 4714 12530 4738 12531
rect 4766 12530 4790 12531
rect 4818 12557 4842 12558
rect 4870 12557 4894 12558
rect 4818 12531 4822 12557
rect 4870 12531 4884 12557
rect 4818 12530 4842 12531
rect 4870 12530 4894 12531
rect 4922 12530 4946 12558
rect 4974 12530 4998 12558
rect 5026 12557 5035 12558
rect 5034 12531 5035 12557
rect 5026 12530 5035 12531
rect 4573 12525 5035 12530
rect 5110 12474 5138 12614
rect 4494 12391 4495 12417
rect 4521 12391 4522 12417
rect 4494 12361 4522 12391
rect 4494 12335 4495 12361
rect 4521 12335 4522 12361
rect 4494 11633 4522 12335
rect 4998 12446 5138 12474
rect 4998 11969 5026 12446
rect 4998 11943 4999 11969
rect 5025 11943 5026 11969
rect 4998 11913 5026 11943
rect 5558 11970 5586 11975
rect 5614 11970 5642 13426
rect 6118 13145 6146 13903
rect 6118 13119 6119 13145
rect 6145 13119 6146 13145
rect 6118 12754 6146 13119
rect 6118 12362 6146 12726
rect 6118 12315 6146 12334
rect 6454 13538 6482 14295
rect 6454 12753 6482 13510
rect 6454 12727 6455 12753
rect 6481 12727 6482 12753
rect 6454 12698 6482 12727
rect 5558 11969 5642 11970
rect 5558 11943 5559 11969
rect 5585 11943 5642 11969
rect 5558 11942 5642 11943
rect 5558 11937 5586 11942
rect 4998 11887 4999 11913
rect 5025 11887 5026 11913
rect 4998 11858 5026 11887
rect 4998 11830 5138 11858
rect 4573 11774 5035 11779
rect 4573 11773 4582 11774
rect 4573 11747 4574 11773
rect 4573 11746 4582 11747
rect 4610 11746 4634 11774
rect 4662 11746 4686 11774
rect 4714 11773 4738 11774
rect 4766 11773 4790 11774
rect 4724 11747 4738 11773
rect 4786 11747 4790 11773
rect 4714 11746 4738 11747
rect 4766 11746 4790 11747
rect 4818 11773 4842 11774
rect 4870 11773 4894 11774
rect 4818 11747 4822 11773
rect 4870 11747 4884 11773
rect 4818 11746 4842 11747
rect 4870 11746 4894 11747
rect 4922 11746 4946 11774
rect 4974 11746 4998 11774
rect 5026 11773 5035 11774
rect 5034 11747 5035 11773
rect 5026 11746 5035 11747
rect 4573 11741 5035 11746
rect 5110 11690 5138 11830
rect 4494 11607 4495 11633
rect 4521 11607 4522 11633
rect 4494 11577 4522 11607
rect 4494 11551 4495 11577
rect 4521 11551 4522 11577
rect 4494 10849 4522 11551
rect 4998 11662 5138 11690
rect 4998 11185 5026 11662
rect 5614 11578 5642 11942
rect 6454 11969 6482 12670
rect 6454 11943 6455 11969
rect 6481 11943 6482 11969
rect 6454 11913 6482 11943
rect 6454 11887 6455 11913
rect 6481 11887 6482 11913
rect 6454 11774 6482 11887
rect 6398 11746 6482 11774
rect 5838 11578 5866 11583
rect 5614 11577 5866 11578
rect 5614 11551 5839 11577
rect 5865 11551 5866 11577
rect 5614 11550 5866 11551
rect 4998 11159 4999 11185
rect 5025 11159 5026 11185
rect 4998 11129 5026 11159
rect 4998 11103 4999 11129
rect 5025 11103 5026 11129
rect 4998 11074 5026 11103
rect 5558 11186 5586 11191
rect 5614 11186 5642 11550
rect 5558 11185 5642 11186
rect 5558 11159 5559 11185
rect 5585 11159 5642 11185
rect 5558 11158 5642 11159
rect 4998 11046 5138 11074
rect 4573 10990 5035 10995
rect 4573 10989 4582 10990
rect 4573 10963 4574 10989
rect 4573 10962 4582 10963
rect 4610 10962 4634 10990
rect 4662 10962 4686 10990
rect 4714 10989 4738 10990
rect 4766 10989 4790 10990
rect 4724 10963 4738 10989
rect 4786 10963 4790 10989
rect 4714 10962 4738 10963
rect 4766 10962 4790 10963
rect 4818 10989 4842 10990
rect 4870 10989 4894 10990
rect 4818 10963 4822 10989
rect 4870 10963 4884 10989
rect 4818 10962 4842 10963
rect 4870 10962 4894 10963
rect 4922 10962 4946 10990
rect 4974 10962 4998 10990
rect 5026 10989 5035 10990
rect 5034 10963 5035 10989
rect 5026 10962 5035 10963
rect 4573 10957 5035 10962
rect 5110 10906 5138 11046
rect 4494 10823 4495 10849
rect 4521 10823 4522 10849
rect 4494 10793 4522 10823
rect 4494 10767 4495 10793
rect 4521 10767 4522 10793
rect 3598 9983 3599 10009
rect 3625 9983 3626 10009
rect 3598 9225 3626 9983
rect 4494 10065 4522 10767
rect 4998 10878 5138 10906
rect 4998 10401 5026 10878
rect 4998 10375 4999 10401
rect 5025 10375 5026 10401
rect 4998 10345 5026 10375
rect 4998 10319 4999 10345
rect 5025 10319 5026 10345
rect 4998 10290 5026 10319
rect 5558 10401 5586 11158
rect 5558 10375 5559 10401
rect 5585 10375 5586 10401
rect 4998 10262 5138 10290
rect 4573 10206 5035 10211
rect 4573 10205 4582 10206
rect 4573 10179 4574 10205
rect 4573 10178 4582 10179
rect 4610 10178 4634 10206
rect 4662 10178 4686 10206
rect 4714 10205 4738 10206
rect 4766 10205 4790 10206
rect 4724 10179 4738 10205
rect 4786 10179 4790 10205
rect 4714 10178 4738 10179
rect 4766 10178 4790 10179
rect 4818 10205 4842 10206
rect 4870 10205 4894 10206
rect 4818 10179 4822 10205
rect 4870 10179 4884 10205
rect 4818 10178 4842 10179
rect 4870 10178 4894 10179
rect 4922 10178 4946 10206
rect 4974 10178 4998 10206
rect 5026 10205 5035 10206
rect 5034 10179 5035 10205
rect 5026 10178 5035 10179
rect 4573 10173 5035 10178
rect 5110 10122 5138 10262
rect 4494 10039 4495 10065
rect 4521 10039 4522 10065
rect 4494 10010 4522 10039
rect 4998 10094 5138 10122
rect 4998 10010 5026 10094
rect 4494 10009 5026 10010
rect 4494 9983 4495 10009
rect 4521 9983 5026 10009
rect 4494 9982 5026 9983
rect 3598 9199 3599 9225
rect 3625 9199 3626 9225
rect 3598 8442 3626 9199
rect 3934 9617 3962 9623
rect 3934 9591 3935 9617
rect 3961 9591 3962 9617
rect 3598 7657 3626 8414
rect 3598 7631 3599 7657
rect 3625 7631 3626 7657
rect 3038 6873 3066 6879
rect 3038 6847 3039 6873
rect 3065 6847 3066 6873
rect 3038 6090 3066 6847
rect 3598 6873 3626 7631
rect 3598 6847 3599 6873
rect 3625 6847 3626 6873
rect 3598 6818 3626 6847
rect 3598 6785 3626 6790
rect 3710 8890 3738 8895
rect 3038 5305 3066 6062
rect 3598 6090 3626 6095
rect 3598 6043 3626 6062
rect 3038 5279 3039 5305
rect 3065 5279 3066 5305
rect 3038 5273 3066 5279
rect 3430 5305 3458 5311
rect 3430 5279 3431 5305
rect 3457 5279 3458 5305
rect 3038 4521 3066 4527
rect 3038 4495 3039 4521
rect 3065 4495 3066 4521
rect 3038 4186 3066 4495
rect 3430 4521 3458 5279
rect 3430 4495 3431 4521
rect 3457 4495 3458 4521
rect 3430 4354 3458 4495
rect 3430 4326 3626 4354
rect 3038 3737 3066 4158
rect 3542 4242 3570 4247
rect 3038 3711 3039 3737
rect 3065 3711 3066 3737
rect 3038 3346 3066 3711
rect 3038 2953 3066 3318
rect 3038 2927 3039 2953
rect 3065 2927 3066 2953
rect 3038 2562 3066 2927
rect 3038 2170 3066 2534
rect 3038 2123 3066 2142
rect 3486 3737 3514 3743
rect 3486 3711 3487 3737
rect 3513 3711 3514 3737
rect 3486 2953 3514 3711
rect 3486 2927 3487 2953
rect 3513 2927 3514 2953
rect 3486 2170 3514 2927
rect 3486 1834 3514 2142
rect 3486 1777 3514 1806
rect 3486 1751 3487 1777
rect 3513 1751 3514 1777
rect 3486 1745 3514 1751
rect 2926 1689 2954 1694
rect 2534 1465 2562 1470
rect 1008 0 1064 400
rect 2464 0 2520 400
rect 3542 378 3570 4214
rect 3598 4130 3626 4326
rect 3710 4242 3738 8862
rect 3934 8833 3962 9591
rect 3934 8807 3935 8833
rect 3961 8807 3962 8833
rect 3934 8049 3962 8807
rect 4270 9281 4298 9287
rect 4270 9255 4271 9281
rect 4297 9255 4298 9281
rect 4270 9225 4298 9255
rect 4270 9199 4271 9225
rect 4297 9199 4298 9225
rect 4270 8834 4298 9199
rect 4494 9226 4522 9982
rect 4998 9617 5026 9982
rect 4998 9591 4999 9617
rect 5025 9591 5026 9617
rect 4998 9562 5026 9591
rect 4998 9515 5026 9534
rect 5558 9617 5586 10375
rect 5558 9591 5559 9617
rect 5585 9591 5586 9617
rect 4573 9422 5035 9427
rect 4573 9421 4582 9422
rect 4573 9395 4574 9421
rect 4573 9394 4582 9395
rect 4610 9394 4634 9422
rect 4662 9394 4686 9422
rect 4714 9421 4738 9422
rect 4766 9421 4790 9422
rect 4724 9395 4738 9421
rect 4786 9395 4790 9421
rect 4714 9394 4738 9395
rect 4766 9394 4790 9395
rect 4818 9421 4842 9422
rect 4870 9421 4894 9422
rect 4818 9395 4822 9421
rect 4870 9395 4884 9421
rect 4818 9394 4842 9395
rect 4870 9394 4894 9395
rect 4922 9394 4946 9422
rect 4974 9394 4998 9422
rect 5026 9421 5035 9422
rect 5034 9395 5035 9421
rect 5026 9394 5035 9395
rect 4573 9389 5035 9394
rect 4494 9193 4522 9198
rect 4494 8834 4522 8839
rect 4270 8833 4494 8834
rect 4270 8807 4271 8833
rect 4297 8807 4494 8833
rect 4270 8806 4494 8807
rect 3934 8023 3935 8049
rect 3961 8023 3962 8049
rect 3934 7574 3962 8023
rect 4214 8498 4242 8503
rect 4270 8498 4298 8806
rect 4494 8768 4522 8806
rect 5558 8833 5586 9591
rect 5558 8807 5559 8833
rect 5585 8807 5586 8833
rect 4573 8638 5035 8643
rect 4573 8637 4582 8638
rect 4573 8611 4574 8637
rect 4573 8610 4582 8611
rect 4610 8610 4634 8638
rect 4662 8610 4686 8638
rect 4714 8637 4738 8638
rect 4766 8637 4790 8638
rect 4724 8611 4738 8637
rect 4786 8611 4790 8637
rect 4714 8610 4738 8611
rect 4766 8610 4790 8611
rect 4818 8637 4842 8638
rect 4870 8637 4894 8638
rect 4818 8611 4822 8637
rect 4870 8611 4884 8637
rect 4818 8610 4842 8611
rect 4870 8610 4894 8611
rect 4922 8610 4946 8638
rect 4974 8610 4998 8638
rect 5026 8637 5035 8638
rect 5034 8611 5035 8637
rect 5026 8610 5035 8611
rect 4573 8605 5035 8610
rect 4242 8497 4298 8498
rect 4242 8471 4271 8497
rect 4297 8471 4298 8497
rect 4242 8470 4298 8471
rect 4214 8441 4242 8470
rect 4270 8465 4298 8470
rect 4214 8415 4215 8441
rect 4241 8415 4242 8441
rect 4214 8050 4242 8415
rect 4270 8050 4298 8055
rect 4214 8049 4298 8050
rect 4214 8023 4271 8049
rect 4297 8023 4298 8049
rect 4214 8022 4298 8023
rect 4214 7714 4242 8022
rect 4270 8017 4298 8022
rect 4494 8049 4522 8055
rect 4494 8023 4495 8049
rect 4521 8023 4522 8049
rect 4270 7714 4298 7719
rect 4214 7713 4298 7714
rect 4214 7687 4271 7713
rect 4297 7687 4298 7713
rect 4214 7686 4298 7687
rect 4214 7657 4242 7686
rect 4214 7631 4215 7657
rect 4241 7631 4242 7657
rect 4214 7625 4242 7631
rect 4270 7574 4298 7686
rect 4494 7574 4522 8023
rect 5558 8049 5586 8807
rect 5558 8023 5559 8049
rect 5585 8023 5586 8049
rect 4573 7854 5035 7859
rect 4573 7853 4582 7854
rect 4573 7827 4574 7853
rect 4573 7826 4582 7827
rect 4610 7826 4634 7854
rect 4662 7826 4686 7854
rect 4714 7853 4738 7854
rect 4766 7853 4790 7854
rect 4724 7827 4738 7853
rect 4786 7827 4790 7853
rect 4714 7826 4738 7827
rect 4766 7826 4790 7827
rect 4818 7853 4842 7854
rect 4870 7853 4894 7854
rect 4818 7827 4822 7853
rect 4870 7827 4884 7853
rect 4818 7826 4842 7827
rect 4870 7826 4894 7827
rect 4922 7826 4946 7854
rect 4974 7826 4998 7854
rect 5026 7853 5035 7854
rect 5034 7827 5035 7853
rect 5026 7826 5035 7827
rect 4573 7821 5035 7826
rect 5558 7574 5586 8023
rect 3934 7546 4130 7574
rect 4270 7546 5026 7574
rect 4102 7265 4130 7546
rect 4102 7239 4103 7265
rect 4129 7239 4130 7265
rect 4102 6818 4130 7239
rect 4494 6929 4522 7546
rect 4998 7265 5026 7546
rect 4998 7239 4999 7265
rect 5025 7239 5026 7265
rect 4998 7209 5026 7239
rect 4998 7183 4999 7209
rect 5025 7183 5026 7209
rect 4998 7177 5026 7183
rect 5278 7546 5586 7574
rect 5838 10793 5866 11550
rect 5838 10767 5839 10793
rect 5865 10767 5866 10793
rect 5838 10009 5866 10767
rect 6398 11578 6426 11746
rect 6510 11578 6538 11583
rect 6398 11577 6538 11578
rect 6398 11551 6399 11577
rect 6425 11551 6511 11577
rect 6537 11551 6538 11577
rect 6398 11550 6538 11551
rect 6398 11185 6426 11550
rect 6510 11545 6538 11550
rect 6398 11159 6399 11185
rect 6425 11159 6426 11185
rect 6398 11129 6426 11159
rect 6398 11103 6399 11129
rect 6425 11103 6426 11129
rect 6398 10794 6426 11103
rect 6510 10794 6538 10799
rect 6398 10793 6538 10794
rect 6398 10767 6399 10793
rect 6425 10767 6511 10793
rect 6537 10767 6538 10793
rect 6398 10766 6538 10767
rect 6398 10761 6426 10766
rect 5838 9983 5839 10009
rect 5865 9983 5866 10009
rect 5838 9225 5866 9983
rect 6454 10401 6482 10766
rect 6510 10761 6538 10766
rect 6454 10375 6455 10401
rect 6481 10375 6482 10401
rect 6454 10345 6482 10375
rect 6454 10319 6455 10345
rect 6481 10319 6482 10345
rect 5838 9199 5839 9225
rect 5865 9199 5866 9225
rect 5838 8441 5866 9199
rect 5838 8415 5839 8441
rect 5865 8415 5866 8441
rect 5838 7657 5866 8415
rect 5894 9954 5922 9959
rect 5894 7994 5922 9926
rect 6454 9617 6482 10319
rect 6454 9591 6455 9617
rect 6481 9591 6482 9617
rect 6454 9562 6482 9591
rect 6454 9515 6482 9534
rect 5950 8834 5978 8839
rect 5950 8787 5978 8806
rect 6230 8834 6258 8839
rect 6230 8778 6258 8806
rect 6790 8834 6818 19614
rect 7350 19530 7378 19614
rect 7504 19600 7560 20000
rect 12488 19600 12544 20000
rect 17472 19600 17528 20000
rect 22456 19600 22512 20000
rect 27440 19600 27496 20000
rect 31934 19614 32298 19642
rect 7518 19530 7546 19600
rect 7350 19502 7546 19530
rect 12502 18522 12530 19600
rect 17486 18522 17514 19600
rect 22470 18522 22498 19600
rect 27454 18522 27482 19600
rect 12502 18494 12642 18522
rect 17486 18494 17626 18522
rect 22470 18494 22610 18522
rect 27454 18494 27594 18522
rect 7073 18438 7535 18443
rect 7073 18437 7082 18438
rect 7073 18411 7074 18437
rect 7073 18410 7082 18411
rect 7110 18410 7134 18438
rect 7162 18410 7186 18438
rect 7214 18437 7238 18438
rect 7266 18437 7290 18438
rect 7224 18411 7238 18437
rect 7286 18411 7290 18437
rect 7214 18410 7238 18411
rect 7266 18410 7290 18411
rect 7318 18437 7342 18438
rect 7370 18437 7394 18438
rect 7318 18411 7322 18437
rect 7370 18411 7384 18437
rect 7318 18410 7342 18411
rect 7370 18410 7394 18411
rect 7422 18410 7446 18438
rect 7474 18410 7498 18438
rect 7526 18437 7535 18438
rect 7534 18411 7535 18437
rect 7526 18410 7535 18411
rect 7073 18405 7535 18410
rect 12073 18438 12535 18443
rect 12073 18437 12082 18438
rect 12073 18411 12074 18437
rect 12073 18410 12082 18411
rect 12110 18410 12134 18438
rect 12162 18410 12186 18438
rect 12214 18437 12238 18438
rect 12266 18437 12290 18438
rect 12224 18411 12238 18437
rect 12286 18411 12290 18437
rect 12214 18410 12238 18411
rect 12266 18410 12290 18411
rect 12318 18437 12342 18438
rect 12370 18437 12394 18438
rect 12318 18411 12322 18437
rect 12370 18411 12384 18437
rect 12318 18410 12342 18411
rect 12370 18410 12394 18411
rect 12422 18410 12446 18438
rect 12474 18410 12498 18438
rect 12526 18437 12535 18438
rect 12534 18411 12535 18437
rect 12526 18410 12535 18411
rect 12073 18405 12535 18410
rect 12614 18354 12642 18494
rect 17073 18438 17535 18443
rect 17073 18437 17082 18438
rect 17073 18411 17074 18437
rect 17073 18410 17082 18411
rect 17110 18410 17134 18438
rect 17162 18410 17186 18438
rect 17214 18437 17238 18438
rect 17266 18437 17290 18438
rect 17224 18411 17238 18437
rect 17286 18411 17290 18437
rect 17214 18410 17238 18411
rect 17266 18410 17290 18411
rect 17318 18437 17342 18438
rect 17370 18437 17394 18438
rect 17318 18411 17322 18437
rect 17370 18411 17384 18437
rect 17318 18410 17342 18411
rect 17370 18410 17394 18411
rect 17422 18410 17446 18438
rect 17474 18410 17498 18438
rect 17526 18437 17535 18438
rect 17534 18411 17535 18437
rect 17526 18410 17535 18411
rect 17073 18405 17535 18410
rect 12558 18326 12642 18354
rect 11102 18241 11130 18247
rect 11102 18215 11103 18241
rect 11129 18215 11130 18241
rect 9573 18046 10035 18051
rect 9573 18045 9582 18046
rect 9573 18019 9574 18045
rect 9573 18018 9582 18019
rect 9610 18018 9634 18046
rect 9662 18018 9686 18046
rect 9714 18045 9738 18046
rect 9766 18045 9790 18046
rect 9724 18019 9738 18045
rect 9786 18019 9790 18045
rect 9714 18018 9738 18019
rect 9766 18018 9790 18019
rect 9818 18045 9842 18046
rect 9870 18045 9894 18046
rect 9818 18019 9822 18045
rect 9870 18019 9884 18045
rect 9818 18018 9842 18019
rect 9870 18018 9894 18019
rect 9922 18018 9946 18046
rect 9974 18018 9998 18046
rect 10026 18045 10035 18046
rect 10034 18019 10035 18045
rect 10026 18018 10035 18019
rect 9573 18013 10035 18018
rect 9254 17850 9282 17855
rect 7073 17654 7535 17659
rect 7073 17653 7082 17654
rect 7073 17627 7074 17653
rect 7073 17626 7082 17627
rect 7110 17626 7134 17654
rect 7162 17626 7186 17654
rect 7214 17653 7238 17654
rect 7266 17653 7290 17654
rect 7224 17627 7238 17653
rect 7286 17627 7290 17653
rect 7214 17626 7238 17627
rect 7266 17626 7290 17627
rect 7318 17653 7342 17654
rect 7370 17653 7394 17654
rect 7318 17627 7322 17653
rect 7370 17627 7384 17653
rect 7318 17626 7342 17627
rect 7370 17626 7394 17627
rect 7422 17626 7446 17654
rect 7474 17626 7498 17654
rect 7526 17653 7535 17654
rect 7534 17627 7535 17653
rect 7526 17626 7535 17627
rect 7073 17621 7535 17626
rect 9254 17457 9282 17822
rect 9814 17850 9842 17855
rect 10262 17850 10290 17855
rect 10486 17850 10514 17855
rect 9814 17803 9842 17822
rect 10206 17849 10514 17850
rect 10206 17823 10263 17849
rect 10289 17823 10487 17849
rect 10513 17823 10514 17849
rect 10206 17822 10514 17823
rect 9254 17431 9255 17457
rect 9281 17431 9282 17457
rect 7073 16870 7535 16875
rect 7073 16869 7082 16870
rect 7073 16843 7074 16869
rect 7073 16842 7082 16843
rect 7110 16842 7134 16870
rect 7162 16842 7186 16870
rect 7214 16869 7238 16870
rect 7266 16869 7290 16870
rect 7224 16843 7238 16869
rect 7286 16843 7290 16869
rect 7214 16842 7238 16843
rect 7266 16842 7290 16843
rect 7318 16869 7342 16870
rect 7370 16869 7394 16870
rect 7318 16843 7322 16869
rect 7370 16843 7384 16869
rect 7318 16842 7342 16843
rect 7370 16842 7394 16843
rect 7422 16842 7446 16870
rect 7474 16842 7498 16870
rect 7526 16869 7535 16870
rect 7534 16843 7535 16869
rect 7526 16842 7535 16843
rect 7073 16837 7535 16842
rect 7798 16674 7826 16679
rect 7073 16086 7535 16091
rect 7073 16085 7082 16086
rect 7073 16059 7074 16085
rect 7073 16058 7082 16059
rect 7110 16058 7134 16086
rect 7162 16058 7186 16086
rect 7214 16085 7238 16086
rect 7266 16085 7290 16086
rect 7224 16059 7238 16085
rect 7286 16059 7290 16085
rect 7214 16058 7238 16059
rect 7266 16058 7290 16059
rect 7318 16085 7342 16086
rect 7370 16085 7394 16086
rect 7318 16059 7322 16085
rect 7370 16059 7384 16085
rect 7318 16058 7342 16059
rect 7370 16058 7394 16059
rect 7422 16058 7446 16086
rect 7474 16058 7498 16086
rect 7526 16085 7535 16086
rect 7534 16059 7535 16085
rect 7526 16058 7535 16059
rect 7073 16053 7535 16058
rect 7014 15553 7042 15559
rect 7014 15527 7015 15553
rect 7041 15527 7042 15553
rect 7014 15497 7042 15527
rect 7014 15471 7015 15497
rect 7041 15471 7042 15497
rect 6790 8801 6818 8806
rect 6902 14826 6930 14831
rect 6902 14658 6930 14798
rect 6230 8777 6314 8778
rect 6230 8751 6231 8777
rect 6257 8751 6314 8777
rect 6230 8750 6314 8751
rect 6230 8745 6258 8750
rect 6286 8442 6314 8750
rect 6510 8442 6538 8447
rect 6286 8441 6538 8442
rect 6286 8415 6287 8441
rect 6313 8415 6511 8441
rect 6537 8415 6538 8441
rect 6286 8414 6538 8415
rect 5894 7961 5922 7966
rect 6230 8049 6258 8055
rect 6230 8023 6231 8049
rect 6257 8023 6258 8049
rect 6230 7993 6258 8023
rect 6230 7967 6231 7993
rect 6257 7967 6258 7993
rect 5838 7631 5839 7657
rect 5865 7631 5866 7657
rect 5838 7574 5866 7631
rect 6230 7658 6258 7967
rect 6230 7625 6258 7630
rect 6286 7658 6314 8414
rect 6510 8409 6538 8414
rect 6510 7658 6538 7663
rect 6286 7657 6538 7658
rect 6286 7631 6287 7657
rect 6313 7631 6511 7657
rect 6537 7631 6538 7657
rect 6286 7630 6538 7631
rect 6286 7625 6314 7630
rect 5838 7546 6146 7574
rect 5278 7265 5306 7546
rect 5278 7239 5279 7265
rect 5305 7239 5306 7265
rect 4573 7070 5035 7075
rect 4573 7069 4582 7070
rect 4573 7043 4574 7069
rect 4573 7042 4582 7043
rect 4610 7042 4634 7070
rect 4662 7042 4686 7070
rect 4714 7069 4738 7070
rect 4766 7069 4790 7070
rect 4724 7043 4738 7069
rect 4786 7043 4790 7069
rect 4714 7042 4738 7043
rect 4766 7042 4790 7043
rect 4818 7069 4842 7070
rect 4870 7069 4894 7070
rect 4818 7043 4822 7069
rect 4870 7043 4884 7069
rect 4818 7042 4842 7043
rect 4870 7042 4894 7043
rect 4922 7042 4946 7070
rect 4974 7042 4998 7070
rect 5026 7069 5035 7070
rect 5034 7043 5035 7069
rect 5026 7042 5035 7043
rect 4573 7037 5035 7042
rect 4494 6903 4495 6929
rect 4521 6903 4522 6929
rect 4494 6873 4522 6903
rect 4494 6847 4495 6873
rect 4521 6847 4522 6873
rect 4494 6841 4522 6847
rect 4102 6481 4130 6790
rect 5278 6818 5306 7239
rect 4102 6455 4103 6481
rect 4129 6455 4130 6481
rect 4102 6449 4130 6455
rect 4382 6482 4410 6487
rect 4494 6482 4522 6487
rect 4382 6481 4522 6482
rect 4382 6455 4383 6481
rect 4409 6455 4495 6481
rect 4521 6455 4522 6481
rect 4382 6454 4522 6455
rect 4382 6449 4410 6454
rect 4494 6145 4522 6454
rect 5278 6481 5306 6790
rect 5278 6455 5279 6481
rect 5305 6455 5306 6481
rect 4573 6286 5035 6291
rect 4573 6285 4582 6286
rect 4573 6259 4574 6285
rect 4573 6258 4582 6259
rect 4610 6258 4634 6286
rect 4662 6258 4686 6286
rect 4714 6285 4738 6286
rect 4766 6285 4790 6286
rect 4724 6259 4738 6285
rect 4786 6259 4790 6285
rect 4714 6258 4738 6259
rect 4766 6258 4790 6259
rect 4818 6285 4842 6286
rect 4870 6285 4894 6286
rect 4818 6259 4822 6285
rect 4870 6259 4884 6285
rect 4818 6258 4842 6259
rect 4870 6258 4894 6259
rect 4922 6258 4946 6286
rect 4974 6258 4998 6286
rect 5026 6285 5035 6286
rect 5034 6259 5035 6285
rect 5026 6258 5035 6259
rect 4573 6253 5035 6258
rect 4494 6119 4495 6145
rect 4521 6119 4522 6145
rect 3710 4209 3738 4214
rect 4102 6090 4130 6095
rect 4102 5697 4130 6062
rect 4102 5671 4103 5697
rect 4129 5671 4130 5697
rect 4102 4913 4130 5671
rect 4494 6089 4522 6119
rect 4494 6063 4495 6089
rect 4521 6063 4522 6089
rect 4494 5361 4522 6063
rect 4998 5698 5026 5703
rect 4998 5641 5026 5670
rect 4998 5615 4999 5641
rect 5025 5615 5026 5641
rect 4998 5609 5026 5615
rect 5278 5697 5306 6455
rect 6118 6873 6146 7546
rect 6118 6847 6119 6873
rect 6145 6847 6146 6873
rect 6118 6089 6146 6847
rect 6118 6063 6119 6089
rect 6145 6063 6146 6089
rect 5278 5671 5279 5697
rect 5305 5671 5306 5697
rect 4573 5502 5035 5507
rect 4573 5501 4582 5502
rect 4573 5475 4574 5501
rect 4573 5474 4582 5475
rect 4610 5474 4634 5502
rect 4662 5474 4686 5502
rect 4714 5501 4738 5502
rect 4766 5501 4790 5502
rect 4724 5475 4738 5501
rect 4786 5475 4790 5501
rect 4714 5474 4738 5475
rect 4766 5474 4790 5475
rect 4818 5501 4842 5502
rect 4870 5501 4894 5502
rect 4818 5475 4822 5501
rect 4870 5475 4884 5501
rect 4818 5474 4842 5475
rect 4870 5474 4894 5475
rect 4922 5474 4946 5502
rect 4974 5474 4998 5502
rect 5026 5501 5035 5502
rect 5034 5475 5035 5501
rect 5026 5474 5035 5475
rect 4573 5469 5035 5474
rect 4494 5335 4495 5361
rect 4521 5335 4522 5361
rect 4494 5305 4522 5335
rect 4494 5279 4495 5305
rect 4521 5279 4522 5305
rect 4494 5082 4522 5279
rect 4494 5049 4522 5054
rect 4998 5082 5026 5087
rect 4102 4887 4103 4913
rect 4129 4887 4130 4913
rect 3598 4097 3626 4102
rect 4102 4130 4130 4887
rect 4998 4913 5026 5054
rect 4998 4887 4999 4913
rect 5025 4887 5026 4913
rect 4998 4857 5026 4887
rect 5278 4913 5306 5671
rect 5838 5698 5866 5703
rect 5950 5698 5978 5703
rect 5866 5697 5978 5698
rect 5866 5671 5951 5697
rect 5977 5671 5978 5697
rect 5866 5670 5978 5671
rect 5838 5632 5866 5670
rect 5278 4887 5279 4913
rect 5305 4887 5306 4913
rect 5278 4881 5306 4887
rect 5950 5082 5978 5670
rect 4998 4831 4999 4857
rect 5025 4831 5026 4857
rect 4998 4825 5026 4831
rect 4573 4718 5035 4723
rect 4573 4717 4582 4718
rect 4573 4691 4574 4717
rect 4573 4690 4582 4691
rect 4610 4690 4634 4718
rect 4662 4690 4686 4718
rect 4714 4717 4738 4718
rect 4766 4717 4790 4718
rect 4724 4691 4738 4717
rect 4786 4691 4790 4717
rect 4714 4690 4738 4691
rect 4766 4690 4790 4691
rect 4818 4717 4842 4718
rect 4870 4717 4894 4718
rect 4818 4691 4822 4717
rect 4870 4691 4884 4717
rect 4818 4690 4842 4691
rect 4870 4690 4894 4691
rect 4922 4690 4946 4718
rect 4974 4690 4998 4718
rect 5026 4717 5035 4718
rect 5034 4691 5035 4717
rect 5026 4690 5035 4691
rect 4573 4685 5035 4690
rect 4494 4577 4522 4583
rect 4494 4551 4495 4577
rect 4521 4551 4522 4577
rect 4494 4522 4522 4551
rect 4494 4475 4522 4494
rect 4774 4522 4802 4527
rect 4102 4064 4130 4102
rect 4774 4129 4802 4494
rect 4774 4103 4775 4129
rect 4801 4103 4802 4129
rect 4774 4073 4802 4103
rect 4774 4047 4775 4073
rect 4801 4047 4802 4073
rect 4774 4041 4802 4047
rect 5278 4130 5306 4135
rect 4573 3934 5035 3939
rect 4573 3933 4582 3934
rect 4573 3907 4574 3933
rect 4573 3906 4582 3907
rect 4610 3906 4634 3934
rect 4662 3906 4686 3934
rect 4714 3933 4738 3934
rect 4766 3933 4790 3934
rect 4724 3907 4738 3933
rect 4786 3907 4790 3933
rect 4714 3906 4738 3907
rect 4766 3906 4790 3907
rect 4818 3933 4842 3934
rect 4870 3933 4894 3934
rect 4818 3907 4822 3933
rect 4870 3907 4884 3933
rect 4818 3906 4842 3907
rect 4870 3906 4894 3907
rect 4922 3906 4946 3934
rect 4974 3906 4998 3934
rect 5026 3933 5035 3934
rect 5034 3907 5035 3933
rect 5026 3906 5035 3907
rect 4573 3901 5035 3906
rect 4494 3793 4522 3799
rect 4494 3767 4495 3793
rect 4521 3767 4522 3793
rect 4494 3737 4522 3767
rect 4494 3711 4495 3737
rect 4521 3711 4522 3737
rect 3822 3345 3850 3351
rect 3822 3319 3823 3345
rect 3849 3319 3850 3345
rect 3822 2561 3850 3319
rect 4382 3346 4410 3351
rect 4494 3346 4522 3711
rect 4382 3345 4522 3346
rect 4382 3319 4383 3345
rect 4409 3319 4495 3345
rect 4521 3319 4522 3345
rect 4382 3318 4522 3319
rect 4382 3313 4410 3318
rect 3822 2535 3823 2561
rect 3849 2535 3850 2561
rect 3822 1834 3850 2535
rect 4494 3009 4522 3318
rect 5278 3738 5306 4102
rect 5950 4130 5978 5054
rect 6118 5306 6146 6063
rect 6454 7266 6482 7271
rect 6510 7266 6538 7630
rect 6454 7265 6538 7266
rect 6454 7239 6455 7265
rect 6481 7239 6538 7265
rect 6454 7238 6538 7239
rect 6454 7209 6482 7238
rect 6454 7183 6455 7209
rect 6481 7183 6482 7209
rect 6454 6481 6482 7183
rect 6454 6455 6455 6481
rect 6481 6455 6482 6481
rect 6454 6425 6482 6455
rect 6454 6399 6455 6425
rect 6481 6399 6482 6425
rect 6454 6090 6482 6399
rect 6454 6057 6482 6062
rect 6118 4521 6146 5278
rect 6790 5361 6818 5367
rect 6790 5335 6791 5361
rect 6817 5335 6818 5361
rect 6790 5305 6818 5335
rect 6790 5279 6791 5305
rect 6817 5279 6818 5305
rect 6454 4914 6482 4919
rect 6454 4857 6482 4886
rect 6454 4831 6455 4857
rect 6481 4831 6482 4857
rect 6454 4825 6482 4831
rect 6790 4914 6818 5279
rect 6118 4495 6119 4521
rect 6145 4495 6146 4521
rect 6118 4489 6146 4495
rect 6790 4577 6818 4886
rect 6790 4551 6791 4577
rect 6817 4551 6818 4577
rect 6790 4522 6818 4551
rect 6790 4456 6818 4494
rect 6902 4214 6930 14630
rect 7014 14769 7042 15471
rect 7574 15497 7602 15503
rect 7574 15471 7575 15497
rect 7601 15471 7602 15497
rect 7073 15302 7535 15307
rect 7073 15301 7082 15302
rect 7073 15275 7074 15301
rect 7073 15274 7082 15275
rect 7110 15274 7134 15302
rect 7162 15274 7186 15302
rect 7214 15301 7238 15302
rect 7266 15301 7290 15302
rect 7224 15275 7238 15301
rect 7286 15275 7290 15301
rect 7214 15274 7238 15275
rect 7266 15274 7290 15275
rect 7318 15301 7342 15302
rect 7370 15301 7394 15302
rect 7318 15275 7322 15301
rect 7370 15275 7384 15301
rect 7318 15274 7342 15275
rect 7370 15274 7394 15275
rect 7422 15274 7446 15302
rect 7474 15274 7498 15302
rect 7526 15301 7535 15302
rect 7534 15275 7535 15301
rect 7526 15274 7535 15275
rect 7073 15269 7535 15274
rect 7014 14743 7015 14769
rect 7041 14743 7042 14769
rect 7014 14713 7042 14743
rect 7014 14687 7015 14713
rect 7041 14687 7042 14713
rect 7014 13985 7042 14687
rect 7574 14713 7602 15471
rect 7574 14687 7575 14713
rect 7601 14687 7602 14713
rect 7073 14518 7535 14523
rect 7073 14517 7082 14518
rect 7073 14491 7074 14517
rect 7073 14490 7082 14491
rect 7110 14490 7134 14518
rect 7162 14490 7186 14518
rect 7214 14517 7238 14518
rect 7266 14517 7290 14518
rect 7224 14491 7238 14517
rect 7286 14491 7290 14517
rect 7214 14490 7238 14491
rect 7266 14490 7290 14491
rect 7318 14517 7342 14518
rect 7370 14517 7394 14518
rect 7318 14491 7322 14517
rect 7370 14491 7384 14517
rect 7318 14490 7342 14491
rect 7370 14490 7394 14491
rect 7422 14490 7446 14518
rect 7474 14490 7498 14518
rect 7526 14517 7535 14518
rect 7534 14491 7535 14517
rect 7526 14490 7535 14491
rect 7073 14485 7535 14490
rect 7014 13959 7015 13985
rect 7041 13959 7042 13985
rect 7014 13929 7042 13959
rect 7014 13903 7015 13929
rect 7041 13903 7042 13929
rect 7014 13201 7042 13903
rect 7574 13929 7602 14687
rect 7798 14714 7826 16646
rect 8974 16673 9002 16679
rect 8974 16647 8975 16673
rect 9001 16647 9002 16673
rect 8974 16617 9002 16647
rect 9254 16674 9282 17431
rect 10206 17458 10234 17822
rect 10262 17817 10290 17822
rect 10486 17817 10514 17822
rect 11102 17850 11130 18215
rect 11830 18241 11858 18247
rect 11830 18215 11831 18241
rect 11857 18215 11858 18241
rect 11830 18186 11858 18215
rect 12054 18186 12082 18191
rect 11830 18185 12082 18186
rect 11830 18159 12055 18185
rect 12081 18159 12082 18185
rect 11830 18158 12082 18159
rect 11102 17817 11130 17822
rect 11270 17849 11298 17855
rect 11270 17823 11271 17849
rect 11297 17823 11298 17849
rect 10374 17458 10402 17463
rect 10206 17457 10402 17458
rect 10206 17431 10375 17457
rect 10401 17431 10402 17457
rect 10206 17430 10402 17431
rect 10374 17401 10402 17430
rect 10374 17375 10375 17401
rect 10401 17375 10402 17401
rect 9573 17262 10035 17267
rect 9573 17261 9582 17262
rect 9573 17235 9574 17261
rect 9573 17234 9582 17235
rect 9610 17234 9634 17262
rect 9662 17234 9686 17262
rect 9714 17261 9738 17262
rect 9766 17261 9790 17262
rect 9724 17235 9738 17261
rect 9786 17235 9790 17261
rect 9714 17234 9738 17235
rect 9766 17234 9790 17235
rect 9818 17261 9842 17262
rect 9870 17261 9894 17262
rect 9818 17235 9822 17261
rect 9870 17235 9884 17261
rect 9818 17234 9842 17235
rect 9870 17234 9894 17235
rect 9922 17234 9946 17262
rect 9974 17234 9998 17262
rect 10026 17261 10035 17262
rect 10034 17235 10035 17261
rect 10026 17234 10035 17235
rect 9573 17229 10035 17234
rect 10094 17065 10122 17071
rect 10094 17039 10095 17065
rect 10121 17039 10122 17065
rect 9254 16641 9282 16646
rect 9478 16673 9506 16679
rect 9478 16647 9479 16673
rect 9505 16647 9506 16673
rect 8974 16591 8975 16617
rect 9001 16591 9002 16617
rect 7798 14681 7826 14686
rect 8078 15889 8106 15895
rect 8078 15863 8079 15889
rect 8105 15863 8106 15889
rect 8078 15105 8106 15863
rect 8974 15889 9002 16591
rect 8974 15863 8975 15889
rect 9001 15863 9002 15889
rect 8974 15833 9002 15863
rect 8974 15807 8975 15833
rect 9001 15807 9002 15833
rect 8078 15079 8079 15105
rect 8105 15079 8106 15105
rect 7574 13903 7575 13929
rect 7601 13903 7602 13929
rect 7073 13734 7535 13739
rect 7073 13733 7082 13734
rect 7073 13707 7074 13733
rect 7073 13706 7082 13707
rect 7110 13706 7134 13734
rect 7162 13706 7186 13734
rect 7214 13733 7238 13734
rect 7266 13733 7290 13734
rect 7224 13707 7238 13733
rect 7286 13707 7290 13733
rect 7214 13706 7238 13707
rect 7266 13706 7290 13707
rect 7318 13733 7342 13734
rect 7370 13733 7394 13734
rect 7318 13707 7322 13733
rect 7370 13707 7384 13733
rect 7318 13706 7342 13707
rect 7370 13706 7394 13707
rect 7422 13706 7446 13734
rect 7474 13706 7498 13734
rect 7526 13733 7535 13734
rect 7534 13707 7535 13733
rect 7526 13706 7535 13707
rect 7073 13701 7535 13706
rect 7014 13175 7015 13201
rect 7041 13175 7042 13201
rect 7014 13145 7042 13175
rect 7014 13119 7015 13145
rect 7041 13119 7042 13145
rect 7014 12698 7042 13119
rect 7574 13145 7602 13903
rect 7574 13119 7575 13145
rect 7601 13119 7602 13145
rect 7073 12950 7535 12955
rect 7073 12949 7082 12950
rect 7073 12923 7074 12949
rect 7073 12922 7082 12923
rect 7110 12922 7134 12950
rect 7162 12922 7186 12950
rect 7214 12949 7238 12950
rect 7266 12949 7290 12950
rect 7224 12923 7238 12949
rect 7286 12923 7290 12949
rect 7214 12922 7238 12923
rect 7266 12922 7290 12923
rect 7318 12949 7342 12950
rect 7370 12949 7394 12950
rect 7318 12923 7322 12949
rect 7370 12923 7384 12949
rect 7318 12922 7342 12923
rect 7370 12922 7394 12923
rect 7422 12922 7446 12950
rect 7474 12922 7498 12950
rect 7526 12949 7535 12950
rect 7534 12923 7535 12949
rect 7526 12922 7535 12923
rect 7073 12917 7535 12922
rect 7014 12418 7042 12670
rect 7014 12361 7042 12390
rect 7014 12335 7015 12361
rect 7041 12335 7042 12361
rect 7014 12329 7042 12335
rect 7574 12362 7602 13119
rect 7073 12166 7535 12171
rect 7073 12165 7082 12166
rect 7073 12139 7074 12165
rect 7073 12138 7082 12139
rect 7110 12138 7134 12166
rect 7162 12138 7186 12166
rect 7214 12165 7238 12166
rect 7266 12165 7290 12166
rect 7224 12139 7238 12165
rect 7286 12139 7290 12165
rect 7214 12138 7238 12139
rect 7266 12138 7290 12139
rect 7318 12165 7342 12166
rect 7370 12165 7394 12166
rect 7318 12139 7322 12165
rect 7370 12139 7384 12165
rect 7318 12138 7342 12139
rect 7370 12138 7394 12139
rect 7422 12138 7446 12166
rect 7474 12138 7498 12166
rect 7526 12165 7535 12166
rect 7534 12139 7535 12165
rect 7526 12138 7535 12139
rect 7073 12133 7535 12138
rect 7574 11802 7602 12334
rect 7574 11577 7602 11774
rect 7574 11551 7575 11577
rect 7601 11551 7602 11577
rect 7574 11545 7602 11551
rect 8078 14321 8106 15079
rect 8078 14295 8079 14321
rect 8105 14295 8106 14321
rect 8078 13537 8106 14295
rect 8470 15553 8498 15559
rect 8470 15527 8471 15553
rect 8497 15527 8498 15553
rect 8470 15497 8498 15527
rect 8470 15471 8471 15497
rect 8497 15471 8498 15497
rect 8470 14769 8498 15471
rect 8470 14743 8471 14769
rect 8497 14743 8498 14769
rect 8470 14714 8498 14743
rect 8470 13985 8498 14686
rect 8974 15105 9002 15807
rect 8974 15079 8975 15105
rect 9001 15079 9002 15105
rect 8974 15049 9002 15079
rect 8974 15023 8975 15049
rect 9001 15023 9002 15049
rect 8974 14714 9002 15023
rect 8974 14322 9002 14686
rect 8974 14265 9002 14294
rect 8974 14239 8975 14265
rect 9001 14239 9002 14265
rect 8974 14233 9002 14239
rect 9478 15889 9506 16647
rect 9573 16478 10035 16483
rect 9573 16477 9582 16478
rect 9573 16451 9574 16477
rect 9573 16450 9582 16451
rect 9610 16450 9634 16478
rect 9662 16450 9686 16478
rect 9714 16477 9738 16478
rect 9766 16477 9790 16478
rect 9724 16451 9738 16477
rect 9786 16451 9790 16477
rect 9714 16450 9738 16451
rect 9766 16450 9790 16451
rect 9818 16477 9842 16478
rect 9870 16477 9894 16478
rect 9818 16451 9822 16477
rect 9870 16451 9884 16477
rect 9818 16450 9842 16451
rect 9870 16450 9894 16451
rect 9922 16450 9946 16478
rect 9974 16450 9998 16478
rect 10026 16477 10035 16478
rect 10034 16451 10035 16477
rect 10026 16450 10035 16451
rect 9573 16445 10035 16450
rect 10094 16282 10122 17039
rect 10374 17066 10402 17375
rect 10486 17066 10514 17071
rect 10374 17065 10514 17066
rect 10374 17039 10375 17065
rect 10401 17039 10487 17065
rect 10513 17039 10514 17065
rect 10374 17038 10514 17039
rect 10374 16674 10402 17038
rect 10486 17033 10514 17038
rect 11270 17065 11298 17823
rect 11830 17850 11858 18158
rect 12054 18153 12082 18158
rect 11942 17850 11970 17855
rect 11830 17849 11970 17850
rect 11830 17823 11831 17849
rect 11857 17823 11943 17849
rect 11969 17823 11970 17849
rect 11830 17822 11970 17823
rect 11270 17039 11271 17065
rect 11297 17039 11298 17065
rect 10430 16674 10458 16679
rect 10374 16673 10458 16674
rect 10374 16647 10431 16673
rect 10457 16647 10458 16673
rect 10374 16646 10458 16647
rect 10094 16235 10122 16254
rect 10430 16617 10458 16646
rect 10430 16591 10431 16617
rect 10457 16591 10458 16617
rect 9478 15863 9479 15889
rect 9505 15863 9506 15889
rect 9478 15105 9506 15863
rect 10430 15889 10458 16591
rect 10430 15863 10431 15889
rect 10457 15863 10458 15889
rect 10430 15834 10458 15863
rect 9573 15694 10035 15699
rect 9573 15693 9582 15694
rect 9573 15667 9574 15693
rect 9573 15666 9582 15667
rect 9610 15666 9634 15694
rect 9662 15666 9686 15694
rect 9714 15693 9738 15694
rect 9766 15693 9790 15694
rect 9724 15667 9738 15693
rect 9786 15667 9790 15693
rect 9714 15666 9738 15667
rect 9766 15666 9790 15667
rect 9818 15693 9842 15694
rect 9870 15693 9894 15694
rect 9818 15667 9822 15693
rect 9870 15667 9884 15693
rect 9818 15666 9842 15667
rect 9870 15666 9894 15667
rect 9922 15666 9946 15694
rect 9974 15666 9998 15694
rect 10026 15693 10035 15694
rect 10034 15667 10035 15693
rect 10026 15666 10035 15667
rect 9573 15661 10035 15666
rect 10038 15498 10066 15503
rect 10038 15451 10066 15470
rect 9478 15079 9479 15105
rect 9505 15079 9506 15105
rect 9478 14321 9506 15079
rect 10430 15105 10458 15806
rect 10990 16337 11018 16343
rect 10990 16311 10991 16337
rect 11017 16311 11018 16337
rect 10990 16282 11018 16311
rect 10990 15834 11018 16254
rect 10990 15553 11018 15806
rect 10990 15527 10991 15553
rect 11017 15527 11018 15553
rect 10990 15497 11018 15527
rect 10990 15471 10991 15497
rect 11017 15471 11018 15497
rect 10990 15465 11018 15471
rect 11270 16281 11298 17039
rect 11270 16255 11271 16281
rect 11297 16255 11298 16281
rect 11270 15498 11298 16255
rect 10430 15079 10431 15105
rect 10457 15079 10458 15105
rect 10430 15050 10458 15079
rect 10374 15049 10458 15050
rect 10374 15023 10431 15049
rect 10457 15023 10458 15049
rect 10374 15022 10458 15023
rect 9573 14910 10035 14915
rect 9573 14909 9582 14910
rect 9573 14883 9574 14909
rect 9573 14882 9582 14883
rect 9610 14882 9634 14910
rect 9662 14882 9686 14910
rect 9714 14909 9738 14910
rect 9766 14909 9790 14910
rect 9724 14883 9738 14909
rect 9786 14883 9790 14909
rect 9714 14882 9738 14883
rect 9766 14882 9790 14883
rect 9818 14909 9842 14910
rect 9870 14909 9894 14910
rect 9818 14883 9822 14909
rect 9870 14883 9884 14909
rect 9818 14882 9842 14883
rect 9870 14882 9894 14883
rect 9922 14882 9946 14910
rect 9974 14882 9998 14910
rect 10026 14909 10035 14910
rect 10034 14883 10035 14909
rect 10026 14882 10035 14883
rect 9573 14877 10035 14882
rect 9478 14295 9479 14321
rect 9505 14295 9506 14321
rect 8470 13959 8471 13985
rect 8497 13959 8498 13985
rect 8470 13929 8498 13959
rect 8470 13903 8471 13929
rect 8497 13903 8498 13929
rect 8078 13511 8079 13537
rect 8105 13511 8106 13537
rect 8078 12753 8106 13511
rect 8078 12727 8079 12753
rect 8105 12727 8106 12753
rect 8078 11969 8106 12727
rect 8358 13538 8386 13543
rect 8470 13538 8498 13903
rect 8358 13537 8498 13538
rect 8358 13511 8359 13537
rect 8385 13511 8471 13537
rect 8497 13511 8498 13537
rect 8358 13510 8498 13511
rect 8358 13201 8386 13510
rect 8470 13505 8498 13510
rect 8862 13874 8890 13879
rect 8358 13175 8359 13201
rect 8385 13175 8386 13201
rect 8358 13145 8386 13175
rect 8358 13119 8359 13145
rect 8385 13119 8386 13145
rect 8358 12754 8386 13119
rect 8470 12754 8498 12759
rect 8358 12753 8498 12754
rect 8358 12727 8359 12753
rect 8385 12727 8471 12753
rect 8497 12727 8498 12753
rect 8358 12726 8498 12727
rect 8358 12418 8386 12726
rect 8470 12721 8498 12726
rect 8358 12361 8386 12390
rect 8358 12335 8359 12361
rect 8385 12335 8386 12361
rect 8358 12329 8386 12335
rect 8078 11943 8079 11969
rect 8105 11943 8106 11969
rect 8078 11802 8106 11943
rect 7073 11382 7535 11387
rect 7073 11381 7082 11382
rect 7073 11355 7074 11381
rect 7073 11354 7082 11355
rect 7110 11354 7134 11382
rect 7162 11354 7186 11382
rect 7214 11381 7238 11382
rect 7266 11381 7290 11382
rect 7224 11355 7238 11381
rect 7286 11355 7290 11381
rect 7214 11354 7238 11355
rect 7266 11354 7290 11355
rect 7318 11381 7342 11382
rect 7370 11381 7394 11382
rect 7318 11355 7322 11381
rect 7370 11355 7384 11381
rect 7318 11354 7342 11355
rect 7370 11354 7394 11355
rect 7422 11354 7446 11382
rect 7474 11354 7498 11382
rect 7526 11381 7535 11382
rect 7534 11355 7535 11381
rect 7526 11354 7535 11355
rect 7073 11349 7535 11354
rect 8078 11185 8106 11774
rect 8078 11159 8079 11185
rect 8105 11159 8106 11185
rect 8078 11153 8106 11159
rect 8470 11633 8498 11639
rect 8470 11607 8471 11633
rect 8497 11607 8498 11633
rect 8470 11577 8498 11607
rect 8470 11551 8471 11577
rect 8497 11551 8498 11577
rect 8470 11130 8498 11551
rect 8470 11097 8498 11102
rect 8302 10849 8330 10855
rect 8302 10823 8303 10849
rect 8329 10823 8330 10849
rect 7574 10793 7602 10799
rect 7574 10767 7575 10793
rect 7601 10767 7602 10793
rect 7073 10598 7535 10603
rect 7073 10597 7082 10598
rect 7073 10571 7074 10597
rect 7073 10570 7082 10571
rect 7110 10570 7134 10598
rect 7162 10570 7186 10598
rect 7214 10597 7238 10598
rect 7266 10597 7290 10598
rect 7224 10571 7238 10597
rect 7286 10571 7290 10597
rect 7214 10570 7238 10571
rect 7266 10570 7290 10571
rect 7318 10597 7342 10598
rect 7370 10597 7394 10598
rect 7318 10571 7322 10597
rect 7370 10571 7384 10597
rect 7318 10570 7342 10571
rect 7370 10570 7394 10571
rect 7422 10570 7446 10598
rect 7474 10570 7498 10598
rect 7526 10597 7535 10598
rect 7534 10571 7535 10597
rect 7526 10570 7535 10571
rect 7073 10565 7535 10570
rect 7574 10402 7602 10767
rect 8302 10793 8330 10823
rect 8302 10767 8303 10793
rect 8329 10767 8330 10793
rect 7798 10402 7826 10407
rect 7574 10401 7826 10402
rect 7574 10375 7799 10401
rect 7825 10375 7826 10401
rect 7574 10374 7826 10375
rect 7014 10065 7042 10071
rect 7014 10039 7015 10065
rect 7041 10039 7042 10065
rect 7014 10009 7042 10039
rect 7014 9983 7015 10009
rect 7041 9983 7042 10009
rect 7014 9562 7042 9983
rect 7574 10009 7602 10374
rect 7798 10369 7826 10374
rect 8302 10402 8330 10767
rect 8470 10402 8498 10407
rect 8302 10401 8498 10402
rect 8302 10375 8303 10401
rect 8329 10375 8471 10401
rect 8497 10375 8498 10401
rect 8302 10374 8498 10375
rect 8302 10094 8330 10374
rect 8470 10369 8498 10374
rect 8302 10066 8386 10094
rect 7574 9983 7575 10009
rect 7601 9983 7602 10009
rect 7073 9814 7535 9819
rect 7073 9813 7082 9814
rect 7073 9787 7074 9813
rect 7073 9786 7082 9787
rect 7110 9786 7134 9814
rect 7162 9786 7186 9814
rect 7214 9813 7238 9814
rect 7266 9813 7290 9814
rect 7224 9787 7238 9813
rect 7286 9787 7290 9813
rect 7214 9786 7238 9787
rect 7266 9786 7290 9787
rect 7318 9813 7342 9814
rect 7370 9813 7394 9814
rect 7318 9787 7322 9813
rect 7370 9787 7384 9813
rect 7318 9786 7342 9787
rect 7370 9786 7394 9787
rect 7422 9786 7446 9814
rect 7474 9786 7498 9814
rect 7526 9813 7535 9814
rect 7534 9787 7535 9813
rect 7526 9786 7535 9787
rect 7073 9781 7535 9786
rect 7014 9281 7042 9534
rect 7014 9255 7015 9281
rect 7041 9255 7042 9281
rect 7014 9225 7042 9255
rect 7014 9199 7015 9225
rect 7041 9199 7042 9225
rect 7014 7658 7042 9199
rect 7574 9618 7602 9983
rect 8358 10065 8386 10066
rect 8358 10039 8359 10065
rect 8385 10039 8386 10065
rect 8358 10009 8386 10039
rect 8358 9983 8359 10009
rect 8385 9983 8386 10009
rect 7798 9618 7826 9623
rect 7574 9617 7826 9618
rect 7574 9591 7799 9617
rect 7825 9591 7826 9617
rect 7574 9590 7826 9591
rect 7574 9225 7602 9590
rect 7798 9585 7826 9590
rect 8358 9618 8386 9983
rect 8470 9618 8498 9623
rect 8358 9617 8498 9618
rect 8358 9591 8359 9617
rect 8385 9591 8471 9617
rect 8497 9591 8498 9617
rect 8358 9590 8498 9591
rect 7574 9199 7575 9225
rect 7601 9199 7602 9225
rect 7073 9030 7535 9035
rect 7073 9029 7082 9030
rect 7073 9003 7074 9029
rect 7073 9002 7082 9003
rect 7110 9002 7134 9030
rect 7162 9002 7186 9030
rect 7214 9029 7238 9030
rect 7266 9029 7290 9030
rect 7224 9003 7238 9029
rect 7286 9003 7290 9029
rect 7214 9002 7238 9003
rect 7266 9002 7290 9003
rect 7318 9029 7342 9030
rect 7370 9029 7394 9030
rect 7318 9003 7322 9029
rect 7370 9003 7384 9029
rect 7318 9002 7342 9003
rect 7370 9002 7394 9003
rect 7422 9002 7446 9030
rect 7474 9002 7498 9030
rect 7526 9029 7535 9030
rect 7534 9003 7535 9029
rect 7526 9002 7535 9003
rect 7073 8997 7535 9002
rect 7574 8834 7602 9199
rect 8358 9281 8386 9590
rect 8470 9585 8498 9590
rect 8358 9255 8359 9281
rect 8385 9255 8386 9281
rect 8358 9225 8386 9255
rect 8358 9199 8359 9225
rect 8385 9199 8386 9225
rect 7798 8834 7826 8839
rect 7574 8833 7826 8834
rect 7574 8807 7799 8833
rect 7825 8807 7826 8833
rect 7574 8806 7826 8807
rect 7574 8441 7602 8806
rect 7798 8801 7826 8806
rect 8358 8834 8386 9199
rect 8470 8834 8498 8839
rect 8358 8833 8498 8834
rect 8358 8807 8359 8833
rect 8385 8807 8471 8833
rect 8497 8807 8498 8833
rect 8358 8806 8498 8807
rect 7574 8415 7575 8441
rect 7601 8415 7602 8441
rect 7073 8246 7535 8251
rect 7073 8245 7082 8246
rect 7073 8219 7074 8245
rect 7073 8218 7082 8219
rect 7110 8218 7134 8246
rect 7162 8218 7186 8246
rect 7214 8245 7238 8246
rect 7266 8245 7290 8246
rect 7224 8219 7238 8245
rect 7286 8219 7290 8245
rect 7214 8218 7238 8219
rect 7266 8218 7290 8219
rect 7318 8245 7342 8246
rect 7370 8245 7394 8246
rect 7318 8219 7322 8245
rect 7370 8219 7384 8245
rect 7318 8218 7342 8219
rect 7370 8218 7394 8219
rect 7422 8218 7446 8246
rect 7474 8218 7498 8246
rect 7526 8245 7535 8246
rect 7534 8219 7535 8245
rect 7526 8218 7535 8219
rect 7073 8213 7535 8218
rect 7014 6929 7042 7630
rect 7574 8050 7602 8415
rect 8358 8498 8386 8806
rect 8470 8801 8498 8806
rect 8358 8441 8386 8470
rect 8358 8415 8359 8441
rect 8385 8415 8386 8441
rect 7798 8050 7826 8055
rect 7574 8049 7826 8050
rect 7574 8023 7799 8049
rect 7825 8023 7826 8049
rect 7574 8022 7826 8023
rect 7574 7657 7602 8022
rect 7798 8017 7826 8022
rect 8358 8050 8386 8415
rect 8470 8050 8498 8055
rect 8358 8049 8498 8050
rect 8358 8023 8359 8049
rect 8385 8023 8471 8049
rect 8497 8023 8498 8049
rect 8358 8022 8498 8023
rect 8358 8017 8386 8022
rect 7574 7631 7575 7657
rect 7601 7631 7602 7657
rect 7073 7462 7535 7467
rect 7073 7461 7082 7462
rect 7073 7435 7074 7461
rect 7073 7434 7082 7435
rect 7110 7434 7134 7462
rect 7162 7434 7186 7462
rect 7214 7461 7238 7462
rect 7266 7461 7290 7462
rect 7224 7435 7238 7461
rect 7286 7435 7290 7461
rect 7214 7434 7238 7435
rect 7266 7434 7290 7435
rect 7318 7461 7342 7462
rect 7370 7461 7394 7462
rect 7318 7435 7322 7461
rect 7370 7435 7384 7461
rect 7318 7434 7342 7435
rect 7370 7434 7394 7435
rect 7422 7434 7446 7462
rect 7474 7434 7498 7462
rect 7526 7461 7535 7462
rect 7534 7435 7535 7461
rect 7526 7434 7535 7435
rect 7073 7429 7535 7434
rect 7014 6903 7015 6929
rect 7041 6903 7042 6929
rect 7014 6873 7042 6903
rect 7014 6847 7015 6873
rect 7041 6847 7042 6873
rect 7014 6841 7042 6847
rect 7574 6873 7602 7631
rect 7742 7658 7770 7663
rect 7742 7611 7770 7630
rect 7966 7658 7994 7663
rect 7966 7611 7994 7630
rect 8470 7658 8498 8022
rect 8470 7574 8498 7630
rect 8470 7546 8778 7574
rect 7574 6847 7575 6873
rect 7601 6847 7602 6873
rect 7073 6678 7535 6683
rect 7073 6677 7082 6678
rect 7073 6651 7074 6677
rect 7073 6650 7082 6651
rect 7110 6650 7134 6678
rect 7162 6650 7186 6678
rect 7214 6677 7238 6678
rect 7266 6677 7290 6678
rect 7224 6651 7238 6677
rect 7286 6651 7290 6677
rect 7214 6650 7238 6651
rect 7266 6650 7290 6651
rect 7318 6677 7342 6678
rect 7370 6677 7394 6678
rect 7318 6651 7322 6677
rect 7370 6651 7384 6677
rect 7318 6650 7342 6651
rect 7370 6650 7394 6651
rect 7422 6650 7446 6678
rect 7474 6650 7498 6678
rect 7526 6677 7535 6678
rect 7534 6651 7535 6677
rect 7526 6650 7535 6651
rect 7073 6645 7535 6650
rect 7014 6145 7042 6151
rect 7014 6119 7015 6145
rect 7041 6119 7042 6145
rect 7014 6090 7042 6119
rect 7014 6043 7042 6062
rect 7574 6089 7602 6847
rect 7574 6063 7575 6089
rect 7601 6063 7602 6089
rect 7073 5894 7535 5899
rect 7073 5893 7082 5894
rect 7073 5867 7074 5893
rect 7073 5866 7082 5867
rect 7110 5866 7134 5894
rect 7162 5866 7186 5894
rect 7214 5893 7238 5894
rect 7266 5893 7290 5894
rect 7224 5867 7238 5893
rect 7286 5867 7290 5893
rect 7214 5866 7238 5867
rect 7266 5866 7290 5867
rect 7318 5893 7342 5894
rect 7370 5893 7394 5894
rect 7318 5867 7322 5893
rect 7370 5867 7384 5893
rect 7318 5866 7342 5867
rect 7370 5866 7394 5867
rect 7422 5866 7446 5894
rect 7474 5866 7498 5894
rect 7526 5893 7535 5894
rect 7534 5867 7535 5893
rect 7526 5866 7535 5867
rect 7073 5861 7535 5866
rect 7574 5866 7602 6063
rect 7574 5833 7602 5838
rect 8078 7265 8106 7271
rect 8078 7239 8079 7265
rect 8105 7239 8106 7265
rect 8078 6481 8106 7239
rect 8750 7265 8778 7546
rect 8750 7239 8751 7265
rect 8777 7239 8778 7265
rect 8750 7209 8778 7239
rect 8750 7183 8751 7209
rect 8777 7183 8778 7209
rect 8750 7177 8778 7183
rect 8078 6455 8079 6481
rect 8105 6455 8106 6481
rect 8078 5866 8106 6455
rect 8358 6929 8386 6935
rect 8358 6903 8359 6929
rect 8385 6903 8386 6929
rect 8358 6873 8386 6903
rect 8358 6847 8359 6873
rect 8385 6847 8386 6873
rect 8358 6146 8386 6847
rect 8470 6146 8498 6151
rect 8358 6145 8498 6146
rect 8358 6119 8471 6145
rect 8497 6119 8498 6145
rect 8358 6118 8498 6119
rect 8358 6090 8386 6118
rect 8358 6057 8386 6062
rect 8470 6089 8498 6118
rect 8470 6063 8471 6089
rect 8497 6063 8498 6089
rect 8078 5697 8106 5838
rect 8078 5671 8079 5697
rect 8105 5671 8106 5697
rect 7294 5306 7322 5311
rect 7294 5259 7322 5278
rect 8078 5306 8106 5671
rect 7073 5110 7535 5115
rect 7073 5109 7082 5110
rect 7073 5083 7074 5109
rect 7073 5082 7082 5083
rect 7110 5082 7134 5110
rect 7162 5082 7186 5110
rect 7214 5109 7238 5110
rect 7266 5109 7290 5110
rect 7224 5083 7238 5109
rect 7286 5083 7290 5109
rect 7214 5082 7238 5083
rect 7266 5082 7290 5083
rect 7318 5109 7342 5110
rect 7370 5109 7394 5110
rect 7318 5083 7322 5109
rect 7370 5083 7384 5109
rect 7318 5082 7342 5083
rect 7370 5082 7394 5083
rect 7422 5082 7446 5110
rect 7474 5082 7498 5110
rect 7526 5109 7535 5110
rect 7534 5083 7535 5109
rect 7526 5082 7535 5083
rect 7073 5077 7535 5082
rect 8078 4913 8106 5278
rect 8078 4887 8079 4913
rect 8105 4887 8106 4913
rect 6846 4186 6930 4214
rect 7014 4522 7042 4527
rect 7014 4186 7042 4494
rect 7574 4521 7602 4527
rect 7574 4495 7575 4521
rect 7601 4495 7602 4521
rect 7073 4326 7535 4331
rect 7073 4325 7082 4326
rect 7073 4299 7074 4325
rect 7073 4298 7082 4299
rect 7110 4298 7134 4326
rect 7162 4298 7186 4326
rect 7214 4325 7238 4326
rect 7266 4325 7290 4326
rect 7224 4299 7238 4325
rect 7286 4299 7290 4325
rect 7214 4298 7238 4299
rect 7266 4298 7290 4299
rect 7318 4325 7342 4326
rect 7370 4325 7394 4326
rect 7318 4299 7322 4325
rect 7370 4299 7384 4325
rect 7318 4298 7342 4299
rect 7370 4298 7394 4299
rect 7422 4298 7446 4326
rect 7474 4298 7498 4326
rect 7526 4325 7535 4326
rect 7534 4299 7535 4325
rect 7526 4298 7535 4299
rect 7073 4293 7535 4298
rect 5950 4097 5978 4102
rect 6454 4130 6482 4135
rect 6454 4073 6482 4102
rect 6454 4047 6455 4073
rect 6481 4047 6482 4073
rect 5278 3345 5306 3710
rect 5838 3738 5866 3743
rect 5278 3319 5279 3345
rect 5305 3319 5306 3345
rect 4573 3150 5035 3155
rect 4573 3149 4582 3150
rect 4573 3123 4574 3149
rect 4573 3122 4582 3123
rect 4610 3122 4634 3150
rect 4662 3122 4686 3150
rect 4714 3149 4738 3150
rect 4766 3149 4790 3150
rect 4724 3123 4738 3149
rect 4786 3123 4790 3149
rect 4714 3122 4738 3123
rect 4766 3122 4790 3123
rect 4818 3149 4842 3150
rect 4870 3149 4894 3150
rect 4818 3123 4822 3149
rect 4870 3123 4884 3149
rect 4818 3122 4842 3123
rect 4870 3122 4894 3123
rect 4922 3122 4946 3150
rect 4974 3122 4998 3150
rect 5026 3149 5035 3150
rect 5034 3123 5035 3149
rect 5026 3122 5035 3123
rect 4573 3117 5035 3122
rect 4494 2983 4495 3009
rect 4521 2983 4522 3009
rect 4494 2953 4522 2983
rect 4494 2927 4495 2953
rect 4521 2927 4522 2953
rect 4494 2506 4522 2927
rect 4494 2473 4522 2478
rect 4998 2561 5026 2567
rect 4998 2535 4999 2561
rect 5025 2535 5026 2561
rect 4998 2506 5026 2535
rect 5278 2561 5306 3319
rect 5278 2535 5279 2561
rect 5305 2535 5306 2561
rect 5278 2529 5306 2535
rect 5390 3458 5418 3463
rect 4998 2459 5026 2478
rect 4573 2366 5035 2371
rect 4573 2365 4582 2366
rect 4573 2339 4574 2365
rect 4573 2338 4582 2339
rect 4610 2338 4634 2366
rect 4662 2338 4686 2366
rect 4714 2365 4738 2366
rect 4766 2365 4790 2366
rect 4724 2339 4738 2365
rect 4786 2339 4790 2365
rect 4714 2338 4738 2339
rect 4766 2338 4790 2339
rect 4818 2365 4842 2366
rect 4870 2365 4894 2366
rect 4818 2339 4822 2365
rect 4870 2339 4884 2365
rect 4818 2338 4842 2339
rect 4870 2338 4894 2339
rect 4922 2338 4946 2366
rect 4974 2338 4998 2366
rect 5026 2365 5035 2366
rect 5034 2339 5035 2365
rect 5026 2338 5035 2339
rect 4573 2333 5035 2338
rect 3822 1801 3850 1806
rect 4438 2226 4466 2231
rect 4438 2169 4466 2198
rect 4438 2143 4439 2169
rect 4465 2143 4466 2169
rect 4438 1777 4466 2143
rect 4438 1751 4439 1777
rect 4465 1751 4466 1777
rect 4438 1722 4466 1751
rect 4438 1675 4466 1694
rect 4573 1582 5035 1587
rect 4573 1581 4582 1582
rect 4573 1555 4574 1581
rect 4573 1554 4582 1555
rect 4610 1554 4634 1582
rect 4662 1554 4686 1582
rect 4714 1581 4738 1582
rect 4766 1581 4790 1582
rect 4724 1555 4738 1581
rect 4786 1555 4790 1581
rect 4714 1554 4738 1555
rect 4766 1554 4790 1555
rect 4818 1581 4842 1582
rect 4870 1581 4894 1582
rect 4818 1555 4822 1581
rect 4870 1555 4884 1581
rect 4818 1554 4842 1555
rect 4870 1554 4894 1555
rect 4922 1554 4946 1582
rect 4974 1554 4998 1582
rect 5026 1581 5035 1582
rect 5034 1555 5035 1581
rect 5026 1554 5035 1555
rect 4573 1549 5035 1554
rect 3766 462 3962 490
rect 3766 378 3794 462
rect 3934 400 3962 462
rect 5390 400 5418 3430
rect 5838 2954 5866 3710
rect 6454 3738 6482 4047
rect 6454 3705 6482 3710
rect 6454 3345 6482 3351
rect 6454 3319 6455 3345
rect 6481 3319 6482 3345
rect 6454 3290 6482 3319
rect 5838 2953 5922 2954
rect 5838 2927 5839 2953
rect 5865 2927 5922 2953
rect 5838 2926 5922 2927
rect 5838 2921 5866 2926
rect 5894 2170 5922 2926
rect 6454 2561 6482 3262
rect 6454 2535 6455 2561
rect 6481 2535 6482 2561
rect 5894 2104 5922 2142
rect 6342 2506 6370 2511
rect 5502 1834 5530 1839
rect 5502 1777 5530 1806
rect 5502 1751 5503 1777
rect 5529 1751 5530 1777
rect 5502 1745 5530 1751
rect 6342 1778 6370 2478
rect 6454 2505 6482 2535
rect 6454 2479 6455 2505
rect 6481 2479 6482 2505
rect 6398 2170 6426 2175
rect 6454 2170 6482 2479
rect 6510 2170 6538 2175
rect 6398 2169 6538 2170
rect 6398 2143 6399 2169
rect 6425 2143 6511 2169
rect 6537 2143 6538 2169
rect 6398 2142 6538 2143
rect 6398 2137 6426 2142
rect 6398 1778 6426 1783
rect 6342 1777 6426 1778
rect 6342 1751 6399 1777
rect 6425 1751 6426 1777
rect 6342 1750 6426 1751
rect 6398 1721 6426 1750
rect 6510 1778 6538 2142
rect 6510 1745 6538 1750
rect 6398 1695 6399 1721
rect 6425 1695 6426 1721
rect 6398 1442 6426 1695
rect 6398 1409 6426 1414
rect 6846 400 6874 4186
rect 6958 3793 6986 3799
rect 6958 3767 6959 3793
rect 6985 3767 6986 3793
rect 6958 3738 6986 3767
rect 6958 3691 6986 3710
rect 7014 3290 7042 4158
rect 7574 3738 7602 4495
rect 8078 4129 8106 4887
rect 8470 5361 8498 6063
rect 8470 5335 8471 5361
rect 8497 5335 8498 5361
rect 8470 5305 8498 5335
rect 8470 5279 8471 5305
rect 8497 5279 8498 5305
rect 8470 4577 8498 5279
rect 8470 4551 8471 4577
rect 8497 4551 8498 4577
rect 8470 4522 8498 4551
rect 8470 4186 8498 4494
rect 8470 4153 8498 4158
rect 8078 4103 8079 4129
rect 8105 4103 8106 4129
rect 8078 3738 8106 4103
rect 7574 3737 8106 3738
rect 7574 3711 7575 3737
rect 7601 3711 8106 3737
rect 7574 3710 8106 3711
rect 7574 3705 7602 3710
rect 7073 3542 7535 3547
rect 7073 3541 7082 3542
rect 7073 3515 7074 3541
rect 7073 3514 7082 3515
rect 7110 3514 7134 3542
rect 7162 3514 7186 3542
rect 7214 3541 7238 3542
rect 7266 3541 7290 3542
rect 7224 3515 7238 3541
rect 7286 3515 7290 3541
rect 7214 3514 7238 3515
rect 7266 3514 7290 3515
rect 7318 3541 7342 3542
rect 7370 3541 7394 3542
rect 7318 3515 7322 3541
rect 7370 3515 7384 3541
rect 7318 3514 7342 3515
rect 7370 3514 7394 3515
rect 7422 3514 7446 3542
rect 7474 3514 7498 3542
rect 7526 3541 7535 3542
rect 7534 3515 7535 3541
rect 7526 3514 7535 3515
rect 7073 3509 7535 3514
rect 8078 3402 8106 3710
rect 8078 3345 8106 3374
rect 8078 3319 8079 3345
rect 8105 3319 8106 3345
rect 8078 3313 8106 3319
rect 8358 3793 8386 3799
rect 8358 3767 8359 3793
rect 8385 3767 8386 3793
rect 8358 3738 8386 3767
rect 7014 3009 7042 3262
rect 7014 2983 7015 3009
rect 7041 2983 7042 3009
rect 7014 2953 7042 2983
rect 8358 3010 8386 3710
rect 8862 3458 8890 13846
rect 9478 13537 9506 14295
rect 10038 14713 10066 14719
rect 10038 14687 10039 14713
rect 10065 14687 10066 14713
rect 10038 14210 10066 14687
rect 10374 14714 10402 15022
rect 10430 15017 10458 15022
rect 10486 14714 10514 14719
rect 10374 14713 10514 14714
rect 10374 14687 10375 14713
rect 10401 14687 10487 14713
rect 10513 14687 10514 14713
rect 10374 14686 10514 14687
rect 10374 14322 10402 14686
rect 10486 14681 10514 14686
rect 11270 14713 11298 15470
rect 11270 14687 11271 14713
rect 11297 14687 11298 14713
rect 10374 14265 10402 14294
rect 10374 14239 10375 14265
rect 10401 14239 10402 14265
rect 10374 14233 10402 14239
rect 10038 14182 10122 14210
rect 9573 14126 10035 14131
rect 9573 14125 9582 14126
rect 9573 14099 9574 14125
rect 9573 14098 9582 14099
rect 9610 14098 9634 14126
rect 9662 14098 9686 14126
rect 9714 14125 9738 14126
rect 9766 14125 9790 14126
rect 9724 14099 9738 14125
rect 9786 14099 9790 14125
rect 9714 14098 9738 14099
rect 9766 14098 9790 14099
rect 9818 14125 9842 14126
rect 9870 14125 9894 14126
rect 9818 14099 9822 14125
rect 9870 14099 9884 14125
rect 9818 14098 9842 14099
rect 9870 14098 9894 14099
rect 9922 14098 9946 14126
rect 9974 14098 9998 14126
rect 10026 14125 10035 14126
rect 10034 14099 10035 14125
rect 10026 14098 10035 14099
rect 9573 14093 10035 14098
rect 9478 13511 9479 13537
rect 9505 13511 9506 13537
rect 9478 12753 9506 13511
rect 10094 13929 10122 14182
rect 10094 13903 10095 13929
rect 10121 13903 10122 13929
rect 9573 13342 10035 13347
rect 9573 13341 9582 13342
rect 9573 13315 9574 13341
rect 9573 13314 9582 13315
rect 9610 13314 9634 13342
rect 9662 13314 9686 13342
rect 9714 13341 9738 13342
rect 9766 13341 9790 13342
rect 9724 13315 9738 13341
rect 9786 13315 9790 13341
rect 9714 13314 9738 13315
rect 9766 13314 9790 13315
rect 9818 13341 9842 13342
rect 9870 13341 9894 13342
rect 9818 13315 9822 13341
rect 9870 13315 9884 13341
rect 9818 13314 9842 13315
rect 9870 13314 9894 13315
rect 9922 13314 9946 13342
rect 9974 13314 9998 13342
rect 10026 13341 10035 13342
rect 10034 13315 10035 13341
rect 10026 13314 10035 13315
rect 9573 13309 10035 13314
rect 9478 12727 9479 12753
rect 9505 12727 9506 12753
rect 9478 12362 9506 12727
rect 10094 13145 10122 13903
rect 10766 13985 10794 13991
rect 10766 13959 10767 13985
rect 10793 13959 10794 13985
rect 10766 13929 10794 13959
rect 10766 13903 10767 13929
rect 10793 13903 10794 13929
rect 10094 13119 10095 13145
rect 10121 13119 10122 13145
rect 9573 12558 10035 12563
rect 9573 12557 9582 12558
rect 9573 12531 9574 12557
rect 9573 12530 9582 12531
rect 9610 12530 9634 12558
rect 9662 12530 9686 12558
rect 9714 12557 9738 12558
rect 9766 12557 9790 12558
rect 9724 12531 9738 12557
rect 9786 12531 9790 12557
rect 9714 12530 9738 12531
rect 9766 12530 9790 12531
rect 9818 12557 9842 12558
rect 9870 12557 9894 12558
rect 9818 12531 9822 12557
rect 9870 12531 9884 12557
rect 9818 12530 9842 12531
rect 9870 12530 9894 12531
rect 9922 12530 9946 12558
rect 9974 12530 9998 12558
rect 10026 12557 10035 12558
rect 10034 12531 10035 12557
rect 10026 12530 10035 12531
rect 9573 12525 10035 12530
rect 9534 12362 9562 12367
rect 9478 12334 9534 12362
rect 8974 11970 9002 11975
rect 9534 11970 9562 12334
rect 10094 12362 10122 13119
rect 10430 13538 10458 13543
rect 10430 13481 10458 13510
rect 10430 13455 10431 13481
rect 10457 13455 10458 13481
rect 10430 12753 10458 13455
rect 10766 13538 10794 13903
rect 10766 13201 10794 13510
rect 10766 13175 10767 13201
rect 10793 13175 10794 13201
rect 10766 13145 10794 13175
rect 10766 13119 10767 13145
rect 10793 13119 10794 13145
rect 10766 13113 10794 13119
rect 11270 13929 11298 14687
rect 11270 13903 11271 13929
rect 11297 13903 11298 13929
rect 11270 13145 11298 13903
rect 11270 13119 11271 13145
rect 11297 13119 11298 13145
rect 10430 12727 10431 12753
rect 10457 12727 10458 12753
rect 10430 12697 10458 12727
rect 10430 12671 10431 12697
rect 10457 12671 10458 12697
rect 10094 12315 10122 12334
rect 10374 12362 10402 12367
rect 10430 12362 10458 12671
rect 10486 12362 10514 12367
rect 10374 12361 10514 12362
rect 10374 12335 10375 12361
rect 10401 12335 10487 12361
rect 10513 12335 10514 12361
rect 10374 12334 10514 12335
rect 8974 11913 9002 11942
rect 8974 11887 8975 11913
rect 9001 11887 9002 11913
rect 8974 11881 9002 11887
rect 9478 11969 9562 11970
rect 9478 11943 9535 11969
rect 9561 11943 9562 11969
rect 9478 11942 9562 11943
rect 9478 11802 9506 11942
rect 9534 11937 9562 11942
rect 9702 11970 9730 11975
rect 9702 11923 9730 11942
rect 10374 11970 10402 12334
rect 10486 12329 10514 12334
rect 11270 12362 11298 13119
rect 9478 11578 9506 11774
rect 9573 11774 10035 11779
rect 9573 11773 9582 11774
rect 9573 11747 9574 11773
rect 9573 11746 9582 11747
rect 9610 11746 9634 11774
rect 9662 11746 9686 11774
rect 9714 11773 9738 11774
rect 9766 11773 9790 11774
rect 9724 11747 9738 11773
rect 9786 11747 9790 11773
rect 9714 11746 9738 11747
rect 9766 11746 9790 11747
rect 9818 11773 9842 11774
rect 9870 11773 9894 11774
rect 9818 11747 9822 11773
rect 9870 11747 9884 11773
rect 9818 11746 9842 11747
rect 9870 11746 9894 11747
rect 9922 11746 9946 11774
rect 9974 11746 9998 11774
rect 10026 11773 10035 11774
rect 10034 11747 10035 11773
rect 10026 11746 10035 11747
rect 9573 11741 10035 11746
rect 9814 11578 9842 11583
rect 9478 11577 9842 11578
rect 9478 11551 9815 11577
rect 9841 11551 9842 11577
rect 9478 11550 9842 11551
rect 8974 11185 9002 11191
rect 8974 11159 8975 11185
rect 9001 11159 9002 11185
rect 8974 11130 9002 11159
rect 8974 11083 9002 11102
rect 9478 11185 9506 11550
rect 9814 11545 9842 11550
rect 10374 11578 10402 11942
rect 11270 11970 11298 12334
rect 11774 17457 11802 17463
rect 11774 17431 11775 17457
rect 11801 17431 11802 17457
rect 11774 16673 11802 17431
rect 11774 16647 11775 16673
rect 11801 16647 11802 16673
rect 11774 15889 11802 16647
rect 11774 15863 11775 15889
rect 11801 15863 11802 15889
rect 11774 15105 11802 15863
rect 11830 17458 11858 17822
rect 11942 17817 11970 17822
rect 12558 17738 12586 18326
rect 13342 18242 13370 18247
rect 13398 18242 13426 18247
rect 13342 18241 13398 18242
rect 13342 18215 13343 18241
rect 13369 18215 13398 18241
rect 13342 18214 13398 18215
rect 13342 18209 13370 18214
rect 13398 17849 13426 18214
rect 13398 17823 13399 17849
rect 13425 17823 13426 17849
rect 12558 17710 12642 17738
rect 12073 17654 12535 17659
rect 12073 17653 12082 17654
rect 12073 17627 12074 17653
rect 12073 17626 12082 17627
rect 12110 17626 12134 17654
rect 12162 17626 12186 17654
rect 12214 17653 12238 17654
rect 12266 17653 12290 17654
rect 12224 17627 12238 17653
rect 12286 17627 12290 17653
rect 12214 17626 12238 17627
rect 12266 17626 12290 17627
rect 12318 17653 12342 17654
rect 12370 17653 12394 17654
rect 12318 17627 12322 17653
rect 12370 17627 12384 17653
rect 12318 17626 12342 17627
rect 12370 17626 12394 17627
rect 12422 17626 12446 17654
rect 12474 17626 12498 17654
rect 12526 17653 12535 17654
rect 12534 17627 12535 17653
rect 12526 17626 12535 17627
rect 12073 17621 12535 17626
rect 12222 17458 12250 17463
rect 12446 17458 12474 17463
rect 11830 17457 12474 17458
rect 11830 17431 12223 17457
rect 12249 17431 12447 17457
rect 12473 17431 12474 17457
rect 11830 17430 12474 17431
rect 11830 17066 11858 17430
rect 12222 17425 12250 17430
rect 12446 17425 12474 17430
rect 12614 17346 12642 17710
rect 12614 17313 12642 17318
rect 13286 17458 13314 17463
rect 13398 17458 13426 17823
rect 13286 17457 13426 17458
rect 13286 17431 13287 17457
rect 13313 17431 13426 17457
rect 13286 17430 13426 17431
rect 14238 18241 14266 18247
rect 14238 18215 14239 18241
rect 14265 18215 14266 18241
rect 14238 18185 14266 18215
rect 14630 18242 14658 18247
rect 14630 18195 14658 18214
rect 15078 18242 15106 18247
rect 14238 18159 14239 18185
rect 14265 18159 14266 18185
rect 14238 17850 14266 18159
rect 14573 18046 15035 18051
rect 14573 18045 14582 18046
rect 14573 18019 14574 18045
rect 14573 18018 14582 18019
rect 14610 18018 14634 18046
rect 14662 18018 14686 18046
rect 14714 18045 14738 18046
rect 14766 18045 14790 18046
rect 14724 18019 14738 18045
rect 14786 18019 14790 18045
rect 14714 18018 14738 18019
rect 14766 18018 14790 18019
rect 14818 18045 14842 18046
rect 14870 18045 14894 18046
rect 14818 18019 14822 18045
rect 14870 18019 14884 18045
rect 14818 18018 14842 18019
rect 14870 18018 14894 18019
rect 14922 18018 14946 18046
rect 14974 18018 14998 18046
rect 15026 18045 15035 18046
rect 15034 18019 15035 18045
rect 15026 18018 15035 18019
rect 14573 18013 15035 18018
rect 14238 17457 14266 17822
rect 14574 17905 14602 17911
rect 14574 17879 14575 17905
rect 14601 17879 14602 17905
rect 14574 17850 14602 17879
rect 14574 17803 14602 17822
rect 15078 17849 15106 18214
rect 15078 17823 15079 17849
rect 15105 17823 15106 17849
rect 14238 17431 14239 17457
rect 14265 17431 14266 17457
rect 11942 17066 11970 17071
rect 11830 17065 11970 17066
rect 11830 17039 11831 17065
rect 11857 17039 11943 17065
rect 11969 17039 11970 17065
rect 11830 17038 11970 17039
rect 11830 16674 11858 17038
rect 11942 17033 11970 17038
rect 12073 16870 12535 16875
rect 12073 16869 12082 16870
rect 12073 16843 12074 16869
rect 12073 16842 12082 16843
rect 12110 16842 12134 16870
rect 12162 16842 12186 16870
rect 12214 16869 12238 16870
rect 12266 16869 12290 16870
rect 12224 16843 12238 16869
rect 12286 16843 12290 16869
rect 12214 16842 12238 16843
rect 12266 16842 12290 16843
rect 12318 16869 12342 16870
rect 12370 16869 12394 16870
rect 12318 16843 12322 16869
rect 12370 16843 12384 16869
rect 12318 16842 12342 16843
rect 12370 16842 12394 16843
rect 12422 16842 12446 16870
rect 12474 16842 12498 16870
rect 12526 16869 12535 16870
rect 12534 16843 12535 16869
rect 12526 16842 12535 16843
rect 12073 16837 12535 16842
rect 11830 16282 11858 16646
rect 12222 16674 12250 16679
rect 12222 16627 12250 16646
rect 12446 16674 12474 16679
rect 12446 16627 12474 16646
rect 13286 16673 13314 17430
rect 14238 17401 14266 17431
rect 14238 17375 14239 17401
rect 14265 17375 14266 17401
rect 13286 16647 13287 16673
rect 13313 16647 13314 16673
rect 11830 16002 11858 16254
rect 11942 16282 11970 16287
rect 11942 16235 11970 16254
rect 12073 16086 12535 16091
rect 12073 16085 12082 16086
rect 12073 16059 12074 16085
rect 12073 16058 12082 16059
rect 12110 16058 12134 16086
rect 12162 16058 12186 16086
rect 12214 16085 12238 16086
rect 12266 16085 12290 16086
rect 12224 16059 12238 16085
rect 12286 16059 12290 16085
rect 12214 16058 12238 16059
rect 12266 16058 12290 16059
rect 12318 16085 12342 16086
rect 12370 16085 12394 16086
rect 12318 16059 12322 16085
rect 12370 16059 12384 16085
rect 12318 16058 12342 16059
rect 12370 16058 12394 16059
rect 12422 16058 12446 16086
rect 12474 16058 12498 16086
rect 12526 16085 12535 16086
rect 12534 16059 12535 16085
rect 12526 16058 12535 16059
rect 12073 16053 12535 16058
rect 11830 15498 11858 15974
rect 12222 16002 12250 16007
rect 12222 15889 12250 15974
rect 12222 15863 12223 15889
rect 12249 15863 12250 15889
rect 12222 15857 12250 15863
rect 12446 16002 12474 16007
rect 12446 15889 12474 15974
rect 12446 15863 12447 15889
rect 12473 15863 12474 15889
rect 12446 15857 12474 15863
rect 13286 15946 13314 16647
rect 13286 15889 13314 15918
rect 13286 15863 13287 15889
rect 13313 15863 13314 15889
rect 11942 15498 11970 15503
rect 11830 15497 11970 15498
rect 11830 15471 11831 15497
rect 11857 15471 11943 15497
rect 11969 15471 11970 15497
rect 11830 15470 11970 15471
rect 11830 15465 11858 15470
rect 11942 15465 11970 15470
rect 12073 15302 12535 15307
rect 12073 15301 12082 15302
rect 12073 15275 12074 15301
rect 12073 15274 12082 15275
rect 12110 15274 12134 15302
rect 12162 15274 12186 15302
rect 12214 15301 12238 15302
rect 12266 15301 12290 15302
rect 12224 15275 12238 15301
rect 12286 15275 12290 15301
rect 12214 15274 12238 15275
rect 12266 15274 12290 15275
rect 12318 15301 12342 15302
rect 12370 15301 12394 15302
rect 12318 15275 12322 15301
rect 12370 15275 12384 15301
rect 12318 15274 12342 15275
rect 12370 15274 12394 15275
rect 12422 15274 12446 15302
rect 12474 15274 12498 15302
rect 12526 15301 12535 15302
rect 12534 15275 12535 15301
rect 12526 15274 12535 15275
rect 12073 15269 12535 15274
rect 11774 15079 11775 15105
rect 11801 15079 11802 15105
rect 11774 14321 11802 15079
rect 12726 15105 12754 15111
rect 12726 15079 12727 15105
rect 12753 15079 12754 15105
rect 12726 15050 12754 15079
rect 12446 15049 12754 15050
rect 12446 15023 12727 15049
rect 12753 15023 12754 15049
rect 12446 15022 12754 15023
rect 12446 14769 12474 15022
rect 12446 14743 12447 14769
rect 12473 14743 12474 14769
rect 12446 14713 12474 14743
rect 12446 14687 12447 14713
rect 12473 14687 12474 14713
rect 12446 14681 12474 14687
rect 12073 14518 12535 14523
rect 12073 14517 12082 14518
rect 12073 14491 12074 14517
rect 12073 14490 12082 14491
rect 12110 14490 12134 14518
rect 12162 14490 12186 14518
rect 12214 14517 12238 14518
rect 12266 14517 12290 14518
rect 12224 14491 12238 14517
rect 12286 14491 12290 14517
rect 12214 14490 12238 14491
rect 12266 14490 12290 14491
rect 12318 14517 12342 14518
rect 12370 14517 12394 14518
rect 12318 14491 12322 14517
rect 12370 14491 12384 14517
rect 12318 14490 12342 14491
rect 12370 14490 12394 14491
rect 12422 14490 12446 14518
rect 12474 14490 12498 14518
rect 12526 14517 12535 14518
rect 12534 14491 12535 14517
rect 12526 14490 12535 14491
rect 12073 14485 12535 14490
rect 12614 14322 12642 15022
rect 12726 15017 12754 15022
rect 13286 15105 13314 15863
rect 13734 17065 13762 17071
rect 13734 17039 13735 17065
rect 13761 17039 13762 17065
rect 13734 16281 13762 17039
rect 14238 16674 14266 17375
rect 15078 17457 15106 17823
rect 15806 18241 15834 18247
rect 15806 18215 15807 18241
rect 15833 18215 15834 18241
rect 15806 18185 15834 18215
rect 15806 18159 15807 18185
rect 15833 18159 15834 18185
rect 15806 17906 15834 18159
rect 15918 17906 15946 17911
rect 15806 17905 15946 17906
rect 15806 17879 15919 17905
rect 15945 17879 15946 17905
rect 15806 17878 15946 17879
rect 15806 17850 15834 17878
rect 15806 17817 15834 17822
rect 15918 17849 15946 17878
rect 15918 17823 15919 17849
rect 15945 17823 15946 17849
rect 15078 17431 15079 17457
rect 15105 17431 15106 17457
rect 14573 17262 15035 17267
rect 14573 17261 14582 17262
rect 14573 17235 14574 17261
rect 14573 17234 14582 17235
rect 14610 17234 14634 17262
rect 14662 17234 14686 17262
rect 14714 17261 14738 17262
rect 14766 17261 14790 17262
rect 14724 17235 14738 17261
rect 14786 17235 14790 17261
rect 14714 17234 14738 17235
rect 14766 17234 14790 17235
rect 14818 17261 14842 17262
rect 14870 17261 14894 17262
rect 14818 17235 14822 17261
rect 14870 17235 14884 17261
rect 14818 17234 14842 17235
rect 14870 17234 14894 17235
rect 14922 17234 14946 17262
rect 14974 17234 14998 17262
rect 15026 17261 15035 17262
rect 15034 17235 15035 17261
rect 15026 17234 15035 17235
rect 14573 17229 15035 17234
rect 14294 17066 14322 17071
rect 14462 17066 14490 17071
rect 14294 17065 14490 17066
rect 14294 17039 14295 17065
rect 14321 17039 14463 17065
rect 14489 17039 14490 17065
rect 14294 17038 14490 17039
rect 14294 17033 14322 17038
rect 14238 16617 14266 16646
rect 14238 16591 14239 16617
rect 14265 16591 14266 16617
rect 14238 16585 14266 16591
rect 13734 16255 13735 16281
rect 13761 16255 13762 16281
rect 13734 15946 13762 16255
rect 13734 15497 13762 15918
rect 14406 16282 14434 16287
rect 14462 16282 14490 17038
rect 15078 17066 15106 17431
rect 15918 17458 15946 17823
rect 17073 17654 17535 17659
rect 17073 17653 17082 17654
rect 17073 17627 17074 17653
rect 17073 17626 17082 17627
rect 17110 17626 17134 17654
rect 17162 17626 17186 17654
rect 17214 17653 17238 17654
rect 17266 17653 17290 17654
rect 17224 17627 17238 17653
rect 17286 17627 17290 17653
rect 17214 17626 17238 17627
rect 17266 17626 17290 17627
rect 17318 17653 17342 17654
rect 17370 17653 17394 17654
rect 17318 17627 17322 17653
rect 17370 17627 17384 17653
rect 17318 17626 17342 17627
rect 17370 17626 17394 17627
rect 17422 17626 17446 17654
rect 17474 17626 17498 17654
rect 17526 17653 17535 17654
rect 17534 17627 17535 17653
rect 17526 17626 17535 17627
rect 17073 17621 17535 17626
rect 15974 17458 16002 17463
rect 15918 17457 16002 17458
rect 15918 17431 15975 17457
rect 16001 17431 16002 17457
rect 15918 17430 16002 17431
rect 15974 17401 16002 17430
rect 15974 17375 15975 17401
rect 16001 17375 16002 17401
rect 15190 17066 15218 17071
rect 15078 17065 15218 17066
rect 15078 17039 15191 17065
rect 15217 17039 15218 17065
rect 15078 17038 15218 17039
rect 15078 16673 15106 17038
rect 15190 17033 15218 17038
rect 15974 17066 16002 17375
rect 16254 17457 16282 17463
rect 16254 17431 16255 17457
rect 16281 17431 16282 17457
rect 16142 17121 16170 17127
rect 16142 17095 16143 17121
rect 16169 17095 16170 17121
rect 16142 17066 16170 17095
rect 15974 17065 16170 17066
rect 15974 17039 15975 17065
rect 16001 17039 16170 17065
rect 15974 17038 16170 17039
rect 15078 16647 15079 16673
rect 15105 16647 15106 16673
rect 14573 16478 15035 16483
rect 14573 16477 14582 16478
rect 14573 16451 14574 16477
rect 14573 16450 14582 16451
rect 14610 16450 14634 16478
rect 14662 16450 14686 16478
rect 14714 16477 14738 16478
rect 14766 16477 14790 16478
rect 14724 16451 14738 16477
rect 14786 16451 14790 16477
rect 14714 16450 14738 16451
rect 14766 16450 14790 16451
rect 14818 16477 14842 16478
rect 14870 16477 14894 16478
rect 14818 16451 14822 16477
rect 14870 16451 14884 16477
rect 14818 16450 14842 16451
rect 14870 16450 14894 16451
rect 14922 16450 14946 16478
rect 14974 16450 14998 16478
rect 15026 16477 15035 16478
rect 15034 16451 15035 16477
rect 15026 16450 15035 16451
rect 14573 16445 15035 16450
rect 14630 16337 14658 16343
rect 14630 16311 14631 16337
rect 14657 16311 14658 16337
rect 14630 16282 14658 16311
rect 14406 16281 14658 16282
rect 14406 16255 14407 16281
rect 14433 16255 14658 16281
rect 14406 16254 14658 16255
rect 15078 16282 15106 16647
rect 15974 16673 16002 17038
rect 15974 16647 15975 16673
rect 16001 16647 16002 16673
rect 15974 16617 16002 16647
rect 15974 16591 15975 16617
rect 16001 16591 16002 16617
rect 15134 16282 15162 16287
rect 15078 16281 15162 16282
rect 15078 16255 15135 16281
rect 15161 16255 15162 16281
rect 15078 16254 15162 16255
rect 14406 15889 14434 16254
rect 14406 15863 14407 15889
rect 14433 15863 14434 15889
rect 14406 15834 14434 15863
rect 15078 15889 15106 16254
rect 15134 16249 15162 16254
rect 15974 16170 16002 16591
rect 15974 16137 16002 16142
rect 16254 16673 16282 17431
rect 16254 16647 16255 16673
rect 16281 16647 16282 16673
rect 16254 16282 16282 16647
rect 16758 17457 16786 17463
rect 16758 17431 16759 17457
rect 16785 17431 16786 17457
rect 16758 16674 16786 17431
rect 16926 17457 16954 17463
rect 16926 17431 16927 17457
rect 16953 17431 16954 17457
rect 15078 15863 15079 15889
rect 15105 15863 15106 15889
rect 14406 15833 14490 15834
rect 14406 15807 14407 15833
rect 14433 15807 14490 15833
rect 14406 15806 14490 15807
rect 14406 15801 14434 15806
rect 13734 15471 13735 15497
rect 13761 15471 13762 15497
rect 13734 15465 13762 15471
rect 14294 15498 14322 15503
rect 14462 15498 14490 15806
rect 14573 15694 15035 15699
rect 14573 15693 14582 15694
rect 14573 15667 14574 15693
rect 14573 15666 14582 15667
rect 14610 15666 14634 15694
rect 14662 15666 14686 15694
rect 14714 15693 14738 15694
rect 14766 15693 14790 15694
rect 14724 15667 14738 15693
rect 14786 15667 14790 15693
rect 14714 15666 14738 15667
rect 14766 15666 14790 15667
rect 14818 15693 14842 15694
rect 14870 15693 14894 15694
rect 14818 15667 14822 15693
rect 14870 15667 14884 15693
rect 14818 15666 14842 15667
rect 14870 15666 14894 15667
rect 14922 15666 14946 15694
rect 14974 15666 14998 15694
rect 15026 15693 15035 15694
rect 15034 15667 15035 15693
rect 15026 15666 15035 15667
rect 14573 15661 15035 15666
rect 14294 15497 14490 15498
rect 14294 15471 14295 15497
rect 14321 15471 14463 15497
rect 14489 15471 14490 15497
rect 14294 15470 14490 15471
rect 14294 15465 14322 15470
rect 13286 15079 13287 15105
rect 13313 15079 13314 15105
rect 11774 14295 11775 14321
rect 11801 14295 11802 14321
rect 11774 13537 11802 14295
rect 12446 14321 12754 14322
rect 12446 14295 12615 14321
rect 12641 14295 12754 14321
rect 12446 14294 12754 14295
rect 12446 13985 12474 14294
rect 12614 14289 12642 14294
rect 12726 14265 12754 14294
rect 12726 14239 12727 14265
rect 12753 14239 12754 14265
rect 12726 14233 12754 14239
rect 13286 14321 13314 15079
rect 14406 15105 14434 15111
rect 14406 15079 14407 15105
rect 14433 15079 14434 15105
rect 14406 15050 14434 15079
rect 14462 15050 14490 15470
rect 15078 15498 15106 15863
rect 15974 15889 16002 15895
rect 15974 15863 15975 15889
rect 16001 15863 16002 15889
rect 15974 15833 16002 15863
rect 15974 15807 15975 15833
rect 16001 15807 16002 15833
rect 15190 15498 15218 15503
rect 15078 15497 15218 15498
rect 15078 15471 15191 15497
rect 15217 15471 15218 15497
rect 15078 15470 15218 15471
rect 15078 15106 15106 15470
rect 15190 15465 15218 15470
rect 15974 15498 16002 15807
rect 16254 15889 16282 16254
rect 16310 16337 16338 16343
rect 16310 16311 16311 16337
rect 16337 16311 16338 16337
rect 16310 16281 16338 16311
rect 16310 16255 16311 16281
rect 16337 16255 16338 16281
rect 16310 16170 16338 16255
rect 16758 16170 16786 16646
rect 16814 17065 16842 17071
rect 16814 17039 16815 17065
rect 16841 17039 16842 17065
rect 16814 16282 16842 17039
rect 16926 16674 16954 17431
rect 17073 16870 17535 16875
rect 17073 16869 17082 16870
rect 17073 16843 17074 16869
rect 17073 16842 17082 16843
rect 17110 16842 17134 16870
rect 17162 16842 17186 16870
rect 17214 16869 17238 16870
rect 17266 16869 17290 16870
rect 17224 16843 17238 16869
rect 17286 16843 17290 16869
rect 17214 16842 17238 16843
rect 17266 16842 17290 16843
rect 17318 16869 17342 16870
rect 17370 16869 17394 16870
rect 17318 16843 17322 16869
rect 17370 16843 17384 16869
rect 17318 16842 17342 16843
rect 17370 16842 17394 16843
rect 17422 16842 17446 16870
rect 17474 16842 17498 16870
rect 17526 16869 17535 16870
rect 17534 16843 17535 16869
rect 17526 16842 17535 16843
rect 17073 16837 17535 16842
rect 16926 16627 16954 16646
rect 16814 16249 16842 16254
rect 16814 16170 16842 16175
rect 16758 16142 16814 16170
rect 16310 16137 16338 16142
rect 16254 15863 16255 15889
rect 16281 15863 16282 15889
rect 16142 15553 16170 15559
rect 16142 15527 16143 15553
rect 16169 15527 16170 15553
rect 16142 15498 16170 15527
rect 15974 15497 16170 15498
rect 15974 15471 15975 15497
rect 16001 15471 16170 15497
rect 15974 15470 16170 15471
rect 15078 15105 15218 15106
rect 15078 15079 15079 15105
rect 15105 15079 15218 15105
rect 15078 15078 15218 15079
rect 15078 15073 15106 15078
rect 14406 15049 14490 15050
rect 14406 15023 14407 15049
rect 14433 15023 14490 15049
rect 14406 15022 14490 15023
rect 14406 15017 14434 15022
rect 13286 14295 13287 14321
rect 13313 14295 13314 14321
rect 12446 13959 12447 13985
rect 12473 13959 12474 13985
rect 11774 13511 11775 13537
rect 11801 13511 11802 13537
rect 11774 12754 11802 13511
rect 11998 13930 12026 13935
rect 11830 13146 11858 13151
rect 11998 13146 12026 13902
rect 12446 13930 12474 13959
rect 12446 13864 12474 13902
rect 12073 13734 12535 13739
rect 12073 13733 12082 13734
rect 12073 13707 12074 13733
rect 12073 13706 12082 13707
rect 12110 13706 12134 13734
rect 12162 13706 12186 13734
rect 12214 13733 12238 13734
rect 12266 13733 12290 13734
rect 12224 13707 12238 13733
rect 12286 13707 12290 13733
rect 12214 13706 12238 13707
rect 12266 13706 12290 13707
rect 12318 13733 12342 13734
rect 12370 13733 12394 13734
rect 12318 13707 12322 13733
rect 12370 13707 12384 13733
rect 12318 13706 12342 13707
rect 12370 13706 12394 13707
rect 12422 13706 12446 13734
rect 12474 13706 12498 13734
rect 12526 13733 12535 13734
rect 12534 13707 12535 13733
rect 12526 13706 12535 13707
rect 12073 13701 12535 13706
rect 12222 13538 12250 13543
rect 12222 13146 12250 13510
rect 12950 13538 12978 13543
rect 12950 13481 12978 13510
rect 12950 13455 12951 13481
rect 12977 13455 12978 13481
rect 12950 13449 12978 13455
rect 13286 13537 13314 14295
rect 13734 14713 13762 14719
rect 13734 14687 13735 14713
rect 13761 14687 13762 14713
rect 13734 13929 13762 14687
rect 14294 14714 14322 14719
rect 14462 14714 14490 15022
rect 14573 14910 15035 14915
rect 14573 14909 14582 14910
rect 14573 14883 14574 14909
rect 14573 14882 14582 14883
rect 14610 14882 14634 14910
rect 14662 14882 14686 14910
rect 14714 14909 14738 14910
rect 14766 14909 14790 14910
rect 14724 14883 14738 14909
rect 14786 14883 14790 14909
rect 14714 14882 14738 14883
rect 14766 14882 14790 14883
rect 14818 14909 14842 14910
rect 14870 14909 14894 14910
rect 14818 14883 14822 14909
rect 14870 14883 14884 14909
rect 14818 14882 14842 14883
rect 14870 14882 14894 14883
rect 14922 14882 14946 14910
rect 14974 14882 14998 14910
rect 15026 14909 15035 14910
rect 15034 14883 15035 14909
rect 15026 14882 15035 14883
rect 14573 14877 15035 14882
rect 15190 14714 15218 15078
rect 14294 14713 14490 14714
rect 14294 14687 14295 14713
rect 14321 14687 14463 14713
rect 14489 14687 14490 14713
rect 14294 14686 14490 14687
rect 14294 14681 14322 14686
rect 14406 14322 14434 14327
rect 14462 14322 14490 14686
rect 14406 14321 14490 14322
rect 14406 14295 14407 14321
rect 14433 14295 14490 14321
rect 14406 14294 14490 14295
rect 14406 14265 14434 14294
rect 14406 14239 14407 14265
rect 14433 14239 14434 14265
rect 14406 14233 14434 14239
rect 14462 13930 14490 14294
rect 15078 14713 15218 14714
rect 15078 14687 15191 14713
rect 15217 14687 15218 14713
rect 15078 14686 15218 14687
rect 15078 14322 15106 14686
rect 15190 14681 15218 14686
rect 15974 15105 16002 15470
rect 15974 15079 15975 15105
rect 16001 15079 16002 15105
rect 15974 15049 16002 15079
rect 15974 15023 15975 15049
rect 16001 15023 16002 15049
rect 15190 14322 15218 14327
rect 15078 14321 15190 14322
rect 15078 14295 15079 14321
rect 15105 14295 15190 14321
rect 15078 14294 15190 14295
rect 15078 14289 15106 14294
rect 14573 14126 15035 14131
rect 14573 14125 14582 14126
rect 14573 14099 14574 14125
rect 14573 14098 14582 14099
rect 14610 14098 14634 14126
rect 14662 14098 14686 14126
rect 14714 14125 14738 14126
rect 14766 14125 14790 14126
rect 14724 14099 14738 14125
rect 14786 14099 14790 14125
rect 14714 14098 14738 14099
rect 14766 14098 14790 14099
rect 14818 14125 14842 14126
rect 14870 14125 14894 14126
rect 14818 14099 14822 14125
rect 14870 14099 14884 14125
rect 14818 14098 14842 14099
rect 14870 14098 14894 14099
rect 14922 14098 14946 14126
rect 14974 14098 14998 14126
rect 15026 14125 15035 14126
rect 15034 14099 15035 14125
rect 15026 14098 15035 14099
rect 14573 14093 15035 14098
rect 13734 13903 13735 13929
rect 13761 13903 13762 13929
rect 13286 13511 13287 13537
rect 13313 13511 13314 13537
rect 13286 13454 13314 13511
rect 11830 13145 12250 13146
rect 11830 13119 11831 13145
rect 11857 13119 11999 13145
rect 12025 13119 12250 13145
rect 11830 13118 12250 13119
rect 13230 13426 13314 13454
rect 13678 13538 13706 13543
rect 13230 13146 13258 13398
rect 13678 13314 13706 13510
rect 13734 13426 13762 13903
rect 14406 13902 14462 13930
rect 14126 13537 14154 13543
rect 14126 13511 14127 13537
rect 14153 13511 14154 13537
rect 13734 13393 13762 13398
rect 13790 13482 13818 13487
rect 13790 13314 13818 13454
rect 14126 13482 14154 13511
rect 14406 13538 14434 13902
rect 14462 13897 14490 13902
rect 14910 13985 14938 13991
rect 14910 13959 14911 13985
rect 14937 13959 14938 13985
rect 14910 13930 14938 13959
rect 14910 13883 14938 13902
rect 15190 13929 15218 14294
rect 15190 13903 15191 13929
rect 15217 13903 15218 13929
rect 15190 13897 15218 13903
rect 15974 14321 16002 15023
rect 15974 14295 15975 14321
rect 16001 14295 16002 14321
rect 15974 14266 16002 14295
rect 16254 15105 16282 15863
rect 16814 15890 16842 16142
rect 17073 16086 17535 16091
rect 17073 16085 17082 16086
rect 17073 16059 17074 16085
rect 17073 16058 17082 16059
rect 17110 16058 17134 16086
rect 17162 16058 17186 16086
rect 17214 16085 17238 16086
rect 17266 16085 17290 16086
rect 17224 16059 17238 16085
rect 17286 16059 17290 16085
rect 17214 16058 17238 16059
rect 17266 16058 17290 16059
rect 17318 16085 17342 16086
rect 17370 16085 17394 16086
rect 17318 16059 17322 16085
rect 17370 16059 17384 16085
rect 17318 16058 17342 16059
rect 17370 16058 17394 16059
rect 17422 16058 17446 16086
rect 17474 16058 17498 16086
rect 17526 16085 17535 16086
rect 17534 16059 17535 16085
rect 17526 16058 17535 16059
rect 17073 16053 17535 16058
rect 16926 15890 16954 15895
rect 16814 15889 16954 15890
rect 16814 15863 16815 15889
rect 16841 15863 16927 15889
rect 16953 15863 16954 15889
rect 16814 15862 16954 15863
rect 16814 15857 16842 15862
rect 16814 15497 16842 15503
rect 16814 15471 16815 15497
rect 16841 15471 16842 15497
rect 16254 15079 16255 15105
rect 16281 15079 16282 15105
rect 16254 14322 16282 15079
rect 16254 14275 16282 14294
rect 16310 15162 16338 15167
rect 15974 13930 16002 14238
rect 15974 13897 16002 13902
rect 14406 13481 14434 13510
rect 14406 13455 14407 13481
rect 14433 13455 14434 13481
rect 14126 13426 14210 13454
rect 14406 13449 14434 13455
rect 15470 13537 15498 13543
rect 15470 13511 15471 13537
rect 15497 13511 15498 13537
rect 13678 13286 13818 13314
rect 13398 13146 13426 13151
rect 13230 13145 13426 13146
rect 13230 13119 13399 13145
rect 13425 13119 13426 13145
rect 13230 13118 13426 13119
rect 11830 13113 11858 13118
rect 11270 11774 11298 11942
rect 11718 11970 11746 11975
rect 11774 11970 11802 12726
rect 11830 12362 11858 12367
rect 11998 12362 12026 13118
rect 12073 12950 12535 12955
rect 12073 12949 12082 12950
rect 12073 12923 12074 12949
rect 12073 12922 12082 12923
rect 12110 12922 12134 12950
rect 12162 12922 12186 12950
rect 12214 12949 12238 12950
rect 12266 12949 12290 12950
rect 12224 12923 12238 12949
rect 12286 12923 12290 12949
rect 12214 12922 12238 12923
rect 12266 12922 12290 12923
rect 12318 12949 12342 12950
rect 12370 12949 12394 12950
rect 12318 12923 12322 12949
rect 12370 12923 12384 12949
rect 12318 12922 12342 12923
rect 12370 12922 12394 12923
rect 12422 12922 12446 12950
rect 12474 12922 12498 12950
rect 12526 12949 12535 12950
rect 12534 12923 12535 12949
rect 12526 12922 12535 12923
rect 12073 12917 12535 12922
rect 12222 12754 12250 12759
rect 12446 12754 12474 12759
rect 12222 12753 12474 12754
rect 12222 12727 12223 12753
rect 12249 12727 12447 12753
rect 12473 12727 12474 12753
rect 12222 12726 12474 12727
rect 12222 12362 12250 12726
rect 12446 12721 12474 12726
rect 13230 12754 13258 13118
rect 13398 13113 13426 13118
rect 14182 13146 14210 13426
rect 14573 13342 15035 13347
rect 14573 13341 14582 13342
rect 14573 13315 14574 13341
rect 14573 13314 14582 13315
rect 14610 13314 14634 13342
rect 14662 13314 14686 13342
rect 14714 13341 14738 13342
rect 14766 13341 14790 13342
rect 14724 13315 14738 13341
rect 14786 13315 14790 13341
rect 14714 13314 14738 13315
rect 14766 13314 14790 13315
rect 14818 13341 14842 13342
rect 14870 13341 14894 13342
rect 14818 13315 14822 13341
rect 14870 13315 14884 13341
rect 14818 13314 14842 13315
rect 14870 13314 14894 13315
rect 14922 13314 14946 13342
rect 14974 13314 14998 13342
rect 15026 13341 15035 13342
rect 15034 13315 15035 13341
rect 15026 13314 15035 13315
rect 14573 13309 15035 13314
rect 14350 13201 14378 13207
rect 14350 13175 14351 13201
rect 14377 13175 14378 13201
rect 14350 13146 14378 13175
rect 14182 13145 14378 13146
rect 14182 13119 14183 13145
rect 14209 13119 14378 13145
rect 14182 13118 14378 13119
rect 15134 13146 15162 13151
rect 13230 12707 13258 12726
rect 14182 12753 14210 13118
rect 15134 13099 15162 13118
rect 15470 13146 15498 13511
rect 16254 13538 16282 13543
rect 16310 13538 16338 15134
rect 16366 14769 16394 14775
rect 16366 14743 16367 14769
rect 16393 14743 16394 14769
rect 16366 14713 16394 14743
rect 16366 14687 16367 14713
rect 16393 14687 16394 14713
rect 16366 14266 16394 14687
rect 16366 13985 16394 14238
rect 16366 13959 16367 13985
rect 16393 13959 16394 13985
rect 16366 13929 16394 13959
rect 16366 13903 16367 13929
rect 16393 13903 16394 13929
rect 16366 13897 16394 13903
rect 16814 14713 16842 15471
rect 16926 15162 16954 15862
rect 17073 15302 17535 15307
rect 17073 15301 17082 15302
rect 17073 15275 17074 15301
rect 17073 15274 17082 15275
rect 17110 15274 17134 15302
rect 17162 15274 17186 15302
rect 17214 15301 17238 15302
rect 17266 15301 17290 15302
rect 17224 15275 17238 15301
rect 17286 15275 17290 15301
rect 17214 15274 17238 15275
rect 17266 15274 17290 15275
rect 17318 15301 17342 15302
rect 17370 15301 17394 15302
rect 17318 15275 17322 15301
rect 17370 15275 17384 15301
rect 17318 15274 17342 15275
rect 17370 15274 17394 15275
rect 17422 15274 17446 15302
rect 17474 15274 17498 15302
rect 17526 15301 17535 15302
rect 17534 15275 17535 15301
rect 17526 15274 17535 15275
rect 17073 15269 17535 15274
rect 16926 15129 16954 15134
rect 16814 14687 16815 14713
rect 16841 14687 16842 14713
rect 16814 14322 16842 14687
rect 16814 13929 16842 14294
rect 16982 15105 17010 15111
rect 16982 15079 16983 15105
rect 17009 15079 17010 15105
rect 16982 15050 17010 15079
rect 17206 15050 17234 15055
rect 16982 15049 17234 15050
rect 16982 15023 17207 15049
rect 17233 15023 17234 15049
rect 16982 15022 17234 15023
rect 16982 14266 17010 15022
rect 17206 15017 17234 15022
rect 17073 14518 17535 14523
rect 17073 14517 17082 14518
rect 17073 14491 17074 14517
rect 17073 14490 17082 14491
rect 17110 14490 17134 14518
rect 17162 14490 17186 14518
rect 17214 14517 17238 14518
rect 17266 14517 17290 14518
rect 17224 14491 17238 14517
rect 17286 14491 17290 14517
rect 17214 14490 17238 14491
rect 17266 14490 17290 14491
rect 17318 14517 17342 14518
rect 17370 14517 17394 14518
rect 17318 14491 17322 14517
rect 17370 14491 17384 14517
rect 17318 14490 17342 14491
rect 17370 14490 17394 14491
rect 17422 14490 17446 14518
rect 17474 14490 17498 14518
rect 17526 14517 17535 14518
rect 17534 14491 17535 14517
rect 17526 14490 17535 14491
rect 17073 14485 17535 14490
rect 16982 14233 17010 14238
rect 17430 14321 17458 14327
rect 17430 14295 17431 14321
rect 17457 14295 17458 14321
rect 17430 14266 17458 14295
rect 17430 14219 17458 14238
rect 16814 13903 16815 13929
rect 16841 13903 16842 13929
rect 16254 13537 16338 13538
rect 16254 13511 16255 13537
rect 16281 13511 16338 13537
rect 16254 13510 16338 13511
rect 16814 13538 16842 13903
rect 17073 13734 17535 13739
rect 17073 13733 17082 13734
rect 17073 13707 17074 13733
rect 17073 13706 17082 13707
rect 17110 13706 17134 13734
rect 17162 13706 17186 13734
rect 17214 13733 17238 13734
rect 17266 13733 17290 13734
rect 17224 13707 17238 13733
rect 17286 13707 17290 13733
rect 17214 13706 17238 13707
rect 17266 13706 17290 13707
rect 17318 13733 17342 13734
rect 17370 13733 17394 13734
rect 17318 13707 17322 13733
rect 17370 13707 17384 13733
rect 17318 13706 17342 13707
rect 17370 13706 17394 13707
rect 17422 13706 17446 13734
rect 17474 13706 17498 13734
rect 17526 13733 17535 13734
rect 17534 13707 17535 13733
rect 17526 13706 17535 13707
rect 17073 13701 17535 13706
rect 16814 13537 17010 13538
rect 16814 13511 16815 13537
rect 16841 13511 17010 13537
rect 16814 13510 17010 13511
rect 16254 13481 16282 13510
rect 16814 13505 16842 13510
rect 16254 13455 16255 13481
rect 16281 13455 16282 13481
rect 16254 13454 16282 13455
rect 16030 13426 16282 13454
rect 16814 13454 16842 13459
rect 16030 13201 16058 13426
rect 16030 13175 16031 13201
rect 16057 13175 16058 13201
rect 15470 13113 15498 13118
rect 15750 13146 15778 13151
rect 14182 12727 14183 12753
rect 14209 12727 14210 12753
rect 14182 12697 14210 12727
rect 15750 12754 15778 13118
rect 16030 13145 16058 13175
rect 16030 13119 16031 13145
rect 16057 13119 16058 13145
rect 15750 12753 15890 12754
rect 15750 12727 15751 12753
rect 15777 12727 15890 12753
rect 15750 12726 15890 12727
rect 15750 12721 15778 12726
rect 14182 12671 14183 12697
rect 14209 12671 14210 12697
rect 14182 12665 14210 12671
rect 14573 12558 15035 12563
rect 14573 12557 14582 12558
rect 14573 12531 14574 12557
rect 14573 12530 14582 12531
rect 14610 12530 14634 12558
rect 14662 12530 14686 12558
rect 14714 12557 14738 12558
rect 14766 12557 14790 12558
rect 14724 12531 14738 12557
rect 14786 12531 14790 12557
rect 14714 12530 14738 12531
rect 14766 12530 14790 12531
rect 14818 12557 14842 12558
rect 14870 12557 14894 12558
rect 14818 12531 14822 12557
rect 14870 12531 14884 12557
rect 14818 12530 14842 12531
rect 14870 12530 14894 12531
rect 14922 12530 14946 12558
rect 14974 12530 14998 12558
rect 15026 12557 15035 12558
rect 15034 12531 15035 12557
rect 15026 12530 15035 12531
rect 14573 12525 15035 12530
rect 14966 12417 14994 12423
rect 14966 12391 14967 12417
rect 14993 12391 14994 12417
rect 11830 12361 12250 12362
rect 11830 12335 11831 12361
rect 11857 12335 11999 12361
rect 12025 12335 12250 12361
rect 11830 12334 12250 12335
rect 14070 12361 14098 12367
rect 14070 12335 14071 12361
rect 14097 12335 14098 12361
rect 11830 12329 11858 12334
rect 11746 11969 11802 11970
rect 11746 11943 11775 11969
rect 11801 11943 11802 11969
rect 11746 11942 11802 11943
rect 11718 11937 11746 11942
rect 11774 11937 11802 11942
rect 11998 11970 12026 12334
rect 12073 12166 12535 12171
rect 12073 12165 12082 12166
rect 12073 12139 12074 12165
rect 12073 12138 12082 12139
rect 12110 12138 12134 12166
rect 12162 12138 12186 12166
rect 12214 12165 12238 12166
rect 12266 12165 12290 12166
rect 12224 12139 12238 12165
rect 12286 12139 12290 12165
rect 12214 12138 12238 12139
rect 12266 12138 12290 12139
rect 12318 12165 12342 12166
rect 12370 12165 12394 12166
rect 12318 12139 12322 12165
rect 12370 12139 12384 12165
rect 12318 12138 12342 12139
rect 12370 12138 12394 12139
rect 12422 12138 12446 12166
rect 12474 12138 12498 12166
rect 12526 12165 12535 12166
rect 12534 12139 12535 12165
rect 12526 12138 12535 12139
rect 12073 12133 12535 12138
rect 12222 11970 12250 11975
rect 12446 11970 12474 11975
rect 11998 11969 12474 11970
rect 11998 11943 12223 11969
rect 12249 11943 12447 11969
rect 12473 11943 12474 11969
rect 11998 11942 12474 11943
rect 11270 11746 11354 11774
rect 10486 11578 10514 11583
rect 10374 11577 10514 11578
rect 10374 11551 10375 11577
rect 10401 11551 10487 11577
rect 10513 11551 10514 11577
rect 10374 11550 10514 11551
rect 9478 11159 9479 11185
rect 9505 11159 9506 11185
rect 9478 10794 9506 11159
rect 10374 11185 10402 11550
rect 10486 11545 10514 11550
rect 11326 11577 11354 11746
rect 11326 11551 11327 11577
rect 11353 11551 11354 11577
rect 10374 11159 10375 11185
rect 10401 11159 10402 11185
rect 10374 11130 10402 11159
rect 9573 10990 10035 10995
rect 9573 10989 9582 10990
rect 9573 10963 9574 10989
rect 9573 10962 9582 10963
rect 9610 10962 9634 10990
rect 9662 10962 9686 10990
rect 9714 10989 9738 10990
rect 9766 10989 9790 10990
rect 9724 10963 9738 10989
rect 9786 10963 9790 10989
rect 9714 10962 9738 10963
rect 9766 10962 9790 10963
rect 9818 10989 9842 10990
rect 9870 10989 9894 10990
rect 9818 10963 9822 10989
rect 9870 10963 9884 10989
rect 9818 10962 9842 10963
rect 9870 10962 9894 10963
rect 9922 10962 9946 10990
rect 9974 10962 9998 10990
rect 10026 10989 10035 10990
rect 10034 10963 10035 10989
rect 10026 10962 10035 10963
rect 9573 10957 10035 10962
rect 9814 10794 9842 10799
rect 9478 10793 9842 10794
rect 9478 10767 9815 10793
rect 9841 10767 9842 10793
rect 9478 10766 9842 10767
rect 9478 10401 9506 10766
rect 9814 10761 9842 10766
rect 10374 10794 10402 11102
rect 10486 10794 10514 10799
rect 10374 10793 10514 10794
rect 10374 10767 10375 10793
rect 10401 10767 10487 10793
rect 10513 10767 10514 10793
rect 10374 10766 10514 10767
rect 9478 10375 9479 10401
rect 9505 10375 9506 10401
rect 9478 10010 9506 10375
rect 10374 10401 10402 10766
rect 10486 10761 10514 10766
rect 11326 10793 11354 11551
rect 11830 11578 11858 11583
rect 11998 11578 12026 11942
rect 12222 11937 12250 11942
rect 12446 11937 12474 11942
rect 13230 11969 13258 11975
rect 13230 11943 13231 11969
rect 13257 11943 13258 11969
rect 11830 11577 12026 11578
rect 11830 11551 11831 11577
rect 11857 11551 11999 11577
rect 12025 11551 12026 11577
rect 11830 11550 12026 11551
rect 11830 11545 11858 11550
rect 11326 10767 11327 10793
rect 11353 10767 11354 10793
rect 10374 10375 10375 10401
rect 10401 10375 10402 10401
rect 10374 10345 10402 10375
rect 10374 10319 10375 10345
rect 10401 10319 10402 10345
rect 9573 10206 10035 10211
rect 9573 10205 9582 10206
rect 9573 10179 9574 10205
rect 9573 10178 9582 10179
rect 9610 10178 9634 10206
rect 9662 10178 9686 10206
rect 9714 10205 9738 10206
rect 9766 10205 9790 10206
rect 9724 10179 9738 10205
rect 9786 10179 9790 10205
rect 9714 10178 9738 10179
rect 9766 10178 9790 10179
rect 9818 10205 9842 10206
rect 9870 10205 9894 10206
rect 9818 10179 9822 10205
rect 9870 10179 9884 10205
rect 9818 10178 9842 10179
rect 9870 10178 9894 10179
rect 9922 10178 9946 10206
rect 9974 10178 9998 10206
rect 10026 10205 10035 10206
rect 10034 10179 10035 10205
rect 10026 10178 10035 10179
rect 9573 10173 10035 10178
rect 9814 10010 9842 10015
rect 9478 10009 9842 10010
rect 9478 9983 9815 10009
rect 9841 9983 9842 10009
rect 9478 9982 9842 9983
rect 9478 9617 9506 9982
rect 9814 9977 9842 9982
rect 10374 10010 10402 10319
rect 11326 10094 11354 10767
rect 11774 11185 11802 11191
rect 11774 11159 11775 11185
rect 11801 11159 11802 11185
rect 11774 10402 11802 11159
rect 11830 10794 11858 10799
rect 11998 10794 12026 11550
rect 12073 11382 12535 11387
rect 12073 11381 12082 11382
rect 12073 11355 12074 11381
rect 12073 11354 12082 11355
rect 12110 11354 12134 11382
rect 12162 11354 12186 11382
rect 12214 11381 12238 11382
rect 12266 11381 12290 11382
rect 12224 11355 12238 11381
rect 12286 11355 12290 11381
rect 12214 11354 12238 11355
rect 12266 11354 12290 11355
rect 12318 11381 12342 11382
rect 12370 11381 12394 11382
rect 12318 11355 12322 11381
rect 12370 11355 12384 11381
rect 12318 11354 12342 11355
rect 12370 11354 12394 11355
rect 12422 11354 12446 11382
rect 12474 11354 12498 11382
rect 12526 11381 12535 11382
rect 12534 11355 12535 11381
rect 12526 11354 12535 11355
rect 12073 11349 12535 11354
rect 11830 10793 12026 10794
rect 11830 10767 11831 10793
rect 11857 10767 11999 10793
rect 12025 10767 12026 10793
rect 11830 10766 12026 10767
rect 11830 10761 11858 10766
rect 11998 10514 12026 10766
rect 12950 11185 12978 11191
rect 12950 11159 12951 11185
rect 12977 11159 12978 11185
rect 12950 11129 12978 11159
rect 13230 11186 13258 11943
rect 14070 11577 14098 12335
rect 14966 12362 14994 12391
rect 15526 12362 15554 12367
rect 15862 12362 15890 12726
rect 16030 12418 16058 13119
rect 16646 12753 16674 12759
rect 16646 12727 16647 12753
rect 16673 12727 16674 12753
rect 16646 12697 16674 12727
rect 16646 12671 16647 12697
rect 16673 12671 16674 12697
rect 16030 12385 16058 12390
rect 16422 12418 16450 12423
rect 14966 12361 15106 12362
rect 14966 12335 14967 12361
rect 14993 12335 15106 12361
rect 14966 12334 15106 12335
rect 14966 12329 14994 12334
rect 14070 11551 14071 11577
rect 14097 11551 14098 11577
rect 13230 11153 13258 11158
rect 13510 11186 13538 11191
rect 12950 11103 12951 11129
rect 12977 11103 12978 11129
rect 12073 10598 12535 10603
rect 12073 10597 12082 10598
rect 12073 10571 12074 10597
rect 12073 10570 12082 10571
rect 12110 10570 12134 10598
rect 12162 10570 12186 10598
rect 12214 10597 12238 10598
rect 12266 10597 12290 10598
rect 12224 10571 12238 10597
rect 12286 10571 12290 10597
rect 12214 10570 12238 10571
rect 12266 10570 12290 10571
rect 12318 10597 12342 10598
rect 12370 10597 12394 10598
rect 12318 10571 12322 10597
rect 12370 10571 12384 10597
rect 12318 10570 12342 10571
rect 12370 10570 12394 10571
rect 12422 10570 12446 10598
rect 12474 10570 12498 10598
rect 12526 10597 12535 10598
rect 12534 10571 12535 10597
rect 12526 10570 12535 10571
rect 12073 10565 12535 10570
rect 11998 10486 12082 10514
rect 11886 10402 11914 10407
rect 11774 10401 11914 10402
rect 11774 10375 11887 10401
rect 11913 10375 11914 10401
rect 11774 10374 11914 10375
rect 11326 10066 11578 10094
rect 10486 10010 10514 10015
rect 10374 10009 10514 10010
rect 10374 9983 10375 10009
rect 10401 9983 10487 10009
rect 10513 9983 10514 10009
rect 10374 9982 10514 9983
rect 10374 9977 10402 9982
rect 9478 9591 9479 9617
rect 9505 9591 9506 9617
rect 9478 9226 9506 9591
rect 10430 9618 10458 9623
rect 10486 9618 10514 9982
rect 10430 9617 10514 9618
rect 10430 9591 10431 9617
rect 10457 9591 10514 9617
rect 10430 9590 10514 9591
rect 11270 10009 11298 10015
rect 11270 9983 11271 10009
rect 11297 9983 11298 10009
rect 10430 9561 10458 9590
rect 10430 9535 10431 9561
rect 10457 9535 10458 9561
rect 9573 9422 10035 9427
rect 9573 9421 9582 9422
rect 9573 9395 9574 9421
rect 9573 9394 9582 9395
rect 9610 9394 9634 9422
rect 9662 9394 9686 9422
rect 9714 9421 9738 9422
rect 9766 9421 9790 9422
rect 9724 9395 9738 9421
rect 9786 9395 9790 9421
rect 9714 9394 9738 9395
rect 9766 9394 9790 9395
rect 9818 9421 9842 9422
rect 9870 9421 9894 9422
rect 9818 9395 9822 9421
rect 9870 9395 9884 9421
rect 9818 9394 9842 9395
rect 9870 9394 9894 9395
rect 9922 9394 9946 9422
rect 9974 9394 9998 9422
rect 10026 9421 10035 9422
rect 10034 9395 10035 9421
rect 10026 9394 10035 9395
rect 9573 9389 10035 9394
rect 10430 9282 10458 9535
rect 10878 9282 10906 9287
rect 10430 9281 10906 9282
rect 10430 9255 10879 9281
rect 10905 9255 10906 9281
rect 10430 9254 10906 9255
rect 9254 8833 9282 8839
rect 9254 8807 9255 8833
rect 9281 8807 9282 8833
rect 9254 8442 9282 8807
rect 9254 8049 9282 8414
rect 9254 8023 9255 8049
rect 9281 8023 9282 8049
rect 9254 7658 9282 8023
rect 9254 7574 9282 7630
rect 9254 7546 9450 7574
rect 9422 7265 9450 7546
rect 9422 7239 9423 7265
rect 9449 7239 9450 7265
rect 8862 3425 8890 3430
rect 8974 6481 9002 6487
rect 8974 6455 8975 6481
rect 9001 6455 9002 6481
rect 8974 6425 9002 6455
rect 8974 6399 8975 6425
rect 9001 6399 9002 6425
rect 8974 5697 9002 6399
rect 8974 5671 8975 5697
rect 9001 5671 9002 5697
rect 8974 5641 9002 5671
rect 8974 5615 8975 5641
rect 9001 5615 9002 5641
rect 8974 4913 9002 5615
rect 8974 4887 8975 4913
rect 9001 4887 9002 4913
rect 8974 4857 9002 4887
rect 8974 4831 8975 4857
rect 9001 4831 9002 4857
rect 8974 4522 9002 4831
rect 8974 4129 9002 4494
rect 8974 4103 8975 4129
rect 9001 4103 9002 4129
rect 8974 4073 9002 4103
rect 9422 6481 9450 7239
rect 9422 6455 9423 6481
rect 9449 6455 9450 6481
rect 9422 5697 9450 6455
rect 9422 5671 9423 5697
rect 9449 5671 9450 5697
rect 9422 4913 9450 5671
rect 9422 4887 9423 4913
rect 9449 4887 9450 4913
rect 9422 4130 9450 4887
rect 9422 4097 9450 4102
rect 8974 4047 8975 4073
rect 9001 4047 9002 4073
rect 8974 3346 9002 4047
rect 8974 3289 9002 3318
rect 8974 3263 8975 3289
rect 9001 3263 9002 3289
rect 8974 3257 9002 3263
rect 8470 3010 8498 3015
rect 8358 3009 8498 3010
rect 8358 2983 8471 3009
rect 8497 2983 8498 3009
rect 8358 2982 8498 2983
rect 7014 2927 7015 2953
rect 7041 2927 7042 2953
rect 7014 2921 7042 2927
rect 7574 2953 7602 2959
rect 7574 2927 7575 2953
rect 7601 2927 7602 2953
rect 7073 2758 7535 2763
rect 7073 2757 7082 2758
rect 7073 2731 7074 2757
rect 7073 2730 7082 2731
rect 7110 2730 7134 2758
rect 7162 2730 7186 2758
rect 7214 2757 7238 2758
rect 7266 2757 7290 2758
rect 7224 2731 7238 2757
rect 7286 2731 7290 2757
rect 7214 2730 7238 2731
rect 7266 2730 7290 2731
rect 7318 2757 7342 2758
rect 7370 2757 7394 2758
rect 7318 2731 7322 2757
rect 7370 2731 7384 2757
rect 7318 2730 7342 2731
rect 7370 2730 7394 2731
rect 7422 2730 7446 2758
rect 7474 2730 7498 2758
rect 7526 2757 7535 2758
rect 7534 2731 7535 2757
rect 7526 2730 7535 2731
rect 7073 2725 7535 2730
rect 7294 2170 7322 2175
rect 7294 2123 7322 2142
rect 7574 2170 7602 2927
rect 8470 2953 8498 2982
rect 8470 2927 8471 2953
rect 8497 2927 8498 2953
rect 7073 1974 7535 1979
rect 7073 1973 7082 1974
rect 7073 1947 7074 1973
rect 7073 1946 7082 1947
rect 7110 1946 7134 1974
rect 7162 1946 7186 1974
rect 7214 1973 7238 1974
rect 7266 1973 7290 1974
rect 7224 1947 7238 1973
rect 7286 1947 7290 1973
rect 7214 1946 7238 1947
rect 7266 1946 7290 1947
rect 7318 1973 7342 1974
rect 7370 1973 7394 1974
rect 7318 1947 7322 1973
rect 7370 1947 7384 1973
rect 7318 1946 7342 1947
rect 7370 1946 7394 1947
rect 7422 1946 7446 1974
rect 7474 1946 7498 1974
rect 7526 1973 7535 1974
rect 7534 1947 7535 1973
rect 7526 1946 7535 1947
rect 7073 1941 7535 1946
rect 7574 1890 7602 2142
rect 7798 2561 7826 2567
rect 7798 2535 7799 2561
rect 7825 2535 7826 2561
rect 7798 2170 7826 2535
rect 7798 2137 7826 2142
rect 8470 2506 8498 2927
rect 8470 2225 8498 2478
rect 8974 2561 9002 2567
rect 8974 2535 8975 2561
rect 9001 2535 9002 2561
rect 8974 2506 9002 2535
rect 8974 2459 9002 2478
rect 8470 2199 8471 2225
rect 8497 2199 8498 2225
rect 8470 2169 8498 2199
rect 8470 2143 8471 2169
rect 8497 2143 8498 2169
rect 8470 2137 8498 2143
rect 7462 1778 7490 1783
rect 7574 1778 7602 1862
rect 8302 1890 8330 1895
rect 7462 1777 7602 1778
rect 7462 1751 7463 1777
rect 7489 1751 7602 1777
rect 7462 1750 7602 1751
rect 8134 1778 8162 1783
rect 7462 1745 7490 1750
rect 8134 1721 8162 1750
rect 8134 1695 8135 1721
rect 8161 1695 8162 1721
rect 8134 1689 8162 1695
rect 8302 400 8330 1862
rect 9422 1890 9450 1895
rect 9422 1777 9450 1862
rect 9422 1751 9423 1777
rect 9449 1751 9450 1777
rect 9422 1745 9450 1751
rect 9478 1498 9506 9198
rect 9814 9226 9842 9231
rect 9814 9179 9842 9198
rect 10878 9225 10906 9254
rect 10878 9199 10879 9225
rect 10905 9199 10906 9225
rect 10262 8833 10290 8839
rect 10262 8807 10263 8833
rect 10289 8807 10290 8833
rect 10262 8777 10290 8807
rect 10262 8751 10263 8777
rect 10289 8751 10290 8777
rect 9573 8638 10035 8643
rect 9573 8637 9582 8638
rect 9573 8611 9574 8637
rect 9573 8610 9582 8611
rect 9610 8610 9634 8638
rect 9662 8610 9686 8638
rect 9714 8637 9738 8638
rect 9766 8637 9790 8638
rect 9724 8611 9738 8637
rect 9786 8611 9790 8637
rect 9714 8610 9738 8611
rect 9766 8610 9790 8611
rect 9818 8637 9842 8638
rect 9870 8637 9894 8638
rect 9818 8611 9822 8637
rect 9870 8611 9884 8637
rect 9818 8610 9842 8611
rect 9870 8610 9894 8611
rect 9922 8610 9946 8638
rect 9974 8610 9998 8638
rect 10026 8637 10035 8638
rect 10034 8611 10035 8637
rect 10026 8610 10035 8611
rect 9573 8605 10035 8610
rect 10262 8498 10290 8751
rect 9814 8442 9842 8447
rect 9814 8395 9842 8414
rect 10262 8442 10290 8470
rect 10486 8442 10514 8447
rect 10262 8441 10514 8442
rect 10262 8415 10263 8441
rect 10289 8415 10487 8441
rect 10513 8415 10514 8441
rect 10262 8414 10514 8415
rect 10262 8049 10290 8414
rect 10486 8409 10514 8414
rect 10262 8023 10263 8049
rect 10289 8023 10290 8049
rect 10262 7993 10290 8023
rect 10262 7967 10263 7993
rect 10289 7967 10290 7993
rect 9573 7854 10035 7859
rect 9573 7853 9582 7854
rect 9573 7827 9574 7853
rect 9573 7826 9582 7827
rect 9610 7826 9634 7854
rect 9662 7826 9686 7854
rect 9714 7853 9738 7854
rect 9766 7853 9790 7854
rect 9724 7827 9738 7853
rect 9786 7827 9790 7853
rect 9714 7826 9738 7827
rect 9766 7826 9790 7827
rect 9818 7853 9842 7854
rect 9870 7853 9894 7854
rect 9818 7827 9822 7853
rect 9870 7827 9884 7853
rect 9818 7826 9842 7827
rect 9870 7826 9894 7827
rect 9922 7826 9946 7854
rect 9974 7826 9998 7854
rect 10026 7853 10035 7854
rect 10034 7827 10035 7853
rect 10026 7826 10035 7827
rect 9573 7821 10035 7826
rect 9814 7658 9842 7663
rect 9814 7611 9842 7630
rect 10262 7658 10290 7967
rect 10486 7658 10514 7663
rect 10262 7657 10514 7658
rect 10262 7631 10263 7657
rect 10289 7631 10487 7657
rect 10513 7631 10514 7657
rect 10262 7630 10514 7631
rect 10206 7546 10234 7551
rect 10206 7265 10234 7518
rect 10206 7239 10207 7265
rect 10233 7239 10234 7265
rect 10206 7209 10234 7239
rect 10206 7183 10207 7209
rect 10233 7183 10234 7209
rect 9573 7070 10035 7075
rect 9573 7069 9582 7070
rect 9573 7043 9574 7069
rect 9573 7042 9582 7043
rect 9610 7042 9634 7070
rect 9662 7042 9686 7070
rect 9714 7069 9738 7070
rect 9766 7069 9790 7070
rect 9724 7043 9738 7069
rect 9786 7043 9790 7069
rect 9714 7042 9738 7043
rect 9766 7042 9790 7043
rect 9818 7069 9842 7070
rect 9870 7069 9894 7070
rect 9818 7043 9822 7069
rect 9870 7043 9884 7069
rect 9818 7042 9842 7043
rect 9870 7042 9894 7043
rect 9922 7042 9946 7070
rect 9974 7042 9998 7070
rect 10026 7069 10035 7070
rect 10034 7043 10035 7069
rect 10026 7042 10035 7043
rect 9573 7037 10035 7042
rect 10038 6873 10066 6879
rect 10038 6847 10039 6873
rect 10065 6847 10066 6873
rect 10038 6370 10066 6847
rect 10206 6482 10234 7183
rect 10206 6449 10234 6454
rect 10262 6986 10290 7630
rect 10486 7625 10514 7630
rect 10878 7602 10906 9199
rect 10878 7569 10906 7574
rect 11270 7657 11298 9983
rect 11550 9225 11578 10066
rect 11886 9674 11914 10374
rect 12054 10010 12082 10486
rect 12950 10401 12978 11103
rect 12950 10375 12951 10401
rect 12977 10375 12978 10401
rect 12950 10345 12978 10375
rect 12950 10319 12951 10345
rect 12977 10319 12978 10345
rect 11886 9641 11914 9646
rect 11942 9982 12082 10010
rect 12446 10065 12474 10071
rect 12446 10039 12447 10065
rect 12473 10039 12474 10065
rect 12446 10010 12474 10039
rect 11550 9199 11551 9225
rect 11577 9199 11578 9225
rect 11550 8442 11578 9199
rect 11550 8395 11578 8414
rect 11774 9226 11802 9231
rect 11942 9226 11970 9982
rect 12446 9963 12474 9982
rect 12950 10010 12978 10319
rect 12073 9814 12535 9819
rect 12073 9813 12082 9814
rect 12073 9787 12074 9813
rect 12073 9786 12082 9787
rect 12110 9786 12134 9814
rect 12162 9786 12186 9814
rect 12214 9813 12238 9814
rect 12266 9813 12290 9814
rect 12224 9787 12238 9813
rect 12286 9787 12290 9813
rect 12214 9786 12238 9787
rect 12266 9786 12290 9787
rect 12318 9813 12342 9814
rect 12370 9813 12394 9814
rect 12318 9787 12322 9813
rect 12370 9787 12384 9813
rect 12318 9786 12342 9787
rect 12370 9786 12394 9787
rect 12422 9786 12446 9814
rect 12474 9786 12498 9814
rect 12526 9813 12535 9814
rect 12534 9787 12535 9813
rect 12526 9786 12535 9787
rect 12073 9781 12535 9786
rect 12054 9674 12082 9679
rect 12054 9617 12082 9646
rect 12054 9591 12055 9617
rect 12081 9591 12082 9617
rect 12054 9585 12082 9591
rect 12950 9617 12978 9982
rect 12950 9591 12951 9617
rect 12977 9591 12978 9617
rect 12950 9562 12978 9591
rect 12950 9515 12978 9534
rect 13510 10401 13538 11158
rect 13510 10375 13511 10401
rect 13537 10375 13538 10401
rect 13510 9674 13538 10375
rect 13510 9617 13538 9646
rect 13510 9591 13511 9617
rect 13537 9591 13538 9617
rect 11774 9225 11970 9226
rect 11774 9199 11775 9225
rect 11801 9199 11943 9225
rect 11969 9199 11970 9225
rect 11774 9198 11970 9199
rect 11774 8442 11802 9198
rect 11942 9193 11970 9198
rect 12073 9030 12535 9035
rect 12073 9029 12082 9030
rect 12073 9003 12074 9029
rect 12073 9002 12082 9003
rect 12110 9002 12134 9030
rect 12162 9002 12186 9030
rect 12214 9029 12238 9030
rect 12266 9029 12290 9030
rect 12224 9003 12238 9029
rect 12286 9003 12290 9029
rect 12214 9002 12238 9003
rect 12266 9002 12290 9003
rect 12318 9029 12342 9030
rect 12370 9029 12394 9030
rect 12318 9003 12322 9029
rect 12370 9003 12384 9029
rect 12318 9002 12342 9003
rect 12370 9002 12394 9003
rect 12422 9002 12446 9030
rect 12474 9002 12498 9030
rect 12526 9029 12535 9030
rect 12534 9003 12535 9029
rect 12526 9002 12535 9003
rect 12073 8997 12535 9002
rect 11998 8833 12026 8839
rect 11998 8807 11999 8833
rect 12025 8807 12026 8833
rect 11942 8442 11970 8447
rect 11774 8441 11970 8442
rect 11774 8415 11775 8441
rect 11801 8415 11943 8441
rect 11969 8415 11970 8441
rect 11774 8414 11970 8415
rect 11270 7631 11271 7657
rect 11297 7631 11298 7657
rect 11270 7574 11298 7631
rect 11774 7657 11802 8414
rect 11942 8386 11970 8414
rect 11942 8353 11970 8358
rect 11998 8442 12026 8807
rect 11998 8050 12026 8414
rect 12222 8834 12250 8839
rect 12446 8834 12474 8839
rect 12222 8833 12474 8834
rect 12222 8807 12223 8833
rect 12249 8807 12447 8833
rect 12473 8807 12474 8833
rect 12222 8806 12474 8807
rect 12222 8386 12250 8806
rect 12446 8801 12474 8806
rect 13510 8834 13538 9591
rect 13510 8787 13538 8806
rect 14070 10793 14098 11551
rect 14406 11969 14434 11975
rect 14406 11943 14407 11969
rect 14433 11943 14434 11969
rect 14406 11913 14434 11943
rect 14406 11887 14407 11913
rect 14433 11887 14434 11913
rect 14406 11185 14434 11887
rect 14573 11774 15035 11779
rect 14573 11773 14582 11774
rect 14573 11747 14574 11773
rect 14573 11746 14582 11747
rect 14610 11746 14634 11774
rect 14662 11746 14686 11774
rect 14714 11773 14738 11774
rect 14766 11773 14790 11774
rect 14724 11747 14738 11773
rect 14786 11747 14790 11773
rect 14714 11746 14738 11747
rect 14766 11746 14790 11747
rect 14818 11773 14842 11774
rect 14870 11773 14894 11774
rect 14818 11747 14822 11773
rect 14870 11747 14884 11773
rect 14818 11746 14842 11747
rect 14870 11746 14894 11747
rect 14922 11746 14946 11774
rect 14974 11746 14998 11774
rect 15026 11773 15035 11774
rect 15034 11747 15035 11773
rect 15026 11746 15035 11747
rect 14573 11741 15035 11746
rect 14966 11633 14994 11639
rect 14966 11607 14967 11633
rect 14993 11607 14994 11633
rect 14966 11578 14994 11607
rect 15078 11634 15106 12334
rect 15526 12361 15890 12362
rect 15526 12335 15527 12361
rect 15553 12335 15890 12361
rect 15526 12334 15890 12335
rect 15526 11774 15554 12334
rect 15862 11970 15890 12334
rect 16422 12362 16450 12390
rect 16646 12362 16674 12671
rect 16422 12361 16674 12362
rect 16422 12335 16423 12361
rect 16449 12335 16674 12361
rect 16422 12334 16674 12335
rect 16422 12329 16450 12334
rect 16646 11970 16674 12334
rect 16758 11970 16786 11975
rect 16646 11969 16786 11970
rect 16646 11943 16759 11969
rect 16785 11943 16786 11969
rect 16646 11942 16786 11943
rect 15862 11923 15890 11942
rect 15078 11578 15106 11606
rect 14966 11577 15106 11578
rect 14966 11551 14967 11577
rect 14993 11551 15106 11577
rect 14966 11550 15106 11551
rect 15470 11746 15554 11774
rect 16758 11913 16786 11942
rect 16758 11887 16759 11913
rect 16785 11887 16786 11913
rect 15470 11577 15498 11746
rect 15470 11551 15471 11577
rect 15497 11551 15498 11577
rect 14966 11545 14994 11550
rect 14406 11159 14407 11185
rect 14433 11159 14434 11185
rect 14406 11129 14434 11159
rect 14406 11103 14407 11129
rect 14433 11103 14434 11129
rect 14070 10767 14071 10793
rect 14097 10767 14098 10793
rect 14070 10009 14098 10767
rect 14350 10794 14378 10799
rect 14406 10794 14434 11103
rect 14573 10990 15035 10995
rect 14573 10989 14582 10990
rect 14573 10963 14574 10989
rect 14573 10962 14582 10963
rect 14610 10962 14634 10990
rect 14662 10962 14686 10990
rect 14714 10989 14738 10990
rect 14766 10989 14790 10990
rect 14724 10963 14738 10989
rect 14786 10963 14790 10989
rect 14714 10962 14738 10963
rect 14766 10962 14790 10963
rect 14818 10989 14842 10990
rect 14870 10989 14894 10990
rect 14818 10963 14822 10989
rect 14870 10963 14884 10989
rect 14818 10962 14842 10963
rect 14870 10962 14894 10963
rect 14922 10962 14946 10990
rect 14974 10962 14998 10990
rect 15026 10989 15035 10990
rect 15034 10963 15035 10989
rect 15026 10962 15035 10963
rect 14573 10957 15035 10962
rect 14462 10794 14490 10799
rect 14350 10793 14490 10794
rect 14350 10767 14351 10793
rect 14377 10767 14463 10793
rect 14489 10767 14490 10793
rect 14350 10766 14490 10767
rect 14350 10761 14378 10766
rect 14406 10401 14434 10766
rect 14462 10761 14490 10766
rect 15470 10793 15498 11551
rect 16198 11634 16226 11639
rect 16198 11577 16226 11606
rect 16758 11634 16786 11887
rect 16758 11601 16786 11606
rect 16198 11551 16199 11577
rect 16225 11551 16226 11577
rect 15470 10767 15471 10793
rect 15497 10767 15498 10793
rect 14406 10375 14407 10401
rect 14433 10375 14434 10401
rect 14406 10345 14434 10375
rect 14406 10319 14407 10345
rect 14433 10319 14434 10345
rect 14070 9983 14071 10009
rect 14097 9983 14098 10009
rect 14070 9225 14098 9983
rect 14350 10010 14378 10015
rect 14406 10010 14434 10319
rect 14573 10206 15035 10211
rect 14573 10205 14582 10206
rect 14573 10179 14574 10205
rect 14573 10178 14582 10179
rect 14610 10178 14634 10206
rect 14662 10178 14686 10206
rect 14714 10205 14738 10206
rect 14766 10205 14790 10206
rect 14724 10179 14738 10205
rect 14786 10179 14790 10205
rect 14714 10178 14738 10179
rect 14766 10178 14790 10179
rect 14818 10205 14842 10206
rect 14870 10205 14894 10206
rect 14818 10179 14822 10205
rect 14870 10179 14884 10205
rect 14818 10178 14842 10179
rect 14870 10178 14894 10179
rect 14922 10178 14946 10206
rect 14974 10178 14998 10206
rect 15026 10205 15035 10206
rect 15034 10179 15035 10205
rect 15026 10178 15035 10179
rect 14573 10173 15035 10178
rect 14462 10010 14490 10015
rect 14350 10009 14490 10010
rect 14350 9983 14351 10009
rect 14377 9983 14463 10009
rect 14489 9983 14490 10009
rect 14350 9982 14490 9983
rect 14350 9977 14378 9982
rect 14406 9618 14434 9623
rect 14462 9618 14490 9982
rect 14406 9617 14490 9618
rect 14406 9591 14407 9617
rect 14433 9591 14490 9617
rect 14406 9590 14490 9591
rect 15470 10010 15498 10767
rect 15694 11185 15722 11191
rect 15694 11159 15695 11185
rect 15721 11159 15722 11185
rect 15694 10401 15722 11159
rect 16198 11186 16226 11551
rect 16310 11186 16338 11191
rect 16198 11185 16338 11186
rect 16198 11159 16199 11185
rect 16225 11159 16311 11185
rect 16337 11159 16338 11185
rect 16198 11158 16338 11159
rect 16198 10849 16226 11158
rect 16310 11153 16338 11158
rect 16198 10823 16199 10849
rect 16225 10823 16226 10849
rect 15694 10375 15695 10401
rect 15721 10375 15722 10401
rect 15694 10010 15722 10375
rect 16142 10794 16170 10799
rect 16198 10794 16226 10823
rect 16142 10793 16226 10794
rect 16142 10767 16143 10793
rect 16169 10767 16226 10793
rect 16142 10766 16226 10767
rect 16142 10402 16170 10766
rect 16366 10402 16394 10407
rect 16142 10401 16366 10402
rect 16142 10375 16143 10401
rect 16169 10375 16366 10401
rect 16142 10374 16366 10375
rect 15470 10009 15722 10010
rect 15470 9983 15471 10009
rect 15497 9983 15722 10009
rect 15470 9982 15722 9983
rect 15806 10010 15834 10015
rect 15918 10010 15946 10015
rect 15806 10009 15946 10010
rect 15806 9983 15807 10009
rect 15833 9983 15919 10009
rect 15945 9983 15946 10009
rect 15806 9982 15946 9983
rect 15470 9618 15498 9982
rect 15806 9977 15834 9982
rect 15526 9618 15554 9623
rect 15470 9617 15554 9618
rect 15470 9591 15527 9617
rect 15553 9591 15554 9617
rect 15470 9590 15554 9591
rect 14406 9562 14434 9590
rect 14070 9199 14071 9225
rect 14097 9199 14098 9225
rect 14070 8834 14098 9199
rect 14350 9226 14378 9231
rect 14406 9226 14434 9534
rect 14573 9422 15035 9427
rect 14573 9421 14582 9422
rect 14573 9395 14574 9421
rect 14573 9394 14582 9395
rect 14610 9394 14634 9422
rect 14662 9394 14686 9422
rect 14714 9421 14738 9422
rect 14766 9421 14790 9422
rect 14724 9395 14738 9421
rect 14786 9395 14790 9421
rect 14714 9394 14738 9395
rect 14766 9394 14790 9395
rect 14818 9421 14842 9422
rect 14870 9421 14894 9422
rect 14818 9395 14822 9421
rect 14870 9395 14884 9421
rect 14818 9394 14842 9395
rect 14870 9394 14894 9395
rect 14922 9394 14946 9422
rect 14974 9394 14998 9422
rect 15026 9421 15035 9422
rect 15034 9395 15035 9421
rect 15026 9394 15035 9395
rect 14573 9389 15035 9394
rect 14462 9226 14490 9231
rect 14350 9225 14490 9226
rect 14350 9199 14351 9225
rect 14377 9199 14463 9225
rect 14489 9199 14490 9225
rect 14350 9198 14490 9199
rect 14350 9193 14378 9198
rect 12222 8353 12250 8358
rect 14070 8441 14098 8806
rect 14070 8415 14071 8441
rect 14097 8415 14098 8441
rect 12073 8246 12535 8251
rect 12073 8245 12082 8246
rect 12073 8219 12074 8245
rect 12073 8218 12082 8219
rect 12110 8218 12134 8246
rect 12162 8218 12186 8246
rect 12214 8245 12238 8246
rect 12266 8245 12290 8246
rect 12224 8219 12238 8245
rect 12286 8219 12290 8245
rect 12214 8218 12238 8219
rect 12266 8218 12290 8219
rect 12318 8245 12342 8246
rect 12370 8245 12394 8246
rect 12318 8219 12322 8245
rect 12370 8219 12384 8245
rect 12318 8218 12342 8219
rect 12370 8218 12394 8219
rect 12422 8218 12446 8246
rect 12474 8218 12498 8246
rect 12526 8245 12535 8246
rect 12534 8219 12535 8245
rect 12526 8218 12535 8219
rect 12073 8213 12535 8218
rect 12054 8050 12082 8055
rect 11998 8022 12054 8050
rect 12054 8003 12082 8022
rect 12222 8050 12250 8055
rect 12446 8050 12474 8055
rect 12222 8049 12474 8050
rect 12222 8023 12223 8049
rect 12249 8023 12447 8049
rect 12473 8023 12474 8049
rect 12222 8022 12474 8023
rect 11774 7631 11775 7657
rect 11801 7631 11802 7657
rect 11774 7602 11802 7631
rect 11270 7546 11578 7574
rect 11774 7569 11802 7574
rect 11942 7657 11970 7663
rect 11942 7631 11943 7657
rect 11969 7631 11970 7657
rect 11942 7602 11970 7631
rect 11942 7569 11970 7574
rect 12222 7602 12250 8022
rect 12446 7994 12474 8022
rect 12446 7961 12474 7966
rect 13398 8050 13426 8055
rect 12222 7569 12250 7574
rect 10262 6958 10570 6986
rect 10262 6873 10290 6958
rect 10262 6847 10263 6873
rect 10289 6847 10290 6873
rect 10038 6342 10122 6370
rect 9573 6286 10035 6291
rect 9573 6285 9582 6286
rect 9573 6259 9574 6285
rect 9573 6258 9582 6259
rect 9610 6258 9634 6286
rect 9662 6258 9686 6286
rect 9714 6285 9738 6286
rect 9766 6285 9790 6286
rect 9724 6259 9738 6285
rect 9786 6259 9790 6285
rect 9714 6258 9738 6259
rect 9766 6258 9790 6259
rect 9818 6285 9842 6286
rect 9870 6285 9894 6286
rect 9818 6259 9822 6285
rect 9870 6259 9884 6285
rect 9818 6258 9842 6259
rect 9870 6258 9894 6259
rect 9922 6258 9946 6286
rect 9974 6258 9998 6286
rect 10026 6285 10035 6286
rect 10034 6259 10035 6285
rect 10026 6258 10035 6259
rect 9573 6253 10035 6258
rect 10094 6202 10122 6342
rect 10038 6174 10122 6202
rect 10038 6089 10066 6174
rect 10038 6063 10039 6089
rect 10065 6063 10066 6089
rect 10038 5586 10066 6063
rect 10262 5697 10290 6847
rect 10542 6873 10570 6958
rect 10542 6847 10543 6873
rect 10569 6847 10570 6873
rect 10542 6841 10570 6847
rect 11550 6873 11578 7546
rect 12073 7462 12535 7467
rect 12073 7461 12082 7462
rect 12073 7435 12074 7461
rect 12073 7434 12082 7435
rect 12110 7434 12134 7462
rect 12162 7434 12186 7462
rect 12214 7461 12238 7462
rect 12266 7461 12290 7462
rect 12224 7435 12238 7461
rect 12286 7435 12290 7461
rect 12214 7434 12238 7435
rect 12266 7434 12290 7435
rect 12318 7461 12342 7462
rect 12370 7461 12394 7462
rect 12318 7435 12322 7461
rect 12370 7435 12384 7461
rect 12318 7434 12342 7435
rect 12370 7434 12394 7435
rect 12422 7434 12446 7462
rect 12474 7434 12498 7462
rect 12526 7461 12535 7462
rect 12534 7435 12535 7461
rect 12526 7434 12535 7435
rect 12073 7429 12535 7434
rect 11830 7265 11858 7271
rect 11830 7239 11831 7265
rect 11857 7239 11858 7265
rect 11550 6847 11551 6873
rect 11577 6847 11578 6873
rect 10262 5671 10263 5697
rect 10289 5671 10290 5697
rect 10262 5641 10290 5671
rect 10262 5615 10263 5641
rect 10289 5615 10290 5641
rect 10038 5558 10122 5586
rect 9573 5502 10035 5507
rect 9573 5501 9582 5502
rect 9573 5475 9574 5501
rect 9573 5474 9582 5475
rect 9610 5474 9634 5502
rect 9662 5474 9686 5502
rect 9714 5501 9738 5502
rect 9766 5501 9790 5502
rect 9724 5475 9738 5501
rect 9786 5475 9790 5501
rect 9714 5474 9738 5475
rect 9766 5474 9790 5475
rect 9818 5501 9842 5502
rect 9870 5501 9894 5502
rect 9818 5475 9822 5501
rect 9870 5475 9884 5501
rect 9818 5474 9842 5475
rect 9870 5474 9894 5475
rect 9922 5474 9946 5502
rect 9974 5474 9998 5502
rect 10026 5501 10035 5502
rect 10034 5475 10035 5501
rect 10026 5474 10035 5475
rect 9573 5469 10035 5474
rect 10094 5418 10122 5558
rect 10038 5390 10122 5418
rect 10038 5305 10066 5390
rect 10038 5279 10039 5305
rect 10065 5279 10066 5305
rect 10038 4802 10066 5279
rect 10038 4774 10122 4802
rect 9573 4718 10035 4723
rect 9573 4717 9582 4718
rect 9573 4691 9574 4717
rect 9573 4690 9582 4691
rect 9610 4690 9634 4718
rect 9662 4690 9686 4718
rect 9714 4717 9738 4718
rect 9766 4717 9790 4718
rect 9724 4691 9738 4717
rect 9786 4691 9790 4717
rect 9714 4690 9738 4691
rect 9766 4690 9790 4691
rect 9818 4717 9842 4718
rect 9870 4717 9894 4718
rect 9818 4691 9822 4717
rect 9870 4691 9884 4717
rect 9818 4690 9842 4691
rect 9870 4690 9894 4691
rect 9922 4690 9946 4718
rect 9974 4690 9998 4718
rect 10026 4717 10035 4718
rect 10034 4691 10035 4717
rect 10026 4690 10035 4691
rect 9573 4685 10035 4690
rect 10094 4634 10122 4774
rect 10038 4606 10122 4634
rect 10038 4521 10066 4606
rect 10038 4495 10039 4521
rect 10065 4495 10066 4521
rect 9534 4130 9562 4135
rect 9534 4083 9562 4102
rect 10038 4130 10066 4495
rect 10038 4018 10066 4102
rect 10038 3990 10122 4018
rect 9573 3934 10035 3939
rect 9573 3933 9582 3934
rect 9573 3907 9574 3933
rect 9573 3906 9582 3907
rect 9610 3906 9634 3934
rect 9662 3906 9686 3934
rect 9714 3933 9738 3934
rect 9766 3933 9790 3934
rect 9724 3907 9738 3933
rect 9786 3907 9790 3933
rect 9714 3906 9738 3907
rect 9766 3906 9790 3907
rect 9818 3933 9842 3934
rect 9870 3933 9894 3934
rect 9818 3907 9822 3933
rect 9870 3907 9884 3933
rect 9818 3906 9842 3907
rect 9870 3906 9894 3907
rect 9922 3906 9946 3934
rect 9974 3906 9998 3934
rect 10026 3933 10035 3934
rect 10034 3907 10035 3933
rect 10026 3906 10035 3907
rect 9573 3901 10035 3906
rect 10094 3850 10122 3990
rect 10038 3822 10122 3850
rect 10038 3737 10066 3822
rect 10038 3711 10039 3737
rect 10065 3711 10066 3737
rect 9534 3402 9562 3407
rect 9534 3345 9562 3374
rect 9534 3319 9535 3345
rect 9561 3319 9562 3345
rect 9534 3313 9562 3319
rect 10038 3402 10066 3711
rect 10038 3234 10066 3374
rect 10262 3738 10290 5615
rect 10038 3206 10122 3234
rect 9573 3150 10035 3155
rect 9573 3149 9582 3150
rect 9573 3123 9574 3149
rect 9573 3122 9582 3123
rect 9610 3122 9634 3150
rect 9662 3122 9686 3150
rect 9714 3149 9738 3150
rect 9766 3149 9790 3150
rect 9724 3123 9738 3149
rect 9786 3123 9790 3149
rect 9714 3122 9738 3123
rect 9766 3122 9790 3123
rect 9818 3149 9842 3150
rect 9870 3149 9894 3150
rect 9818 3123 9822 3149
rect 9870 3123 9884 3149
rect 9818 3122 9842 3123
rect 9870 3122 9894 3123
rect 9922 3122 9946 3150
rect 9974 3122 9998 3150
rect 10026 3149 10035 3150
rect 10034 3123 10035 3149
rect 10026 3122 10035 3123
rect 9573 3117 10035 3122
rect 10094 3066 10122 3206
rect 10038 3038 10122 3066
rect 10038 2953 10066 3038
rect 10038 2927 10039 2953
rect 10065 2927 10066 2953
rect 9534 2562 9562 2567
rect 10038 2562 10066 2927
rect 9534 2561 10066 2562
rect 9534 2535 9535 2561
rect 9561 2535 10066 2561
rect 9534 2534 10066 2535
rect 9534 2529 9562 2534
rect 10038 2450 10066 2534
rect 10262 2561 10290 3710
rect 10318 6482 10346 6487
rect 10318 6425 10346 6454
rect 10318 6399 10319 6425
rect 10345 6399 10346 6425
rect 10318 6090 10346 6399
rect 10486 6090 10514 6095
rect 10318 6089 10514 6090
rect 10318 6063 10319 6089
rect 10345 6063 10487 6089
rect 10513 6063 10514 6089
rect 10318 6062 10514 6063
rect 10318 5306 10346 6062
rect 10486 6057 10514 6062
rect 11550 6089 11578 6847
rect 11774 6874 11802 6879
rect 11774 6827 11802 6846
rect 11550 6063 11551 6089
rect 11577 6063 11578 6089
rect 10486 5306 10514 5311
rect 10318 5305 10514 5306
rect 10318 5279 10319 5305
rect 10345 5279 10487 5305
rect 10513 5279 10514 5305
rect 10318 5278 10514 5279
rect 10318 4913 10346 5278
rect 10486 5273 10514 5278
rect 11550 5305 11578 6063
rect 11830 6481 11858 7239
rect 12222 7266 12250 7271
rect 12446 7266 12474 7271
rect 12222 7265 12474 7266
rect 12222 7239 12223 7265
rect 12249 7239 12447 7265
rect 12473 7239 12474 7265
rect 12222 7238 12474 7239
rect 13398 7266 13426 8022
rect 14070 7658 14098 8415
rect 14406 8833 14434 9198
rect 14462 9193 14490 9198
rect 15246 9225 15274 9231
rect 15246 9199 15247 9225
rect 15273 9199 15274 9225
rect 14406 8807 14407 8833
rect 14433 8807 14434 8833
rect 14406 8777 14434 8807
rect 14406 8751 14407 8777
rect 14433 8751 14434 8777
rect 14406 8442 14434 8751
rect 15246 8834 15274 9199
rect 15470 8834 15498 9590
rect 15526 9585 15554 9590
rect 15918 9618 15946 9982
rect 15974 9618 16002 9623
rect 16142 9618 16170 10374
rect 16366 10336 16394 10374
rect 16198 9618 16226 9623
rect 15918 9617 16226 9618
rect 15918 9591 15975 9617
rect 16001 9591 16199 9617
rect 16225 9591 16226 9617
rect 15918 9590 16226 9591
rect 15806 9226 15834 9231
rect 15918 9226 15946 9590
rect 15974 9585 16002 9590
rect 16198 9585 16226 9590
rect 15806 9225 15946 9226
rect 15806 9199 15807 9225
rect 15833 9199 15919 9225
rect 15945 9199 15946 9225
rect 15806 9198 15946 9199
rect 15806 9193 15834 9198
rect 15246 8833 15498 8834
rect 15246 8807 15471 8833
rect 15497 8807 15498 8833
rect 15246 8806 15498 8807
rect 14573 8638 15035 8643
rect 14573 8637 14582 8638
rect 14573 8611 14574 8637
rect 14573 8610 14582 8611
rect 14610 8610 14634 8638
rect 14662 8610 14686 8638
rect 14714 8637 14738 8638
rect 14766 8637 14790 8638
rect 14724 8611 14738 8637
rect 14786 8611 14790 8637
rect 14714 8610 14738 8611
rect 14766 8610 14790 8611
rect 14818 8637 14842 8638
rect 14870 8637 14894 8638
rect 14818 8611 14822 8637
rect 14870 8611 14884 8637
rect 14818 8610 14842 8611
rect 14870 8610 14894 8611
rect 14922 8610 14946 8638
rect 14974 8610 14998 8638
rect 15026 8637 15035 8638
rect 15034 8611 15035 8637
rect 15026 8610 15035 8611
rect 14573 8605 15035 8610
rect 14406 8409 14434 8414
rect 14966 8497 14994 8503
rect 14966 8471 14967 8497
rect 14993 8471 14994 8497
rect 14966 8442 14994 8471
rect 14966 8395 14994 8414
rect 15246 8441 15274 8806
rect 15470 8801 15498 8806
rect 15526 9170 15554 9175
rect 15246 8415 15247 8441
rect 15273 8415 15274 8441
rect 14182 8049 14210 8055
rect 14182 8023 14183 8049
rect 14209 8023 14210 8049
rect 14182 7994 14210 8023
rect 14182 7928 14210 7966
rect 15246 8050 15274 8415
rect 15302 8050 15330 8055
rect 15246 8049 15330 8050
rect 15246 8023 15303 8049
rect 15329 8023 15330 8049
rect 15246 8022 15330 8023
rect 14573 7854 15035 7859
rect 14573 7853 14582 7854
rect 14573 7827 14574 7853
rect 14573 7826 14582 7827
rect 14610 7826 14634 7854
rect 14662 7826 14686 7854
rect 14714 7853 14738 7854
rect 14766 7853 14790 7854
rect 14724 7827 14738 7853
rect 14786 7827 14790 7853
rect 14714 7826 14738 7827
rect 14766 7826 14790 7827
rect 14818 7853 14842 7854
rect 14870 7853 14894 7854
rect 14818 7827 14822 7853
rect 14870 7827 14884 7853
rect 14818 7826 14842 7827
rect 14870 7826 14894 7827
rect 14922 7826 14946 7854
rect 14974 7826 14998 7854
rect 15026 7853 15035 7854
rect 15034 7827 15035 7853
rect 15026 7826 15035 7827
rect 14573 7821 15035 7826
rect 14070 7611 14098 7630
rect 14966 7713 14994 7719
rect 14966 7687 14967 7713
rect 14993 7687 14994 7713
rect 14966 7658 14994 7687
rect 15190 7658 15218 7663
rect 15246 7658 15274 8022
rect 15302 8017 15330 8022
rect 14966 7657 15106 7658
rect 14966 7631 14967 7657
rect 14993 7631 15106 7657
rect 14966 7630 15106 7631
rect 14966 7625 14994 7630
rect 13510 7266 13538 7271
rect 13398 7265 13762 7266
rect 13398 7239 13511 7265
rect 13537 7239 13762 7265
rect 13398 7238 13762 7239
rect 11830 6455 11831 6481
rect 11857 6455 11858 6481
rect 11830 5894 11858 6455
rect 11998 6874 12026 6879
rect 11998 6482 12026 6846
rect 12222 6874 12250 7238
rect 12446 7233 12474 7238
rect 13510 7233 13538 7238
rect 12222 6841 12250 6846
rect 13734 6873 13762 7238
rect 14406 7265 14434 7271
rect 14406 7239 14407 7265
rect 14433 7239 14434 7265
rect 14406 7209 14434 7239
rect 14406 7183 14407 7209
rect 14433 7183 14434 7209
rect 14294 6874 14322 6879
rect 13734 6847 13735 6873
rect 13761 6847 13762 6873
rect 13734 6841 13762 6847
rect 14238 6846 14294 6874
rect 12073 6678 12535 6683
rect 12073 6677 12082 6678
rect 12073 6651 12074 6677
rect 12073 6650 12082 6651
rect 12110 6650 12134 6678
rect 12162 6650 12186 6678
rect 12214 6677 12238 6678
rect 12266 6677 12290 6678
rect 12224 6651 12238 6677
rect 12286 6651 12290 6677
rect 12214 6650 12238 6651
rect 12266 6650 12290 6651
rect 12318 6677 12342 6678
rect 12370 6677 12394 6678
rect 12318 6651 12322 6677
rect 12370 6651 12384 6677
rect 12318 6650 12342 6651
rect 12370 6650 12394 6651
rect 12422 6650 12446 6678
rect 12474 6650 12498 6678
rect 12526 6677 12535 6678
rect 12534 6651 12535 6677
rect 12526 6650 12535 6651
rect 12073 6645 12535 6650
rect 11998 6449 12026 6454
rect 12334 6482 12362 6487
rect 12446 6482 12474 6487
rect 12362 6481 12474 6482
rect 12362 6455 12447 6481
rect 12473 6455 12474 6481
rect 12362 6454 12474 6455
rect 12334 6416 12362 6454
rect 12446 6145 12474 6454
rect 12446 6119 12447 6145
rect 12473 6119 12474 6145
rect 12446 6090 12474 6119
rect 13510 6481 13538 6487
rect 13510 6455 13511 6481
rect 13537 6455 13538 6481
rect 12446 6043 12474 6062
rect 12950 6090 12978 6095
rect 12073 5894 12535 5899
rect 11830 5866 12026 5894
rect 11550 5279 11551 5305
rect 11577 5279 11578 5305
rect 10318 4887 10319 4913
rect 10345 4887 10346 4913
rect 10318 4857 10346 4887
rect 10318 4831 10319 4857
rect 10345 4831 10346 4857
rect 10318 4522 10346 4831
rect 10486 4522 10514 4527
rect 10318 4521 10514 4522
rect 10318 4495 10319 4521
rect 10345 4495 10487 4521
rect 10513 4495 10514 4521
rect 10318 4494 10514 4495
rect 10318 4129 10346 4494
rect 10486 4489 10514 4494
rect 11550 4521 11578 5279
rect 11550 4495 11551 4521
rect 11577 4495 11578 4521
rect 10318 4103 10319 4129
rect 10345 4103 10346 4129
rect 10318 4073 10346 4103
rect 10318 4047 10319 4073
rect 10345 4047 10346 4073
rect 10318 3346 10346 4047
rect 10486 3738 10514 3743
rect 10486 3691 10514 3710
rect 11550 3737 11578 4495
rect 11550 3711 11551 3737
rect 11577 3711 11578 3737
rect 10430 3346 10458 3351
rect 10346 3345 10458 3346
rect 10346 3319 10431 3345
rect 10457 3319 10458 3345
rect 10346 3318 10458 3319
rect 10318 3280 10346 3318
rect 10430 3289 10458 3318
rect 10430 3263 10431 3289
rect 10457 3263 10458 3289
rect 10430 3010 10458 3263
rect 10766 3010 10794 3015
rect 10430 3009 10794 3010
rect 10430 2983 10767 3009
rect 10793 2983 10794 3009
rect 10430 2982 10794 2983
rect 10262 2535 10263 2561
rect 10289 2535 10290 2561
rect 10262 2506 10290 2535
rect 10038 2422 10122 2450
rect 9573 2366 10035 2371
rect 9573 2365 9582 2366
rect 9573 2339 9574 2365
rect 9573 2338 9582 2339
rect 9610 2338 9634 2366
rect 9662 2338 9686 2366
rect 9714 2365 9738 2366
rect 9766 2365 9790 2366
rect 9724 2339 9738 2365
rect 9786 2339 9790 2365
rect 9714 2338 9738 2339
rect 9766 2338 9790 2339
rect 9818 2365 9842 2366
rect 9870 2365 9894 2366
rect 9818 2339 9822 2365
rect 9870 2339 9884 2365
rect 9818 2338 9842 2339
rect 9870 2338 9894 2339
rect 9922 2338 9946 2366
rect 9974 2338 9998 2366
rect 10026 2365 10035 2366
rect 10034 2339 10035 2365
rect 10026 2338 10035 2339
rect 9573 2333 10035 2338
rect 10094 2282 10122 2422
rect 10038 2254 10122 2282
rect 10038 2170 10066 2254
rect 10038 2123 10066 2142
rect 10262 1777 10290 2478
rect 10766 2953 10794 2982
rect 10766 2927 10767 2953
rect 10793 2927 10794 2953
rect 10766 2225 10794 2927
rect 10766 2199 10767 2225
rect 10793 2199 10794 2225
rect 10766 2169 10794 2199
rect 11550 2953 11578 3711
rect 11998 5697 12026 5866
rect 12073 5893 12082 5894
rect 12073 5867 12074 5893
rect 12073 5866 12082 5867
rect 12110 5866 12134 5894
rect 12162 5866 12186 5894
rect 12214 5893 12238 5894
rect 12266 5893 12290 5894
rect 12224 5867 12238 5893
rect 12286 5867 12290 5893
rect 12214 5866 12238 5867
rect 12266 5866 12290 5867
rect 12318 5893 12342 5894
rect 12370 5893 12394 5894
rect 12318 5867 12322 5893
rect 12370 5867 12384 5893
rect 12318 5866 12342 5867
rect 12370 5866 12394 5867
rect 12422 5866 12446 5894
rect 12474 5866 12498 5894
rect 12526 5893 12535 5894
rect 12534 5867 12535 5893
rect 12526 5866 12535 5867
rect 12073 5861 12535 5866
rect 11998 5671 11999 5697
rect 12025 5671 12026 5697
rect 11998 4913 12026 5671
rect 12950 5697 12978 6062
rect 12950 5671 12951 5697
rect 12977 5671 12978 5697
rect 12950 5641 12978 5671
rect 12950 5615 12951 5641
rect 12977 5615 12978 5641
rect 12446 5361 12474 5367
rect 12446 5335 12447 5361
rect 12473 5335 12474 5361
rect 12446 5306 12474 5335
rect 12446 5259 12474 5278
rect 12950 5306 12978 5615
rect 12073 5110 12535 5115
rect 12073 5109 12082 5110
rect 12073 5083 12074 5109
rect 12073 5082 12082 5083
rect 12110 5082 12134 5110
rect 12162 5082 12186 5110
rect 12214 5109 12238 5110
rect 12266 5109 12290 5110
rect 12224 5083 12238 5109
rect 12286 5083 12290 5109
rect 12214 5082 12238 5083
rect 12266 5082 12290 5083
rect 12318 5109 12342 5110
rect 12370 5109 12394 5110
rect 12318 5083 12322 5109
rect 12370 5083 12384 5109
rect 12318 5082 12342 5083
rect 12370 5082 12394 5083
rect 12422 5082 12446 5110
rect 12474 5082 12498 5110
rect 12526 5109 12535 5110
rect 12534 5083 12535 5109
rect 12526 5082 12535 5083
rect 12073 5077 12535 5082
rect 11998 4887 11999 4913
rect 12025 4887 12026 4913
rect 11998 4129 12026 4887
rect 12950 4913 12978 5278
rect 12950 4887 12951 4913
rect 12977 4887 12978 4913
rect 12950 4858 12978 4887
rect 12670 4634 12698 4639
rect 12446 4577 12474 4583
rect 12446 4551 12447 4577
rect 12473 4551 12474 4577
rect 12446 4522 12474 4551
rect 12446 4456 12474 4494
rect 12073 4326 12535 4331
rect 12073 4325 12082 4326
rect 12073 4299 12074 4325
rect 12073 4298 12082 4299
rect 12110 4298 12134 4326
rect 12162 4298 12186 4326
rect 12214 4325 12238 4326
rect 12266 4325 12290 4326
rect 12224 4299 12238 4325
rect 12286 4299 12290 4325
rect 12214 4298 12238 4299
rect 12266 4298 12290 4299
rect 12318 4325 12342 4326
rect 12370 4325 12394 4326
rect 12318 4299 12322 4325
rect 12370 4299 12384 4325
rect 12318 4298 12342 4299
rect 12370 4298 12394 4299
rect 12422 4298 12446 4326
rect 12474 4298 12498 4326
rect 12526 4325 12535 4326
rect 12534 4299 12535 4325
rect 12526 4298 12535 4299
rect 12073 4293 12535 4298
rect 11998 4103 11999 4129
rect 12025 4103 12026 4129
rect 11998 3402 12026 4103
rect 12446 3793 12474 3799
rect 12446 3767 12447 3793
rect 12473 3767 12474 3793
rect 12446 3738 12474 3767
rect 12446 3691 12474 3710
rect 12073 3542 12535 3547
rect 12073 3541 12082 3542
rect 12073 3515 12074 3541
rect 12073 3514 12082 3515
rect 12110 3514 12134 3542
rect 12162 3514 12186 3542
rect 12214 3541 12238 3542
rect 12266 3541 12290 3542
rect 12224 3515 12238 3541
rect 12286 3515 12290 3541
rect 12214 3514 12238 3515
rect 12266 3514 12290 3515
rect 12318 3541 12342 3542
rect 12370 3541 12394 3542
rect 12318 3515 12322 3541
rect 12370 3515 12384 3541
rect 12318 3514 12342 3515
rect 12370 3514 12394 3515
rect 12422 3514 12446 3542
rect 12474 3514 12498 3542
rect 12526 3541 12535 3542
rect 12534 3515 12535 3541
rect 12526 3514 12535 3515
rect 12073 3509 12535 3514
rect 12054 3402 12082 3407
rect 11550 2927 11551 2953
rect 11577 2927 11578 2953
rect 11550 2562 11578 2927
rect 11886 3374 12054 3402
rect 11886 2562 11914 3374
rect 12054 3345 12082 3374
rect 12054 3319 12055 3345
rect 12081 3319 12082 3345
rect 12054 3313 12082 3319
rect 12446 3010 12474 3015
rect 12446 2953 12474 2982
rect 12446 2927 12447 2953
rect 12473 2927 12474 2953
rect 12446 2921 12474 2927
rect 12073 2758 12535 2763
rect 12073 2757 12082 2758
rect 12073 2731 12074 2757
rect 12073 2730 12082 2731
rect 12110 2730 12134 2758
rect 12162 2730 12186 2758
rect 12214 2757 12238 2758
rect 12266 2757 12290 2758
rect 12224 2731 12238 2757
rect 12286 2731 12290 2757
rect 12214 2730 12238 2731
rect 12266 2730 12290 2731
rect 12318 2757 12342 2758
rect 12370 2757 12394 2758
rect 12318 2731 12322 2757
rect 12370 2731 12384 2757
rect 12318 2730 12342 2731
rect 12370 2730 12394 2731
rect 12422 2730 12446 2758
rect 12474 2730 12498 2758
rect 12526 2757 12535 2758
rect 12534 2731 12535 2757
rect 12526 2730 12535 2731
rect 12073 2725 12535 2730
rect 11550 2561 11914 2562
rect 11550 2535 11887 2561
rect 11913 2535 11914 2561
rect 11550 2534 11914 2535
rect 10766 2143 10767 2169
rect 10793 2143 10794 2169
rect 10766 2137 10794 2143
rect 11214 2170 11242 2175
rect 10262 1751 10263 1777
rect 10289 1751 10290 1777
rect 10262 1721 10290 1751
rect 10262 1695 10263 1721
rect 10289 1695 10290 1721
rect 10262 1689 10290 1695
rect 11214 1694 11242 2142
rect 11550 2169 11578 2534
rect 11886 2529 11914 2534
rect 11550 2143 11551 2169
rect 11577 2143 11578 2169
rect 11382 1778 11410 1783
rect 11550 1778 11578 2143
rect 11382 1777 11578 1778
rect 11382 1751 11383 1777
rect 11409 1751 11578 1777
rect 11382 1750 11578 1751
rect 11998 2226 12026 2231
rect 11998 1777 12026 2198
rect 12446 2226 12474 2231
rect 12446 2169 12474 2198
rect 12446 2143 12447 2169
rect 12473 2143 12474 2169
rect 12446 2137 12474 2143
rect 12073 1974 12535 1979
rect 12073 1973 12082 1974
rect 12073 1947 12074 1973
rect 12073 1946 12082 1947
rect 12110 1946 12134 1974
rect 12162 1946 12186 1974
rect 12214 1973 12238 1974
rect 12266 1973 12290 1974
rect 12224 1947 12238 1973
rect 12286 1947 12290 1973
rect 12214 1946 12238 1947
rect 12266 1946 12290 1947
rect 12318 1973 12342 1974
rect 12370 1973 12394 1974
rect 12318 1947 12322 1973
rect 12370 1947 12384 1973
rect 12318 1946 12342 1947
rect 12370 1946 12394 1947
rect 12422 1946 12446 1974
rect 12474 1946 12498 1974
rect 12526 1973 12535 1974
rect 12534 1947 12535 1973
rect 12526 1946 12535 1947
rect 12073 1941 12535 1946
rect 11998 1751 11999 1777
rect 12025 1751 12026 1777
rect 11382 1694 11410 1750
rect 11998 1722 12026 1751
rect 12054 1722 12082 1727
rect 11998 1721 12082 1722
rect 11998 1695 12055 1721
rect 12081 1695 12082 1721
rect 11998 1694 12082 1695
rect 11214 1666 11410 1694
rect 12054 1689 12082 1694
rect 9573 1582 10035 1587
rect 9573 1581 9582 1582
rect 9573 1555 9574 1581
rect 9573 1554 9582 1555
rect 9610 1554 9634 1582
rect 9662 1554 9686 1582
rect 9714 1581 9738 1582
rect 9766 1581 9790 1582
rect 9724 1555 9738 1581
rect 9786 1555 9790 1581
rect 9714 1554 9738 1555
rect 9766 1554 9790 1555
rect 9818 1581 9842 1582
rect 9870 1581 9894 1582
rect 9818 1555 9822 1581
rect 9870 1555 9884 1581
rect 9818 1554 9842 1555
rect 9870 1554 9894 1555
rect 9922 1554 9946 1582
rect 9974 1554 9998 1582
rect 10026 1581 10035 1582
rect 10034 1555 10035 1581
rect 10026 1554 10035 1555
rect 9573 1549 10035 1554
rect 9478 1470 9786 1498
rect 9758 400 9786 1470
rect 11214 400 11242 1666
rect 12670 400 12698 4606
rect 12726 4522 12754 4527
rect 12726 4129 12754 4494
rect 12726 4103 12727 4129
rect 12753 4103 12754 4129
rect 12726 4073 12754 4103
rect 12726 4047 12727 4073
rect 12753 4047 12754 4073
rect 12726 3346 12754 4047
rect 12950 3738 12978 4830
rect 12950 3705 12978 3710
rect 13342 6090 13370 6095
rect 13342 5697 13370 6062
rect 13510 6090 13538 6455
rect 14238 6481 14266 6846
rect 14294 6827 14322 6846
rect 14406 6874 14434 7183
rect 14573 7070 15035 7075
rect 14573 7069 14582 7070
rect 14573 7043 14574 7069
rect 14573 7042 14582 7043
rect 14610 7042 14634 7070
rect 14662 7042 14686 7070
rect 14714 7069 14738 7070
rect 14766 7069 14790 7070
rect 14724 7043 14738 7069
rect 14786 7043 14790 7069
rect 14714 7042 14738 7043
rect 14766 7042 14790 7043
rect 14818 7069 14842 7070
rect 14870 7069 14894 7070
rect 14818 7043 14822 7069
rect 14870 7043 14884 7069
rect 14818 7042 14842 7043
rect 14870 7042 14894 7043
rect 14922 7042 14946 7070
rect 14974 7042 14998 7070
rect 15026 7069 15035 7070
rect 15034 7043 15035 7069
rect 15026 7042 15035 7043
rect 14573 7037 15035 7042
rect 14406 6827 14434 6846
rect 15078 6874 15106 7630
rect 15078 6841 15106 6846
rect 15218 7657 15274 7658
rect 15218 7631 15247 7657
rect 15273 7631 15274 7657
rect 15218 7630 15274 7631
rect 15190 7265 15218 7630
rect 15246 7625 15274 7630
rect 15190 7239 15191 7265
rect 15217 7239 15218 7265
rect 15190 6874 15218 7239
rect 15246 6874 15274 6879
rect 15190 6873 15274 6874
rect 15190 6847 15247 6873
rect 15273 6847 15274 6873
rect 15190 6846 15274 6847
rect 14238 6455 14239 6481
rect 14265 6455 14266 6481
rect 14238 6425 14266 6455
rect 14238 6399 14239 6425
rect 14265 6399 14266 6425
rect 14238 6393 14266 6399
rect 14573 6286 15035 6291
rect 14573 6285 14582 6286
rect 14573 6259 14574 6285
rect 14573 6258 14582 6259
rect 14610 6258 14634 6286
rect 14662 6258 14686 6286
rect 14714 6285 14738 6286
rect 14766 6285 14790 6286
rect 14724 6259 14738 6285
rect 14786 6259 14790 6285
rect 14714 6258 14738 6259
rect 14766 6258 14790 6259
rect 14818 6285 14842 6286
rect 14870 6285 14894 6286
rect 14818 6259 14822 6285
rect 14870 6259 14884 6285
rect 14818 6258 14842 6259
rect 14870 6258 14894 6259
rect 14922 6258 14946 6286
rect 14974 6258 14998 6286
rect 15026 6285 15035 6286
rect 15034 6259 15035 6285
rect 15026 6258 15035 6259
rect 14573 6253 15035 6258
rect 14462 6146 14490 6151
rect 13510 6057 13538 6062
rect 13958 6090 13986 6095
rect 13958 6043 13986 6062
rect 13342 5671 13343 5697
rect 13369 5671 13370 5697
rect 13342 4913 13370 5671
rect 14406 5698 14434 5703
rect 14462 5698 14490 6118
rect 14854 6146 14882 6151
rect 14854 6089 14882 6118
rect 14854 6063 14855 6089
rect 14881 6063 14882 6089
rect 14854 6057 14882 6063
rect 15190 6090 15218 6846
rect 15246 6841 15274 6846
rect 14406 5697 14490 5698
rect 14406 5671 14407 5697
rect 14433 5671 14490 5697
rect 14406 5670 14490 5671
rect 14406 5641 14434 5670
rect 14406 5615 14407 5641
rect 14433 5615 14434 5641
rect 14406 5609 14434 5615
rect 14462 5361 14490 5670
rect 15190 5697 15218 6062
rect 15190 5671 15191 5697
rect 15217 5671 15218 5697
rect 14573 5502 15035 5507
rect 14573 5501 14582 5502
rect 14573 5475 14574 5501
rect 14573 5474 14582 5475
rect 14610 5474 14634 5502
rect 14662 5474 14686 5502
rect 14714 5501 14738 5502
rect 14766 5501 14790 5502
rect 14724 5475 14738 5501
rect 14786 5475 14790 5501
rect 14714 5474 14738 5475
rect 14766 5474 14790 5475
rect 14818 5501 14842 5502
rect 14870 5501 14894 5502
rect 14818 5475 14822 5501
rect 14870 5475 14884 5501
rect 14818 5474 14842 5475
rect 14870 5474 14894 5475
rect 14922 5474 14946 5502
rect 14974 5474 14998 5502
rect 15026 5501 15035 5502
rect 15034 5475 15035 5501
rect 15026 5474 15035 5475
rect 14573 5469 15035 5474
rect 14462 5335 14463 5361
rect 14489 5335 14490 5361
rect 13342 4887 13343 4913
rect 13369 4887 13370 4913
rect 13342 4129 13370 4887
rect 13342 4103 13343 4129
rect 13369 4103 13370 4129
rect 13342 3738 13370 4103
rect 12726 3289 12754 3318
rect 12726 3263 12727 3289
rect 12753 3263 12754 3289
rect 12726 3010 12754 3263
rect 12726 2561 12754 2982
rect 12726 2535 12727 2561
rect 12753 2535 12754 2561
rect 12726 2505 12754 2535
rect 12726 2479 12727 2505
rect 12753 2479 12754 2505
rect 12726 2226 12754 2479
rect 12726 2193 12754 2198
rect 13342 3402 13370 3710
rect 13566 5305 13594 5311
rect 13566 5279 13567 5305
rect 13593 5279 13594 5305
rect 13566 4521 13594 5279
rect 14182 5306 14210 5311
rect 14182 4913 14210 5278
rect 14462 5306 14490 5335
rect 14462 5240 14490 5278
rect 15190 5305 15218 5671
rect 15190 5279 15191 5305
rect 15217 5279 15218 5305
rect 15190 5273 15218 5279
rect 14182 4887 14183 4913
rect 14209 4887 14210 4913
rect 14182 4858 14210 4887
rect 13566 4495 13567 4521
rect 13593 4495 13594 4521
rect 13566 3738 13594 4495
rect 14126 4522 14154 4527
rect 14182 4522 14210 4830
rect 14573 4718 15035 4723
rect 14573 4717 14582 4718
rect 14573 4691 14574 4717
rect 14573 4690 14582 4691
rect 14610 4690 14634 4718
rect 14662 4690 14686 4718
rect 14714 4717 14738 4718
rect 14766 4717 14790 4718
rect 14724 4691 14738 4717
rect 14786 4691 14790 4717
rect 14714 4690 14738 4691
rect 14766 4690 14790 4691
rect 14818 4717 14842 4718
rect 14870 4717 14894 4718
rect 14818 4691 14822 4717
rect 14870 4691 14884 4717
rect 14818 4690 14842 4691
rect 14870 4690 14894 4691
rect 14922 4690 14946 4718
rect 14974 4690 14998 4718
rect 15026 4717 15035 4718
rect 15034 4691 15035 4717
rect 15026 4690 15035 4691
rect 14573 4685 15035 4690
rect 15526 4634 15554 9142
rect 15918 8834 15946 9198
rect 16142 8834 16170 8839
rect 15918 8833 16170 8834
rect 15918 8807 15919 8833
rect 15945 8807 16143 8833
rect 16169 8807 16170 8833
rect 15918 8806 16170 8807
rect 15694 8442 15722 8447
rect 15694 7266 15722 8414
rect 15918 8442 15946 8806
rect 16142 8801 16170 8806
rect 15918 8395 15946 8414
rect 16422 8049 16450 8055
rect 16422 8023 16423 8049
rect 16449 8023 16450 8049
rect 16422 7993 16450 8023
rect 16422 7967 16423 7993
rect 16449 7967 16450 7993
rect 16422 7713 16450 7967
rect 16422 7687 16423 7713
rect 16449 7687 16450 7713
rect 16422 7657 16450 7687
rect 16422 7631 16423 7657
rect 16449 7631 16450 7657
rect 15806 7266 15834 7271
rect 15694 7265 15834 7266
rect 15694 7239 15695 7265
rect 15721 7239 15807 7265
rect 15833 7239 15834 7265
rect 15694 7238 15834 7239
rect 15694 6146 15722 7238
rect 15806 7233 15834 7238
rect 16198 6929 16226 6935
rect 16198 6903 16199 6929
rect 16225 6903 16226 6929
rect 16198 6874 16226 6903
rect 16198 6827 16226 6846
rect 16422 6874 16450 7631
rect 16758 7658 16786 7663
rect 16758 7266 16786 7630
rect 16814 7546 16842 13426
rect 16982 13145 17010 13510
rect 17598 13482 17626 18494
rect 22073 18438 22535 18443
rect 22073 18437 22082 18438
rect 22073 18411 22074 18437
rect 22073 18410 22082 18411
rect 22110 18410 22134 18438
rect 22162 18410 22186 18438
rect 22214 18437 22238 18438
rect 22266 18437 22290 18438
rect 22224 18411 22238 18437
rect 22286 18411 22290 18437
rect 22214 18410 22238 18411
rect 22266 18410 22290 18411
rect 22318 18437 22342 18438
rect 22370 18437 22394 18438
rect 22318 18411 22322 18437
rect 22370 18411 22384 18437
rect 22318 18410 22342 18411
rect 22370 18410 22394 18411
rect 22422 18410 22446 18438
rect 22474 18410 22498 18438
rect 22526 18437 22535 18438
rect 22534 18411 22535 18437
rect 22526 18410 22535 18411
rect 22073 18405 22535 18410
rect 19573 18046 20035 18051
rect 19573 18045 19582 18046
rect 19573 18019 19574 18045
rect 19573 18018 19582 18019
rect 19610 18018 19634 18046
rect 19662 18018 19686 18046
rect 19714 18045 19738 18046
rect 19766 18045 19790 18046
rect 19724 18019 19738 18045
rect 19786 18019 19790 18045
rect 19714 18018 19738 18019
rect 19766 18018 19790 18019
rect 19818 18045 19842 18046
rect 19870 18045 19894 18046
rect 19818 18019 19822 18045
rect 19870 18019 19884 18045
rect 19818 18018 19842 18019
rect 19870 18018 19894 18019
rect 19922 18018 19946 18046
rect 19974 18018 19998 18046
rect 20026 18045 20035 18046
rect 20034 18019 20035 18045
rect 20026 18018 20035 18019
rect 19573 18013 20035 18018
rect 22073 17654 22535 17659
rect 22073 17653 22082 17654
rect 22073 17627 22074 17653
rect 22073 17626 22082 17627
rect 22110 17626 22134 17654
rect 22162 17626 22186 17654
rect 22214 17653 22238 17654
rect 22266 17653 22290 17654
rect 22224 17627 22238 17653
rect 22286 17627 22290 17653
rect 22214 17626 22238 17627
rect 22266 17626 22290 17627
rect 22318 17653 22342 17654
rect 22370 17653 22394 17654
rect 22318 17627 22322 17653
rect 22370 17627 22384 17653
rect 22318 17626 22342 17627
rect 22370 17626 22394 17627
rect 22422 17626 22446 17654
rect 22474 17626 22498 17654
rect 22526 17653 22535 17654
rect 22534 17627 22535 17653
rect 22526 17626 22535 17627
rect 22073 17621 22535 17626
rect 18494 17346 18522 17351
rect 17598 13449 17626 13454
rect 17878 17121 17906 17127
rect 17878 17095 17879 17121
rect 17905 17095 17906 17121
rect 17878 17065 17906 17095
rect 17878 17039 17879 17065
rect 17905 17039 17906 17065
rect 17878 16337 17906 17039
rect 18494 16394 18522 17318
rect 19573 17262 20035 17267
rect 19573 17261 19582 17262
rect 19573 17235 19574 17261
rect 19573 17234 19582 17235
rect 19610 17234 19634 17262
rect 19662 17234 19686 17262
rect 19714 17261 19738 17262
rect 19766 17261 19790 17262
rect 19724 17235 19738 17261
rect 19786 17235 19790 17261
rect 19714 17234 19738 17235
rect 19766 17234 19790 17235
rect 19818 17261 19842 17262
rect 19870 17261 19894 17262
rect 19818 17235 19822 17261
rect 19870 17235 19884 17261
rect 19818 17234 19842 17235
rect 19870 17234 19894 17235
rect 19922 17234 19946 17262
rect 19974 17234 19998 17262
rect 20026 17261 20035 17262
rect 20034 17235 20035 17261
rect 20026 17234 20035 17235
rect 19573 17229 20035 17234
rect 22073 16870 22535 16875
rect 22073 16869 22082 16870
rect 22073 16843 22074 16869
rect 22073 16842 22082 16843
rect 22110 16842 22134 16870
rect 22162 16842 22186 16870
rect 22214 16869 22238 16870
rect 22266 16869 22290 16870
rect 22224 16843 22238 16869
rect 22286 16843 22290 16869
rect 22214 16842 22238 16843
rect 22266 16842 22290 16843
rect 22318 16869 22342 16870
rect 22370 16869 22394 16870
rect 22318 16843 22322 16869
rect 22370 16843 22384 16869
rect 22318 16842 22342 16843
rect 22370 16842 22394 16843
rect 22422 16842 22446 16870
rect 22474 16842 22498 16870
rect 22526 16869 22535 16870
rect 22534 16843 22535 16869
rect 22526 16842 22535 16843
rect 22073 16837 22535 16842
rect 19573 16478 20035 16483
rect 19573 16477 19582 16478
rect 19573 16451 19574 16477
rect 19573 16450 19582 16451
rect 19610 16450 19634 16478
rect 19662 16450 19686 16478
rect 19714 16477 19738 16478
rect 19766 16477 19790 16478
rect 19724 16451 19738 16477
rect 19786 16451 19790 16477
rect 19714 16450 19738 16451
rect 19766 16450 19790 16451
rect 19818 16477 19842 16478
rect 19870 16477 19894 16478
rect 19818 16451 19822 16477
rect 19870 16451 19884 16477
rect 19818 16450 19842 16451
rect 19870 16450 19894 16451
rect 19922 16450 19946 16478
rect 19974 16450 19998 16478
rect 20026 16477 20035 16478
rect 20034 16451 20035 16477
rect 20026 16450 20035 16451
rect 19573 16445 20035 16450
rect 18494 16361 18522 16366
rect 17878 16311 17879 16337
rect 17905 16311 17906 16337
rect 17878 16281 17906 16311
rect 17878 16255 17879 16281
rect 17905 16255 17906 16281
rect 17878 16002 17906 16255
rect 17878 15553 17906 15974
rect 17878 15527 17879 15553
rect 17905 15527 17906 15553
rect 17878 15497 17906 15527
rect 17878 15471 17879 15497
rect 17905 15471 17906 15497
rect 16982 13119 16983 13145
rect 17009 13119 17010 13145
rect 16982 13113 17010 13119
rect 17073 12950 17535 12955
rect 17073 12949 17082 12950
rect 17073 12923 17074 12949
rect 17073 12922 17082 12923
rect 17110 12922 17134 12950
rect 17162 12922 17186 12950
rect 17214 12949 17238 12950
rect 17266 12949 17290 12950
rect 17224 12923 17238 12949
rect 17286 12923 17290 12949
rect 17214 12922 17238 12923
rect 17266 12922 17290 12923
rect 17318 12949 17342 12950
rect 17370 12949 17394 12950
rect 17318 12923 17322 12949
rect 17370 12923 17384 12949
rect 17318 12922 17342 12923
rect 17370 12922 17394 12923
rect 17422 12922 17446 12950
rect 17474 12922 17498 12950
rect 17526 12949 17535 12950
rect 17534 12923 17535 12949
rect 17526 12922 17535 12923
rect 17073 12917 17535 12922
rect 16926 12753 16954 12759
rect 16926 12727 16927 12753
rect 16953 12727 16954 12753
rect 16926 12361 16954 12727
rect 16926 12335 16927 12361
rect 16953 12335 16954 12361
rect 16926 11970 16954 12335
rect 17878 12753 17906 15471
rect 18270 16281 18298 16287
rect 18270 16255 18271 16281
rect 18297 16255 18298 16281
rect 18270 15890 18298 16255
rect 18270 15497 18298 15862
rect 18270 15471 18271 15497
rect 18297 15471 18298 15497
rect 17934 14769 17962 14775
rect 17934 14743 17935 14769
rect 17961 14743 17962 14769
rect 17934 14713 17962 14743
rect 17934 14687 17935 14713
rect 17961 14687 17962 14713
rect 17934 14266 17962 14687
rect 17934 13985 17962 14238
rect 17934 13959 17935 13985
rect 17961 13959 17962 13985
rect 17934 13929 17962 13959
rect 17934 13903 17935 13929
rect 17961 13903 17962 13929
rect 17934 13537 17962 13903
rect 17934 13511 17935 13537
rect 17961 13511 17962 13537
rect 17934 13482 17962 13511
rect 18270 14713 18298 15471
rect 18718 16282 18746 16287
rect 18942 16282 18970 16287
rect 18718 16281 18970 16282
rect 18718 16255 18719 16281
rect 18745 16255 18943 16281
rect 18969 16255 18970 16281
rect 18718 16254 18970 16255
rect 18718 16002 18746 16254
rect 18942 16249 18970 16254
rect 22582 16282 22610 18494
rect 27073 18438 27535 18443
rect 27073 18437 27082 18438
rect 27073 18411 27074 18437
rect 27073 18410 27082 18411
rect 27110 18410 27134 18438
rect 27162 18410 27186 18438
rect 27214 18437 27238 18438
rect 27266 18437 27290 18438
rect 27224 18411 27238 18437
rect 27286 18411 27290 18437
rect 27214 18410 27238 18411
rect 27266 18410 27290 18411
rect 27318 18437 27342 18438
rect 27370 18437 27394 18438
rect 27318 18411 27322 18437
rect 27370 18411 27384 18437
rect 27318 18410 27342 18411
rect 27370 18410 27394 18411
rect 27422 18410 27446 18438
rect 27474 18410 27498 18438
rect 27526 18437 27535 18438
rect 27534 18411 27535 18437
rect 27526 18410 27535 18411
rect 27073 18405 27535 18410
rect 24573 18046 25035 18051
rect 24573 18045 24582 18046
rect 24573 18019 24574 18045
rect 24573 18018 24582 18019
rect 24610 18018 24634 18046
rect 24662 18018 24686 18046
rect 24714 18045 24738 18046
rect 24766 18045 24790 18046
rect 24724 18019 24738 18045
rect 24786 18019 24790 18045
rect 24714 18018 24738 18019
rect 24766 18018 24790 18019
rect 24818 18045 24842 18046
rect 24870 18045 24894 18046
rect 24818 18019 24822 18045
rect 24870 18019 24884 18045
rect 24818 18018 24842 18019
rect 24870 18018 24894 18019
rect 24922 18018 24946 18046
rect 24974 18018 24998 18046
rect 25026 18045 25035 18046
rect 25034 18019 25035 18045
rect 25026 18018 25035 18019
rect 24573 18013 25035 18018
rect 27073 17654 27535 17659
rect 27073 17653 27082 17654
rect 27073 17627 27074 17653
rect 27073 17626 27082 17627
rect 27110 17626 27134 17654
rect 27162 17626 27186 17654
rect 27214 17653 27238 17654
rect 27266 17653 27290 17654
rect 27224 17627 27238 17653
rect 27286 17627 27290 17653
rect 27214 17626 27238 17627
rect 27266 17626 27290 17627
rect 27318 17653 27342 17654
rect 27370 17653 27394 17654
rect 27318 17627 27322 17653
rect 27370 17627 27384 17653
rect 27318 17626 27342 17627
rect 27370 17626 27394 17627
rect 27422 17626 27446 17654
rect 27474 17626 27498 17654
rect 27526 17653 27535 17654
rect 27534 17627 27535 17653
rect 27526 17626 27535 17627
rect 27073 17621 27535 17626
rect 24573 17262 25035 17267
rect 24573 17261 24582 17262
rect 24573 17235 24574 17261
rect 24573 17234 24582 17235
rect 24610 17234 24634 17262
rect 24662 17234 24686 17262
rect 24714 17261 24738 17262
rect 24766 17261 24790 17262
rect 24724 17235 24738 17261
rect 24786 17235 24790 17261
rect 24714 17234 24738 17235
rect 24766 17234 24790 17235
rect 24818 17261 24842 17262
rect 24870 17261 24894 17262
rect 24818 17235 24822 17261
rect 24870 17235 24884 17261
rect 24818 17234 24842 17235
rect 24870 17234 24894 17235
rect 24922 17234 24946 17262
rect 24974 17234 24998 17262
rect 25026 17261 25035 17262
rect 25034 17235 25035 17261
rect 25026 17234 25035 17235
rect 24573 17229 25035 17234
rect 27073 16870 27535 16875
rect 27073 16869 27082 16870
rect 27073 16843 27074 16869
rect 27073 16842 27082 16843
rect 27110 16842 27134 16870
rect 27162 16842 27186 16870
rect 27214 16869 27238 16870
rect 27266 16869 27290 16870
rect 27224 16843 27238 16869
rect 27286 16843 27290 16869
rect 27214 16842 27238 16843
rect 27266 16842 27290 16843
rect 27318 16869 27342 16870
rect 27370 16869 27394 16870
rect 27318 16843 27322 16869
rect 27370 16843 27384 16869
rect 27318 16842 27342 16843
rect 27370 16842 27394 16843
rect 27422 16842 27446 16870
rect 27474 16842 27498 16870
rect 27526 16869 27535 16870
rect 27534 16843 27535 16869
rect 27526 16842 27535 16843
rect 27073 16837 27535 16842
rect 24573 16478 25035 16483
rect 24573 16477 24582 16478
rect 24573 16451 24574 16477
rect 24573 16450 24582 16451
rect 24610 16450 24634 16478
rect 24662 16450 24686 16478
rect 24714 16477 24738 16478
rect 24766 16477 24790 16478
rect 24724 16451 24738 16477
rect 24786 16451 24790 16477
rect 24714 16450 24738 16451
rect 24766 16450 24790 16451
rect 24818 16477 24842 16478
rect 24870 16477 24894 16478
rect 24818 16451 24822 16477
rect 24870 16451 24884 16477
rect 24818 16450 24842 16451
rect 24870 16450 24894 16451
rect 24922 16450 24946 16478
rect 24974 16450 24998 16478
rect 25026 16477 25035 16478
rect 25034 16451 25035 16477
rect 25026 16450 25035 16451
rect 24573 16445 25035 16450
rect 22582 16249 22610 16254
rect 24094 16394 24122 16399
rect 22073 16086 22535 16091
rect 22073 16085 22082 16086
rect 22073 16059 22074 16085
rect 22073 16058 22082 16059
rect 22110 16058 22134 16086
rect 22162 16058 22186 16086
rect 22214 16085 22238 16086
rect 22266 16085 22290 16086
rect 22224 16059 22238 16085
rect 22286 16059 22290 16085
rect 22214 16058 22238 16059
rect 22266 16058 22290 16059
rect 22318 16085 22342 16086
rect 22370 16085 22394 16086
rect 22318 16059 22322 16085
rect 22370 16059 22384 16085
rect 22318 16058 22342 16059
rect 22370 16058 22394 16059
rect 22422 16058 22446 16086
rect 22474 16058 22498 16086
rect 22526 16085 22535 16086
rect 22534 16059 22535 16085
rect 22526 16058 22535 16059
rect 22073 16053 22535 16058
rect 18718 15498 18746 15974
rect 19222 16002 19250 16007
rect 18774 15890 18802 15895
rect 18774 15843 18802 15862
rect 19222 15890 19250 15974
rect 19446 15890 19474 15895
rect 19222 15889 19474 15890
rect 19222 15863 19223 15889
rect 19249 15863 19447 15889
rect 19473 15863 19474 15889
rect 19222 15862 19474 15863
rect 19222 15857 19250 15862
rect 18942 15498 18970 15503
rect 18718 15497 18970 15498
rect 18718 15471 18719 15497
rect 18745 15471 18943 15497
rect 18969 15471 18970 15497
rect 18718 15470 18970 15471
rect 18718 15465 18746 15470
rect 18942 15465 18970 15470
rect 18270 14687 18271 14713
rect 18297 14687 18298 14713
rect 18270 14322 18298 14687
rect 18270 13929 18298 14294
rect 18270 13903 18271 13929
rect 18297 13903 18298 13929
rect 17934 13481 18018 13482
rect 17934 13455 17935 13481
rect 17961 13455 18018 13481
rect 17934 13454 18018 13455
rect 17934 13449 17962 13454
rect 17990 13201 18018 13454
rect 18270 13454 18298 13903
rect 18830 15105 18858 15111
rect 18830 15079 18831 15105
rect 18857 15079 18858 15105
rect 18830 14321 18858 15079
rect 19334 15106 19362 15111
rect 19446 15106 19474 15862
rect 19573 15694 20035 15699
rect 19573 15693 19582 15694
rect 19573 15667 19574 15693
rect 19573 15666 19582 15667
rect 19610 15666 19634 15694
rect 19662 15666 19686 15694
rect 19714 15693 19738 15694
rect 19766 15693 19790 15694
rect 19724 15667 19738 15693
rect 19786 15667 19790 15693
rect 19714 15666 19738 15667
rect 19766 15666 19790 15667
rect 19818 15693 19842 15694
rect 19870 15693 19894 15694
rect 19818 15667 19822 15693
rect 19870 15667 19884 15693
rect 19818 15666 19842 15667
rect 19870 15666 19894 15667
rect 19922 15666 19946 15694
rect 19974 15666 19998 15694
rect 20026 15693 20035 15694
rect 20034 15667 20035 15693
rect 20026 15666 20035 15667
rect 19573 15661 20035 15666
rect 23422 15553 23450 15559
rect 23422 15527 23423 15553
rect 23449 15527 23450 15553
rect 20790 15497 20818 15503
rect 20790 15471 20791 15497
rect 20817 15471 20818 15497
rect 19334 15105 19474 15106
rect 19334 15079 19335 15105
rect 19361 15079 19447 15105
rect 19473 15079 19474 15105
rect 19334 15078 19474 15079
rect 19334 15073 19362 15078
rect 19446 14769 19474 15078
rect 20510 15105 20538 15111
rect 20510 15079 20511 15105
rect 20537 15079 20538 15105
rect 19573 14910 20035 14915
rect 19573 14909 19582 14910
rect 19573 14883 19574 14909
rect 19573 14882 19582 14883
rect 19610 14882 19634 14910
rect 19662 14882 19686 14910
rect 19714 14909 19738 14910
rect 19766 14909 19790 14910
rect 19724 14883 19738 14909
rect 19786 14883 19790 14909
rect 19714 14882 19738 14883
rect 19766 14882 19790 14883
rect 19818 14909 19842 14910
rect 19870 14909 19894 14910
rect 19818 14883 19822 14909
rect 19870 14883 19884 14909
rect 19818 14882 19842 14883
rect 19870 14882 19894 14883
rect 19922 14882 19946 14910
rect 19974 14882 19998 14910
rect 20026 14909 20035 14910
rect 20034 14883 20035 14909
rect 20026 14882 20035 14883
rect 19573 14877 20035 14882
rect 19446 14743 19447 14769
rect 19473 14743 19474 14769
rect 19446 14713 19474 14743
rect 19446 14687 19447 14713
rect 19473 14687 19474 14713
rect 18830 14295 18831 14321
rect 18857 14295 18858 14321
rect 18830 13537 18858 14295
rect 19334 14322 19362 14327
rect 19446 14322 19474 14687
rect 19334 14321 19446 14322
rect 19334 14295 19335 14321
rect 19361 14295 19446 14321
rect 19334 14294 19446 14295
rect 19334 14289 19362 14294
rect 19446 13985 19474 14294
rect 20510 14321 20538 15079
rect 20790 14713 20818 15471
rect 21238 15498 21266 15503
rect 21462 15498 21490 15503
rect 21238 15497 21490 15498
rect 21238 15471 21239 15497
rect 21265 15471 21463 15497
rect 21489 15471 21490 15497
rect 21238 15470 21490 15471
rect 20790 14687 20791 14713
rect 20817 14687 20818 14713
rect 20790 14658 20818 14687
rect 20790 14625 20818 14630
rect 21014 15105 21042 15111
rect 21014 15079 21015 15105
rect 21041 15079 21042 15105
rect 21014 15050 21042 15079
rect 21182 15050 21210 15055
rect 21238 15050 21266 15470
rect 21462 15465 21490 15470
rect 22526 15498 22554 15503
rect 22526 15497 22610 15498
rect 22526 15471 22527 15497
rect 22553 15471 22610 15497
rect 22526 15470 22610 15471
rect 22526 15465 22554 15470
rect 22073 15302 22535 15307
rect 22073 15301 22082 15302
rect 22073 15275 22074 15301
rect 22073 15274 22082 15275
rect 22110 15274 22134 15302
rect 22162 15274 22186 15302
rect 22214 15301 22238 15302
rect 22266 15301 22290 15302
rect 22224 15275 22238 15301
rect 22286 15275 22290 15301
rect 22214 15274 22238 15275
rect 22266 15274 22290 15275
rect 22318 15301 22342 15302
rect 22370 15301 22394 15302
rect 22318 15275 22322 15301
rect 22370 15275 22384 15301
rect 22318 15274 22342 15275
rect 22370 15274 22394 15275
rect 22422 15274 22446 15302
rect 22474 15274 22498 15302
rect 22526 15301 22535 15302
rect 22534 15275 22535 15301
rect 22526 15274 22535 15275
rect 22073 15269 22535 15274
rect 21014 15049 21266 15050
rect 21014 15023 21183 15049
rect 21209 15023 21266 15049
rect 21014 15022 21266 15023
rect 20510 14295 20511 14321
rect 20537 14295 20538 14321
rect 19573 14126 20035 14131
rect 19573 14125 19582 14126
rect 19573 14099 19574 14125
rect 19573 14098 19582 14099
rect 19610 14098 19634 14126
rect 19662 14098 19686 14126
rect 19714 14125 19738 14126
rect 19766 14125 19790 14126
rect 19724 14099 19738 14125
rect 19786 14099 19790 14125
rect 19714 14098 19738 14099
rect 19766 14098 19790 14099
rect 19818 14125 19842 14126
rect 19870 14125 19894 14126
rect 19818 14099 19822 14125
rect 19870 14099 19884 14125
rect 19818 14098 19842 14099
rect 19870 14098 19894 14099
rect 19922 14098 19946 14126
rect 19974 14098 19998 14126
rect 20026 14125 20035 14126
rect 20034 14099 20035 14125
rect 20026 14098 20035 14099
rect 19573 14093 20035 14098
rect 19446 13959 19447 13985
rect 19473 13959 19474 13985
rect 19446 13929 19474 13959
rect 19446 13903 19447 13929
rect 19473 13903 19474 13929
rect 18830 13511 18831 13537
rect 18857 13511 18858 13537
rect 18830 13454 18858 13511
rect 19334 13538 19362 13543
rect 19446 13538 19474 13903
rect 19334 13537 19474 13538
rect 19334 13511 19335 13537
rect 19361 13511 19447 13537
rect 19473 13511 19474 13537
rect 19334 13510 19474 13511
rect 19334 13505 19362 13510
rect 19446 13505 19474 13510
rect 20510 13537 20538 14295
rect 20678 14322 20706 14327
rect 20678 14275 20706 14294
rect 21014 14322 21042 15022
rect 21182 15017 21210 15022
rect 21238 14714 21266 15022
rect 21462 14714 21490 14719
rect 21238 14713 21490 14714
rect 21238 14687 21239 14713
rect 21265 14687 21463 14713
rect 21489 14687 21490 14713
rect 21238 14686 21490 14687
rect 21238 14681 21266 14686
rect 21462 14681 21490 14686
rect 22526 14714 22554 14719
rect 22582 14714 22610 15470
rect 23422 15497 23450 15527
rect 23422 15471 23423 15497
rect 23449 15471 23450 15497
rect 22526 14713 22610 14714
rect 22526 14687 22527 14713
rect 22553 14687 22610 14713
rect 22526 14686 22610 14687
rect 22526 14681 22554 14686
rect 22582 14658 22610 14686
rect 22073 14518 22535 14523
rect 22073 14517 22082 14518
rect 22073 14491 22074 14517
rect 22073 14490 22082 14491
rect 22110 14490 22134 14518
rect 22162 14490 22186 14518
rect 22214 14517 22238 14518
rect 22266 14517 22290 14518
rect 22224 14491 22238 14517
rect 22286 14491 22290 14517
rect 22214 14490 22238 14491
rect 22266 14490 22290 14491
rect 22318 14517 22342 14518
rect 22370 14517 22394 14518
rect 22318 14491 22322 14517
rect 22370 14491 22384 14517
rect 22318 14490 22342 14491
rect 22370 14490 22394 14491
rect 22422 14490 22446 14518
rect 22474 14490 22498 14518
rect 22526 14517 22535 14518
rect 22534 14491 22535 14517
rect 22526 14490 22535 14491
rect 22073 14485 22535 14490
rect 20510 13511 20511 13537
rect 20537 13511 20538 13537
rect 18270 13426 18578 13454
rect 18830 13426 19082 13454
rect 17990 13175 17991 13201
rect 18017 13175 18018 13201
rect 17990 13146 18018 13175
rect 17990 13099 18018 13118
rect 18550 13145 18578 13398
rect 19054 13393 19082 13398
rect 19573 13342 20035 13347
rect 19573 13341 19582 13342
rect 19573 13315 19574 13341
rect 19573 13314 19582 13315
rect 19610 13314 19634 13342
rect 19662 13314 19686 13342
rect 19714 13341 19738 13342
rect 19766 13341 19790 13342
rect 19724 13315 19738 13341
rect 19786 13315 19790 13341
rect 19714 13314 19738 13315
rect 19766 13314 19790 13315
rect 19818 13341 19842 13342
rect 19870 13341 19894 13342
rect 19818 13315 19822 13341
rect 19870 13315 19884 13341
rect 19818 13314 19842 13315
rect 19870 13314 19894 13315
rect 19922 13314 19946 13342
rect 19974 13314 19998 13342
rect 20026 13341 20035 13342
rect 20034 13315 20035 13341
rect 20026 13314 20035 13315
rect 19573 13309 20035 13314
rect 18550 13119 18551 13145
rect 18577 13119 18578 13145
rect 17878 12727 17879 12753
rect 17905 12727 17906 12753
rect 17878 12697 17906 12727
rect 17878 12671 17879 12697
rect 17905 12671 17906 12697
rect 17878 12417 17906 12671
rect 17878 12391 17879 12417
rect 17905 12391 17906 12417
rect 17878 12361 17906 12391
rect 17878 12335 17879 12361
rect 17905 12335 17906 12361
rect 17073 12166 17535 12171
rect 17073 12165 17082 12166
rect 17073 12139 17074 12165
rect 17073 12138 17082 12139
rect 17110 12138 17134 12166
rect 17162 12138 17186 12166
rect 17214 12165 17238 12166
rect 17266 12165 17290 12166
rect 17224 12139 17238 12165
rect 17286 12139 17290 12165
rect 17214 12138 17238 12139
rect 17266 12138 17290 12139
rect 17318 12165 17342 12166
rect 17370 12165 17394 12166
rect 17318 12139 17322 12165
rect 17370 12139 17384 12165
rect 17318 12138 17342 12139
rect 17370 12138 17394 12139
rect 17422 12138 17446 12166
rect 17474 12138 17498 12166
rect 17526 12165 17535 12166
rect 17534 12139 17535 12165
rect 17526 12138 17535 12139
rect 17073 12133 17535 12138
rect 17038 11970 17066 11975
rect 16954 11969 17066 11970
rect 16954 11943 17039 11969
rect 17065 11943 17066 11969
rect 16954 11942 17066 11943
rect 16926 11904 16954 11942
rect 17038 11937 17066 11942
rect 17878 11970 17906 12335
rect 18550 12362 18578 13119
rect 19446 13201 19474 13207
rect 19446 13175 19447 13201
rect 19473 13175 19474 13201
rect 19446 13146 19474 13175
rect 18774 12753 18802 12759
rect 18774 12727 18775 12753
rect 18801 12727 18802 12753
rect 18774 12642 18802 12727
rect 18774 12362 18802 12614
rect 18550 12361 18802 12362
rect 18550 12335 18551 12361
rect 18577 12335 18802 12361
rect 18550 12334 18802 12335
rect 18550 12329 18578 12334
rect 17878 11969 18018 11970
rect 17878 11943 17879 11969
rect 17905 11943 18018 11969
rect 17878 11942 18018 11943
rect 17878 11937 17906 11942
rect 17990 11913 18018 11942
rect 18774 11969 18802 12334
rect 19446 12698 19474 13118
rect 19446 12417 19474 12670
rect 19950 12753 19978 12759
rect 19950 12727 19951 12753
rect 19977 12727 19978 12753
rect 19950 12698 19978 12727
rect 19950 12642 19978 12670
rect 20510 12753 20538 13511
rect 20510 12727 20511 12753
rect 20537 12727 20538 12753
rect 20510 12642 20538 12727
rect 19950 12614 20146 12642
rect 19573 12558 20035 12563
rect 19573 12557 19582 12558
rect 19573 12531 19574 12557
rect 19573 12530 19582 12531
rect 19610 12530 19634 12558
rect 19662 12530 19686 12558
rect 19714 12557 19738 12558
rect 19766 12557 19790 12558
rect 19724 12531 19738 12557
rect 19786 12531 19790 12557
rect 19714 12530 19738 12531
rect 19766 12530 19790 12531
rect 19818 12557 19842 12558
rect 19870 12557 19894 12558
rect 19818 12531 19822 12557
rect 19870 12531 19884 12557
rect 19818 12530 19842 12531
rect 19870 12530 19894 12531
rect 19922 12530 19946 12558
rect 19974 12530 19998 12558
rect 20026 12557 20035 12558
rect 20034 12531 20035 12557
rect 20026 12530 20035 12531
rect 19573 12525 20035 12530
rect 19446 12391 19447 12417
rect 19473 12391 19474 12417
rect 19446 12361 19474 12391
rect 19446 12335 19447 12361
rect 19473 12335 19474 12361
rect 19446 12329 19474 12335
rect 18774 11943 18775 11969
rect 18801 11943 18802 11969
rect 18774 11937 18802 11943
rect 19950 11970 19978 11975
rect 17990 11887 17991 11913
rect 18017 11887 18018 11913
rect 17990 11633 18018 11887
rect 19950 11913 19978 11942
rect 20118 11970 20146 12614
rect 20118 11937 20146 11942
rect 20510 11969 20538 12614
rect 20510 11943 20511 11969
rect 20537 11943 20538 11969
rect 19950 11887 19951 11913
rect 19977 11887 19978 11913
rect 19950 11881 19978 11887
rect 19573 11774 20035 11779
rect 19573 11773 19582 11774
rect 19573 11747 19574 11773
rect 19573 11746 19582 11747
rect 19610 11746 19634 11774
rect 19662 11746 19686 11774
rect 19714 11773 19738 11774
rect 19766 11773 19790 11774
rect 19724 11747 19738 11773
rect 19786 11747 19790 11773
rect 19714 11746 19738 11747
rect 19766 11746 19790 11747
rect 19818 11773 19842 11774
rect 19870 11773 19894 11774
rect 19818 11747 19822 11773
rect 19870 11747 19884 11773
rect 19818 11746 19842 11747
rect 19870 11746 19894 11747
rect 19922 11746 19946 11774
rect 19974 11746 19998 11774
rect 20026 11773 20035 11774
rect 20034 11747 20035 11773
rect 20026 11746 20035 11747
rect 19573 11741 20035 11746
rect 17990 11607 17991 11633
rect 18017 11607 18018 11633
rect 16982 11577 17010 11583
rect 16982 11551 16983 11577
rect 17009 11551 17010 11577
rect 16982 11186 17010 11551
rect 17990 11577 18018 11607
rect 19334 11633 19362 11639
rect 19334 11607 19335 11633
rect 19361 11607 19362 11633
rect 17990 11551 17991 11577
rect 18017 11551 18018 11577
rect 17073 11382 17535 11387
rect 17073 11381 17082 11382
rect 17073 11355 17074 11381
rect 17073 11354 17082 11355
rect 17110 11354 17134 11382
rect 17162 11354 17186 11382
rect 17214 11381 17238 11382
rect 17266 11381 17290 11382
rect 17224 11355 17238 11381
rect 17286 11355 17290 11381
rect 17214 11354 17238 11355
rect 17266 11354 17290 11355
rect 17318 11381 17342 11382
rect 17370 11381 17394 11382
rect 17318 11355 17322 11381
rect 17370 11355 17384 11381
rect 17318 11354 17342 11355
rect 17370 11354 17394 11355
rect 17422 11354 17446 11382
rect 17474 11354 17498 11382
rect 17526 11381 17535 11382
rect 17534 11355 17535 11381
rect 17526 11354 17535 11355
rect 17073 11349 17535 11354
rect 17094 11186 17122 11191
rect 16982 11185 17122 11186
rect 16982 11159 17095 11185
rect 17121 11159 17122 11185
rect 16982 11158 17122 11159
rect 16982 10793 17010 11158
rect 17094 11153 17122 11158
rect 17990 11186 18018 11551
rect 18550 11577 18578 11583
rect 18550 11551 18551 11577
rect 18577 11551 18578 11577
rect 17990 11185 18074 11186
rect 17990 11159 17991 11185
rect 18017 11159 18074 11185
rect 17990 11158 18074 11159
rect 16982 10767 16983 10793
rect 17009 10767 17010 10793
rect 16982 10010 17010 10767
rect 17990 10849 18018 11158
rect 18046 11129 18074 11158
rect 18046 11103 18047 11129
rect 18073 11103 18074 11129
rect 18046 11097 18074 11103
rect 17990 10823 17991 10849
rect 18017 10823 18018 10849
rect 17990 10793 18018 10823
rect 17990 10767 17991 10793
rect 18017 10767 18018 10793
rect 17654 10738 17682 10743
rect 17073 10598 17535 10603
rect 17073 10597 17082 10598
rect 17073 10571 17074 10597
rect 17073 10570 17082 10571
rect 17110 10570 17134 10598
rect 17162 10570 17186 10598
rect 17214 10597 17238 10598
rect 17266 10597 17290 10598
rect 17224 10571 17238 10597
rect 17286 10571 17290 10597
rect 17214 10570 17238 10571
rect 17266 10570 17290 10571
rect 17318 10597 17342 10598
rect 17370 10597 17394 10598
rect 17318 10571 17322 10597
rect 17370 10571 17384 10597
rect 17318 10570 17342 10571
rect 17370 10570 17394 10571
rect 17422 10570 17446 10598
rect 17474 10570 17498 10598
rect 17526 10597 17535 10598
rect 17534 10571 17535 10597
rect 17526 10570 17535 10571
rect 17073 10565 17535 10570
rect 17150 10401 17178 10407
rect 17150 10375 17151 10401
rect 17177 10375 17178 10401
rect 17150 10010 17178 10375
rect 16982 10009 17178 10010
rect 16982 9983 16983 10009
rect 17009 9983 17178 10009
rect 16982 9982 17178 9983
rect 16982 9618 17010 9982
rect 17073 9814 17535 9819
rect 17073 9813 17082 9814
rect 17073 9787 17074 9813
rect 17073 9786 17082 9787
rect 17110 9786 17134 9814
rect 17162 9786 17186 9814
rect 17214 9813 17238 9814
rect 17266 9813 17290 9814
rect 17224 9787 17238 9813
rect 17286 9787 17290 9813
rect 17214 9786 17238 9787
rect 17266 9786 17290 9787
rect 17318 9813 17342 9814
rect 17370 9813 17394 9814
rect 17318 9787 17322 9813
rect 17370 9787 17384 9813
rect 17318 9786 17342 9787
rect 17370 9786 17394 9787
rect 17422 9786 17446 9814
rect 17474 9786 17498 9814
rect 17526 9813 17535 9814
rect 17534 9787 17535 9813
rect 17526 9786 17535 9787
rect 17073 9781 17535 9786
rect 17094 9618 17122 9623
rect 16982 9617 17122 9618
rect 16982 9591 17095 9617
rect 17121 9591 17122 9617
rect 16982 9590 17122 9591
rect 17094 9226 17122 9590
rect 17206 9226 17234 9231
rect 16982 9225 17234 9226
rect 16982 9199 17207 9225
rect 17233 9199 17234 9225
rect 16982 9198 17234 9199
rect 16982 8834 17010 9198
rect 17206 9193 17234 9198
rect 17654 9170 17682 10710
rect 17990 10402 18018 10767
rect 18550 10793 18578 11551
rect 19334 11577 19362 11607
rect 19334 11551 19335 11577
rect 19361 11551 19362 11577
rect 18886 11242 18914 11247
rect 18550 10767 18551 10793
rect 18577 10767 18578 10793
rect 18018 10374 18130 10402
rect 17990 10065 18018 10374
rect 18102 10346 18130 10374
rect 18102 10280 18130 10318
rect 17990 10039 17991 10065
rect 18017 10039 18018 10065
rect 17990 10009 18018 10039
rect 17990 9983 17991 10009
rect 18017 9983 18018 10009
rect 17990 9977 18018 9983
rect 18550 10009 18578 10767
rect 18774 11185 18802 11191
rect 18774 11159 18775 11185
rect 18801 11159 18802 11185
rect 18774 10401 18802 11159
rect 18774 10375 18775 10401
rect 18801 10375 18802 10401
rect 18550 9983 18551 10009
rect 18577 9983 18578 10009
rect 18270 9618 18298 9623
rect 18270 9561 18298 9590
rect 18270 9535 18271 9561
rect 18297 9535 18298 9561
rect 18270 9281 18298 9535
rect 18550 9506 18578 9983
rect 18718 10010 18746 10015
rect 18718 9618 18746 9982
rect 18718 9585 18746 9590
rect 18774 9617 18802 10375
rect 18774 9591 18775 9617
rect 18801 9591 18802 9617
rect 18774 9506 18802 9591
rect 18550 9478 18802 9506
rect 18270 9255 18271 9281
rect 18297 9255 18298 9281
rect 18270 9225 18298 9255
rect 18270 9199 18271 9225
rect 18297 9199 18298 9225
rect 17654 9137 17682 9142
rect 18214 9170 18242 9175
rect 17073 9030 17535 9035
rect 17073 9029 17082 9030
rect 17073 9003 17074 9029
rect 17073 9002 17082 9003
rect 17110 9002 17134 9030
rect 17162 9002 17186 9030
rect 17214 9029 17238 9030
rect 17266 9029 17290 9030
rect 17224 9003 17238 9029
rect 17286 9003 17290 9029
rect 17214 9002 17238 9003
rect 17266 9002 17290 9003
rect 17318 9029 17342 9030
rect 17370 9029 17394 9030
rect 17318 9003 17322 9029
rect 17370 9003 17384 9029
rect 17318 9002 17342 9003
rect 17370 9002 17394 9003
rect 17422 9002 17446 9030
rect 17474 9002 17498 9030
rect 17526 9029 17535 9030
rect 17534 9003 17535 9029
rect 17526 9002 17535 9003
rect 17073 8997 17535 9002
rect 17206 8834 17234 8839
rect 16982 8806 17206 8834
rect 17094 8442 17122 8806
rect 17206 8768 17234 8806
rect 16870 8441 17122 8442
rect 16870 8415 17095 8441
rect 17121 8415 17122 8441
rect 16870 8414 17122 8415
rect 16870 8049 16898 8414
rect 17094 8409 17122 8414
rect 17073 8246 17535 8251
rect 17073 8245 17082 8246
rect 17073 8219 17074 8245
rect 17073 8218 17082 8219
rect 17110 8218 17134 8246
rect 17162 8218 17186 8246
rect 17214 8245 17238 8246
rect 17266 8245 17290 8246
rect 17224 8219 17238 8245
rect 17286 8219 17290 8245
rect 17214 8218 17238 8219
rect 17266 8218 17290 8219
rect 17318 8245 17342 8246
rect 17370 8245 17394 8246
rect 17318 8219 17322 8245
rect 17370 8219 17384 8245
rect 17318 8218 17342 8219
rect 17370 8218 17394 8219
rect 17422 8218 17446 8246
rect 17474 8218 17498 8246
rect 17526 8245 17535 8246
rect 17534 8219 17535 8245
rect 17526 8218 17535 8219
rect 17073 8213 17535 8218
rect 16870 8023 16871 8049
rect 16897 8023 16898 8049
rect 16870 7658 16898 8023
rect 16870 7611 16898 7630
rect 17710 8049 17738 8055
rect 17710 8023 17711 8049
rect 17737 8023 17738 8049
rect 17710 7993 17738 8023
rect 17710 7967 17711 7993
rect 17737 7967 17738 7993
rect 17710 7714 17738 7967
rect 17766 7714 17794 7719
rect 17710 7713 17794 7714
rect 17710 7687 17767 7713
rect 17793 7687 17794 7713
rect 17710 7686 17794 7687
rect 17710 7657 17738 7686
rect 17766 7681 17794 7686
rect 17710 7631 17711 7657
rect 17737 7631 17738 7657
rect 16814 7518 16898 7546
rect 16814 7266 16842 7271
rect 16758 7265 16842 7266
rect 16758 7239 16815 7265
rect 16841 7239 16842 7265
rect 16758 7238 16842 7239
rect 16422 6841 16450 6846
rect 16814 6873 16842 7238
rect 16814 6847 16815 6873
rect 16841 6847 16842 6873
rect 15694 6090 15722 6118
rect 16366 6481 16394 6487
rect 16366 6455 16367 6481
rect 16393 6455 16394 6481
rect 15862 6090 15890 6095
rect 15694 6089 15890 6090
rect 15694 6063 15695 6089
rect 15721 6063 15863 6089
rect 15889 6063 15890 6089
rect 15694 6062 15890 6063
rect 15694 6057 15722 6062
rect 15862 5697 15890 6062
rect 16366 5894 16394 6455
rect 16814 6089 16842 6847
rect 16814 6063 16815 6089
rect 16841 6063 16842 6089
rect 16366 5866 16450 5894
rect 16422 5833 16450 5838
rect 16814 5866 16842 6063
rect 16870 5894 16898 7518
rect 17073 7462 17535 7467
rect 17073 7461 17082 7462
rect 17073 7435 17074 7461
rect 17073 7434 17082 7435
rect 17110 7434 17134 7462
rect 17162 7434 17186 7462
rect 17214 7461 17238 7462
rect 17266 7461 17290 7462
rect 17224 7435 17238 7461
rect 17286 7435 17290 7461
rect 17214 7434 17238 7435
rect 17266 7434 17290 7435
rect 17318 7461 17342 7462
rect 17370 7461 17394 7462
rect 17318 7435 17322 7461
rect 17370 7435 17384 7461
rect 17318 7434 17342 7435
rect 17370 7434 17394 7435
rect 17422 7434 17446 7462
rect 17474 7434 17498 7462
rect 17526 7461 17535 7462
rect 17534 7435 17535 7461
rect 17526 7434 17535 7435
rect 17073 7429 17535 7434
rect 17262 7266 17290 7271
rect 17374 7266 17402 7271
rect 17262 7265 17402 7266
rect 17262 7239 17263 7265
rect 17289 7239 17375 7265
rect 17401 7239 17402 7265
rect 17262 7238 17402 7239
rect 17262 7233 17290 7238
rect 17374 6874 17402 7238
rect 17598 6874 17626 6879
rect 17710 6874 17738 7631
rect 17402 6873 17738 6874
rect 17402 6847 17599 6873
rect 17625 6847 17738 6873
rect 17402 6846 17738 6847
rect 17374 6808 17402 6846
rect 17073 6678 17535 6683
rect 17073 6677 17082 6678
rect 17073 6651 17074 6677
rect 17073 6650 17082 6651
rect 17110 6650 17134 6678
rect 17162 6650 17186 6678
rect 17214 6677 17238 6678
rect 17266 6677 17290 6678
rect 17224 6651 17238 6677
rect 17286 6651 17290 6677
rect 17214 6650 17238 6651
rect 17266 6650 17290 6651
rect 17318 6677 17342 6678
rect 17370 6677 17394 6678
rect 17318 6651 17322 6677
rect 17370 6651 17384 6677
rect 17318 6650 17342 6651
rect 17370 6650 17394 6651
rect 17422 6650 17446 6678
rect 17474 6650 17498 6678
rect 17526 6677 17535 6678
rect 17534 6651 17535 6677
rect 17526 6650 17535 6651
rect 17073 6645 17535 6650
rect 17318 6481 17346 6487
rect 17318 6455 17319 6481
rect 17345 6455 17346 6481
rect 17318 6425 17346 6455
rect 17318 6399 17319 6425
rect 17345 6399 17346 6425
rect 17318 6090 17346 6399
rect 17598 6090 17626 6846
rect 17766 6145 17794 6151
rect 17766 6119 17767 6145
rect 17793 6119 17794 6145
rect 17710 6090 17738 6095
rect 17766 6090 17794 6119
rect 17318 6089 17794 6090
rect 17318 6063 17711 6089
rect 17737 6063 17794 6089
rect 17318 6062 17794 6063
rect 17073 5894 17535 5899
rect 16870 5866 17010 5894
rect 15862 5671 15863 5697
rect 15889 5671 15890 5697
rect 15862 5642 15890 5671
rect 16814 5697 16842 5838
rect 16814 5671 16815 5697
rect 16841 5671 16842 5697
rect 16030 5642 16058 5647
rect 15862 5641 16058 5642
rect 15862 5615 16031 5641
rect 16057 5615 16058 5641
rect 15862 5614 16058 5615
rect 15862 5361 15890 5614
rect 16030 5609 16058 5614
rect 15862 5335 15863 5361
rect 15889 5335 15890 5361
rect 15862 5305 15890 5335
rect 15862 5279 15863 5305
rect 15889 5279 15890 5305
rect 15862 5273 15890 5279
rect 16814 5305 16842 5671
rect 16982 5362 17010 5866
rect 17073 5893 17082 5894
rect 17073 5867 17074 5893
rect 17073 5866 17082 5867
rect 17110 5866 17134 5894
rect 17162 5866 17186 5894
rect 17214 5893 17238 5894
rect 17266 5893 17290 5894
rect 17224 5867 17238 5893
rect 17286 5867 17290 5893
rect 17214 5866 17238 5867
rect 17266 5866 17290 5867
rect 17318 5893 17342 5894
rect 17370 5893 17394 5894
rect 17318 5867 17322 5893
rect 17370 5867 17384 5893
rect 17318 5866 17342 5867
rect 17370 5866 17394 5867
rect 17422 5866 17446 5894
rect 17474 5866 17498 5894
rect 17526 5893 17535 5894
rect 17534 5867 17535 5893
rect 17526 5866 17535 5867
rect 17073 5861 17535 5866
rect 17710 5697 17738 6062
rect 17710 5671 17711 5697
rect 17737 5671 17738 5697
rect 17710 5642 17738 5671
rect 17710 5641 17794 5642
rect 17710 5615 17711 5641
rect 17737 5615 17794 5641
rect 17710 5614 17794 5615
rect 17710 5609 17738 5614
rect 16982 5329 17010 5334
rect 17766 5361 17794 5614
rect 17766 5335 17767 5361
rect 17793 5335 17794 5361
rect 16814 5279 16815 5305
rect 16841 5279 16842 5305
rect 15414 4606 15554 4634
rect 15582 4913 15610 4919
rect 15806 4914 15834 4919
rect 16030 4914 16058 4919
rect 15582 4887 15583 4913
rect 15609 4887 15610 4913
rect 14238 4522 14266 4527
rect 14126 4521 14266 4522
rect 14126 4495 14127 4521
rect 14153 4495 14239 4521
rect 14265 4495 14266 4521
rect 14126 4494 14266 4495
rect 14126 4489 14154 4494
rect 14238 4129 14266 4494
rect 14238 4103 14239 4129
rect 14265 4103 14266 4129
rect 14238 4073 14266 4103
rect 14238 4047 14239 4073
rect 14265 4047 14266 4073
rect 13678 3738 13706 3743
rect 13594 3737 13706 3738
rect 13594 3711 13679 3737
rect 13705 3711 13706 3737
rect 13594 3710 13706 3711
rect 13566 3672 13594 3710
rect 13678 3705 13706 3710
rect 14126 3738 14154 3743
rect 13342 3345 13370 3374
rect 13342 3319 13343 3345
rect 13369 3319 13370 3345
rect 13342 2953 13370 3319
rect 13678 3346 13706 3351
rect 13678 3299 13706 3318
rect 13902 3346 13930 3351
rect 13902 3299 13930 3318
rect 14126 3346 14154 3710
rect 14126 3313 14154 3318
rect 14238 3009 14266 4047
rect 15134 4521 15162 4527
rect 15134 4495 15135 4521
rect 15161 4495 15162 4521
rect 14573 3934 15035 3939
rect 14573 3933 14582 3934
rect 14573 3907 14574 3933
rect 14573 3906 14582 3907
rect 14610 3906 14634 3934
rect 14662 3906 14686 3934
rect 14714 3933 14738 3934
rect 14766 3933 14790 3934
rect 14724 3907 14738 3933
rect 14786 3907 14790 3933
rect 14714 3906 14738 3907
rect 14766 3906 14790 3907
rect 14818 3933 14842 3934
rect 14870 3933 14894 3934
rect 14818 3907 14822 3933
rect 14870 3907 14884 3933
rect 14818 3906 14842 3907
rect 14870 3906 14894 3907
rect 14922 3906 14946 3934
rect 14974 3906 14998 3934
rect 15026 3933 15035 3934
rect 15034 3907 15035 3933
rect 15026 3906 15035 3907
rect 14573 3901 15035 3906
rect 14350 3738 14378 3743
rect 14350 3691 14378 3710
rect 15134 3737 15162 4495
rect 15134 3711 15135 3737
rect 15161 3711 15162 3737
rect 15134 3346 15162 3711
rect 14573 3150 15035 3155
rect 14573 3149 14582 3150
rect 14573 3123 14574 3149
rect 14573 3122 14582 3123
rect 14610 3122 14634 3150
rect 14662 3122 14686 3150
rect 14714 3149 14738 3150
rect 14766 3149 14790 3150
rect 14724 3123 14738 3149
rect 14786 3123 14790 3149
rect 14714 3122 14738 3123
rect 14766 3122 14790 3123
rect 14818 3149 14842 3150
rect 14870 3149 14894 3150
rect 14818 3123 14822 3149
rect 14870 3123 14884 3149
rect 14818 3122 14842 3123
rect 14870 3122 14894 3123
rect 14922 3122 14946 3150
rect 14974 3122 14998 3150
rect 15026 3149 15035 3150
rect 15034 3123 15035 3149
rect 15026 3122 15035 3123
rect 14573 3117 15035 3122
rect 14238 2983 14239 3009
rect 14265 2983 14266 3009
rect 13342 2927 13343 2953
rect 13369 2927 13370 2953
rect 13342 2561 13370 2927
rect 13342 2535 13343 2561
rect 13369 2535 13370 2561
rect 13342 2170 13370 2535
rect 14126 2954 14154 2959
rect 13342 1777 13370 2142
rect 13342 1751 13343 1777
rect 13369 1751 13370 1777
rect 13342 1745 13370 1751
rect 13510 2226 13538 2231
rect 13510 1778 13538 2198
rect 14070 2226 14098 2231
rect 13622 2170 13650 2175
rect 13622 2123 13650 2142
rect 14070 2169 14098 2198
rect 14070 2143 14071 2169
rect 14097 2143 14098 2169
rect 14070 2137 14098 2143
rect 13734 1778 13762 1783
rect 13510 1777 13762 1778
rect 13510 1751 13511 1777
rect 13537 1751 13735 1777
rect 13761 1751 13762 1777
rect 13510 1750 13762 1751
rect 13510 1745 13538 1750
rect 13734 1745 13762 1750
rect 14126 400 14154 2926
rect 14238 2953 14266 2983
rect 14238 2927 14239 2953
rect 14265 2927 14266 2953
rect 14238 2618 14266 2927
rect 15078 2954 15106 2959
rect 15134 2954 15162 3318
rect 15078 2953 15162 2954
rect 15078 2927 15079 2953
rect 15105 2927 15162 2953
rect 15078 2926 15162 2927
rect 15078 2921 15106 2926
rect 14238 2561 14266 2590
rect 14238 2535 14239 2561
rect 14265 2535 14266 2561
rect 14238 2505 14266 2535
rect 14238 2479 14239 2505
rect 14265 2479 14266 2505
rect 14238 2473 14266 2479
rect 15134 2562 15162 2926
rect 15246 3290 15274 3295
rect 15246 2954 15274 3262
rect 15246 2953 15330 2954
rect 15246 2927 15247 2953
rect 15273 2927 15330 2953
rect 15246 2926 15330 2927
rect 15246 2921 15274 2926
rect 15302 2898 15330 2926
rect 15246 2562 15274 2567
rect 15134 2561 15274 2562
rect 15134 2535 15247 2561
rect 15273 2535 15274 2561
rect 15134 2534 15274 2535
rect 14573 2366 15035 2371
rect 14573 2365 14582 2366
rect 14573 2339 14574 2365
rect 14573 2338 14582 2339
rect 14610 2338 14634 2366
rect 14662 2338 14686 2366
rect 14714 2365 14738 2366
rect 14766 2365 14790 2366
rect 14724 2339 14738 2365
rect 14786 2339 14790 2365
rect 14714 2338 14738 2339
rect 14766 2338 14790 2339
rect 14818 2365 14842 2366
rect 14870 2365 14894 2366
rect 14818 2339 14822 2365
rect 14870 2339 14884 2365
rect 14818 2338 14842 2339
rect 14870 2338 14894 2339
rect 14922 2338 14946 2366
rect 14974 2338 14998 2366
rect 15026 2365 15035 2366
rect 15034 2339 15035 2365
rect 15026 2338 15035 2339
rect 14573 2333 15035 2338
rect 14294 2226 14322 2231
rect 14294 2169 14322 2198
rect 14294 2143 14295 2169
rect 14321 2143 14322 2169
rect 14294 2137 14322 2143
rect 15134 2170 15162 2534
rect 15246 2506 15274 2534
rect 15246 2473 15274 2478
rect 15134 1777 15162 2142
rect 15134 1751 15135 1777
rect 15161 1751 15162 1777
rect 15134 1745 15162 1751
rect 15302 1834 15330 2870
rect 15302 1777 15330 1806
rect 15302 1751 15303 1777
rect 15329 1751 15330 1777
rect 15302 1745 15330 1751
rect 15414 1694 15442 4606
rect 15470 4522 15498 4527
rect 15470 3738 15498 4494
rect 15470 2953 15498 3710
rect 15526 4130 15554 4135
rect 15582 4130 15610 4887
rect 15694 4913 16058 4914
rect 15694 4887 15807 4913
rect 15833 4887 16031 4913
rect 16057 4887 16058 4913
rect 15694 4886 16058 4887
rect 15694 4522 15722 4886
rect 15806 4881 15834 4886
rect 16030 4881 16058 4886
rect 16814 4913 16842 5279
rect 17766 5305 17794 5335
rect 17766 5279 17767 5305
rect 17793 5279 17794 5305
rect 17073 5110 17535 5115
rect 17073 5109 17082 5110
rect 17073 5083 17074 5109
rect 17073 5082 17082 5083
rect 17110 5082 17134 5110
rect 17162 5082 17186 5110
rect 17214 5109 17238 5110
rect 17266 5109 17290 5110
rect 17224 5083 17238 5109
rect 17286 5083 17290 5109
rect 17214 5082 17238 5083
rect 17266 5082 17290 5083
rect 17318 5109 17342 5110
rect 17370 5109 17394 5110
rect 17318 5083 17322 5109
rect 17370 5083 17384 5109
rect 17318 5082 17342 5083
rect 17370 5082 17394 5083
rect 17422 5082 17446 5110
rect 17474 5082 17498 5110
rect 17526 5109 17535 5110
rect 17534 5083 17535 5109
rect 17526 5082 17535 5083
rect 17073 5077 17535 5082
rect 16814 4887 16815 4913
rect 16841 4887 16842 4913
rect 15694 4475 15722 4494
rect 16814 4521 16842 4887
rect 16814 4495 16815 4521
rect 16841 4495 16842 4521
rect 15526 4129 15610 4130
rect 15526 4103 15527 4129
rect 15553 4103 15610 4129
rect 15526 4102 15610 4103
rect 15806 4129 15834 4135
rect 15806 4103 15807 4129
rect 15833 4103 15834 4129
rect 15526 3346 15554 4102
rect 15582 3738 15610 3743
rect 15582 3691 15610 3710
rect 15806 3738 15834 4103
rect 16030 4129 16058 4135
rect 16030 4103 16031 4129
rect 16057 4103 16058 4129
rect 15806 3691 15834 3710
rect 15974 3738 16002 3743
rect 16030 3738 16058 4103
rect 16002 3710 16058 3738
rect 16814 4129 16842 4495
rect 17766 4913 17794 5279
rect 17766 4887 17767 4913
rect 17793 4887 17794 4913
rect 17766 4857 17794 4887
rect 17766 4831 17767 4857
rect 17793 4831 17794 4857
rect 17766 4577 17794 4831
rect 18214 4690 18242 9142
rect 18270 8833 18298 9199
rect 18270 8807 18271 8833
rect 18297 8807 18298 8833
rect 18270 8777 18298 8807
rect 18270 8751 18271 8777
rect 18297 8751 18298 8777
rect 18270 8497 18298 8751
rect 18270 8471 18271 8497
rect 18297 8471 18298 8497
rect 18270 8441 18298 8471
rect 18270 8415 18271 8441
rect 18297 8415 18298 8441
rect 18270 8409 18298 8415
rect 18774 9225 18802 9478
rect 18774 9199 18775 9225
rect 18801 9199 18802 9225
rect 18774 8834 18802 9199
rect 18774 8441 18802 8806
rect 18774 8415 18775 8441
rect 18801 8415 18802 8441
rect 18774 8049 18802 8415
rect 18774 8023 18775 8049
rect 18801 8023 18802 8049
rect 18550 7657 18578 7663
rect 18550 7631 18551 7657
rect 18577 7631 18578 7657
rect 18550 7574 18578 7631
rect 18774 7574 18802 8023
rect 18550 7546 18802 7574
rect 18774 7265 18802 7546
rect 18774 7239 18775 7265
rect 18801 7239 18802 7265
rect 18214 4657 18242 4662
rect 18550 6873 18578 6879
rect 18550 6847 18551 6873
rect 18577 6847 18578 6873
rect 18550 6089 18578 6847
rect 18550 6063 18551 6089
rect 18577 6063 18578 6089
rect 18550 5305 18578 6063
rect 18550 5279 18551 5305
rect 18577 5279 18578 5305
rect 17766 4551 17767 4577
rect 17793 4551 17794 4577
rect 17766 4521 17794 4551
rect 17766 4495 17767 4521
rect 17793 4495 17794 4521
rect 17073 4326 17535 4331
rect 17073 4325 17082 4326
rect 17073 4299 17074 4325
rect 17073 4298 17082 4299
rect 17110 4298 17134 4326
rect 17162 4298 17186 4326
rect 17214 4325 17238 4326
rect 17266 4325 17290 4326
rect 17224 4299 17238 4325
rect 17286 4299 17290 4325
rect 17214 4298 17238 4299
rect 17266 4298 17290 4299
rect 17318 4325 17342 4326
rect 17370 4325 17394 4326
rect 17318 4299 17322 4325
rect 17370 4299 17384 4325
rect 17318 4298 17342 4299
rect 17370 4298 17394 4299
rect 17422 4298 17446 4326
rect 17474 4298 17498 4326
rect 17526 4325 17535 4326
rect 17534 4299 17535 4325
rect 17526 4298 17535 4299
rect 17073 4293 17535 4298
rect 16814 4103 16815 4129
rect 16841 4103 16842 4129
rect 16814 3737 16842 4103
rect 16814 3711 16815 3737
rect 16841 3711 16842 3737
rect 15526 3299 15554 3318
rect 15974 3346 16002 3710
rect 16198 3346 16226 3351
rect 15974 3345 16226 3346
rect 15974 3319 15975 3345
rect 16001 3319 16199 3345
rect 16225 3319 16226 3345
rect 15974 3318 16226 3319
rect 15974 3313 16002 3318
rect 16198 3313 16226 3318
rect 16814 3346 16842 3711
rect 17766 4129 17794 4495
rect 17766 4103 17767 4129
rect 17793 4103 17794 4129
rect 17766 4073 17794 4103
rect 17766 4047 17767 4073
rect 17793 4047 17794 4073
rect 17766 3793 17794 4047
rect 17766 3767 17767 3793
rect 17793 3767 17794 3793
rect 17766 3737 17794 3767
rect 17766 3711 17767 3737
rect 17793 3711 17794 3737
rect 17073 3542 17535 3547
rect 17073 3541 17082 3542
rect 17073 3515 17074 3541
rect 17073 3514 17082 3515
rect 17110 3514 17134 3542
rect 17162 3514 17186 3542
rect 17214 3541 17238 3542
rect 17266 3541 17290 3542
rect 17224 3515 17238 3541
rect 17286 3515 17290 3541
rect 17214 3514 17238 3515
rect 17266 3514 17290 3515
rect 17318 3541 17342 3542
rect 17370 3541 17394 3542
rect 17318 3515 17322 3541
rect 17370 3515 17384 3541
rect 17318 3514 17342 3515
rect 17370 3514 17394 3515
rect 17422 3514 17446 3542
rect 17474 3514 17498 3542
rect 17526 3541 17535 3542
rect 17534 3515 17535 3541
rect 17526 3514 17535 3515
rect 17073 3509 17535 3514
rect 16982 3346 17010 3351
rect 16814 3345 17010 3346
rect 16814 3319 16983 3345
rect 17009 3319 17010 3345
rect 16814 3318 17010 3319
rect 15470 2927 15471 2953
rect 15497 2927 15498 2953
rect 15470 2898 15498 2927
rect 15470 2865 15498 2870
rect 16814 2953 16842 3318
rect 16982 3313 17010 3318
rect 17766 3345 17794 3711
rect 17990 4634 18018 4639
rect 17766 3319 17767 3345
rect 17793 3319 17794 3345
rect 17766 3290 17794 3319
rect 17934 3346 17962 3351
rect 17934 3290 17962 3318
rect 17766 3289 17962 3290
rect 17766 3263 17935 3289
rect 17961 3263 17962 3289
rect 17766 3262 17962 3263
rect 17766 3009 17794 3262
rect 17934 3257 17962 3262
rect 17766 2983 17767 3009
rect 17793 2983 17794 3009
rect 16814 2927 16815 2953
rect 16841 2927 16842 2953
rect 15694 2562 15722 2567
rect 15918 2562 15946 2567
rect 15694 2561 15918 2562
rect 15694 2535 15695 2561
rect 15721 2535 15918 2561
rect 15694 2534 15918 2535
rect 15582 2170 15610 2175
rect 15694 2170 15722 2534
rect 15918 2496 15946 2534
rect 16814 2561 16842 2927
rect 17654 2954 17682 2959
rect 17766 2954 17794 2983
rect 17654 2953 17794 2954
rect 17654 2927 17655 2953
rect 17681 2927 17794 2953
rect 17654 2926 17794 2927
rect 17073 2758 17535 2763
rect 17073 2757 17082 2758
rect 17073 2731 17074 2757
rect 17073 2730 17082 2731
rect 17110 2730 17134 2758
rect 17162 2730 17186 2758
rect 17214 2757 17238 2758
rect 17266 2757 17290 2758
rect 17224 2731 17238 2757
rect 17286 2731 17290 2757
rect 17214 2730 17238 2731
rect 17266 2730 17290 2731
rect 17318 2757 17342 2758
rect 17370 2757 17394 2758
rect 17318 2731 17322 2757
rect 17370 2731 17384 2757
rect 17318 2730 17342 2731
rect 17370 2730 17394 2731
rect 17422 2730 17446 2758
rect 17474 2730 17498 2758
rect 17526 2757 17535 2758
rect 17534 2731 17535 2757
rect 17526 2730 17535 2731
rect 17073 2725 17535 2730
rect 17598 2618 17626 2623
rect 16814 2535 16815 2561
rect 16841 2535 16842 2561
rect 16814 2506 16842 2535
rect 17150 2562 17178 2567
rect 17150 2515 17178 2534
rect 17374 2562 17402 2567
rect 17374 2515 17402 2534
rect 15806 2170 15834 2175
rect 15526 2169 15834 2170
rect 15526 2143 15583 2169
rect 15609 2143 15807 2169
rect 15833 2143 15834 2169
rect 15526 2142 15834 2143
rect 15526 1834 15554 2142
rect 15582 2137 15610 2142
rect 15806 2137 15834 2142
rect 16590 2170 16618 2175
rect 15526 1777 15554 1806
rect 15526 1751 15527 1777
rect 15553 1751 15554 1777
rect 15526 1745 15554 1751
rect 16590 1890 16618 2142
rect 16814 2169 16842 2478
rect 16814 2143 16815 2169
rect 16841 2143 16842 2169
rect 16814 2137 16842 2143
rect 17073 1974 17535 1979
rect 17073 1973 17082 1974
rect 17073 1947 17074 1973
rect 17073 1946 17082 1947
rect 17110 1946 17134 1974
rect 17162 1946 17186 1974
rect 17214 1973 17238 1974
rect 17266 1973 17290 1974
rect 17224 1947 17238 1973
rect 17286 1947 17290 1973
rect 17214 1946 17238 1947
rect 17266 1946 17290 1947
rect 17318 1973 17342 1974
rect 17370 1973 17394 1974
rect 17318 1947 17322 1973
rect 17370 1947 17384 1973
rect 17318 1946 17342 1947
rect 17370 1946 17394 1947
rect 17422 1946 17446 1974
rect 17474 1946 17498 1974
rect 17526 1973 17535 1974
rect 17534 1947 17535 1973
rect 17526 1946 17535 1947
rect 17073 1941 17535 1946
rect 16590 1777 16618 1862
rect 16590 1751 16591 1777
rect 16617 1751 16618 1777
rect 16590 1745 16618 1751
rect 17038 1890 17066 1895
rect 15414 1666 15498 1694
rect 14573 1582 15035 1587
rect 14573 1581 14582 1582
rect 14573 1555 14574 1581
rect 14573 1554 14582 1555
rect 14610 1554 14634 1582
rect 14662 1554 14686 1582
rect 14714 1581 14738 1582
rect 14766 1581 14790 1582
rect 14724 1555 14738 1581
rect 14786 1555 14790 1581
rect 14714 1554 14738 1555
rect 14766 1554 14790 1555
rect 14818 1581 14842 1582
rect 14870 1581 14894 1582
rect 14818 1555 14822 1581
rect 14870 1555 14884 1581
rect 14818 1554 14842 1555
rect 14870 1554 14894 1555
rect 14922 1554 14946 1582
rect 14974 1554 14998 1582
rect 15026 1581 15035 1582
rect 15034 1555 15035 1581
rect 15026 1554 15035 1555
rect 14573 1549 15035 1554
rect 15470 490 15498 1666
rect 15470 462 15610 490
rect 15582 400 15610 462
rect 17038 400 17066 1862
rect 17542 1778 17570 1783
rect 17598 1778 17626 2590
rect 17654 2562 17682 2926
rect 17654 2226 17682 2534
rect 17766 2226 17794 2231
rect 17654 2225 17794 2226
rect 17654 2199 17767 2225
rect 17793 2199 17794 2225
rect 17654 2198 17794 2199
rect 17654 2169 17682 2198
rect 17766 2193 17794 2198
rect 17654 2143 17655 2169
rect 17681 2143 17682 2169
rect 17654 2137 17682 2143
rect 17990 1890 18018 4606
rect 18550 4521 18578 5279
rect 18550 4495 18551 4521
rect 18577 4495 18578 4521
rect 18550 4130 18578 4495
rect 18774 6481 18802 7239
rect 18774 6455 18775 6481
rect 18801 6455 18802 6481
rect 18774 5697 18802 6455
rect 18774 5671 18775 5697
rect 18801 5671 18802 5697
rect 18774 5082 18802 5671
rect 18774 4913 18802 5054
rect 18774 4887 18775 4913
rect 18801 4887 18802 4913
rect 18774 4130 18802 4887
rect 18550 4129 18802 4130
rect 18550 4103 18775 4129
rect 18801 4103 18802 4129
rect 18550 4102 18802 4103
rect 18550 3737 18578 4102
rect 18774 4097 18802 4102
rect 18550 3711 18551 3737
rect 18577 3711 18578 3737
rect 18550 3705 18578 3711
rect 18494 3402 18522 3407
rect 18270 2953 18298 2959
rect 18270 2927 18271 2953
rect 18297 2927 18298 2953
rect 18270 2170 18298 2927
rect 18270 2123 18298 2142
rect 17990 1857 18018 1862
rect 17542 1777 17626 1778
rect 17542 1751 17543 1777
rect 17569 1751 17626 1777
rect 17542 1750 17626 1751
rect 17542 1721 17570 1750
rect 17542 1695 17543 1721
rect 17569 1695 17570 1721
rect 17542 1689 17570 1695
rect 18494 1498 18522 3374
rect 18774 3345 18802 3351
rect 18774 3319 18775 3345
rect 18801 3319 18802 3345
rect 18774 2506 18802 3319
rect 18886 2954 18914 11214
rect 19334 11186 19362 11551
rect 19502 11186 19530 11191
rect 19334 11185 19530 11186
rect 19334 11159 19335 11185
rect 19361 11159 19503 11185
rect 19529 11159 19530 11185
rect 19334 11158 19530 11159
rect 19334 11153 19362 11158
rect 19446 10850 19474 10855
rect 19502 10850 19530 11158
rect 20510 11185 20538 11943
rect 20958 13929 20986 13935
rect 20958 13903 20959 13929
rect 20985 13903 20986 13929
rect 20958 13145 20986 13903
rect 21014 13538 21042 14294
rect 22526 14322 22554 14327
rect 22582 14322 22610 14630
rect 22554 14294 22610 14322
rect 23030 15105 23058 15111
rect 23030 15079 23031 15105
rect 23057 15079 23058 15105
rect 23030 14322 23058 15079
rect 23422 14769 23450 15471
rect 23422 14743 23423 14769
rect 23449 14743 23450 14769
rect 23422 14714 23450 14743
rect 23422 14667 23450 14686
rect 23926 15105 23954 15111
rect 23926 15079 23927 15105
rect 23953 15079 23954 15105
rect 23926 15049 23954 15079
rect 23926 15023 23927 15049
rect 23953 15023 23954 15049
rect 23926 14714 23954 15023
rect 21238 13930 21266 13935
rect 21462 13930 21490 13935
rect 21182 13929 21462 13930
rect 21182 13903 21239 13929
rect 21265 13903 21462 13929
rect 21182 13902 21462 13903
rect 21182 13538 21210 13902
rect 21238 13897 21266 13902
rect 21462 13864 21490 13902
rect 22526 13929 22554 14294
rect 22526 13903 22527 13929
rect 22553 13903 22554 13929
rect 22526 13897 22554 13903
rect 22073 13734 22535 13739
rect 22073 13733 22082 13734
rect 22073 13707 22074 13733
rect 22073 13706 22082 13707
rect 22110 13706 22134 13734
rect 22162 13706 22186 13734
rect 22214 13733 22238 13734
rect 22266 13733 22290 13734
rect 22224 13707 22238 13733
rect 22286 13707 22290 13733
rect 22214 13706 22238 13707
rect 22266 13706 22290 13707
rect 22318 13733 22342 13734
rect 22370 13733 22394 13734
rect 22318 13707 22322 13733
rect 22370 13707 22384 13733
rect 22318 13706 22342 13707
rect 22370 13706 22394 13707
rect 22422 13706 22446 13734
rect 22474 13706 22498 13734
rect 22526 13733 22535 13734
rect 22534 13707 22535 13733
rect 22526 13706 22535 13707
rect 22073 13701 22535 13706
rect 21014 13537 21210 13538
rect 21014 13511 21015 13537
rect 21041 13511 21210 13537
rect 21014 13510 21210 13511
rect 21014 13505 21042 13510
rect 20958 13119 20959 13145
rect 20985 13119 20986 13145
rect 20958 12642 20986 13119
rect 20958 12361 20986 12614
rect 20958 12335 20959 12361
rect 20985 12335 20986 12361
rect 20958 11577 20986 12335
rect 21182 13481 21210 13510
rect 23030 13537 23058 14294
rect 23926 14321 23954 14686
rect 23926 14295 23927 14321
rect 23953 14295 23954 14321
rect 23926 14266 23954 14295
rect 23926 14219 23954 14238
rect 23030 13511 23031 13537
rect 23057 13511 23058 13537
rect 23030 13505 23058 13511
rect 23422 13985 23450 13991
rect 23422 13959 23423 13985
rect 23449 13959 23450 13985
rect 23422 13930 23450 13959
rect 21182 13455 21183 13481
rect 21209 13455 21210 13481
rect 21182 13146 21210 13455
rect 23422 13482 23450 13902
rect 23422 13201 23450 13454
rect 23926 13537 23954 13543
rect 23926 13511 23927 13537
rect 23953 13511 23954 13537
rect 23926 13482 23954 13511
rect 23926 13435 23954 13454
rect 23422 13175 23423 13201
rect 23449 13175 23450 13201
rect 21238 13146 21266 13151
rect 21462 13146 21490 13151
rect 21182 13145 21490 13146
rect 21182 13119 21239 13145
rect 21265 13119 21463 13145
rect 21489 13119 21490 13145
rect 21182 13118 21490 13119
rect 21182 12753 21210 13118
rect 21238 13113 21266 13118
rect 21462 13113 21490 13118
rect 22526 13146 22554 13151
rect 22526 13145 22610 13146
rect 22526 13119 22527 13145
rect 22553 13119 22610 13145
rect 22526 13118 22610 13119
rect 22526 13113 22554 13118
rect 22073 12950 22535 12955
rect 22073 12949 22082 12950
rect 22073 12923 22074 12949
rect 22073 12922 22082 12923
rect 22110 12922 22134 12950
rect 22162 12922 22186 12950
rect 22214 12949 22238 12950
rect 22266 12949 22290 12950
rect 22224 12923 22238 12949
rect 22286 12923 22290 12949
rect 22214 12922 22238 12923
rect 22266 12922 22290 12923
rect 22318 12949 22342 12950
rect 22370 12949 22394 12950
rect 22318 12923 22322 12949
rect 22370 12923 22384 12949
rect 22318 12922 22342 12923
rect 22370 12922 22394 12923
rect 22422 12922 22446 12950
rect 22474 12922 22498 12950
rect 22526 12949 22535 12950
rect 22534 12923 22535 12949
rect 22526 12922 22535 12923
rect 22073 12917 22535 12922
rect 22582 12754 22610 13118
rect 23422 13145 23450 13175
rect 23422 13119 23423 13145
rect 23449 13119 23450 13145
rect 22750 12754 22778 12759
rect 21182 12727 21183 12753
rect 21209 12727 21210 12753
rect 21182 12697 21210 12727
rect 21182 12671 21183 12697
rect 21209 12671 21210 12697
rect 21182 12362 21210 12671
rect 22526 12753 22778 12754
rect 22526 12727 22751 12753
rect 22777 12727 22778 12753
rect 22526 12726 22778 12727
rect 22526 12642 22554 12726
rect 22750 12721 22778 12726
rect 23310 12754 23338 12759
rect 23422 12754 23450 13119
rect 23310 12753 23450 12754
rect 23310 12727 23311 12753
rect 23337 12727 23423 12753
rect 23449 12727 23450 12753
rect 23310 12726 23450 12727
rect 23310 12721 23338 12726
rect 21238 12362 21266 12367
rect 21462 12362 21490 12367
rect 21182 12361 21490 12362
rect 21182 12335 21239 12361
rect 21265 12335 21463 12361
rect 21489 12335 21490 12361
rect 21182 12334 21490 12335
rect 21238 12329 21266 12334
rect 21462 12329 21490 12334
rect 22526 12361 22554 12614
rect 22526 12335 22527 12361
rect 22553 12335 22554 12361
rect 22526 12329 22554 12335
rect 23422 12417 23450 12726
rect 23422 12391 23423 12417
rect 23449 12391 23450 12417
rect 23422 12361 23450 12391
rect 23422 12335 23423 12361
rect 23449 12335 23450 12361
rect 23422 12329 23450 12335
rect 22073 12166 22535 12171
rect 22073 12165 22082 12166
rect 22073 12139 22074 12165
rect 22073 12138 22082 12139
rect 22110 12138 22134 12166
rect 22162 12138 22186 12166
rect 22214 12165 22238 12166
rect 22266 12165 22290 12166
rect 22224 12139 22238 12165
rect 22286 12139 22290 12165
rect 22214 12138 22238 12139
rect 22266 12138 22290 12139
rect 22318 12165 22342 12166
rect 22370 12165 22394 12166
rect 22318 12139 22322 12165
rect 22370 12139 22384 12165
rect 22318 12138 22342 12139
rect 22370 12138 22394 12139
rect 22422 12138 22446 12166
rect 22474 12138 22498 12166
rect 22526 12165 22535 12166
rect 22534 12139 22535 12165
rect 22526 12138 22535 12139
rect 22073 12133 22535 12138
rect 20958 11551 20959 11577
rect 20985 11551 20986 11577
rect 20958 11545 20986 11551
rect 21182 11970 21210 11975
rect 21182 11913 21210 11942
rect 21182 11887 21183 11913
rect 21209 11887 21210 11913
rect 21182 11578 21210 11887
rect 22806 11969 22834 11975
rect 22806 11943 22807 11969
rect 22833 11943 22834 11969
rect 21238 11578 21266 11583
rect 21462 11578 21490 11583
rect 21182 11577 21490 11578
rect 21182 11551 21239 11577
rect 21265 11551 21463 11577
rect 21489 11551 21490 11577
rect 21182 11550 21490 11551
rect 20510 11159 20511 11185
rect 20537 11159 20538 11185
rect 20510 11153 20538 11159
rect 21014 11185 21042 11191
rect 21014 11159 21015 11185
rect 21041 11159 21042 11185
rect 21014 11130 21042 11159
rect 21182 11130 21210 11550
rect 21238 11545 21266 11550
rect 21462 11545 21490 11550
rect 22526 11578 22554 11583
rect 22526 11577 22610 11578
rect 22526 11551 22527 11577
rect 22553 11551 22610 11577
rect 22526 11550 22610 11551
rect 22526 11545 22554 11550
rect 22073 11382 22535 11387
rect 22073 11381 22082 11382
rect 22073 11355 22074 11381
rect 22073 11354 22082 11355
rect 22110 11354 22134 11382
rect 22162 11354 22186 11382
rect 22214 11381 22238 11382
rect 22266 11381 22290 11382
rect 22224 11355 22238 11381
rect 22286 11355 22290 11381
rect 22214 11354 22238 11355
rect 22266 11354 22290 11355
rect 22318 11381 22342 11382
rect 22370 11381 22394 11382
rect 22318 11355 22322 11381
rect 22370 11355 22384 11381
rect 22318 11354 22342 11355
rect 22370 11354 22394 11355
rect 22422 11354 22446 11382
rect 22474 11354 22498 11382
rect 22526 11381 22535 11382
rect 22534 11355 22535 11381
rect 22526 11354 22535 11355
rect 22073 11349 22535 11354
rect 21014 11129 21210 11130
rect 21014 11103 21183 11129
rect 21209 11103 21210 11129
rect 21014 11102 21210 11103
rect 19573 10990 20035 10995
rect 19573 10989 19582 10990
rect 19573 10963 19574 10989
rect 19573 10962 19582 10963
rect 19610 10962 19634 10990
rect 19662 10962 19686 10990
rect 19714 10989 19738 10990
rect 19766 10989 19790 10990
rect 19724 10963 19738 10989
rect 19786 10963 19790 10989
rect 19714 10962 19738 10963
rect 19766 10962 19790 10963
rect 19818 10989 19842 10990
rect 19870 10989 19894 10990
rect 19818 10963 19822 10989
rect 19870 10963 19884 10989
rect 19818 10962 19842 10963
rect 19870 10962 19894 10963
rect 19922 10962 19946 10990
rect 19974 10962 19998 10990
rect 20026 10989 20035 10990
rect 20034 10963 20035 10989
rect 20026 10962 20035 10963
rect 19573 10957 20035 10962
rect 19446 10849 19530 10850
rect 19446 10823 19447 10849
rect 19473 10823 19530 10849
rect 19446 10822 19530 10823
rect 19446 10793 19474 10822
rect 19446 10767 19447 10793
rect 19473 10767 19474 10793
rect 19446 10761 19474 10767
rect 19502 10346 19530 10822
rect 20790 10793 20818 10799
rect 20790 10767 20791 10793
rect 20817 10767 20818 10793
rect 19502 10313 19530 10318
rect 19950 10401 19978 10407
rect 19950 10375 19951 10401
rect 19977 10375 19978 10401
rect 19950 10346 19978 10375
rect 19950 10299 19978 10318
rect 20230 10401 20258 10407
rect 20230 10375 20231 10401
rect 20257 10375 20258 10401
rect 19573 10206 20035 10211
rect 19573 10205 19582 10206
rect 19573 10179 19574 10205
rect 19573 10178 19582 10179
rect 19610 10178 19634 10206
rect 19662 10178 19686 10206
rect 19714 10205 19738 10206
rect 19766 10205 19790 10206
rect 19724 10179 19738 10205
rect 19786 10179 19790 10205
rect 19714 10178 19738 10179
rect 19766 10178 19790 10179
rect 19818 10205 19842 10206
rect 19870 10205 19894 10206
rect 19818 10179 19822 10205
rect 19870 10179 19884 10205
rect 19818 10178 19842 10179
rect 19870 10178 19894 10179
rect 19922 10178 19946 10206
rect 19974 10178 19998 10206
rect 20026 10205 20035 10206
rect 20034 10179 20035 10205
rect 20026 10178 20035 10179
rect 19573 10173 20035 10178
rect 18942 10010 18970 10015
rect 18942 9963 18970 9982
rect 19222 9618 19250 9623
rect 19446 9618 19474 9623
rect 19250 9617 19474 9618
rect 19250 9591 19447 9617
rect 19473 9591 19474 9617
rect 19250 9590 19474 9591
rect 19222 9226 19250 9590
rect 19446 9585 19474 9590
rect 20230 9617 20258 10375
rect 20230 9591 20231 9617
rect 20257 9591 20258 9617
rect 19573 9422 20035 9427
rect 19573 9421 19582 9422
rect 19573 9395 19574 9421
rect 19573 9394 19582 9395
rect 19610 9394 19634 9422
rect 19662 9394 19686 9422
rect 19714 9421 19738 9422
rect 19766 9421 19790 9422
rect 19724 9395 19738 9421
rect 19786 9395 19790 9421
rect 19714 9394 19738 9395
rect 19766 9394 19790 9395
rect 19818 9421 19842 9422
rect 19870 9421 19894 9422
rect 19818 9395 19822 9421
rect 19870 9395 19884 9421
rect 19818 9394 19842 9395
rect 19870 9394 19894 9395
rect 19922 9394 19946 9422
rect 19974 9394 19998 9422
rect 20026 9421 20035 9422
rect 20034 9395 20035 9421
rect 20026 9394 20035 9395
rect 19573 9389 20035 9394
rect 19334 9226 19362 9231
rect 19222 9225 19362 9226
rect 19222 9199 19223 9225
rect 19249 9199 19335 9225
rect 19361 9199 19362 9225
rect 19222 9198 19362 9199
rect 19222 9193 19250 9198
rect 19334 8833 19362 9198
rect 19334 8807 19335 8833
rect 19361 8807 19362 8833
rect 19334 8442 19362 8807
rect 19502 8833 19530 8839
rect 19502 8807 19503 8833
rect 19529 8807 19530 8833
rect 19502 8497 19530 8807
rect 20230 8833 20258 9591
rect 20230 8807 20231 8833
rect 20257 8807 20258 8833
rect 19573 8638 20035 8643
rect 19573 8637 19582 8638
rect 19573 8611 19574 8637
rect 19573 8610 19582 8611
rect 19610 8610 19634 8638
rect 19662 8610 19686 8638
rect 19714 8637 19738 8638
rect 19766 8637 19790 8638
rect 19724 8611 19738 8637
rect 19786 8611 19790 8637
rect 19714 8610 19738 8611
rect 19766 8610 19790 8611
rect 19818 8637 19842 8638
rect 19870 8637 19894 8638
rect 19818 8611 19822 8637
rect 19870 8611 19884 8637
rect 19818 8610 19842 8611
rect 19870 8610 19894 8611
rect 19922 8610 19946 8638
rect 19974 8610 19998 8638
rect 20026 8637 20035 8638
rect 20034 8611 20035 8637
rect 20026 8610 20035 8611
rect 19573 8605 20035 8610
rect 19502 8471 19503 8497
rect 19529 8471 19530 8497
rect 19502 8442 19530 8471
rect 19334 8441 19530 8442
rect 19334 8415 19335 8441
rect 19361 8415 19530 8441
rect 19334 8414 19530 8415
rect 19334 8050 19362 8414
rect 19446 8050 19474 8055
rect 19334 8049 19474 8050
rect 19334 8023 19335 8049
rect 19361 8023 19447 8049
rect 19473 8023 19474 8049
rect 19334 8022 19474 8023
rect 19334 7713 19362 8022
rect 19446 8017 19474 8022
rect 20230 8049 20258 8807
rect 20230 8023 20231 8049
rect 20257 8023 20258 8049
rect 19573 7854 20035 7859
rect 19573 7853 19582 7854
rect 19573 7827 19574 7853
rect 19573 7826 19582 7827
rect 19610 7826 19634 7854
rect 19662 7826 19686 7854
rect 19714 7853 19738 7854
rect 19766 7853 19790 7854
rect 19724 7827 19738 7853
rect 19786 7827 19790 7853
rect 19714 7826 19738 7827
rect 19766 7826 19790 7827
rect 19818 7853 19842 7854
rect 19870 7853 19894 7854
rect 19818 7827 19822 7853
rect 19870 7827 19884 7853
rect 19818 7826 19842 7827
rect 19870 7826 19894 7827
rect 19922 7826 19946 7854
rect 19974 7826 19998 7854
rect 20026 7853 20035 7854
rect 20034 7827 20035 7853
rect 20026 7826 20035 7827
rect 19573 7821 20035 7826
rect 19334 7687 19335 7713
rect 19361 7687 19362 7713
rect 19334 7657 19362 7687
rect 19334 7631 19335 7657
rect 19361 7631 19362 7657
rect 19334 7266 19362 7631
rect 19446 7266 19474 7271
rect 19334 7265 19474 7266
rect 19334 7239 19335 7265
rect 19361 7239 19447 7265
rect 19473 7239 19474 7265
rect 19334 7238 19474 7239
rect 19334 6929 19362 7238
rect 19446 7233 19474 7238
rect 20230 7265 20258 8023
rect 20230 7239 20231 7265
rect 20257 7239 20258 7265
rect 19573 7070 20035 7075
rect 19573 7069 19582 7070
rect 19573 7043 19574 7069
rect 19573 7042 19582 7043
rect 19610 7042 19634 7070
rect 19662 7042 19686 7070
rect 19714 7069 19738 7070
rect 19766 7069 19790 7070
rect 19724 7043 19738 7069
rect 19786 7043 19790 7069
rect 19714 7042 19738 7043
rect 19766 7042 19790 7043
rect 19818 7069 19842 7070
rect 19870 7069 19894 7070
rect 19818 7043 19822 7069
rect 19870 7043 19884 7069
rect 19818 7042 19842 7043
rect 19870 7042 19894 7043
rect 19922 7042 19946 7070
rect 19974 7042 19998 7070
rect 20026 7069 20035 7070
rect 20034 7043 20035 7069
rect 20026 7042 20035 7043
rect 19573 7037 20035 7042
rect 19334 6903 19335 6929
rect 19361 6903 19362 6929
rect 19334 6873 19362 6903
rect 19334 6847 19335 6873
rect 19361 6847 19362 6873
rect 19334 6482 19362 6847
rect 19446 6482 19474 6487
rect 19334 6481 19474 6482
rect 19334 6455 19335 6481
rect 19361 6455 19447 6481
rect 19473 6455 19474 6481
rect 19334 6454 19474 6455
rect 19334 6449 19362 6454
rect 19446 6145 19474 6454
rect 20230 6481 20258 7239
rect 20230 6455 20231 6481
rect 20257 6455 20258 6481
rect 19573 6286 20035 6291
rect 19573 6285 19582 6286
rect 19573 6259 19574 6285
rect 19573 6258 19582 6259
rect 19610 6258 19634 6286
rect 19662 6258 19686 6286
rect 19714 6285 19738 6286
rect 19766 6285 19790 6286
rect 19724 6259 19738 6285
rect 19786 6259 19790 6285
rect 19714 6258 19738 6259
rect 19766 6258 19790 6259
rect 19818 6285 19842 6286
rect 19870 6285 19894 6286
rect 19818 6259 19822 6285
rect 19870 6259 19884 6285
rect 19818 6258 19842 6259
rect 19870 6258 19894 6259
rect 19922 6258 19946 6286
rect 19974 6258 19998 6286
rect 20026 6285 20035 6286
rect 20034 6259 20035 6285
rect 20026 6258 20035 6259
rect 19573 6253 20035 6258
rect 19446 6119 19447 6145
rect 19473 6119 19474 6145
rect 19446 6089 19474 6119
rect 19446 6063 19447 6089
rect 19473 6063 19474 6089
rect 19446 5361 19474 6063
rect 19950 5697 19978 5703
rect 19950 5671 19951 5697
rect 19977 5671 19978 5697
rect 19950 5642 19978 5671
rect 20230 5697 20258 6455
rect 20230 5671 20231 5697
rect 20257 5671 20258 5697
rect 19950 5641 20146 5642
rect 19950 5615 19951 5641
rect 19977 5615 20146 5641
rect 19950 5614 20146 5615
rect 19950 5609 19978 5614
rect 19573 5502 20035 5507
rect 19573 5501 19582 5502
rect 19573 5475 19574 5501
rect 19573 5474 19582 5475
rect 19610 5474 19634 5502
rect 19662 5474 19686 5502
rect 19714 5501 19738 5502
rect 19766 5501 19790 5502
rect 19724 5475 19738 5501
rect 19786 5475 19790 5501
rect 19714 5474 19738 5475
rect 19766 5474 19790 5475
rect 19818 5501 19842 5502
rect 19870 5501 19894 5502
rect 19818 5475 19822 5501
rect 19870 5475 19884 5501
rect 19818 5474 19842 5475
rect 19870 5474 19894 5475
rect 19922 5474 19946 5502
rect 19974 5474 19998 5502
rect 20026 5501 20035 5502
rect 20034 5475 20035 5501
rect 20026 5474 20035 5475
rect 19573 5469 20035 5474
rect 19446 5335 19447 5361
rect 19473 5335 19474 5361
rect 19446 5305 19474 5335
rect 19446 5279 19447 5305
rect 19473 5279 19474 5305
rect 19446 4577 19474 5279
rect 19950 4913 19978 4919
rect 19950 4887 19951 4913
rect 19977 4887 19978 4913
rect 19950 4857 19978 4887
rect 19950 4831 19951 4857
rect 19977 4831 19978 4857
rect 19950 4802 19978 4831
rect 20118 4802 20146 5614
rect 20230 5306 20258 5671
rect 20230 5082 20258 5278
rect 20230 4913 20258 5054
rect 20230 4887 20231 4913
rect 20257 4887 20258 4913
rect 20230 4881 20258 4887
rect 20566 10122 20594 10127
rect 19950 4774 20146 4802
rect 19573 4718 20035 4723
rect 19573 4717 19582 4718
rect 19573 4691 19574 4717
rect 19573 4690 19582 4691
rect 19610 4690 19634 4718
rect 19662 4690 19686 4718
rect 19714 4717 19738 4718
rect 19766 4717 19790 4718
rect 19724 4691 19738 4717
rect 19786 4691 19790 4717
rect 19714 4690 19738 4691
rect 19766 4690 19790 4691
rect 19818 4717 19842 4718
rect 19870 4717 19894 4718
rect 19818 4691 19822 4717
rect 19870 4691 19884 4717
rect 19818 4690 19842 4691
rect 19870 4690 19894 4691
rect 19922 4690 19946 4718
rect 19974 4690 19998 4718
rect 20026 4717 20035 4718
rect 20034 4691 20035 4717
rect 20026 4690 20035 4691
rect 19573 4685 20035 4690
rect 19446 4551 19447 4577
rect 19473 4551 19474 4577
rect 19446 4521 19474 4551
rect 19446 4495 19447 4521
rect 19473 4495 19474 4521
rect 19446 4074 19474 4495
rect 20118 4186 20146 4774
rect 19950 4158 20118 4186
rect 19950 4129 19978 4158
rect 20118 4153 20146 4158
rect 19950 4103 19951 4129
rect 19977 4103 19978 4129
rect 19950 4074 19978 4103
rect 19446 4073 19978 4074
rect 19446 4047 19951 4073
rect 19977 4047 19978 4073
rect 19446 4046 19978 4047
rect 19446 3793 19474 4046
rect 19950 4041 19978 4046
rect 20230 4129 20258 4135
rect 20230 4103 20231 4129
rect 20257 4103 20258 4129
rect 19573 3934 20035 3939
rect 19573 3933 19582 3934
rect 19573 3907 19574 3933
rect 19573 3906 19582 3907
rect 19610 3906 19634 3934
rect 19662 3906 19686 3934
rect 19714 3933 19738 3934
rect 19766 3933 19790 3934
rect 19724 3907 19738 3933
rect 19786 3907 19790 3933
rect 19714 3906 19738 3907
rect 19766 3906 19790 3907
rect 19818 3933 19842 3934
rect 19870 3933 19894 3934
rect 19818 3907 19822 3933
rect 19870 3907 19884 3933
rect 19818 3906 19842 3907
rect 19870 3906 19894 3907
rect 19922 3906 19946 3934
rect 19974 3906 19998 3934
rect 20026 3933 20035 3934
rect 20034 3907 20035 3933
rect 20026 3906 20035 3907
rect 19573 3901 20035 3906
rect 19446 3767 19447 3793
rect 19473 3767 19474 3793
rect 19446 3738 19474 3767
rect 19166 3737 19474 3738
rect 19166 3711 19447 3737
rect 19473 3711 19474 3737
rect 19166 3710 19474 3711
rect 19166 3346 19194 3710
rect 19446 3705 19474 3710
rect 19166 3313 19194 3318
rect 19222 3346 19250 3351
rect 19446 3346 19474 3351
rect 19222 3345 19446 3346
rect 19222 3319 19223 3345
rect 19249 3319 19446 3345
rect 19222 3318 19446 3319
rect 18886 2921 18914 2926
rect 19222 3009 19250 3318
rect 19446 3280 19474 3318
rect 20230 3345 20258 4103
rect 20566 3402 20594 10094
rect 20790 10009 20818 10767
rect 21014 10094 21042 11102
rect 21182 11097 21210 11102
rect 21742 10849 21770 10855
rect 21742 10823 21743 10849
rect 21769 10823 21770 10849
rect 21742 10793 21770 10823
rect 21742 10767 21743 10793
rect 21769 10767 21770 10793
rect 21406 10401 21434 10407
rect 21406 10375 21407 10401
rect 21433 10375 21434 10401
rect 21406 10346 21434 10375
rect 21406 10299 21434 10318
rect 21742 10346 21770 10767
rect 22526 10794 22554 10799
rect 22582 10794 22610 11550
rect 22526 10793 22610 10794
rect 22526 10767 22527 10793
rect 22553 10767 22610 10793
rect 22526 10766 22610 10767
rect 22526 10761 22554 10766
rect 22073 10598 22535 10603
rect 22073 10597 22082 10598
rect 22073 10571 22074 10597
rect 22073 10570 22082 10571
rect 22110 10570 22134 10598
rect 22162 10570 22186 10598
rect 22214 10597 22238 10598
rect 22266 10597 22290 10598
rect 22224 10571 22238 10597
rect 22286 10571 22290 10597
rect 22214 10570 22238 10571
rect 22266 10570 22290 10571
rect 22318 10597 22342 10598
rect 22370 10597 22394 10598
rect 22318 10571 22322 10597
rect 22370 10571 22384 10597
rect 22318 10570 22342 10571
rect 22370 10570 22394 10571
rect 22422 10570 22446 10598
rect 22474 10570 22498 10598
rect 22526 10597 22535 10598
rect 22534 10571 22535 10597
rect 22526 10570 22535 10571
rect 22073 10565 22535 10570
rect 21014 10066 21322 10094
rect 20790 9983 20791 10009
rect 20817 9983 20818 10009
rect 20790 9225 20818 9983
rect 20790 9199 20791 9225
rect 20817 9199 20818 9225
rect 20790 8441 20818 9199
rect 20790 8415 20791 8441
rect 20817 8415 20818 8441
rect 20790 7657 20818 8415
rect 20790 7631 20791 7657
rect 20817 7631 20818 7657
rect 20790 6873 20818 7631
rect 20790 6847 20791 6873
rect 20817 6847 20818 6873
rect 20790 6090 20818 6847
rect 20790 5306 20818 6062
rect 20790 5259 20818 5278
rect 21294 9617 21322 10066
rect 21742 10065 21770 10318
rect 21742 10039 21743 10065
rect 21769 10039 21770 10065
rect 21742 10010 21770 10039
rect 22582 10094 22610 10766
rect 22750 11185 22778 11191
rect 22750 11159 22751 11185
rect 22777 11159 22778 11185
rect 22750 10401 22778 11159
rect 22750 10375 22751 10401
rect 22777 10375 22778 10401
rect 22750 10094 22778 10375
rect 22582 10066 22778 10094
rect 22806 10906 22834 11943
rect 23926 11969 23954 11975
rect 23926 11943 23927 11969
rect 23953 11943 23954 11969
rect 23926 11914 23954 11943
rect 23926 11867 23954 11886
rect 23310 11633 23338 11639
rect 23310 11607 23311 11633
rect 23337 11607 23338 11633
rect 23310 11577 23338 11607
rect 23310 11551 23311 11577
rect 23337 11551 23338 11577
rect 23310 11186 23338 11551
rect 23422 11186 23450 11191
rect 23310 11185 23450 11186
rect 23310 11159 23311 11185
rect 23337 11159 23423 11185
rect 23449 11159 23450 11185
rect 23310 11158 23450 11159
rect 23310 11153 23338 11158
rect 22806 10122 22834 10878
rect 22806 10089 22834 10094
rect 23366 10849 23394 11158
rect 23422 11153 23450 11158
rect 23366 10823 23367 10849
rect 23393 10823 23394 10849
rect 23366 10793 23394 10823
rect 23366 10767 23367 10793
rect 23393 10767 23394 10793
rect 21742 9944 21770 9982
rect 22526 10010 22554 10015
rect 22582 10010 22610 10066
rect 22526 10009 22610 10010
rect 22526 9983 22527 10009
rect 22553 9983 22610 10009
rect 22526 9982 22610 9983
rect 22694 10010 22722 10015
rect 22526 9977 22554 9982
rect 22694 9963 22722 9982
rect 22073 9814 22535 9819
rect 22073 9813 22082 9814
rect 22073 9787 22074 9813
rect 22073 9786 22082 9787
rect 22110 9786 22134 9814
rect 22162 9786 22186 9814
rect 22214 9813 22238 9814
rect 22266 9813 22290 9814
rect 22224 9787 22238 9813
rect 22286 9787 22290 9813
rect 22214 9786 22238 9787
rect 22266 9786 22290 9787
rect 22318 9813 22342 9814
rect 22370 9813 22394 9814
rect 22318 9787 22322 9813
rect 22370 9787 22384 9813
rect 22318 9786 22342 9787
rect 22370 9786 22394 9787
rect 22422 9786 22446 9814
rect 22474 9786 22498 9814
rect 22526 9813 22535 9814
rect 22534 9787 22535 9813
rect 22526 9786 22535 9787
rect 22073 9781 22535 9786
rect 21294 9591 21295 9617
rect 21321 9591 21322 9617
rect 21294 9561 21322 9591
rect 21294 9535 21295 9561
rect 21321 9535 21322 9561
rect 21294 9226 21322 9535
rect 22750 9617 22778 10066
rect 22918 10010 22946 10015
rect 22918 9963 22946 9982
rect 23366 10010 23394 10767
rect 22750 9591 22751 9617
rect 22777 9591 22778 9617
rect 22750 9282 22778 9591
rect 23310 9618 23338 9623
rect 23366 9618 23394 9982
rect 23702 10401 23730 10407
rect 23702 10375 23703 10401
rect 23729 10375 23730 10401
rect 23702 10345 23730 10375
rect 23702 10319 23703 10345
rect 23729 10319 23730 10345
rect 23422 9618 23450 9623
rect 23310 9617 23422 9618
rect 23310 9591 23311 9617
rect 23337 9591 23422 9617
rect 23310 9590 23422 9591
rect 23310 9585 23338 9590
rect 23422 9552 23450 9590
rect 21462 9226 21490 9231
rect 21294 9225 21490 9226
rect 21294 9199 21295 9225
rect 21321 9199 21463 9225
rect 21489 9199 21490 9225
rect 21294 9198 21490 9199
rect 21294 8833 21322 9198
rect 21462 9193 21490 9198
rect 22526 9226 22554 9231
rect 22526 9225 22610 9226
rect 22526 9199 22527 9225
rect 22553 9199 22610 9225
rect 22526 9198 22610 9199
rect 22526 9193 22554 9198
rect 22073 9030 22535 9035
rect 22073 9029 22082 9030
rect 22073 9003 22074 9029
rect 22073 9002 22082 9003
rect 22110 9002 22134 9030
rect 22162 9002 22186 9030
rect 22214 9029 22238 9030
rect 22266 9029 22290 9030
rect 22224 9003 22238 9029
rect 22286 9003 22290 9029
rect 22214 9002 22238 9003
rect 22266 9002 22290 9003
rect 22318 9029 22342 9030
rect 22370 9029 22394 9030
rect 22318 9003 22322 9029
rect 22370 9003 22384 9029
rect 22318 9002 22342 9003
rect 22370 9002 22394 9003
rect 22422 9002 22446 9030
rect 22474 9002 22498 9030
rect 22526 9029 22535 9030
rect 22534 9003 22535 9029
rect 22526 9002 22535 9003
rect 22073 8997 22535 9002
rect 21294 8807 21295 8833
rect 21321 8807 21322 8833
rect 21294 8777 21322 8807
rect 21294 8751 21295 8777
rect 21321 8751 21322 8777
rect 21294 8442 21322 8751
rect 21462 8442 21490 8447
rect 21294 8441 21490 8442
rect 21294 8415 21295 8441
rect 21321 8415 21463 8441
rect 21489 8415 21490 8441
rect 21294 8414 21490 8415
rect 21294 8049 21322 8414
rect 21462 8409 21490 8414
rect 22526 8442 22554 8447
rect 22582 8442 22610 9198
rect 22526 8441 22610 8442
rect 22526 8415 22527 8441
rect 22553 8415 22610 8441
rect 22526 8414 22610 8415
rect 22526 8409 22554 8414
rect 22073 8246 22535 8251
rect 22073 8245 22082 8246
rect 22073 8219 22074 8245
rect 22073 8218 22082 8219
rect 22110 8218 22134 8246
rect 22162 8218 22186 8246
rect 22214 8245 22238 8246
rect 22266 8245 22290 8246
rect 22224 8219 22238 8245
rect 22286 8219 22290 8245
rect 22214 8218 22238 8219
rect 22266 8218 22290 8219
rect 22318 8245 22342 8246
rect 22370 8245 22394 8246
rect 22318 8219 22322 8245
rect 22370 8219 22384 8245
rect 22318 8218 22342 8219
rect 22370 8218 22394 8219
rect 22422 8218 22446 8246
rect 22474 8218 22498 8246
rect 22526 8245 22535 8246
rect 22534 8219 22535 8245
rect 22526 8218 22535 8219
rect 22073 8213 22535 8218
rect 21294 8023 21295 8049
rect 21321 8023 21322 8049
rect 21294 7993 21322 8023
rect 21294 7967 21295 7993
rect 21321 7967 21322 7993
rect 21294 7658 21322 7967
rect 21462 7658 21490 7663
rect 21294 7657 21490 7658
rect 21294 7631 21295 7657
rect 21321 7631 21463 7657
rect 21489 7631 21490 7657
rect 21294 7630 21490 7631
rect 21294 7265 21322 7630
rect 21462 7625 21490 7630
rect 22526 7658 22554 7663
rect 22582 7658 22610 8414
rect 22526 7657 22610 7658
rect 22526 7631 22527 7657
rect 22553 7631 22610 7657
rect 22526 7630 22610 7631
rect 22526 7625 22554 7630
rect 22073 7462 22535 7467
rect 22073 7461 22082 7462
rect 22073 7435 22074 7461
rect 22073 7434 22082 7435
rect 22110 7434 22134 7462
rect 22162 7434 22186 7462
rect 22214 7461 22238 7462
rect 22266 7461 22290 7462
rect 22224 7435 22238 7461
rect 22286 7435 22290 7461
rect 22214 7434 22238 7435
rect 22266 7434 22290 7435
rect 22318 7461 22342 7462
rect 22370 7461 22394 7462
rect 22318 7435 22322 7461
rect 22370 7435 22384 7461
rect 22318 7434 22342 7435
rect 22370 7434 22394 7435
rect 22422 7434 22446 7462
rect 22474 7434 22498 7462
rect 22526 7461 22535 7462
rect 22534 7435 22535 7461
rect 22526 7434 22535 7435
rect 22073 7429 22535 7434
rect 21294 7239 21295 7265
rect 21321 7239 21322 7265
rect 21294 7209 21322 7239
rect 21294 7183 21295 7209
rect 21321 7183 21322 7209
rect 21294 6874 21322 7183
rect 21462 6874 21490 6879
rect 21294 6873 21490 6874
rect 21294 6847 21295 6873
rect 21321 6847 21463 6873
rect 21489 6847 21490 6873
rect 21294 6846 21490 6847
rect 21294 6481 21322 6846
rect 21462 6841 21490 6846
rect 22526 6874 22554 6879
rect 22582 6874 22610 7630
rect 22526 6873 22610 6874
rect 22526 6847 22527 6873
rect 22553 6847 22610 6873
rect 22526 6846 22610 6847
rect 22526 6841 22554 6846
rect 22073 6678 22535 6683
rect 22073 6677 22082 6678
rect 22073 6651 22074 6677
rect 22073 6650 22082 6651
rect 22110 6650 22134 6678
rect 22162 6650 22186 6678
rect 22214 6677 22238 6678
rect 22266 6677 22290 6678
rect 22224 6651 22238 6677
rect 22286 6651 22290 6677
rect 22214 6650 22238 6651
rect 22266 6650 22290 6651
rect 22318 6677 22342 6678
rect 22370 6677 22394 6678
rect 22318 6651 22322 6677
rect 22370 6651 22384 6677
rect 22318 6650 22342 6651
rect 22370 6650 22394 6651
rect 22422 6650 22446 6678
rect 22474 6650 22498 6678
rect 22526 6677 22535 6678
rect 22534 6651 22535 6677
rect 22526 6650 22535 6651
rect 22073 6645 22535 6650
rect 21294 6455 21295 6481
rect 21321 6455 21322 6481
rect 21294 6425 21322 6455
rect 21294 6399 21295 6425
rect 21321 6399 21322 6425
rect 21294 6090 21322 6399
rect 22582 6482 22610 6846
rect 22750 8833 22778 9254
rect 23422 9281 23450 9287
rect 23422 9255 23423 9281
rect 23449 9255 23450 9281
rect 23422 9226 23450 9255
rect 22750 8807 22751 8833
rect 22777 8807 22778 8833
rect 22750 8049 22778 8807
rect 23310 8834 23338 8839
rect 23422 8834 23450 9198
rect 23702 9226 23730 10319
rect 23702 9193 23730 9198
rect 23310 8833 23450 8834
rect 23310 8807 23311 8833
rect 23337 8807 23423 8833
rect 23449 8807 23450 8833
rect 23310 8806 23450 8807
rect 23310 8801 23338 8806
rect 23422 8497 23450 8806
rect 23422 8471 23423 8497
rect 23449 8471 23450 8497
rect 23422 8442 23450 8471
rect 22750 8023 22751 8049
rect 22777 8023 22778 8049
rect 22750 7265 22778 8023
rect 23310 8050 23338 8055
rect 23422 8050 23450 8414
rect 23310 8049 23450 8050
rect 23310 8023 23311 8049
rect 23337 8023 23423 8049
rect 23449 8023 23450 8049
rect 23310 8022 23450 8023
rect 23310 8017 23338 8022
rect 23422 7713 23450 8022
rect 23422 7687 23423 7713
rect 23449 7687 23450 7713
rect 23422 7657 23450 7687
rect 23422 7631 23423 7657
rect 23449 7631 23450 7657
rect 22750 7239 22751 7265
rect 22777 7239 22778 7265
rect 22750 6482 22778 7239
rect 23310 7266 23338 7271
rect 23422 7266 23450 7631
rect 23310 7265 23450 7266
rect 23310 7239 23311 7265
rect 23337 7239 23423 7265
rect 23449 7239 23450 7265
rect 23310 7238 23450 7239
rect 23310 7233 23338 7238
rect 23422 6929 23450 7238
rect 23422 6903 23423 6929
rect 23449 6903 23450 6929
rect 23422 6873 23450 6903
rect 23422 6847 23423 6873
rect 23449 6847 23450 6873
rect 23198 6482 23226 6487
rect 23422 6482 23450 6847
rect 22582 6481 22778 6482
rect 22582 6455 22751 6481
rect 22777 6455 22778 6481
rect 22582 6454 22778 6455
rect 21462 6090 21490 6095
rect 21294 6089 21490 6090
rect 21294 6063 21295 6089
rect 21321 6063 21463 6089
rect 21489 6063 21490 6089
rect 21294 6062 21490 6063
rect 21294 5697 21322 6062
rect 21462 6034 21490 6062
rect 22246 6090 22274 6095
rect 22246 6043 22274 6062
rect 22582 6090 22610 6454
rect 22750 6449 22778 6454
rect 22918 6481 23450 6482
rect 22918 6455 23199 6481
rect 23225 6455 23423 6481
rect 23449 6455 23450 6481
rect 22918 6454 23450 6455
rect 22582 6057 22610 6062
rect 22694 6090 22722 6095
rect 22918 6090 22946 6454
rect 23198 6449 23226 6454
rect 23422 6449 23450 6454
rect 22694 6089 22946 6090
rect 22694 6063 22695 6089
rect 22721 6063 22919 6089
rect 22945 6063 22946 6089
rect 22694 6062 22946 6063
rect 21462 6001 21490 6006
rect 22694 6034 22722 6062
rect 22918 6057 22946 6062
rect 23086 6370 23114 6375
rect 22694 6001 22722 6006
rect 22073 5894 22535 5899
rect 22073 5893 22082 5894
rect 22073 5867 22074 5893
rect 22073 5866 22082 5867
rect 22110 5866 22134 5894
rect 22162 5866 22186 5894
rect 22214 5893 22238 5894
rect 22266 5893 22290 5894
rect 22224 5867 22238 5893
rect 22286 5867 22290 5893
rect 22214 5866 22238 5867
rect 22266 5866 22290 5867
rect 22318 5893 22342 5894
rect 22370 5893 22394 5894
rect 22318 5867 22322 5893
rect 22370 5867 22384 5893
rect 22318 5866 22342 5867
rect 22370 5866 22394 5867
rect 22422 5866 22446 5894
rect 22474 5866 22498 5894
rect 22526 5893 22535 5894
rect 22534 5867 22535 5893
rect 22526 5866 22535 5867
rect 22073 5861 22535 5866
rect 21294 5671 21295 5697
rect 21321 5671 21322 5697
rect 21294 5641 21322 5671
rect 21294 5615 21295 5641
rect 21321 5615 21322 5641
rect 21294 5306 21322 5615
rect 22750 5697 22778 5703
rect 22750 5671 22751 5697
rect 22777 5671 22778 5697
rect 21462 5306 21490 5311
rect 21294 5305 21490 5306
rect 21294 5279 21295 5305
rect 21321 5279 21463 5305
rect 21489 5279 21490 5305
rect 21294 5278 21490 5279
rect 21294 4913 21322 5278
rect 21462 5273 21490 5278
rect 22526 5306 22554 5311
rect 22526 5305 22610 5306
rect 22526 5279 22527 5305
rect 22553 5279 22610 5305
rect 22526 5278 22610 5279
rect 22526 5273 22554 5278
rect 22073 5110 22535 5115
rect 22073 5109 22082 5110
rect 22073 5083 22074 5109
rect 22073 5082 22082 5083
rect 22110 5082 22134 5110
rect 22162 5082 22186 5110
rect 22214 5109 22238 5110
rect 22266 5109 22290 5110
rect 22224 5083 22238 5109
rect 22286 5083 22290 5109
rect 22214 5082 22238 5083
rect 22266 5082 22290 5083
rect 22318 5109 22342 5110
rect 22370 5109 22394 5110
rect 22318 5083 22322 5109
rect 22370 5083 22384 5109
rect 22318 5082 22342 5083
rect 22370 5082 22394 5083
rect 22422 5082 22446 5110
rect 22474 5082 22498 5110
rect 22526 5109 22535 5110
rect 22534 5083 22535 5109
rect 22526 5082 22535 5083
rect 22073 5077 22535 5082
rect 21294 4887 21295 4913
rect 21321 4887 21322 4913
rect 21294 4857 21322 4887
rect 21294 4831 21295 4857
rect 21321 4831 21322 4857
rect 20566 3369 20594 3374
rect 20790 4521 20818 4527
rect 20790 4495 20791 4521
rect 20817 4495 20818 4521
rect 20790 3737 20818 4495
rect 21294 4214 21322 4831
rect 21798 4577 21826 4583
rect 21798 4551 21799 4577
rect 21825 4551 21826 4577
rect 21406 4522 21434 4527
rect 21294 4186 21378 4214
rect 21406 4186 21434 4494
rect 21798 4522 21826 4551
rect 21798 4214 21826 4494
rect 22526 4522 22554 4527
rect 22582 4522 22610 5278
rect 22750 4913 22778 5671
rect 22750 4887 22751 4913
rect 22777 4887 22778 4913
rect 22526 4521 22610 4522
rect 22526 4495 22527 4521
rect 22553 4495 22610 4521
rect 22526 4494 22610 4495
rect 22526 4489 22554 4494
rect 22073 4326 22535 4331
rect 22073 4325 22082 4326
rect 22073 4299 22074 4325
rect 22073 4298 22082 4299
rect 22110 4298 22134 4326
rect 22162 4298 22186 4326
rect 22214 4325 22238 4326
rect 22266 4325 22290 4326
rect 22224 4299 22238 4325
rect 22286 4299 22290 4325
rect 22214 4298 22238 4299
rect 22266 4298 22290 4299
rect 22318 4325 22342 4326
rect 22370 4325 22394 4326
rect 22318 4299 22322 4325
rect 22370 4299 22384 4325
rect 22318 4298 22342 4299
rect 22370 4298 22394 4299
rect 22422 4298 22446 4326
rect 22474 4298 22498 4326
rect 22526 4325 22535 4326
rect 22534 4299 22535 4325
rect 22526 4298 22535 4299
rect 22073 4293 22535 4298
rect 21686 4186 21714 4191
rect 21406 4158 21490 4186
rect 21350 4153 21378 4158
rect 20790 3711 20791 3737
rect 20817 3711 20818 3737
rect 20230 3319 20231 3345
rect 20257 3319 20258 3345
rect 19573 3150 20035 3155
rect 19573 3149 19582 3150
rect 19573 3123 19574 3149
rect 19573 3122 19582 3123
rect 19610 3122 19634 3150
rect 19662 3122 19686 3150
rect 19714 3149 19738 3150
rect 19766 3149 19790 3150
rect 19724 3123 19738 3149
rect 19786 3123 19790 3149
rect 19714 3122 19738 3123
rect 19766 3122 19790 3123
rect 19818 3149 19842 3150
rect 19870 3149 19894 3150
rect 19818 3123 19822 3149
rect 19870 3123 19884 3149
rect 19818 3122 19842 3123
rect 19870 3122 19894 3123
rect 19922 3122 19946 3150
rect 19974 3122 19998 3150
rect 20026 3149 20035 3150
rect 20034 3123 20035 3149
rect 20026 3122 20035 3123
rect 19573 3117 20035 3122
rect 19222 2983 19223 3009
rect 19249 2983 19250 3009
rect 19222 2953 19250 2983
rect 19222 2927 19223 2953
rect 19249 2927 19250 2953
rect 18550 2170 18578 2175
rect 18550 1777 18578 2142
rect 18774 2170 18802 2478
rect 19222 2618 19250 2927
rect 19222 2225 19250 2590
rect 20118 2562 20146 2567
rect 20118 2515 20146 2534
rect 20230 2506 20258 3319
rect 20230 2473 20258 2478
rect 20790 2954 20818 3711
rect 21182 4129 21210 4135
rect 21182 4103 21183 4129
rect 21209 4103 21210 4129
rect 21182 4073 21210 4103
rect 21182 4047 21183 4073
rect 21209 4047 21210 4073
rect 21182 4018 21210 4047
rect 21462 4018 21490 4158
rect 21182 3990 21490 4018
rect 21014 3346 21042 3351
rect 21014 3299 21042 3318
rect 21182 3346 21210 3990
rect 21686 3402 21714 4158
rect 21742 4186 21826 4214
rect 21742 3793 21770 4186
rect 21742 3767 21743 3793
rect 21769 3767 21770 3793
rect 21742 3737 21770 3767
rect 22582 4130 22610 4494
rect 22694 4522 22722 4527
rect 22694 4475 22722 4494
rect 22750 4130 22778 4887
rect 22918 4522 22946 4527
rect 22918 4475 22946 4494
rect 22582 4102 22750 4130
rect 21742 3711 21743 3737
rect 21769 3711 21770 3737
rect 21742 3705 21770 3711
rect 22526 3738 22554 3743
rect 22582 3738 22610 4102
rect 22750 4064 22778 4102
rect 22526 3737 22610 3738
rect 22526 3711 22527 3737
rect 22553 3711 22610 3737
rect 22526 3710 22610 3711
rect 22526 3705 22554 3710
rect 22073 3542 22535 3547
rect 22073 3541 22082 3542
rect 22073 3515 22074 3541
rect 22073 3514 22082 3515
rect 22110 3514 22134 3542
rect 22162 3514 22186 3542
rect 22214 3541 22238 3542
rect 22266 3541 22290 3542
rect 22224 3515 22238 3541
rect 22286 3515 22290 3541
rect 22214 3514 22238 3515
rect 22266 3514 22290 3515
rect 22318 3541 22342 3542
rect 22370 3541 22394 3542
rect 22318 3515 22322 3541
rect 22370 3515 22384 3541
rect 22318 3514 22342 3515
rect 22370 3514 22394 3515
rect 22422 3514 22446 3542
rect 22474 3514 22498 3542
rect 22526 3541 22535 3542
rect 22534 3515 22535 3541
rect 22526 3514 22535 3515
rect 22073 3509 22535 3514
rect 21742 3402 21770 3407
rect 21686 3374 21742 3402
rect 21182 3289 21210 3318
rect 21182 3263 21183 3289
rect 21209 3263 21210 3289
rect 21182 3257 21210 3263
rect 20790 2506 20818 2926
rect 21406 3066 21434 3071
rect 19573 2366 20035 2371
rect 19573 2365 19582 2366
rect 19573 2339 19574 2365
rect 19573 2338 19582 2339
rect 19610 2338 19634 2366
rect 19662 2338 19686 2366
rect 19714 2365 19738 2366
rect 19766 2365 19790 2366
rect 19724 2339 19738 2365
rect 19786 2339 19790 2365
rect 19714 2338 19738 2339
rect 19766 2338 19790 2339
rect 19818 2365 19842 2366
rect 19870 2365 19894 2366
rect 19818 2339 19822 2365
rect 19870 2339 19884 2365
rect 19818 2338 19842 2339
rect 19870 2338 19894 2339
rect 19922 2338 19946 2366
rect 19974 2338 19998 2366
rect 20026 2365 20035 2366
rect 20034 2339 20035 2365
rect 20026 2338 20035 2339
rect 19573 2333 20035 2338
rect 19222 2199 19223 2225
rect 19249 2199 19250 2225
rect 18774 2137 18802 2142
rect 19110 2170 19138 2175
rect 19222 2170 19250 2199
rect 19110 2169 19250 2170
rect 19110 2143 19111 2169
rect 19137 2143 19250 2169
rect 19110 2142 19250 2143
rect 20790 2169 20818 2478
rect 20958 2618 20986 2623
rect 20958 2561 20986 2590
rect 20958 2535 20959 2561
rect 20985 2535 20986 2561
rect 20958 2505 20986 2535
rect 20958 2479 20959 2505
rect 20985 2479 20986 2505
rect 20958 2473 20986 2479
rect 21406 2562 21434 3038
rect 20790 2143 20791 2169
rect 20817 2143 20818 2169
rect 18550 1751 18551 1777
rect 18577 1751 18578 1777
rect 18550 1745 18578 1751
rect 19110 1778 19138 2142
rect 20790 2137 20818 2143
rect 19222 1778 19250 1783
rect 19110 1777 19250 1778
rect 19110 1751 19111 1777
rect 19137 1751 19223 1777
rect 19249 1751 19250 1777
rect 19110 1750 19250 1751
rect 19110 1745 19138 1750
rect 19222 1745 19250 1750
rect 20118 1778 20146 1783
rect 19573 1582 20035 1587
rect 19573 1581 19582 1582
rect 19573 1555 19574 1581
rect 19573 1554 19582 1555
rect 19610 1554 19634 1582
rect 19662 1554 19686 1582
rect 19714 1581 19738 1582
rect 19766 1581 19790 1582
rect 19724 1555 19738 1581
rect 19786 1555 19790 1581
rect 19714 1554 19738 1555
rect 19766 1554 19790 1555
rect 19818 1581 19842 1582
rect 19870 1581 19894 1582
rect 19818 1555 19822 1581
rect 19870 1555 19884 1581
rect 19818 1554 19842 1555
rect 19870 1554 19894 1555
rect 19922 1554 19946 1582
rect 19974 1554 19998 1582
rect 20026 1581 20035 1582
rect 20034 1555 20035 1581
rect 20026 1554 20035 1555
rect 19573 1549 20035 1554
rect 18494 400 18522 1470
rect 20118 490 20146 1750
rect 21182 1778 21210 1783
rect 21182 1731 21210 1750
rect 19950 462 20146 490
rect 19950 400 19978 462
rect 21406 400 21434 2534
rect 21742 3009 21770 3374
rect 21742 2983 21743 3009
rect 21769 2983 21770 3009
rect 21742 2953 21770 2983
rect 22582 3346 22610 3710
rect 22806 3738 22834 3743
rect 22918 3738 22946 3743
rect 22806 3737 22946 3738
rect 22806 3711 22807 3737
rect 22833 3711 22919 3737
rect 22945 3711 22946 3737
rect 22806 3710 22946 3711
rect 22806 3402 22834 3710
rect 22918 3705 22946 3710
rect 22806 3369 22834 3374
rect 22750 3346 22778 3351
rect 22582 3345 22778 3346
rect 22582 3319 22751 3345
rect 22777 3319 22778 3345
rect 22582 3318 22778 3319
rect 21742 2927 21743 2953
rect 21769 2927 21770 2953
rect 21742 2225 21770 2927
rect 22246 2954 22274 2959
rect 22246 2907 22274 2926
rect 22582 2954 22610 3318
rect 22750 3313 22778 3318
rect 22582 2921 22610 2926
rect 22073 2758 22535 2763
rect 22073 2757 22082 2758
rect 22073 2731 22074 2757
rect 22073 2730 22082 2731
rect 22110 2730 22134 2758
rect 22162 2730 22186 2758
rect 22214 2757 22238 2758
rect 22266 2757 22290 2758
rect 22224 2731 22238 2757
rect 22286 2731 22290 2757
rect 22214 2730 22238 2731
rect 22266 2730 22290 2731
rect 22318 2757 22342 2758
rect 22370 2757 22394 2758
rect 22318 2731 22322 2757
rect 22370 2731 22384 2757
rect 22318 2730 22342 2731
rect 22370 2730 22394 2731
rect 22422 2730 22446 2758
rect 22474 2730 22498 2758
rect 22526 2757 22535 2758
rect 22534 2731 22535 2757
rect 22526 2730 22535 2731
rect 22073 2725 22535 2730
rect 21742 2199 21743 2225
rect 21769 2199 21770 2225
rect 21742 2169 21770 2199
rect 22750 2561 22778 2567
rect 22750 2535 22751 2561
rect 22777 2535 22778 2561
rect 22750 2450 22778 2535
rect 21742 2143 21743 2169
rect 21769 2143 21770 2169
rect 21742 2137 21770 2143
rect 22526 2170 22554 2175
rect 22750 2170 22778 2422
rect 22526 2169 22778 2170
rect 22526 2143 22527 2169
rect 22553 2143 22778 2169
rect 22526 2142 22778 2143
rect 22526 2137 22554 2142
rect 22073 1974 22535 1979
rect 22073 1973 22082 1974
rect 22073 1947 22074 1973
rect 22073 1946 22082 1947
rect 22110 1946 22134 1974
rect 22162 1946 22186 1974
rect 22214 1973 22238 1974
rect 22266 1973 22290 1974
rect 22224 1947 22238 1973
rect 22286 1947 22290 1973
rect 22214 1946 22238 1947
rect 22266 1946 22290 1947
rect 22318 1973 22342 1974
rect 22370 1973 22394 1974
rect 22318 1947 22322 1973
rect 22370 1947 22384 1973
rect 22318 1946 22342 1947
rect 22370 1946 22394 1947
rect 22422 1946 22446 1974
rect 22474 1946 22498 1974
rect 22526 1973 22535 1974
rect 22534 1947 22535 1973
rect 22526 1946 22535 1947
rect 22073 1941 22535 1946
rect 22470 1834 22498 1839
rect 22582 1834 22610 2142
rect 22498 1806 22610 1834
rect 21798 1777 21826 1783
rect 21798 1751 21799 1777
rect 21825 1751 21826 1777
rect 21798 1722 21826 1751
rect 22470 1777 22498 1806
rect 22470 1751 22471 1777
rect 22497 1751 22498 1777
rect 22470 1745 22498 1751
rect 22862 1778 22890 1783
rect 21854 1722 21882 1727
rect 21826 1721 21882 1722
rect 21826 1695 21855 1721
rect 21881 1695 21882 1721
rect 21826 1694 21882 1695
rect 21798 1656 21826 1694
rect 21854 1689 21882 1694
rect 22862 400 22890 1750
rect 22918 1777 22946 1783
rect 22918 1751 22919 1777
rect 22945 1751 22946 1777
rect 22918 1666 22946 1751
rect 23086 1778 23114 6342
rect 23198 5698 23226 5703
rect 23422 5698 23450 5703
rect 23198 5697 23450 5698
rect 23198 5671 23199 5697
rect 23225 5671 23423 5697
rect 23449 5671 23450 5697
rect 23198 5670 23450 5671
rect 23198 5361 23226 5670
rect 23422 5665 23450 5670
rect 23198 5335 23199 5361
rect 23225 5335 23226 5361
rect 23198 5305 23226 5335
rect 23198 5279 23199 5305
rect 23225 5279 23226 5305
rect 23198 4914 23226 5279
rect 23422 4914 23450 4919
rect 23198 4913 23450 4914
rect 23198 4887 23199 4913
rect 23225 4887 23423 4913
rect 23449 4887 23450 4913
rect 23198 4886 23450 4887
rect 23198 4522 23226 4886
rect 23422 4881 23450 4886
rect 23198 4489 23226 4494
rect 23310 4130 23338 4135
rect 23422 4130 23450 4135
rect 23310 4129 23450 4130
rect 23310 4103 23311 4129
rect 23337 4103 23423 4129
rect 23449 4103 23450 4129
rect 23310 4102 23450 4103
rect 23310 4097 23338 4102
rect 23422 4074 23450 4102
rect 23198 3402 23226 3407
rect 23198 3345 23226 3374
rect 23198 3319 23199 3345
rect 23225 3319 23226 3345
rect 23198 3313 23226 3319
rect 23422 3402 23450 4046
rect 23422 3345 23450 3374
rect 23422 3319 23423 3345
rect 23449 3319 23450 3345
rect 23422 3009 23450 3319
rect 23422 2983 23423 3009
rect 23449 2983 23450 3009
rect 23422 2953 23450 2983
rect 23422 2927 23423 2953
rect 23449 2927 23450 2953
rect 23422 2921 23450 2927
rect 23198 2562 23226 2567
rect 23198 2225 23226 2534
rect 23534 2562 23562 2567
rect 23534 2515 23562 2534
rect 23198 2199 23199 2225
rect 23225 2199 23226 2225
rect 23086 1745 23114 1750
rect 23142 2170 23170 2175
rect 23198 2170 23226 2199
rect 24094 2506 24122 16366
rect 24430 16282 24458 16287
rect 24430 12810 24458 16254
rect 27073 16086 27535 16091
rect 27073 16085 27082 16086
rect 27073 16059 27074 16085
rect 27073 16058 27082 16059
rect 27110 16058 27134 16086
rect 27162 16058 27186 16086
rect 27214 16085 27238 16086
rect 27266 16085 27290 16086
rect 27224 16059 27238 16085
rect 27286 16059 27290 16085
rect 27214 16058 27238 16059
rect 27266 16058 27290 16059
rect 27318 16085 27342 16086
rect 27370 16085 27394 16086
rect 27318 16059 27322 16085
rect 27370 16059 27384 16085
rect 27318 16058 27342 16059
rect 27370 16058 27394 16059
rect 27422 16058 27446 16086
rect 27474 16058 27498 16086
rect 27526 16085 27535 16086
rect 27534 16059 27535 16085
rect 27526 16058 27535 16059
rect 27073 16053 27535 16058
rect 24573 15694 25035 15699
rect 24573 15693 24582 15694
rect 24573 15667 24574 15693
rect 24573 15666 24582 15667
rect 24610 15666 24634 15694
rect 24662 15666 24686 15694
rect 24714 15693 24738 15694
rect 24766 15693 24790 15694
rect 24724 15667 24738 15693
rect 24786 15667 24790 15693
rect 24714 15666 24738 15667
rect 24766 15666 24790 15667
rect 24818 15693 24842 15694
rect 24870 15693 24894 15694
rect 24818 15667 24822 15693
rect 24870 15667 24884 15693
rect 24818 15666 24842 15667
rect 24870 15666 24894 15667
rect 24922 15666 24946 15694
rect 24974 15666 24998 15694
rect 25026 15693 25035 15694
rect 25034 15667 25035 15693
rect 25026 15666 25035 15667
rect 24573 15661 25035 15666
rect 27073 15302 27535 15307
rect 27073 15301 27082 15302
rect 27073 15275 27074 15301
rect 27073 15274 27082 15275
rect 27110 15274 27134 15302
rect 27162 15274 27186 15302
rect 27214 15301 27238 15302
rect 27266 15301 27290 15302
rect 27224 15275 27238 15301
rect 27286 15275 27290 15301
rect 27214 15274 27238 15275
rect 27266 15274 27290 15275
rect 27318 15301 27342 15302
rect 27370 15301 27394 15302
rect 27318 15275 27322 15301
rect 27370 15275 27384 15301
rect 27318 15274 27342 15275
rect 27370 15274 27394 15275
rect 27422 15274 27446 15302
rect 27474 15274 27498 15302
rect 27526 15301 27535 15302
rect 27534 15275 27535 15301
rect 27526 15274 27535 15275
rect 27073 15269 27535 15274
rect 24486 15105 24514 15111
rect 24486 15079 24487 15105
rect 24513 15079 24514 15105
rect 24486 14322 24514 15079
rect 25326 15105 25354 15111
rect 25326 15079 25327 15105
rect 25353 15079 25354 15105
rect 25326 15049 25354 15079
rect 25326 15023 25327 15049
rect 25353 15023 25354 15049
rect 24573 14910 25035 14915
rect 24573 14909 24582 14910
rect 24573 14883 24574 14909
rect 24573 14882 24582 14883
rect 24610 14882 24634 14910
rect 24662 14882 24686 14910
rect 24714 14909 24738 14910
rect 24766 14909 24790 14910
rect 24724 14883 24738 14909
rect 24786 14883 24790 14909
rect 24714 14882 24738 14883
rect 24766 14882 24790 14883
rect 24818 14909 24842 14910
rect 24870 14909 24894 14910
rect 24818 14883 24822 14909
rect 24870 14883 24884 14909
rect 24818 14882 24842 14883
rect 24870 14882 24894 14883
rect 24922 14882 24946 14910
rect 24974 14882 24998 14910
rect 25026 14909 25035 14910
rect 25034 14883 25035 14909
rect 25026 14882 25035 14883
rect 24573 14877 25035 14882
rect 25046 14714 25074 14719
rect 25326 14714 25354 15023
rect 25438 14714 25466 14719
rect 25046 14713 25130 14714
rect 25046 14687 25047 14713
rect 25073 14687 25130 14713
rect 25046 14686 25130 14687
rect 25046 14681 25074 14686
rect 24486 13537 24514 14294
rect 24573 14126 25035 14131
rect 24573 14125 24582 14126
rect 24573 14099 24574 14125
rect 24573 14098 24582 14099
rect 24610 14098 24634 14126
rect 24662 14098 24686 14126
rect 24714 14125 24738 14126
rect 24766 14125 24790 14126
rect 24724 14099 24738 14125
rect 24786 14099 24790 14125
rect 24714 14098 24738 14099
rect 24766 14098 24790 14099
rect 24818 14125 24842 14126
rect 24870 14125 24894 14126
rect 24818 14099 24822 14125
rect 24870 14099 24884 14125
rect 24818 14098 24842 14099
rect 24870 14098 24894 14099
rect 24922 14098 24946 14126
rect 24974 14098 24998 14126
rect 25026 14125 25035 14126
rect 25034 14099 25035 14125
rect 25026 14098 25035 14099
rect 24573 14093 25035 14098
rect 25046 13930 25074 13935
rect 25102 13930 25130 14686
rect 25326 14713 25466 14714
rect 25326 14687 25327 14713
rect 25353 14687 25439 14713
rect 25465 14687 25466 14713
rect 25326 14686 25466 14687
rect 25326 14681 25354 14686
rect 25046 13929 25130 13930
rect 25046 13903 25047 13929
rect 25073 13903 25130 13929
rect 25046 13902 25130 13903
rect 25046 13897 25074 13902
rect 24486 13511 24487 13537
rect 24513 13511 24514 13537
rect 24486 13146 24514 13511
rect 24573 13342 25035 13347
rect 24573 13341 24582 13342
rect 24573 13315 24574 13341
rect 24573 13314 24582 13315
rect 24610 13314 24634 13342
rect 24662 13314 24686 13342
rect 24714 13341 24738 13342
rect 24766 13341 24790 13342
rect 24724 13315 24738 13341
rect 24786 13315 24790 13341
rect 24714 13314 24738 13315
rect 24766 13314 24790 13315
rect 24818 13341 24842 13342
rect 24870 13341 24894 13342
rect 24818 13315 24822 13341
rect 24870 13315 24884 13341
rect 24818 13314 24842 13315
rect 24870 13314 24894 13315
rect 24922 13314 24946 13342
rect 24974 13314 24998 13342
rect 25026 13341 25035 13342
rect 25034 13315 25035 13341
rect 25026 13314 25035 13315
rect 24573 13309 25035 13314
rect 24486 13113 24514 13118
rect 25046 13146 25074 13151
rect 25102 13146 25130 13902
rect 25382 14322 25410 14327
rect 25438 14322 25466 14686
rect 27073 14518 27535 14523
rect 27073 14517 27082 14518
rect 27073 14491 27074 14517
rect 27073 14490 27082 14491
rect 27110 14490 27134 14518
rect 27162 14490 27186 14518
rect 27214 14517 27238 14518
rect 27266 14517 27290 14518
rect 27224 14491 27238 14517
rect 27286 14491 27290 14517
rect 27214 14490 27238 14491
rect 27266 14490 27290 14491
rect 27318 14517 27342 14518
rect 27370 14517 27394 14518
rect 27318 14491 27322 14517
rect 27370 14491 27384 14517
rect 27318 14490 27342 14491
rect 27370 14490 27394 14491
rect 27422 14490 27446 14518
rect 27474 14490 27498 14518
rect 27526 14517 27535 14518
rect 27534 14491 27535 14517
rect 27526 14490 27535 14491
rect 27073 14485 27535 14490
rect 25382 14321 25466 14322
rect 25382 14295 25383 14321
rect 25409 14295 25466 14321
rect 25382 14294 25466 14295
rect 26726 14321 26754 14327
rect 26726 14295 26727 14321
rect 26753 14295 26754 14321
rect 25382 14266 25410 14294
rect 25382 13538 25410 14238
rect 25382 13481 25410 13510
rect 25382 13455 25383 13481
rect 25409 13455 25410 13481
rect 25382 13449 25410 13455
rect 25942 13985 25970 13991
rect 25942 13959 25943 13985
rect 25969 13959 25970 13985
rect 25942 13929 25970 13959
rect 25942 13903 25943 13929
rect 25969 13903 25970 13929
rect 25942 13538 25970 13903
rect 26222 13929 26250 13935
rect 26222 13903 26223 13929
rect 26249 13903 26250 13929
rect 26222 13874 26250 13903
rect 26222 13841 26250 13846
rect 26726 13874 26754 14295
rect 27398 13986 27426 13991
rect 27398 13929 27426 13958
rect 27398 13903 27399 13929
rect 27425 13903 27426 13929
rect 27398 13897 27426 13903
rect 25074 13118 25130 13146
rect 25942 13201 25970 13510
rect 26726 13538 26754 13846
rect 27073 13734 27535 13739
rect 27073 13733 27082 13734
rect 27073 13707 27074 13733
rect 27073 13706 27082 13707
rect 27110 13706 27134 13734
rect 27162 13706 27186 13734
rect 27214 13733 27238 13734
rect 27266 13733 27290 13734
rect 27224 13707 27238 13733
rect 27286 13707 27290 13733
rect 27214 13706 27238 13707
rect 27266 13706 27290 13707
rect 27318 13733 27342 13734
rect 27370 13733 27394 13734
rect 27318 13707 27322 13733
rect 27370 13707 27384 13733
rect 27318 13706 27342 13707
rect 27370 13706 27394 13707
rect 27422 13706 27446 13734
rect 27474 13706 27498 13734
rect 27526 13733 27535 13734
rect 27534 13707 27535 13733
rect 27526 13706 27535 13707
rect 27073 13701 27535 13706
rect 26726 13472 26754 13510
rect 25942 13175 25943 13201
rect 25969 13175 25970 13201
rect 25942 13146 25970 13175
rect 26502 13146 26530 13151
rect 25942 13145 26026 13146
rect 25942 13119 25943 13145
rect 25969 13119 26026 13145
rect 25942 13118 26026 13119
rect 25046 13099 25074 13118
rect 25942 13113 25970 13118
rect 24430 12782 24682 12810
rect 24374 12753 24402 12759
rect 24374 12727 24375 12753
rect 24401 12727 24402 12753
rect 24374 11970 24402 12727
rect 24654 12754 24682 12782
rect 24878 12754 24906 12759
rect 24654 12753 25130 12754
rect 24654 12727 24655 12753
rect 24681 12727 24879 12753
rect 24905 12727 25130 12753
rect 24654 12726 25130 12727
rect 24654 12721 24682 12726
rect 24878 12721 24906 12726
rect 24573 12558 25035 12563
rect 24573 12557 24582 12558
rect 24573 12531 24574 12557
rect 24573 12530 24582 12531
rect 24610 12530 24634 12558
rect 24662 12530 24686 12558
rect 24714 12557 24738 12558
rect 24766 12557 24790 12558
rect 24724 12531 24738 12557
rect 24786 12531 24790 12557
rect 24714 12530 24738 12531
rect 24766 12530 24790 12531
rect 24818 12557 24842 12558
rect 24870 12557 24894 12558
rect 24818 12531 24822 12557
rect 24870 12531 24884 12557
rect 24818 12530 24842 12531
rect 24870 12530 24894 12531
rect 24922 12530 24946 12558
rect 24974 12530 24998 12558
rect 25026 12557 25035 12558
rect 25034 12531 25035 12557
rect 25026 12530 25035 12531
rect 24573 12525 25035 12530
rect 24766 12361 24794 12367
rect 24766 12335 24767 12361
rect 24793 12335 24794 12361
rect 24766 11970 24794 12335
rect 25102 12362 25130 12726
rect 25214 12362 25242 12367
rect 25438 12362 25466 12367
rect 25102 12361 25466 12362
rect 25102 12335 25215 12361
rect 25241 12335 25439 12361
rect 25465 12335 25466 12361
rect 25102 12334 25466 12335
rect 25214 12329 25242 12334
rect 24374 11969 24794 11970
rect 24374 11943 24375 11969
rect 24401 11943 24794 11969
rect 24374 11942 24794 11943
rect 25158 11969 25186 11975
rect 25158 11943 25159 11969
rect 25185 11943 25186 11969
rect 24374 11578 24402 11942
rect 25158 11914 25186 11943
rect 25158 11802 25186 11886
rect 24573 11774 25035 11779
rect 24573 11773 24582 11774
rect 24573 11747 24574 11773
rect 24573 11746 24582 11747
rect 24610 11746 24634 11774
rect 24662 11746 24686 11774
rect 24714 11773 24738 11774
rect 24766 11773 24790 11774
rect 24724 11747 24738 11773
rect 24786 11747 24790 11773
rect 24714 11746 24738 11747
rect 24766 11746 24790 11747
rect 24818 11773 24842 11774
rect 24870 11773 24894 11774
rect 24818 11747 24822 11773
rect 24870 11747 24884 11773
rect 24818 11746 24842 11747
rect 24870 11746 24894 11747
rect 24922 11746 24946 11774
rect 24974 11746 24998 11774
rect 25026 11773 25035 11774
rect 25034 11747 25035 11773
rect 25026 11746 25035 11747
rect 24573 11741 25035 11746
rect 24766 11578 24794 11583
rect 24374 11577 24794 11578
rect 24374 11551 24767 11577
rect 24793 11551 24794 11577
rect 24374 11550 24794 11551
rect 24374 11185 24402 11550
rect 24766 11545 24794 11550
rect 24374 11159 24375 11185
rect 24401 11159 24402 11185
rect 24374 10906 24402 11159
rect 25158 11185 25186 11774
rect 25326 11578 25354 11583
rect 25438 11578 25466 12334
rect 25998 12362 26026 13118
rect 25326 11577 25466 11578
rect 25326 11551 25327 11577
rect 25353 11551 25439 11577
rect 25465 11551 25466 11577
rect 25326 11550 25466 11551
rect 25326 11545 25354 11550
rect 25158 11159 25159 11185
rect 25185 11159 25186 11185
rect 25158 11129 25186 11159
rect 25158 11103 25159 11129
rect 25185 11103 25186 11129
rect 25158 11097 25186 11103
rect 24573 10990 25035 10995
rect 24573 10989 24582 10990
rect 24573 10963 24574 10989
rect 24573 10962 24582 10963
rect 24610 10962 24634 10990
rect 24662 10962 24686 10990
rect 24714 10989 24738 10990
rect 24766 10989 24790 10990
rect 24724 10963 24738 10989
rect 24786 10963 24790 10989
rect 24714 10962 24738 10963
rect 24766 10962 24790 10963
rect 24818 10989 24842 10990
rect 24870 10989 24894 10990
rect 24818 10963 24822 10989
rect 24870 10963 24884 10989
rect 24818 10962 24842 10963
rect 24870 10962 24894 10963
rect 24922 10962 24946 10990
rect 24974 10962 24998 10990
rect 25026 10989 25035 10990
rect 25034 10963 25035 10989
rect 25026 10962 25035 10963
rect 24573 10957 25035 10962
rect 24374 10873 24402 10878
rect 24766 10906 24794 10911
rect 24766 10793 24794 10878
rect 24766 10767 24767 10793
rect 24793 10767 24794 10793
rect 24766 10761 24794 10767
rect 24486 10401 24514 10407
rect 24486 10375 24487 10401
rect 24513 10375 24514 10401
rect 24374 9617 24402 9623
rect 24374 9591 24375 9617
rect 24401 9591 24402 9617
rect 24374 9282 24402 9591
rect 24374 8833 24402 9254
rect 24486 9226 24514 10375
rect 25382 10401 25410 11550
rect 25438 11545 25466 11550
rect 25942 11802 25970 11807
rect 25942 10849 25970 11774
rect 25942 10823 25943 10849
rect 25969 10823 25970 10849
rect 25942 10793 25970 10823
rect 25942 10767 25943 10793
rect 25969 10767 25970 10793
rect 25942 10761 25970 10767
rect 25382 10375 25383 10401
rect 25409 10375 25410 10401
rect 25382 10346 25410 10375
rect 25382 10280 25410 10318
rect 25942 10346 25970 10351
rect 24573 10206 25035 10211
rect 24573 10205 24582 10206
rect 24573 10179 24574 10205
rect 24573 10178 24582 10179
rect 24610 10178 24634 10206
rect 24662 10178 24686 10206
rect 24714 10205 24738 10206
rect 24766 10205 24790 10206
rect 24724 10179 24738 10205
rect 24786 10179 24790 10205
rect 24714 10178 24738 10179
rect 24766 10178 24790 10179
rect 24818 10205 24842 10206
rect 24870 10205 24894 10206
rect 24818 10179 24822 10205
rect 24870 10179 24884 10205
rect 24818 10178 24842 10179
rect 24870 10178 24894 10179
rect 24922 10178 24946 10206
rect 24974 10178 24998 10206
rect 25026 10205 25035 10206
rect 25034 10179 25035 10205
rect 25026 10178 25035 10179
rect 24573 10173 25035 10178
rect 25942 10122 25970 10318
rect 25942 10065 25970 10094
rect 25942 10039 25943 10065
rect 25969 10039 25970 10065
rect 25046 10010 25074 10015
rect 25046 10009 25130 10010
rect 25046 9983 25047 10009
rect 25073 9983 25130 10009
rect 25046 9982 25130 9983
rect 25046 9977 25074 9982
rect 24654 9618 24682 9623
rect 24654 9571 24682 9590
rect 24878 9618 24906 9623
rect 24878 9571 24906 9590
rect 24573 9422 25035 9427
rect 24573 9421 24582 9422
rect 24573 9395 24574 9421
rect 24573 9394 24582 9395
rect 24610 9394 24634 9422
rect 24662 9394 24686 9422
rect 24714 9421 24738 9422
rect 24766 9421 24790 9422
rect 24724 9395 24738 9421
rect 24786 9395 24790 9421
rect 24714 9394 24738 9395
rect 24766 9394 24790 9395
rect 24818 9421 24842 9422
rect 24870 9421 24894 9422
rect 24818 9395 24822 9421
rect 24870 9395 24884 9421
rect 24818 9394 24842 9395
rect 24870 9394 24894 9395
rect 24922 9394 24946 9422
rect 24974 9394 24998 9422
rect 25026 9421 25035 9422
rect 25034 9395 25035 9421
rect 25026 9394 25035 9395
rect 24573 9389 25035 9394
rect 24486 9193 24514 9198
rect 24766 9282 24794 9287
rect 24766 9225 24794 9254
rect 24766 9199 24767 9225
rect 24793 9199 24794 9225
rect 24766 9193 24794 9199
rect 25102 9226 25130 9982
rect 25942 10009 25970 10039
rect 25942 9983 25943 10009
rect 25969 9983 25970 10009
rect 25942 9977 25970 9983
rect 25102 9193 25130 9198
rect 25158 9618 25186 9623
rect 25158 8890 25186 9590
rect 24374 8807 24375 8833
rect 24401 8807 24402 8833
rect 24374 8442 24402 8807
rect 25102 8862 25186 8890
rect 25214 9226 25242 9231
rect 25438 9226 25466 9231
rect 25214 9225 25466 9226
rect 25214 9199 25215 9225
rect 25241 9199 25439 9225
rect 25465 9199 25466 9225
rect 25214 9198 25466 9199
rect 24573 8638 25035 8643
rect 24573 8637 24582 8638
rect 24573 8611 24574 8637
rect 24573 8610 24582 8611
rect 24610 8610 24634 8638
rect 24662 8610 24686 8638
rect 24714 8637 24738 8638
rect 24766 8637 24790 8638
rect 24724 8611 24738 8637
rect 24786 8611 24790 8637
rect 24714 8610 24738 8611
rect 24766 8610 24790 8611
rect 24818 8637 24842 8638
rect 24870 8637 24894 8638
rect 24818 8611 24822 8637
rect 24870 8611 24884 8637
rect 24818 8610 24842 8611
rect 24870 8610 24894 8611
rect 24922 8610 24946 8638
rect 24974 8610 24998 8638
rect 25026 8637 25035 8638
rect 25034 8611 25035 8637
rect 25026 8610 25035 8611
rect 24573 8605 25035 8610
rect 24766 8442 24794 8447
rect 24374 8441 24794 8442
rect 24374 8415 24767 8441
rect 24793 8415 24794 8441
rect 24374 8414 24794 8415
rect 24374 8049 24402 8414
rect 24766 8409 24794 8414
rect 24878 8442 24906 8447
rect 24374 8023 24375 8049
rect 24401 8023 24402 8049
rect 24374 8017 24402 8023
rect 24766 8050 24794 8055
rect 24878 8050 24906 8414
rect 24766 8049 24906 8050
rect 24766 8023 24767 8049
rect 24793 8023 24879 8049
rect 24905 8023 24906 8049
rect 24766 8022 24906 8023
rect 24766 8017 24794 8022
rect 24878 8017 24906 8022
rect 24573 7854 25035 7859
rect 24573 7853 24582 7854
rect 24573 7827 24574 7853
rect 24573 7826 24582 7827
rect 24610 7826 24634 7854
rect 24662 7826 24686 7854
rect 24714 7853 24738 7854
rect 24766 7853 24790 7854
rect 24724 7827 24738 7853
rect 24786 7827 24790 7853
rect 24714 7826 24738 7827
rect 24766 7826 24790 7827
rect 24818 7853 24842 7854
rect 24870 7853 24894 7854
rect 24818 7827 24822 7853
rect 24870 7827 24884 7853
rect 24818 7826 24842 7827
rect 24870 7826 24894 7827
rect 24922 7826 24946 7854
rect 24974 7826 24998 7854
rect 25026 7853 25035 7854
rect 25034 7827 25035 7853
rect 25026 7826 25035 7827
rect 24573 7821 25035 7826
rect 24766 7657 24794 7663
rect 24766 7631 24767 7657
rect 24793 7631 24794 7657
rect 24374 7266 24402 7271
rect 24766 7266 24794 7631
rect 24374 7265 24794 7266
rect 24374 7239 24375 7265
rect 24401 7239 24794 7265
rect 24374 7238 24794 7239
rect 25102 7658 25130 8862
rect 25214 8833 25242 9198
rect 25438 9114 25466 9198
rect 25438 9081 25466 9086
rect 25998 9114 26026 12334
rect 26502 12362 26530 13118
rect 26782 13146 26810 13151
rect 26894 13146 26922 13151
rect 26782 13145 26922 13146
rect 26782 13119 26783 13145
rect 26809 13119 26895 13145
rect 26921 13119 26922 13145
rect 26782 13118 26922 13119
rect 26782 13113 26810 13118
rect 26726 12753 26754 12759
rect 26726 12727 26727 12753
rect 26753 12727 26754 12753
rect 26726 12362 26754 12727
rect 26502 12361 26754 12362
rect 26502 12335 26503 12361
rect 26529 12335 26754 12361
rect 26502 12334 26754 12335
rect 26894 12362 26922 13118
rect 27073 12950 27535 12955
rect 27073 12949 27082 12950
rect 27073 12923 27074 12949
rect 27073 12922 27082 12923
rect 27110 12922 27134 12950
rect 27162 12922 27186 12950
rect 27214 12949 27238 12950
rect 27266 12949 27290 12950
rect 27224 12923 27238 12949
rect 27286 12923 27290 12949
rect 27214 12922 27238 12923
rect 27266 12922 27290 12923
rect 27318 12949 27342 12950
rect 27370 12949 27394 12950
rect 27318 12923 27322 12949
rect 27370 12923 27384 12949
rect 27318 12922 27342 12923
rect 27370 12922 27394 12923
rect 27422 12922 27446 12950
rect 27474 12922 27498 12950
rect 27526 12949 27535 12950
rect 27534 12923 27535 12949
rect 27526 12922 27535 12923
rect 27073 12917 27535 12922
rect 26502 12329 26530 12334
rect 26894 12315 26922 12334
rect 27174 12754 27202 12759
rect 27398 12754 27426 12759
rect 27174 12753 27426 12754
rect 27174 12727 27175 12753
rect 27201 12727 27399 12753
rect 27425 12727 27426 12753
rect 27174 12726 27426 12727
rect 27174 12417 27202 12726
rect 27398 12721 27426 12726
rect 27174 12391 27175 12417
rect 27201 12391 27202 12417
rect 27174 12362 27202 12391
rect 27174 12329 27202 12334
rect 27073 12166 27535 12171
rect 27073 12165 27082 12166
rect 27073 12139 27074 12165
rect 27073 12138 27082 12139
rect 27110 12138 27134 12166
rect 27162 12138 27186 12166
rect 27214 12165 27238 12166
rect 27266 12165 27290 12166
rect 27224 12139 27238 12165
rect 27286 12139 27290 12165
rect 27214 12138 27238 12139
rect 27266 12138 27290 12139
rect 27318 12165 27342 12166
rect 27370 12165 27394 12166
rect 27318 12139 27322 12165
rect 27370 12139 27384 12165
rect 27318 12138 27342 12139
rect 27370 12138 27394 12139
rect 27422 12138 27446 12166
rect 27474 12138 27498 12166
rect 27526 12165 27535 12166
rect 27534 12139 27535 12165
rect 27526 12138 27535 12139
rect 27073 12133 27535 12138
rect 27006 11970 27034 11975
rect 27006 11923 27034 11942
rect 27566 11970 27594 18494
rect 29573 18046 30035 18051
rect 29573 18045 29582 18046
rect 29573 18019 29574 18045
rect 29573 18018 29582 18019
rect 29610 18018 29634 18046
rect 29662 18018 29686 18046
rect 29714 18045 29738 18046
rect 29766 18045 29790 18046
rect 29724 18019 29738 18045
rect 29786 18019 29790 18045
rect 29714 18018 29738 18019
rect 29766 18018 29790 18019
rect 29818 18045 29842 18046
rect 29870 18045 29894 18046
rect 29818 18019 29822 18045
rect 29870 18019 29884 18045
rect 29818 18018 29842 18019
rect 29870 18018 29894 18019
rect 29922 18018 29946 18046
rect 29974 18018 29998 18046
rect 30026 18045 30035 18046
rect 30034 18019 30035 18045
rect 30026 18018 30035 18019
rect 29573 18013 30035 18018
rect 29573 17262 30035 17267
rect 29573 17261 29582 17262
rect 29573 17235 29574 17261
rect 29573 17234 29582 17235
rect 29610 17234 29634 17262
rect 29662 17234 29686 17262
rect 29714 17261 29738 17262
rect 29766 17261 29790 17262
rect 29724 17235 29738 17261
rect 29786 17235 29790 17261
rect 29714 17234 29738 17235
rect 29766 17234 29790 17235
rect 29818 17261 29842 17262
rect 29870 17261 29894 17262
rect 29818 17235 29822 17261
rect 29870 17235 29884 17261
rect 29818 17234 29842 17235
rect 29870 17234 29894 17235
rect 29922 17234 29946 17262
rect 29974 17234 29998 17262
rect 30026 17261 30035 17262
rect 30034 17235 30035 17261
rect 30026 17234 30035 17235
rect 29573 17229 30035 17234
rect 29573 16478 30035 16483
rect 29573 16477 29582 16478
rect 29573 16451 29574 16477
rect 29573 16450 29582 16451
rect 29610 16450 29634 16478
rect 29662 16450 29686 16478
rect 29714 16477 29738 16478
rect 29766 16477 29790 16478
rect 29724 16451 29738 16477
rect 29786 16451 29790 16477
rect 29714 16450 29738 16451
rect 29766 16450 29790 16451
rect 29818 16477 29842 16478
rect 29870 16477 29894 16478
rect 29818 16451 29822 16477
rect 29870 16451 29884 16477
rect 29818 16450 29842 16451
rect 29870 16450 29894 16451
rect 29922 16450 29946 16478
rect 29974 16450 29998 16478
rect 30026 16477 30035 16478
rect 30034 16451 30035 16477
rect 30026 16450 30035 16451
rect 29573 16445 30035 16450
rect 29573 15694 30035 15699
rect 29573 15693 29582 15694
rect 29573 15667 29574 15693
rect 29573 15666 29582 15667
rect 29610 15666 29634 15694
rect 29662 15666 29686 15694
rect 29714 15693 29738 15694
rect 29766 15693 29790 15694
rect 29724 15667 29738 15693
rect 29786 15667 29790 15693
rect 29714 15666 29738 15667
rect 29766 15666 29790 15667
rect 29818 15693 29842 15694
rect 29870 15693 29894 15694
rect 29818 15667 29822 15693
rect 29870 15667 29884 15693
rect 29818 15666 29842 15667
rect 29870 15666 29894 15667
rect 29922 15666 29946 15694
rect 29974 15666 29998 15694
rect 30026 15693 30035 15694
rect 30034 15667 30035 15693
rect 30026 15666 30035 15667
rect 29573 15661 30035 15666
rect 29573 14910 30035 14915
rect 29573 14909 29582 14910
rect 29573 14883 29574 14909
rect 29573 14882 29582 14883
rect 29610 14882 29634 14910
rect 29662 14882 29686 14910
rect 29714 14909 29738 14910
rect 29766 14909 29790 14910
rect 29724 14883 29738 14909
rect 29786 14883 29790 14909
rect 29714 14882 29738 14883
rect 29766 14882 29790 14883
rect 29818 14909 29842 14910
rect 29870 14909 29894 14910
rect 29818 14883 29822 14909
rect 29870 14883 29884 14909
rect 29818 14882 29842 14883
rect 29870 14882 29894 14883
rect 29922 14882 29946 14910
rect 29974 14882 29998 14910
rect 30026 14909 30035 14910
rect 30034 14883 30035 14909
rect 30026 14882 30035 14883
rect 29573 14877 30035 14882
rect 27678 14321 27706 14327
rect 27678 14295 27679 14321
rect 27705 14295 27706 14321
rect 27678 14265 27706 14295
rect 27678 14239 27679 14265
rect 27705 14239 27706 14265
rect 27678 13986 27706 14239
rect 27678 13537 27706 13958
rect 27678 13511 27679 13537
rect 27705 13511 27706 13537
rect 27678 13482 27706 13511
rect 27678 13416 27706 13454
rect 28462 14321 28490 14327
rect 28462 14295 28463 14321
rect 28489 14295 28490 14321
rect 28462 13538 28490 14295
rect 29358 14321 29386 14327
rect 29358 14295 29359 14321
rect 29385 14295 29386 14321
rect 29358 14266 29386 14295
rect 28462 12753 28490 13510
rect 29246 14265 29386 14266
rect 29246 14239 29359 14265
rect 29385 14239 29386 14265
rect 29246 14238 29386 14239
rect 28462 12727 28463 12753
rect 28489 12727 28490 12753
rect 28462 12642 28490 12727
rect 28462 12609 28490 12614
rect 29022 13145 29050 13151
rect 29022 13119 29023 13145
rect 29049 13119 29050 13145
rect 29022 12642 29050 13119
rect 27622 12362 27650 12367
rect 27622 12082 27650 12334
rect 29022 12361 29050 12614
rect 29022 12335 29023 12361
rect 29049 12335 29050 12361
rect 29022 12329 29050 12335
rect 29246 12362 29274 14238
rect 29358 14233 29386 14238
rect 29573 14126 30035 14131
rect 29573 14125 29582 14126
rect 29573 14099 29574 14125
rect 29573 14098 29582 14099
rect 29610 14098 29634 14126
rect 29662 14098 29686 14126
rect 29714 14125 29738 14126
rect 29766 14125 29790 14126
rect 29724 14099 29738 14125
rect 29786 14099 29790 14125
rect 29714 14098 29738 14099
rect 29766 14098 29790 14099
rect 29818 14125 29842 14126
rect 29870 14125 29894 14126
rect 29818 14099 29822 14125
rect 29870 14099 29884 14125
rect 29818 14098 29842 14099
rect 29870 14098 29894 14099
rect 29922 14098 29946 14126
rect 29974 14098 29998 14126
rect 30026 14125 30035 14126
rect 30034 14099 30035 14125
rect 30026 14098 30035 14099
rect 29573 14093 30035 14098
rect 29358 13537 29386 13543
rect 29358 13511 29359 13537
rect 29385 13511 29386 13537
rect 29358 13482 29386 13511
rect 29302 13146 29330 13151
rect 29358 13146 29386 13454
rect 29573 13342 30035 13347
rect 29573 13341 29582 13342
rect 29573 13315 29574 13341
rect 29573 13314 29582 13315
rect 29610 13314 29634 13342
rect 29662 13314 29686 13342
rect 29714 13341 29738 13342
rect 29766 13341 29790 13342
rect 29724 13315 29738 13341
rect 29786 13315 29790 13341
rect 29714 13314 29738 13315
rect 29766 13314 29790 13315
rect 29818 13341 29842 13342
rect 29870 13341 29894 13342
rect 29818 13315 29822 13341
rect 29870 13315 29884 13341
rect 29818 13314 29842 13315
rect 29870 13314 29894 13315
rect 29922 13314 29946 13342
rect 29974 13314 29998 13342
rect 30026 13341 30035 13342
rect 30034 13315 30035 13341
rect 30026 13314 30035 13315
rect 29573 13309 30035 13314
rect 29414 13146 29442 13151
rect 29302 13145 29442 13146
rect 29302 13119 29303 13145
rect 29329 13119 29415 13145
rect 29441 13119 29442 13145
rect 29302 13118 29442 13119
rect 29302 13113 29330 13118
rect 29358 12753 29386 12759
rect 29358 12727 29359 12753
rect 29385 12727 29386 12753
rect 29358 12698 29386 12727
rect 29414 12698 29442 13118
rect 29358 12697 29442 12698
rect 29358 12671 29359 12697
rect 29385 12671 29442 12697
rect 29358 12670 29442 12671
rect 29358 12665 29386 12670
rect 29414 12362 29442 12670
rect 30478 12642 30506 12647
rect 29573 12558 30035 12563
rect 29573 12557 29582 12558
rect 29573 12531 29574 12557
rect 29573 12530 29582 12531
rect 29610 12530 29634 12558
rect 29662 12530 29686 12558
rect 29714 12557 29738 12558
rect 29766 12557 29790 12558
rect 29724 12531 29738 12557
rect 29786 12531 29790 12557
rect 29714 12530 29738 12531
rect 29766 12530 29790 12531
rect 29818 12557 29842 12558
rect 29870 12557 29894 12558
rect 29818 12531 29822 12557
rect 29870 12531 29884 12557
rect 29818 12530 29842 12531
rect 29870 12530 29894 12531
rect 29922 12530 29946 12558
rect 29974 12530 29998 12558
rect 30026 12557 30035 12558
rect 30034 12531 30035 12557
rect 30026 12530 30035 12531
rect 29573 12525 30035 12530
rect 29694 12417 29722 12423
rect 29694 12391 29695 12417
rect 29721 12391 29722 12417
rect 29470 12362 29498 12367
rect 29694 12362 29722 12391
rect 29414 12361 29722 12362
rect 29414 12335 29471 12361
rect 29497 12335 29722 12361
rect 29414 12334 29722 12335
rect 30478 12361 30506 12614
rect 31150 12417 31178 12423
rect 31150 12391 31151 12417
rect 31177 12391 31178 12417
rect 30478 12335 30479 12361
rect 30505 12335 30506 12361
rect 27622 12049 27650 12054
rect 29246 12082 29274 12334
rect 29246 12049 29274 12054
rect 28462 11970 28490 11975
rect 27566 11969 27706 11970
rect 27566 11943 27567 11969
rect 27593 11943 27706 11969
rect 27566 11942 27706 11943
rect 27566 11937 27594 11942
rect 27678 11913 27706 11942
rect 27678 11887 27679 11913
rect 27705 11887 27706 11913
rect 27678 11802 27706 11887
rect 26726 11578 26754 11583
rect 26950 11578 26978 11583
rect 26726 11577 26978 11578
rect 26726 11551 26727 11577
rect 26753 11551 26951 11577
rect 26977 11551 26978 11577
rect 26726 11550 26978 11551
rect 26726 11545 26754 11550
rect 26950 11074 26978 11550
rect 27398 11578 27426 11583
rect 27398 11531 27426 11550
rect 27073 11382 27535 11387
rect 27073 11381 27082 11382
rect 27073 11355 27074 11381
rect 27073 11354 27082 11355
rect 27110 11354 27134 11382
rect 27162 11354 27186 11382
rect 27214 11381 27238 11382
rect 27266 11381 27290 11382
rect 27224 11355 27238 11381
rect 27286 11355 27290 11381
rect 27214 11354 27238 11355
rect 27266 11354 27290 11355
rect 27318 11381 27342 11382
rect 27370 11381 27394 11382
rect 27318 11355 27322 11381
rect 27370 11355 27384 11381
rect 27318 11354 27342 11355
rect 27370 11354 27394 11355
rect 27422 11354 27446 11382
rect 27474 11354 27498 11382
rect 27526 11381 27535 11382
rect 27534 11355 27535 11381
rect 27526 11354 27535 11355
rect 27073 11349 27535 11354
rect 26950 11041 26978 11046
rect 27230 11185 27258 11191
rect 27230 11159 27231 11185
rect 27257 11159 27258 11185
rect 27230 11074 27258 11159
rect 27230 11041 27258 11046
rect 27454 11185 27482 11191
rect 27454 11159 27455 11185
rect 27481 11159 27482 11185
rect 27454 11074 27482 11159
rect 27678 11130 27706 11774
rect 27678 11097 27706 11102
rect 27846 11578 27874 11583
rect 27846 11185 27874 11550
rect 27846 11159 27847 11185
rect 27873 11159 27874 11185
rect 27454 11041 27482 11046
rect 26222 10906 26250 10911
rect 26222 10793 26250 10878
rect 26222 10767 26223 10793
rect 26249 10767 26250 10793
rect 26222 10761 26250 10767
rect 26726 10906 26754 10911
rect 26726 10402 26754 10878
rect 27286 10849 27314 10855
rect 27286 10823 27287 10849
rect 27313 10823 27314 10849
rect 27286 10794 27314 10823
rect 27286 10728 27314 10766
rect 27566 10794 27594 10799
rect 27073 10598 27535 10603
rect 27073 10597 27082 10598
rect 27073 10571 27074 10597
rect 27073 10570 27082 10571
rect 27110 10570 27134 10598
rect 27162 10570 27186 10598
rect 27214 10597 27238 10598
rect 27266 10597 27290 10598
rect 27224 10571 27238 10597
rect 27286 10571 27290 10597
rect 27214 10570 27238 10571
rect 27266 10570 27290 10571
rect 27318 10597 27342 10598
rect 27370 10597 27394 10598
rect 27318 10571 27322 10597
rect 27370 10571 27384 10597
rect 27318 10570 27342 10571
rect 27370 10570 27394 10571
rect 27422 10570 27446 10598
rect 27474 10570 27498 10598
rect 27526 10597 27535 10598
rect 27534 10571 27535 10597
rect 27526 10570 27535 10571
rect 27073 10565 27535 10570
rect 26726 10336 26754 10374
rect 27566 10402 27594 10766
rect 27566 10401 27706 10402
rect 27566 10375 27567 10401
rect 27593 10375 27706 10401
rect 27566 10374 27706 10375
rect 27566 10066 27594 10374
rect 27678 10345 27706 10374
rect 27678 10319 27679 10345
rect 27705 10319 27706 10345
rect 27678 10313 27706 10319
rect 27846 10234 27874 11159
rect 28462 11186 28490 11942
rect 28966 11969 28994 11975
rect 28966 11943 28967 11969
rect 28993 11943 28994 11969
rect 28966 11914 28994 11943
rect 29134 11914 29162 11919
rect 28966 11913 29162 11914
rect 28966 11887 29135 11913
rect 29161 11887 29162 11913
rect 28966 11886 29162 11887
rect 28462 11139 28490 11158
rect 28630 11185 28658 11191
rect 28630 11159 28631 11185
rect 28657 11159 28658 11185
rect 28630 11130 28658 11159
rect 28630 11097 28658 11102
rect 28854 11185 28882 11191
rect 28854 11159 28855 11185
rect 28881 11159 28882 11185
rect 28854 11130 28882 11159
rect 28854 11097 28882 11102
rect 28182 10401 28210 10407
rect 28182 10375 28183 10401
rect 28209 10375 28210 10401
rect 28182 10234 28210 10375
rect 27622 10206 28210 10234
rect 28406 10402 28434 10407
rect 27622 10094 27650 10206
rect 28406 10094 28434 10374
rect 28630 10346 28658 10351
rect 28630 10094 28658 10318
rect 27622 10066 27706 10094
rect 28406 10066 28490 10094
rect 26726 10010 26754 10015
rect 26950 10010 26978 10015
rect 26726 10009 26978 10010
rect 26726 9983 26727 10009
rect 26753 9983 26951 10009
rect 26977 9983 26978 10009
rect 26726 9982 26978 9983
rect 26726 9977 26754 9982
rect 26950 9618 26978 9982
rect 27398 10010 27426 10015
rect 27398 9963 27426 9982
rect 27073 9814 27535 9819
rect 27073 9813 27082 9814
rect 27073 9787 27074 9813
rect 27073 9786 27082 9787
rect 27110 9786 27134 9814
rect 27162 9786 27186 9814
rect 27214 9813 27238 9814
rect 27266 9813 27290 9814
rect 27224 9787 27238 9813
rect 27286 9787 27290 9813
rect 27214 9786 27238 9787
rect 27266 9786 27290 9787
rect 27318 9813 27342 9814
rect 27370 9813 27394 9814
rect 27318 9787 27322 9813
rect 27370 9787 27384 9813
rect 27318 9786 27342 9787
rect 27370 9786 27394 9787
rect 27422 9786 27446 9814
rect 27474 9786 27498 9814
rect 27526 9813 27535 9814
rect 27534 9787 27535 9813
rect 27526 9786 27535 9787
rect 27073 9781 27535 9786
rect 26950 9585 26978 9590
rect 27230 9618 27258 9623
rect 27230 9571 27258 9590
rect 27454 9618 27482 9623
rect 27454 9571 27482 9590
rect 27566 9450 27594 10038
rect 27398 9422 27594 9450
rect 27398 9281 27426 9422
rect 27398 9255 27399 9281
rect 27425 9255 27426 9281
rect 26502 9226 26530 9231
rect 26530 9198 26698 9226
rect 26502 9160 26530 9198
rect 25998 9081 26026 9086
rect 25214 8807 25215 8833
rect 25241 8807 25242 8833
rect 25158 8778 25186 8783
rect 25214 8778 25242 8807
rect 25158 8777 25242 8778
rect 25158 8751 25159 8777
rect 25185 8751 25242 8777
rect 25158 8750 25242 8751
rect 26670 8834 26698 9198
rect 27398 9225 27426 9255
rect 27398 9199 27399 9225
rect 27425 9199 27426 9225
rect 27398 9193 27426 9199
rect 27073 9030 27535 9035
rect 27073 9029 27082 9030
rect 27073 9003 27074 9029
rect 27073 9002 27082 9003
rect 27110 9002 27134 9030
rect 27162 9002 27186 9030
rect 27214 9029 27238 9030
rect 27266 9029 27290 9030
rect 27224 9003 27238 9029
rect 27286 9003 27290 9029
rect 27214 9002 27238 9003
rect 27266 9002 27290 9003
rect 27318 9029 27342 9030
rect 27370 9029 27394 9030
rect 27318 9003 27322 9029
rect 27370 9003 27384 9029
rect 27318 9002 27342 9003
rect 27370 9002 27394 9003
rect 27422 9002 27446 9030
rect 27474 9002 27498 9030
rect 27526 9029 27535 9030
rect 27534 9003 27535 9029
rect 27526 9002 27535 9003
rect 27073 8997 27535 9002
rect 27566 8946 27594 9422
rect 27510 8918 27594 8946
rect 26726 8834 26754 8839
rect 26670 8833 26754 8834
rect 26670 8807 26727 8833
rect 26753 8807 26754 8833
rect 26670 8806 26754 8807
rect 25158 8442 25186 8750
rect 25214 8442 25242 8447
rect 25186 8441 25242 8442
rect 25186 8415 25215 8441
rect 25241 8415 25242 8441
rect 25186 8414 25242 8415
rect 25158 8409 25186 8414
rect 25214 8409 25242 8414
rect 25438 8442 25466 8447
rect 25438 8395 25466 8414
rect 26222 8441 26250 8447
rect 26222 8415 26223 8441
rect 26249 8415 26250 8441
rect 25214 7658 25242 7663
rect 25438 7658 25466 7663
rect 25102 7657 25466 7658
rect 25102 7631 25215 7657
rect 25241 7631 25439 7657
rect 25465 7631 25466 7657
rect 25102 7630 25466 7631
rect 25102 7266 25130 7630
rect 25214 7625 25242 7630
rect 25438 7625 25466 7630
rect 26222 7657 26250 8415
rect 26222 7631 26223 7657
rect 26249 7631 26250 7657
rect 25158 7266 25186 7271
rect 25102 7265 25158 7266
rect 25102 7239 25103 7265
rect 25129 7239 25158 7265
rect 25102 7238 25158 7239
rect 24374 6482 24402 7238
rect 25102 7233 25130 7238
rect 25158 7210 25186 7238
rect 25158 7209 25242 7210
rect 25158 7183 25159 7209
rect 25185 7183 25242 7209
rect 25158 7182 25242 7183
rect 25158 7177 25186 7182
rect 24573 7070 25035 7075
rect 24573 7069 24582 7070
rect 24573 7043 24574 7069
rect 24573 7042 24582 7043
rect 24610 7042 24634 7070
rect 24662 7042 24686 7070
rect 24714 7069 24738 7070
rect 24766 7069 24790 7070
rect 24724 7043 24738 7069
rect 24786 7043 24790 7069
rect 24714 7042 24738 7043
rect 24766 7042 24790 7043
rect 24818 7069 24842 7070
rect 24870 7069 24894 7070
rect 24818 7043 24822 7069
rect 24870 7043 24884 7069
rect 24818 7042 24842 7043
rect 24870 7042 24894 7043
rect 24922 7042 24946 7070
rect 24974 7042 24998 7070
rect 25026 7069 25035 7070
rect 25034 7043 25035 7069
rect 25026 7042 25035 7043
rect 24573 7037 25035 7042
rect 24374 6090 24402 6454
rect 24766 6873 24794 6879
rect 24766 6847 24767 6873
rect 24793 6847 24794 6873
rect 24766 6482 24794 6847
rect 24766 6449 24794 6454
rect 25214 6874 25242 7182
rect 25214 6481 25242 6846
rect 25214 6455 25215 6481
rect 25241 6455 25242 6481
rect 25214 6425 25242 6455
rect 25214 6399 25215 6425
rect 25241 6399 25242 6425
rect 24573 6286 25035 6291
rect 24573 6285 24582 6286
rect 24573 6259 24574 6285
rect 24573 6258 24582 6259
rect 24610 6258 24634 6286
rect 24662 6258 24686 6286
rect 24714 6285 24738 6286
rect 24766 6285 24790 6286
rect 24724 6259 24738 6285
rect 24786 6259 24790 6285
rect 24714 6258 24738 6259
rect 24766 6258 24790 6259
rect 24818 6285 24842 6286
rect 24870 6285 24894 6286
rect 24818 6259 24822 6285
rect 24870 6259 24884 6285
rect 24818 6258 24842 6259
rect 24870 6258 24894 6259
rect 24922 6258 24946 6286
rect 24974 6258 24998 6286
rect 25026 6285 25035 6286
rect 25034 6259 25035 6285
rect 25026 6258 25035 6259
rect 24573 6253 25035 6258
rect 24374 5697 24402 6062
rect 24766 6090 24794 6095
rect 25214 6090 25242 6399
rect 24766 6043 24794 6062
rect 25158 6089 25242 6090
rect 25158 6063 25215 6089
rect 25241 6063 25242 6089
rect 25158 6062 25242 6063
rect 24374 5671 24375 5697
rect 24401 5671 24402 5697
rect 24374 5474 24402 5671
rect 25158 5697 25186 6062
rect 25214 6057 25242 6062
rect 25382 7154 25410 7159
rect 25158 5671 25159 5697
rect 25185 5671 25186 5697
rect 25158 5641 25186 5671
rect 25158 5615 25159 5641
rect 25185 5615 25186 5641
rect 25158 5609 25186 5615
rect 24573 5502 25035 5507
rect 24573 5501 24582 5502
rect 24573 5475 24574 5501
rect 24573 5474 24582 5475
rect 24610 5474 24634 5502
rect 24662 5474 24686 5502
rect 24714 5501 24738 5502
rect 24766 5501 24790 5502
rect 24724 5475 24738 5501
rect 24786 5475 24790 5501
rect 24714 5474 24738 5475
rect 24766 5474 24790 5475
rect 24818 5501 24842 5502
rect 24870 5501 24894 5502
rect 24818 5475 24822 5501
rect 24870 5475 24884 5501
rect 24818 5474 24842 5475
rect 24870 5474 24894 5475
rect 24922 5474 24946 5502
rect 24974 5474 24998 5502
rect 25026 5501 25035 5502
rect 25034 5475 25035 5501
rect 25026 5474 25035 5475
rect 24374 5446 24514 5474
rect 24573 5469 25035 5474
rect 24374 4913 24402 5446
rect 24374 4887 24375 4913
rect 24401 4887 24402 4913
rect 24374 4130 24402 4887
rect 24374 4083 24402 4102
rect 24430 5362 24458 5367
rect 24094 2226 24122 2478
rect 24374 3738 24402 3743
rect 24374 3345 24402 3710
rect 24374 3319 24375 3345
rect 24401 3319 24402 3345
rect 24374 2561 24402 3319
rect 24374 2535 24375 2561
rect 24401 2535 24402 2561
rect 24374 2450 24402 2535
rect 24374 2417 24402 2422
rect 24374 2226 24402 2231
rect 24430 2226 24458 5334
rect 24486 5306 24514 5446
rect 24766 5306 24794 5311
rect 24486 5305 24794 5306
rect 24486 5279 24767 5305
rect 24793 5279 24794 5305
rect 24486 5278 24794 5279
rect 24766 5273 24794 5278
rect 25214 5305 25242 5311
rect 25214 5279 25215 5305
rect 25241 5279 25242 5305
rect 25214 4913 25242 5279
rect 25214 4887 25215 4913
rect 25241 4887 25242 4913
rect 25214 4857 25242 4887
rect 25214 4831 25215 4857
rect 25241 4831 25242 4857
rect 24573 4718 25035 4723
rect 24573 4717 24582 4718
rect 24573 4691 24574 4717
rect 24573 4690 24582 4691
rect 24610 4690 24634 4718
rect 24662 4690 24686 4718
rect 24714 4717 24738 4718
rect 24766 4717 24790 4718
rect 24724 4691 24738 4717
rect 24786 4691 24790 4717
rect 24714 4690 24738 4691
rect 24766 4690 24790 4691
rect 24818 4717 24842 4718
rect 24870 4717 24894 4718
rect 24818 4691 24822 4717
rect 24870 4691 24884 4717
rect 24818 4690 24842 4691
rect 24870 4690 24894 4691
rect 24922 4690 24946 4718
rect 24974 4690 24998 4718
rect 25026 4717 25035 4718
rect 25034 4691 25035 4717
rect 25026 4690 25035 4691
rect 24573 4685 25035 4690
rect 24766 4521 24794 4527
rect 24766 4495 24767 4521
rect 24793 4495 24794 4521
rect 24654 4129 24682 4135
rect 24654 4103 24655 4129
rect 24681 4103 24682 4129
rect 24654 4074 24682 4103
rect 24766 4130 24794 4495
rect 25214 4521 25242 4831
rect 25214 4495 25215 4521
rect 25241 4495 25242 4521
rect 24766 4097 24794 4102
rect 24878 4129 24906 4135
rect 24878 4103 24879 4129
rect 24905 4103 24906 4129
rect 24654 4041 24682 4046
rect 24878 4074 24906 4103
rect 24878 4041 24906 4046
rect 25214 4074 25242 4495
rect 25382 4214 25410 7126
rect 25438 6874 25466 6879
rect 25438 6089 25466 6846
rect 25438 6063 25439 6089
rect 25465 6063 25466 6089
rect 25438 6057 25466 6063
rect 26222 6873 26250 7631
rect 26222 6847 26223 6873
rect 26249 6847 26250 6873
rect 26222 6090 26250 6847
rect 25942 5305 25970 5311
rect 25942 5279 25943 5305
rect 25969 5279 25970 5305
rect 25942 5250 25970 5279
rect 25942 4521 25970 5222
rect 25942 4495 25943 4521
rect 25969 4495 25970 4521
rect 25942 4489 25970 4495
rect 26054 5306 26082 5311
rect 26054 5194 26082 5278
rect 26222 5305 26250 6062
rect 26670 5978 26698 8806
rect 26726 8801 26754 8806
rect 27286 8834 27314 8839
rect 27510 8834 27538 8918
rect 27286 8833 27538 8834
rect 27286 8807 27287 8833
rect 27313 8807 27511 8833
rect 27537 8807 27538 8833
rect 27286 8806 27538 8807
rect 27286 8801 27314 8806
rect 27510 8801 27538 8806
rect 27174 8497 27202 8503
rect 27174 8471 27175 8497
rect 27201 8471 27202 8497
rect 26894 8442 26922 8447
rect 26670 5945 26698 5950
rect 26726 8049 26754 8055
rect 26726 8023 26727 8049
rect 26753 8023 26754 8049
rect 26726 7265 26754 8023
rect 26894 8050 26922 8414
rect 27174 8442 27202 8471
rect 27174 8409 27202 8414
rect 27073 8246 27535 8251
rect 27073 8245 27082 8246
rect 27073 8219 27074 8245
rect 27073 8218 27082 8219
rect 27110 8218 27134 8246
rect 27162 8218 27186 8246
rect 27214 8245 27238 8246
rect 27266 8245 27290 8246
rect 27224 8219 27238 8245
rect 27286 8219 27290 8245
rect 27214 8218 27238 8219
rect 27266 8218 27290 8219
rect 27318 8245 27342 8246
rect 27370 8245 27394 8246
rect 27318 8219 27322 8245
rect 27370 8219 27384 8245
rect 27318 8218 27342 8219
rect 27370 8218 27394 8219
rect 27422 8218 27446 8246
rect 27474 8218 27498 8246
rect 27526 8245 27535 8246
rect 27534 8219 27535 8245
rect 27526 8218 27535 8219
rect 27073 8213 27535 8218
rect 27174 8050 27202 8055
rect 27398 8050 27426 8055
rect 26894 8049 27426 8050
rect 26894 8023 27175 8049
rect 27201 8023 27399 8049
rect 27425 8023 27426 8049
rect 26894 8022 27426 8023
rect 26782 7658 26810 7663
rect 26894 7658 26922 8022
rect 27174 8017 27202 8022
rect 27398 8017 27426 8022
rect 26782 7657 26922 7658
rect 26782 7631 26783 7657
rect 26809 7631 26895 7657
rect 26921 7631 26922 7657
rect 26782 7630 26922 7631
rect 26782 7625 26810 7630
rect 26726 7239 26727 7265
rect 26753 7239 26754 7265
rect 26726 6874 26754 7239
rect 26726 6481 26754 6846
rect 26782 6874 26810 6879
rect 26894 6874 26922 7630
rect 27073 7462 27535 7467
rect 27073 7461 27082 7462
rect 27073 7435 27074 7461
rect 27073 7434 27082 7435
rect 27110 7434 27134 7462
rect 27162 7434 27186 7462
rect 27214 7461 27238 7462
rect 27266 7461 27290 7462
rect 27224 7435 27238 7461
rect 27286 7435 27290 7461
rect 27214 7434 27238 7435
rect 27266 7434 27290 7435
rect 27318 7461 27342 7462
rect 27370 7461 27394 7462
rect 27318 7435 27322 7461
rect 27370 7435 27384 7461
rect 27318 7434 27342 7435
rect 27370 7434 27394 7435
rect 27422 7434 27446 7462
rect 27474 7434 27498 7462
rect 27526 7461 27535 7462
rect 27534 7435 27535 7461
rect 27526 7434 27535 7435
rect 27073 7429 27535 7434
rect 27174 7266 27202 7271
rect 27174 7219 27202 7238
rect 27398 7266 27426 7271
rect 27398 7219 27426 7238
rect 26782 6873 26922 6874
rect 26782 6847 26783 6873
rect 26809 6847 26895 6873
rect 26921 6847 26922 6873
rect 26782 6846 26922 6847
rect 26782 6841 26810 6846
rect 26726 6455 26727 6481
rect 26753 6455 26754 6481
rect 26726 6090 26754 6455
rect 26726 5697 26754 6062
rect 26726 5671 26727 5697
rect 26753 5671 26754 5697
rect 26726 5665 26754 5671
rect 26894 6762 26922 6846
rect 26894 6146 26922 6734
rect 27006 7210 27034 7215
rect 27006 6594 27034 7182
rect 27678 7210 27706 10066
rect 27902 10010 27930 10015
rect 27902 9617 27930 9982
rect 27902 9591 27903 9617
rect 27929 9591 27930 9617
rect 27902 9562 27930 9591
rect 28462 9617 28490 10066
rect 28462 9591 28463 9617
rect 28489 9591 28490 9617
rect 27902 9529 27930 9534
rect 28406 9562 28434 9567
rect 28406 8834 28434 9534
rect 28462 9226 28490 9591
rect 28574 10066 28658 10094
rect 28966 10066 28994 11886
rect 29134 11881 29162 11886
rect 29022 11577 29050 11583
rect 29022 11551 29023 11577
rect 29049 11551 29050 11577
rect 29022 11186 29050 11551
rect 29470 11522 29498 12334
rect 29573 11774 30035 11779
rect 29573 11773 29582 11774
rect 29573 11747 29574 11773
rect 29573 11746 29582 11747
rect 29610 11746 29634 11774
rect 29662 11746 29686 11774
rect 29714 11773 29738 11774
rect 29766 11773 29790 11774
rect 29724 11747 29738 11773
rect 29786 11747 29790 11773
rect 29714 11746 29738 11747
rect 29766 11746 29790 11747
rect 29818 11773 29842 11774
rect 29870 11773 29894 11774
rect 29818 11747 29822 11773
rect 29870 11747 29884 11773
rect 29818 11746 29842 11747
rect 29870 11746 29894 11747
rect 29922 11746 29946 11774
rect 29974 11746 29998 11774
rect 30026 11773 30035 11774
rect 30034 11747 30035 11773
rect 30026 11746 30035 11747
rect 29573 11741 30035 11746
rect 29918 11633 29946 11639
rect 29918 11607 29919 11633
rect 29945 11607 29946 11633
rect 29918 11578 29946 11607
rect 30478 11578 30506 12335
rect 31094 12362 31122 12367
rect 31150 12362 31178 12391
rect 31122 12334 31178 12362
rect 31094 12315 31122 12334
rect 29918 11577 30114 11578
rect 29918 11551 29919 11577
rect 29945 11551 30114 11577
rect 29918 11550 30114 11551
rect 29918 11545 29946 11550
rect 29470 11489 29498 11494
rect 29022 10794 29050 11158
rect 29414 11410 29442 11415
rect 29414 11074 29442 11382
rect 29022 10793 29106 10794
rect 29022 10767 29023 10793
rect 29049 10767 29106 10793
rect 29022 10766 29106 10767
rect 29022 10761 29050 10766
rect 28574 10010 28602 10066
rect 28742 10010 28770 10015
rect 28574 9618 28602 9982
rect 28574 9585 28602 9590
rect 28630 10009 28770 10010
rect 28630 9983 28743 10009
rect 28769 9983 28770 10009
rect 28630 9982 28770 9983
rect 28462 9193 28490 9198
rect 28462 8834 28490 8839
rect 28406 8833 28490 8834
rect 28406 8807 28463 8833
rect 28489 8807 28490 8833
rect 28406 8806 28490 8807
rect 28462 8050 28490 8806
rect 28462 8003 28490 8022
rect 27678 7177 27706 7182
rect 28462 7265 28490 7271
rect 28462 7239 28463 7265
rect 28489 7239 28490 7265
rect 28462 6874 28490 7239
rect 27073 6678 27535 6683
rect 27073 6677 27082 6678
rect 27073 6651 27074 6677
rect 27073 6650 27082 6651
rect 27110 6650 27134 6678
rect 27162 6650 27186 6678
rect 27214 6677 27238 6678
rect 27266 6677 27290 6678
rect 27224 6651 27238 6677
rect 27286 6651 27290 6677
rect 27214 6650 27238 6651
rect 27266 6650 27290 6651
rect 27318 6677 27342 6678
rect 27370 6677 27394 6678
rect 27318 6651 27322 6677
rect 27370 6651 27384 6677
rect 27318 6650 27342 6651
rect 27370 6650 27394 6651
rect 27422 6650 27446 6678
rect 27474 6650 27498 6678
rect 27526 6677 27535 6678
rect 27534 6651 27535 6677
rect 27526 6650 27535 6651
rect 27073 6645 27535 6650
rect 27006 6566 27146 6594
rect 26894 6089 26922 6118
rect 26894 6063 26895 6089
rect 26921 6063 26922 6089
rect 26222 5279 26223 5305
rect 26249 5279 26250 5305
rect 26222 5273 26250 5279
rect 26782 5306 26810 5311
rect 26894 5306 26922 6063
rect 27118 6034 27146 6566
rect 27174 6482 27202 6487
rect 27398 6482 27426 6487
rect 27174 6481 27594 6482
rect 27174 6455 27175 6481
rect 27201 6455 27399 6481
rect 27425 6455 27594 6481
rect 27174 6454 27594 6455
rect 27174 6146 27202 6454
rect 27398 6449 27426 6454
rect 27174 6099 27202 6118
rect 26782 5305 26922 5306
rect 26782 5279 26783 5305
rect 26809 5279 26895 5305
rect 26921 5279 26922 5305
rect 26782 5278 26922 5279
rect 26782 5250 26810 5278
rect 26894 5273 26922 5278
rect 27006 6006 27146 6034
rect 26782 5217 26810 5222
rect 25214 4041 25242 4046
rect 25326 4186 25410 4214
rect 24573 3934 25035 3939
rect 24573 3933 24582 3934
rect 24573 3907 24574 3933
rect 24573 3906 24582 3907
rect 24610 3906 24634 3934
rect 24662 3906 24686 3934
rect 24714 3933 24738 3934
rect 24766 3933 24790 3934
rect 24724 3907 24738 3933
rect 24786 3907 24790 3933
rect 24714 3906 24738 3907
rect 24766 3906 24790 3907
rect 24818 3933 24842 3934
rect 24870 3933 24894 3934
rect 24818 3907 24822 3933
rect 24870 3907 24884 3933
rect 24818 3906 24842 3907
rect 24870 3906 24894 3907
rect 24922 3906 24946 3934
rect 24974 3906 24998 3934
rect 25026 3933 25035 3934
rect 25034 3907 25035 3933
rect 25026 3906 25035 3907
rect 24573 3901 25035 3906
rect 24766 3738 24794 3743
rect 24766 3691 24794 3710
rect 25214 3738 25242 3743
rect 25214 3345 25242 3710
rect 25214 3319 25215 3345
rect 25241 3319 25242 3345
rect 25214 3289 25242 3319
rect 25214 3263 25215 3289
rect 25241 3263 25242 3289
rect 24573 3150 25035 3155
rect 24573 3149 24582 3150
rect 24573 3123 24574 3149
rect 24573 3122 24582 3123
rect 24610 3122 24634 3150
rect 24662 3122 24686 3150
rect 24714 3149 24738 3150
rect 24766 3149 24790 3150
rect 24724 3123 24738 3149
rect 24786 3123 24790 3149
rect 24714 3122 24738 3123
rect 24766 3122 24790 3123
rect 24818 3149 24842 3150
rect 24870 3149 24894 3150
rect 24818 3123 24822 3149
rect 24870 3123 24884 3149
rect 24818 3122 24842 3123
rect 24870 3122 24894 3123
rect 24922 3122 24946 3150
rect 24974 3122 24998 3150
rect 25026 3149 25035 3150
rect 25034 3123 25035 3149
rect 25026 3122 25035 3123
rect 24573 3117 25035 3122
rect 24766 2953 24794 2959
rect 24766 2927 24767 2953
rect 24793 2927 24794 2953
rect 24654 2562 24682 2567
rect 24654 2515 24682 2534
rect 24094 2225 24234 2226
rect 24094 2199 24095 2225
rect 24121 2199 24234 2225
rect 24094 2198 24234 2199
rect 24094 2193 24122 2198
rect 23142 2169 23226 2170
rect 23142 2143 23143 2169
rect 23169 2143 23226 2169
rect 23142 2142 23226 2143
rect 24206 2169 24234 2198
rect 24374 2225 24458 2226
rect 24374 2199 24375 2225
rect 24401 2199 24458 2225
rect 24374 2198 24458 2199
rect 24486 2450 24514 2455
rect 24374 2193 24402 2198
rect 24206 2143 24207 2169
rect 24233 2143 24234 2169
rect 23142 1777 23170 2142
rect 24206 2137 24234 2143
rect 24486 2170 24514 2422
rect 24766 2450 24794 2927
rect 25214 2953 25242 3263
rect 25214 2927 25215 2953
rect 25241 2927 25242 2953
rect 24878 2562 24906 2567
rect 24878 2515 24906 2534
rect 25214 2562 25242 2927
rect 24766 2417 24794 2422
rect 24573 2366 25035 2371
rect 24573 2365 24582 2366
rect 24573 2339 24574 2365
rect 24573 2338 24582 2339
rect 24610 2338 24634 2366
rect 24662 2338 24686 2366
rect 24714 2365 24738 2366
rect 24766 2365 24790 2366
rect 24724 2339 24738 2365
rect 24786 2339 24790 2365
rect 24714 2338 24738 2339
rect 24766 2338 24790 2339
rect 24818 2365 24842 2366
rect 24870 2365 24894 2366
rect 24818 2339 24822 2365
rect 24870 2339 24884 2365
rect 24818 2338 24842 2339
rect 24870 2338 24894 2339
rect 24922 2338 24946 2366
rect 24974 2338 24998 2366
rect 25026 2365 25035 2366
rect 25034 2339 25035 2365
rect 25026 2338 25035 2339
rect 24573 2333 25035 2338
rect 23142 1751 23143 1777
rect 23169 1751 23170 1777
rect 23142 1666 23170 1751
rect 22918 1638 23170 1666
rect 24318 1890 24346 1895
rect 22918 1442 22946 1638
rect 22918 1409 22946 1414
rect 24318 400 24346 1862
rect 24486 1777 24514 2142
rect 24766 2170 24794 2175
rect 24766 2123 24794 2142
rect 25214 2169 25242 2534
rect 25214 2143 25215 2169
rect 25241 2143 25242 2169
rect 24486 1751 24487 1777
rect 24513 1751 24514 1777
rect 24486 1745 24514 1751
rect 25214 1778 25242 2143
rect 25326 1834 25354 4186
rect 25438 3738 25466 3743
rect 25438 3691 25466 3710
rect 26054 3346 26082 5166
rect 26726 4913 26754 4919
rect 26726 4887 26727 4913
rect 26753 4887 26754 4913
rect 26278 4521 26306 4527
rect 26278 4495 26279 4521
rect 26305 4495 26306 4521
rect 26278 3737 26306 4495
rect 26278 3711 26279 3737
rect 26305 3711 26306 3737
rect 26166 3346 26194 3351
rect 26054 3345 26194 3346
rect 26054 3319 26055 3345
rect 26081 3319 26167 3345
rect 26193 3319 26194 3345
rect 26054 3318 26194 3319
rect 26054 3313 26082 3318
rect 26166 3313 26194 3318
rect 25438 2953 25466 2959
rect 25438 2927 25439 2953
rect 25465 2927 25466 2953
rect 25438 2562 25466 2927
rect 25438 2169 25466 2534
rect 26278 2953 26306 3711
rect 26334 4522 26362 4527
rect 26334 3345 26362 4494
rect 26334 3319 26335 3345
rect 26361 3319 26362 3345
rect 26334 3313 26362 3319
rect 26726 4129 26754 4887
rect 26726 4103 26727 4129
rect 26753 4103 26754 4129
rect 26726 3345 26754 4103
rect 26726 3319 26727 3345
rect 26753 3319 26754 3345
rect 26278 2927 26279 2953
rect 26305 2927 26306 2953
rect 26278 2562 26306 2927
rect 26054 2506 26082 2511
rect 26054 2459 26082 2478
rect 26222 2506 26250 2511
rect 26222 2459 26250 2478
rect 25438 2143 25439 2169
rect 25465 2143 25466 2169
rect 25438 2137 25466 2143
rect 26222 2170 26250 2175
rect 26278 2170 26306 2534
rect 26726 2562 26754 3319
rect 26894 3738 26922 3743
rect 26894 3402 26922 3710
rect 26782 2954 26810 2959
rect 26894 2954 26922 3374
rect 26782 2953 26922 2954
rect 26782 2927 26783 2953
rect 26809 2927 26895 2953
rect 26921 2927 26922 2953
rect 26782 2926 26922 2927
rect 26782 2921 26810 2926
rect 26726 2515 26754 2534
rect 26894 2674 26922 2926
rect 26334 2505 26362 2511
rect 26334 2479 26335 2505
rect 26361 2479 26362 2505
rect 26334 2450 26362 2479
rect 26334 2417 26362 2422
rect 26250 2142 26306 2170
rect 26222 2123 26250 2142
rect 25326 1806 25466 1834
rect 25214 1777 25410 1778
rect 25214 1751 25215 1777
rect 25241 1751 25410 1777
rect 25214 1750 25410 1751
rect 25214 1745 25242 1750
rect 25382 1721 25410 1750
rect 25382 1695 25383 1721
rect 25409 1695 25410 1721
rect 25382 1689 25410 1695
rect 24573 1582 25035 1587
rect 24573 1581 24582 1582
rect 24573 1555 24574 1581
rect 24573 1554 24582 1555
rect 24610 1554 24634 1582
rect 24662 1554 24686 1582
rect 24714 1581 24738 1582
rect 24766 1581 24790 1582
rect 24724 1555 24738 1581
rect 24786 1555 24790 1581
rect 24714 1554 24738 1555
rect 24766 1554 24790 1555
rect 24818 1581 24842 1582
rect 24870 1581 24894 1582
rect 24818 1555 24822 1581
rect 24870 1555 24884 1581
rect 24818 1554 24842 1555
rect 24870 1554 24894 1555
rect 24922 1554 24946 1582
rect 24974 1554 24998 1582
rect 25026 1581 25035 1582
rect 25034 1555 25035 1581
rect 25026 1554 25035 1555
rect 24573 1549 25035 1554
rect 3542 350 3794 378
rect 3920 0 3976 400
rect 5376 0 5432 400
rect 6832 0 6888 400
rect 8288 0 8344 400
rect 9744 0 9800 400
rect 11200 0 11256 400
rect 12656 0 12712 400
rect 14112 0 14168 400
rect 15568 0 15624 400
rect 17024 0 17080 400
rect 18480 0 18536 400
rect 19936 0 19992 400
rect 21392 0 21448 400
rect 22848 0 22904 400
rect 24304 0 24360 400
rect 25438 378 25466 1806
rect 26278 1778 26306 2142
rect 26782 2170 26810 2175
rect 26894 2170 26922 2646
rect 26782 2169 26922 2170
rect 26782 2143 26783 2169
rect 26809 2143 26895 2169
rect 26921 2143 26922 2169
rect 26782 2142 26922 2143
rect 26782 2137 26810 2142
rect 26390 1778 26418 1783
rect 26278 1777 26418 1778
rect 26278 1751 26391 1777
rect 26417 1751 26418 1777
rect 26278 1750 26418 1751
rect 26390 1745 26418 1750
rect 26894 1777 26922 2142
rect 27006 1890 27034 6006
rect 27073 5894 27535 5899
rect 27073 5893 27082 5894
rect 27073 5867 27074 5893
rect 27073 5866 27082 5867
rect 27110 5866 27134 5894
rect 27162 5866 27186 5894
rect 27214 5893 27238 5894
rect 27266 5893 27290 5894
rect 27224 5867 27238 5893
rect 27286 5867 27290 5893
rect 27214 5866 27238 5867
rect 27266 5866 27290 5867
rect 27318 5893 27342 5894
rect 27370 5893 27394 5894
rect 27318 5867 27322 5893
rect 27370 5867 27384 5893
rect 27318 5866 27342 5867
rect 27370 5866 27394 5867
rect 27422 5866 27446 5894
rect 27474 5866 27498 5894
rect 27526 5893 27535 5894
rect 27534 5867 27535 5893
rect 27526 5866 27535 5867
rect 27073 5861 27535 5866
rect 27566 5698 27594 6454
rect 28462 6481 28490 6846
rect 28462 6455 28463 6481
rect 28489 6455 28490 6481
rect 28462 6449 28490 6455
rect 28070 5810 28098 5815
rect 27566 5697 27706 5698
rect 27566 5671 27567 5697
rect 27593 5671 27706 5697
rect 27566 5670 27706 5671
rect 27566 5665 27594 5670
rect 27678 5641 27706 5670
rect 27678 5615 27679 5641
rect 27705 5615 27706 5641
rect 27678 5609 27706 5615
rect 28070 5362 28098 5782
rect 28014 5306 28042 5311
rect 28070 5296 28098 5334
rect 28238 5697 28266 5703
rect 28238 5671 28239 5697
rect 28265 5671 28266 5697
rect 28182 5306 28210 5311
rect 28014 5194 28042 5278
rect 28182 5259 28210 5278
rect 27073 5110 27535 5115
rect 27073 5109 27082 5110
rect 27073 5083 27074 5109
rect 27073 5082 27082 5083
rect 27110 5082 27134 5110
rect 27162 5082 27186 5110
rect 27214 5109 27238 5110
rect 27266 5109 27290 5110
rect 27224 5083 27238 5109
rect 27286 5083 27290 5109
rect 27214 5082 27238 5083
rect 27266 5082 27290 5083
rect 27318 5109 27342 5110
rect 27370 5109 27394 5110
rect 27318 5083 27322 5109
rect 27370 5083 27384 5109
rect 27318 5082 27342 5083
rect 27370 5082 27394 5083
rect 27422 5082 27446 5110
rect 27474 5082 27498 5110
rect 27526 5109 27535 5110
rect 27534 5083 27535 5109
rect 27526 5082 27535 5083
rect 27073 5077 27535 5082
rect 27286 4914 27314 4919
rect 27398 4914 27426 4919
rect 27286 4913 27426 4914
rect 27286 4887 27287 4913
rect 27313 4887 27399 4913
rect 27425 4887 27426 4913
rect 27286 4886 27426 4887
rect 27286 4881 27314 4886
rect 27398 4577 27426 4886
rect 27398 4551 27399 4577
rect 27425 4551 27426 4577
rect 27398 4522 27426 4551
rect 27398 4521 27706 4522
rect 27398 4495 27399 4521
rect 27425 4495 27706 4521
rect 27398 4494 27706 4495
rect 27398 4489 27426 4494
rect 27073 4326 27535 4331
rect 27073 4325 27082 4326
rect 27073 4299 27074 4325
rect 27073 4298 27082 4299
rect 27110 4298 27134 4326
rect 27162 4298 27186 4326
rect 27214 4325 27238 4326
rect 27266 4325 27290 4326
rect 27224 4299 27238 4325
rect 27286 4299 27290 4325
rect 27214 4298 27238 4299
rect 27266 4298 27290 4299
rect 27318 4325 27342 4326
rect 27370 4325 27394 4326
rect 27318 4299 27322 4325
rect 27370 4299 27384 4325
rect 27318 4298 27342 4299
rect 27370 4298 27394 4299
rect 27422 4298 27446 4326
rect 27474 4298 27498 4326
rect 27526 4325 27535 4326
rect 27534 4299 27535 4325
rect 27526 4298 27535 4299
rect 27073 4293 27535 4298
rect 27174 4130 27202 4135
rect 27398 4130 27426 4135
rect 27174 4129 27398 4130
rect 27174 4103 27175 4129
rect 27201 4103 27398 4129
rect 27174 4102 27398 4103
rect 27174 3793 27202 4102
rect 27398 4064 27426 4102
rect 27678 4130 27706 4494
rect 27678 4097 27706 4102
rect 27174 3767 27175 3793
rect 27201 3767 27202 3793
rect 27174 3738 27202 3767
rect 27174 3705 27202 3710
rect 27073 3542 27535 3547
rect 27073 3541 27082 3542
rect 27073 3515 27074 3541
rect 27073 3514 27082 3515
rect 27110 3514 27134 3542
rect 27162 3514 27186 3542
rect 27214 3541 27238 3542
rect 27266 3541 27290 3542
rect 27224 3515 27238 3541
rect 27286 3515 27290 3541
rect 27214 3514 27238 3515
rect 27266 3514 27290 3515
rect 27318 3541 27342 3542
rect 27370 3541 27394 3542
rect 27318 3515 27322 3541
rect 27370 3515 27384 3541
rect 27318 3514 27342 3515
rect 27370 3514 27394 3515
rect 27422 3514 27446 3542
rect 27474 3514 27498 3542
rect 27526 3541 27535 3542
rect 27534 3515 27535 3541
rect 27526 3514 27535 3515
rect 27073 3509 27535 3514
rect 27174 3402 27202 3407
rect 27174 3345 27202 3374
rect 27174 3319 27175 3345
rect 27201 3319 27202 3345
rect 27174 3313 27202 3319
rect 27398 3402 27426 3407
rect 27398 3345 27426 3374
rect 27398 3319 27399 3345
rect 27425 3319 27426 3345
rect 27398 3313 27426 3319
rect 28014 2954 28042 5166
rect 28238 4914 28266 5671
rect 28406 5306 28434 5311
rect 28406 5259 28434 5278
rect 28238 4913 28434 4914
rect 28238 4887 28239 4913
rect 28265 4887 28434 4913
rect 28238 4886 28434 4887
rect 28238 4881 28266 4886
rect 28182 4606 28378 4634
rect 28182 4577 28210 4606
rect 28182 4551 28183 4577
rect 28209 4551 28210 4577
rect 28182 4545 28210 4551
rect 28126 4522 28154 4527
rect 28126 4475 28154 4494
rect 28350 4521 28378 4606
rect 28350 4495 28351 4521
rect 28377 4495 28378 4521
rect 28350 4298 28378 4495
rect 28182 4270 28378 4298
rect 28070 3738 28098 3743
rect 28182 3738 28210 4270
rect 28406 4214 28434 4886
rect 28238 4186 28434 4214
rect 28238 4130 28266 4186
rect 28462 4130 28490 4135
rect 28238 4129 28490 4130
rect 28238 4103 28463 4129
rect 28489 4103 28490 4129
rect 28238 4102 28490 4103
rect 28350 3794 28378 3799
rect 28294 3766 28350 3794
rect 28238 3738 28266 3743
rect 28070 3737 28266 3738
rect 28070 3711 28071 3737
rect 28097 3711 28239 3737
rect 28265 3711 28266 3737
rect 28070 3710 28266 3711
rect 28070 3705 28098 3710
rect 28182 2954 28210 2959
rect 28014 2953 28210 2954
rect 28014 2927 28015 2953
rect 28041 2927 28183 2953
rect 28209 2927 28210 2953
rect 28014 2926 28210 2927
rect 28014 2921 28042 2926
rect 28182 2921 28210 2926
rect 27073 2758 27535 2763
rect 27073 2757 27082 2758
rect 27073 2731 27074 2757
rect 27073 2730 27082 2731
rect 27110 2730 27134 2758
rect 27162 2730 27186 2758
rect 27214 2757 27238 2758
rect 27266 2757 27290 2758
rect 27224 2731 27238 2757
rect 27286 2731 27290 2757
rect 27214 2730 27238 2731
rect 27266 2730 27290 2731
rect 27318 2757 27342 2758
rect 27370 2757 27394 2758
rect 27318 2731 27322 2757
rect 27370 2731 27384 2757
rect 27318 2730 27342 2731
rect 27370 2730 27394 2731
rect 27422 2730 27446 2758
rect 27474 2730 27498 2758
rect 27526 2757 27535 2758
rect 27534 2731 27535 2757
rect 27526 2730 27535 2731
rect 27073 2725 27535 2730
rect 27174 2674 27202 2679
rect 27174 2562 27202 2646
rect 27398 2562 27426 2567
rect 27174 2561 27426 2562
rect 27174 2535 27175 2561
rect 27201 2535 27399 2561
rect 27425 2535 27426 2561
rect 27174 2534 27426 2535
rect 27174 2529 27202 2534
rect 27398 2529 27426 2534
rect 28238 2506 28266 3710
rect 28070 2226 28098 2231
rect 28238 2226 28266 2478
rect 28070 2225 28266 2226
rect 28070 2199 28071 2225
rect 28097 2199 28239 2225
rect 28265 2199 28266 2225
rect 28070 2198 28266 2199
rect 28070 2193 28098 2198
rect 28238 2193 28266 2198
rect 28294 2169 28322 3766
rect 28350 3747 28378 3766
rect 28462 3345 28490 4102
rect 28462 3319 28463 3345
rect 28489 3319 28490 3345
rect 28350 3290 28378 3295
rect 28350 3009 28378 3262
rect 28350 2983 28351 3009
rect 28377 2983 28378 3009
rect 28350 2977 28378 2983
rect 28462 2562 28490 3319
rect 28630 3066 28658 9982
rect 28742 9977 28770 9982
rect 28742 9618 28770 9623
rect 28966 9618 28994 10038
rect 28742 9617 28966 9618
rect 28742 9591 28743 9617
rect 28769 9591 28966 9617
rect 28742 9590 28966 9591
rect 28742 9585 28770 9590
rect 28966 9552 28994 9590
rect 29022 9226 29050 9231
rect 29022 9179 29050 9198
rect 29078 9114 29106 10766
rect 29134 10401 29162 10407
rect 29134 10375 29135 10401
rect 29161 10375 29162 10401
rect 29134 10346 29162 10375
rect 29134 10280 29162 10318
rect 29414 10094 29442 11046
rect 29573 10990 30035 10995
rect 29573 10989 29582 10990
rect 29573 10963 29574 10989
rect 29573 10962 29582 10963
rect 29610 10962 29634 10990
rect 29662 10962 29686 10990
rect 29714 10989 29738 10990
rect 29766 10989 29790 10990
rect 29724 10963 29738 10989
rect 29786 10963 29790 10989
rect 29714 10962 29738 10963
rect 29766 10962 29790 10963
rect 29818 10989 29842 10990
rect 29870 10989 29894 10990
rect 29818 10963 29822 10989
rect 29870 10963 29884 10989
rect 29818 10962 29842 10963
rect 29870 10962 29894 10963
rect 29922 10962 29946 10990
rect 29974 10962 29998 10990
rect 30026 10989 30035 10990
rect 30034 10963 30035 10989
rect 30026 10962 30035 10963
rect 29573 10957 30035 10962
rect 29918 10849 29946 10855
rect 29918 10823 29919 10849
rect 29945 10823 29946 10849
rect 29918 10794 29946 10823
rect 29918 10747 29946 10766
rect 30086 10794 30114 11550
rect 30478 11531 30506 11550
rect 30982 11969 31010 11975
rect 30982 11943 30983 11969
rect 31009 11943 31010 11969
rect 30982 11578 31010 11943
rect 31150 11970 31178 12334
rect 31374 11970 31402 11975
rect 31150 11969 31374 11970
rect 31150 11943 31151 11969
rect 31177 11943 31374 11969
rect 31150 11942 31374 11943
rect 31150 11937 31178 11942
rect 31374 11904 31402 11942
rect 30702 11242 30730 11247
rect 30702 11185 30730 11214
rect 30702 11159 30703 11185
rect 30729 11159 30730 11185
rect 30702 11153 30730 11159
rect 30982 11186 31010 11550
rect 31374 11633 31402 11639
rect 31374 11607 31375 11633
rect 31401 11607 31402 11633
rect 31374 11577 31402 11607
rect 31374 11551 31375 11577
rect 31401 11551 31402 11577
rect 31374 11522 31402 11551
rect 31374 11489 31402 11494
rect 31934 11410 31962 19614
rect 32270 19530 32298 19614
rect 32424 19600 32480 20000
rect 36974 19614 37282 19642
rect 32438 19530 32466 19600
rect 32270 19502 32466 19530
rect 32073 18438 32535 18443
rect 32073 18437 32082 18438
rect 32073 18411 32074 18437
rect 32073 18410 32082 18411
rect 32110 18410 32134 18438
rect 32162 18410 32186 18438
rect 32214 18437 32238 18438
rect 32266 18437 32290 18438
rect 32224 18411 32238 18437
rect 32286 18411 32290 18437
rect 32214 18410 32238 18411
rect 32266 18410 32290 18411
rect 32318 18437 32342 18438
rect 32370 18437 32394 18438
rect 32318 18411 32322 18437
rect 32370 18411 32384 18437
rect 32318 18410 32342 18411
rect 32370 18410 32394 18411
rect 32422 18410 32446 18438
rect 32474 18410 32498 18438
rect 32526 18437 32535 18438
rect 32534 18411 32535 18437
rect 32526 18410 32535 18411
rect 32073 18405 32535 18410
rect 34573 18046 35035 18051
rect 34573 18045 34582 18046
rect 34573 18019 34574 18045
rect 34573 18018 34582 18019
rect 34610 18018 34634 18046
rect 34662 18018 34686 18046
rect 34714 18045 34738 18046
rect 34766 18045 34790 18046
rect 34724 18019 34738 18045
rect 34786 18019 34790 18045
rect 34714 18018 34738 18019
rect 34766 18018 34790 18019
rect 34818 18045 34842 18046
rect 34870 18045 34894 18046
rect 34818 18019 34822 18045
rect 34870 18019 34884 18045
rect 34818 18018 34842 18019
rect 34870 18018 34894 18019
rect 34922 18018 34946 18046
rect 34974 18018 34998 18046
rect 35026 18045 35035 18046
rect 35034 18019 35035 18045
rect 35026 18018 35035 18019
rect 34573 18013 35035 18018
rect 32073 17654 32535 17659
rect 32073 17653 32082 17654
rect 32073 17627 32074 17653
rect 32073 17626 32082 17627
rect 32110 17626 32134 17654
rect 32162 17626 32186 17654
rect 32214 17653 32238 17654
rect 32266 17653 32290 17654
rect 32224 17627 32238 17653
rect 32286 17627 32290 17653
rect 32214 17626 32238 17627
rect 32266 17626 32290 17627
rect 32318 17653 32342 17654
rect 32370 17653 32394 17654
rect 32318 17627 32322 17653
rect 32370 17627 32384 17653
rect 32318 17626 32342 17627
rect 32370 17626 32394 17627
rect 32422 17626 32446 17654
rect 32474 17626 32498 17654
rect 32526 17653 32535 17654
rect 32534 17627 32535 17653
rect 32526 17626 32535 17627
rect 32073 17621 32535 17626
rect 34573 17262 35035 17267
rect 34573 17261 34582 17262
rect 34573 17235 34574 17261
rect 34573 17234 34582 17235
rect 34610 17234 34634 17262
rect 34662 17234 34686 17262
rect 34714 17261 34738 17262
rect 34766 17261 34790 17262
rect 34724 17235 34738 17261
rect 34786 17235 34790 17261
rect 34714 17234 34738 17235
rect 34766 17234 34790 17235
rect 34818 17261 34842 17262
rect 34870 17261 34894 17262
rect 34818 17235 34822 17261
rect 34870 17235 34884 17261
rect 34818 17234 34842 17235
rect 34870 17234 34894 17235
rect 34922 17234 34946 17262
rect 34974 17234 34998 17262
rect 35026 17261 35035 17262
rect 35034 17235 35035 17261
rect 35026 17234 35035 17235
rect 34573 17229 35035 17234
rect 32073 16870 32535 16875
rect 32073 16869 32082 16870
rect 32073 16843 32074 16869
rect 32073 16842 32082 16843
rect 32110 16842 32134 16870
rect 32162 16842 32186 16870
rect 32214 16869 32238 16870
rect 32266 16869 32290 16870
rect 32224 16843 32238 16869
rect 32286 16843 32290 16869
rect 32214 16842 32238 16843
rect 32266 16842 32290 16843
rect 32318 16869 32342 16870
rect 32370 16869 32394 16870
rect 32318 16843 32322 16869
rect 32370 16843 32384 16869
rect 32318 16842 32342 16843
rect 32370 16842 32394 16843
rect 32422 16842 32446 16870
rect 32474 16842 32498 16870
rect 32526 16869 32535 16870
rect 32534 16843 32535 16869
rect 32526 16842 32535 16843
rect 32073 16837 32535 16842
rect 34573 16478 35035 16483
rect 34573 16477 34582 16478
rect 34573 16451 34574 16477
rect 34573 16450 34582 16451
rect 34610 16450 34634 16478
rect 34662 16450 34686 16478
rect 34714 16477 34738 16478
rect 34766 16477 34790 16478
rect 34724 16451 34738 16477
rect 34786 16451 34790 16477
rect 34714 16450 34738 16451
rect 34766 16450 34790 16451
rect 34818 16477 34842 16478
rect 34870 16477 34894 16478
rect 34818 16451 34822 16477
rect 34870 16451 34884 16477
rect 34818 16450 34842 16451
rect 34870 16450 34894 16451
rect 34922 16450 34946 16478
rect 34974 16450 34998 16478
rect 35026 16477 35035 16478
rect 35034 16451 35035 16477
rect 35026 16450 35035 16451
rect 34573 16445 35035 16450
rect 32073 16086 32535 16091
rect 32073 16085 32082 16086
rect 32073 16059 32074 16085
rect 32073 16058 32082 16059
rect 32110 16058 32134 16086
rect 32162 16058 32186 16086
rect 32214 16085 32238 16086
rect 32266 16085 32290 16086
rect 32224 16059 32238 16085
rect 32286 16059 32290 16085
rect 32214 16058 32238 16059
rect 32266 16058 32290 16059
rect 32318 16085 32342 16086
rect 32370 16085 32394 16086
rect 32318 16059 32322 16085
rect 32370 16059 32384 16085
rect 32318 16058 32342 16059
rect 32370 16058 32394 16059
rect 32422 16058 32446 16086
rect 32474 16058 32498 16086
rect 32526 16085 32535 16086
rect 32534 16059 32535 16085
rect 32526 16058 32535 16059
rect 32073 16053 32535 16058
rect 34573 15694 35035 15699
rect 34573 15693 34582 15694
rect 34573 15667 34574 15693
rect 34573 15666 34582 15667
rect 34610 15666 34634 15694
rect 34662 15666 34686 15694
rect 34714 15693 34738 15694
rect 34766 15693 34790 15694
rect 34724 15667 34738 15693
rect 34786 15667 34790 15693
rect 34714 15666 34738 15667
rect 34766 15666 34790 15667
rect 34818 15693 34842 15694
rect 34870 15693 34894 15694
rect 34818 15667 34822 15693
rect 34870 15667 34884 15693
rect 34818 15666 34842 15667
rect 34870 15666 34894 15667
rect 34922 15666 34946 15694
rect 34974 15666 34998 15694
rect 35026 15693 35035 15694
rect 35034 15667 35035 15693
rect 35026 15666 35035 15667
rect 34573 15661 35035 15666
rect 32073 15302 32535 15307
rect 32073 15301 32082 15302
rect 32073 15275 32074 15301
rect 32073 15274 32082 15275
rect 32110 15274 32134 15302
rect 32162 15274 32186 15302
rect 32214 15301 32238 15302
rect 32266 15301 32290 15302
rect 32224 15275 32238 15301
rect 32286 15275 32290 15301
rect 32214 15274 32238 15275
rect 32266 15274 32290 15275
rect 32318 15301 32342 15302
rect 32370 15301 32394 15302
rect 32318 15275 32322 15301
rect 32370 15275 32384 15301
rect 32318 15274 32342 15275
rect 32370 15274 32394 15275
rect 32422 15274 32446 15302
rect 32474 15274 32498 15302
rect 32526 15301 32535 15302
rect 32534 15275 32535 15301
rect 32526 15274 32535 15275
rect 32073 15269 32535 15274
rect 34573 14910 35035 14915
rect 34573 14909 34582 14910
rect 34573 14883 34574 14909
rect 34573 14882 34582 14883
rect 34610 14882 34634 14910
rect 34662 14882 34686 14910
rect 34714 14909 34738 14910
rect 34766 14909 34790 14910
rect 34724 14883 34738 14909
rect 34786 14883 34790 14909
rect 34714 14882 34738 14883
rect 34766 14882 34790 14883
rect 34818 14909 34842 14910
rect 34870 14909 34894 14910
rect 34818 14883 34822 14909
rect 34870 14883 34884 14909
rect 34818 14882 34842 14883
rect 34870 14882 34894 14883
rect 34922 14882 34946 14910
rect 34974 14882 34998 14910
rect 35026 14909 35035 14910
rect 35034 14883 35035 14909
rect 35026 14882 35035 14883
rect 34573 14877 35035 14882
rect 32073 14518 32535 14523
rect 32073 14517 32082 14518
rect 32073 14491 32074 14517
rect 32073 14490 32082 14491
rect 32110 14490 32134 14518
rect 32162 14490 32186 14518
rect 32214 14517 32238 14518
rect 32266 14517 32290 14518
rect 32224 14491 32238 14517
rect 32286 14491 32290 14517
rect 32214 14490 32238 14491
rect 32266 14490 32290 14491
rect 32318 14517 32342 14518
rect 32370 14517 32394 14518
rect 32318 14491 32322 14517
rect 32370 14491 32384 14517
rect 32318 14490 32342 14491
rect 32370 14490 32394 14491
rect 32422 14490 32446 14518
rect 32474 14490 32498 14518
rect 32526 14517 32535 14518
rect 32534 14491 32535 14517
rect 32526 14490 32535 14491
rect 32073 14485 32535 14490
rect 34573 14126 35035 14131
rect 34573 14125 34582 14126
rect 34573 14099 34574 14125
rect 34573 14098 34582 14099
rect 34610 14098 34634 14126
rect 34662 14098 34686 14126
rect 34714 14125 34738 14126
rect 34766 14125 34790 14126
rect 34724 14099 34738 14125
rect 34786 14099 34790 14125
rect 34714 14098 34738 14099
rect 34766 14098 34790 14099
rect 34818 14125 34842 14126
rect 34870 14125 34894 14126
rect 34818 14099 34822 14125
rect 34870 14099 34884 14125
rect 34818 14098 34842 14099
rect 34870 14098 34894 14099
rect 34922 14098 34946 14126
rect 34974 14098 34998 14126
rect 35026 14125 35035 14126
rect 35034 14099 35035 14125
rect 35026 14098 35035 14099
rect 34573 14093 35035 14098
rect 32073 13734 32535 13739
rect 32073 13733 32082 13734
rect 32073 13707 32074 13733
rect 32073 13706 32082 13707
rect 32110 13706 32134 13734
rect 32162 13706 32186 13734
rect 32214 13733 32238 13734
rect 32266 13733 32290 13734
rect 32224 13707 32238 13733
rect 32286 13707 32290 13733
rect 32214 13706 32238 13707
rect 32266 13706 32290 13707
rect 32318 13733 32342 13734
rect 32370 13733 32394 13734
rect 32318 13707 32322 13733
rect 32370 13707 32384 13733
rect 32318 13706 32342 13707
rect 32370 13706 32394 13707
rect 32422 13706 32446 13734
rect 32474 13706 32498 13734
rect 32526 13733 32535 13734
rect 32534 13707 32535 13733
rect 32526 13706 32535 13707
rect 32073 13701 32535 13706
rect 34573 13342 35035 13347
rect 34573 13341 34582 13342
rect 34573 13315 34574 13341
rect 34573 13314 34582 13315
rect 34610 13314 34634 13342
rect 34662 13314 34686 13342
rect 34714 13341 34738 13342
rect 34766 13341 34790 13342
rect 34724 13315 34738 13341
rect 34786 13315 34790 13341
rect 34714 13314 34738 13315
rect 34766 13314 34790 13315
rect 34818 13341 34842 13342
rect 34870 13341 34894 13342
rect 34818 13315 34822 13341
rect 34870 13315 34884 13341
rect 34818 13314 34842 13315
rect 34870 13314 34894 13315
rect 34922 13314 34946 13342
rect 34974 13314 34998 13342
rect 35026 13341 35035 13342
rect 35034 13315 35035 13341
rect 35026 13314 35035 13315
rect 34573 13309 35035 13314
rect 32073 12950 32535 12955
rect 32073 12949 32082 12950
rect 32073 12923 32074 12949
rect 32073 12922 32082 12923
rect 32110 12922 32134 12950
rect 32162 12922 32186 12950
rect 32214 12949 32238 12950
rect 32266 12949 32290 12950
rect 32224 12923 32238 12949
rect 32286 12923 32290 12949
rect 32214 12922 32238 12923
rect 32266 12922 32290 12923
rect 32318 12949 32342 12950
rect 32370 12949 32394 12950
rect 32318 12923 32322 12949
rect 32370 12923 32384 12949
rect 32318 12922 32342 12923
rect 32370 12922 32394 12923
rect 32422 12922 32446 12950
rect 32474 12922 32498 12950
rect 32526 12949 32535 12950
rect 32534 12923 32535 12949
rect 32526 12922 32535 12923
rect 32073 12917 32535 12922
rect 34573 12558 35035 12563
rect 34573 12557 34582 12558
rect 34573 12531 34574 12557
rect 34573 12530 34582 12531
rect 34610 12530 34634 12558
rect 34662 12530 34686 12558
rect 34714 12557 34738 12558
rect 34766 12557 34790 12558
rect 34724 12531 34738 12557
rect 34786 12531 34790 12557
rect 34714 12530 34738 12531
rect 34766 12530 34790 12531
rect 34818 12557 34842 12558
rect 34870 12557 34894 12558
rect 34818 12531 34822 12557
rect 34870 12531 34884 12557
rect 34818 12530 34842 12531
rect 34870 12530 34894 12531
rect 34922 12530 34946 12558
rect 34974 12530 34998 12558
rect 35026 12557 35035 12558
rect 35034 12531 35035 12557
rect 35026 12530 35035 12531
rect 34573 12525 35035 12530
rect 32073 12166 32535 12171
rect 32073 12165 32082 12166
rect 32073 12139 32074 12165
rect 32073 12138 32082 12139
rect 32110 12138 32134 12166
rect 32162 12138 32186 12166
rect 32214 12165 32238 12166
rect 32266 12165 32290 12166
rect 32224 12139 32238 12165
rect 32286 12139 32290 12165
rect 32214 12138 32238 12139
rect 32266 12138 32290 12139
rect 32318 12165 32342 12166
rect 32370 12165 32394 12166
rect 32318 12139 32322 12165
rect 32370 12139 32384 12165
rect 32318 12138 32342 12139
rect 32370 12138 32394 12139
rect 32422 12138 32446 12166
rect 32474 12138 32498 12166
rect 32526 12165 32535 12166
rect 32534 12139 32535 12165
rect 32526 12138 32535 12139
rect 32073 12133 32535 12138
rect 32158 11970 32186 11975
rect 31934 11377 31962 11382
rect 31990 11969 32186 11970
rect 31990 11943 32159 11969
rect 32185 11943 32186 11969
rect 31990 11942 32186 11943
rect 31990 11578 32018 11942
rect 32158 11937 32186 11942
rect 32830 11970 32858 11975
rect 32830 11923 32858 11942
rect 33110 11970 33138 11975
rect 33110 11913 33138 11942
rect 33110 11887 33111 11913
rect 33137 11887 33138 11913
rect 31934 11242 31962 11247
rect 30982 11153 31010 11158
rect 31262 11186 31290 11191
rect 31374 11186 31402 11191
rect 31262 11185 31402 11186
rect 31262 11159 31263 11185
rect 31289 11159 31375 11185
rect 31401 11159 31402 11185
rect 31262 11158 31402 11159
rect 31262 11153 31290 11158
rect 31094 11130 31122 11135
rect 31094 10850 31122 11102
rect 31150 10850 31178 10855
rect 31094 10849 31178 10850
rect 31094 10823 31151 10849
rect 31177 10823 31178 10849
rect 31094 10822 31178 10823
rect 30086 10761 30114 10766
rect 30254 10793 30282 10799
rect 30254 10767 30255 10793
rect 30281 10767 30282 10793
rect 30254 10738 30282 10767
rect 31094 10793 31122 10822
rect 31094 10767 31095 10793
rect 31121 10767 31122 10793
rect 31094 10761 31122 10767
rect 30254 10705 30282 10710
rect 30702 10738 30730 10743
rect 30702 10402 30730 10710
rect 30702 10336 30730 10374
rect 29573 10206 30035 10211
rect 29573 10205 29582 10206
rect 29573 10179 29574 10205
rect 29573 10178 29582 10179
rect 29610 10178 29634 10206
rect 29662 10178 29686 10206
rect 29714 10205 29738 10206
rect 29766 10205 29790 10206
rect 29724 10179 29738 10205
rect 29786 10179 29790 10205
rect 29714 10178 29738 10179
rect 29766 10178 29790 10179
rect 29818 10205 29842 10206
rect 29870 10205 29894 10206
rect 29818 10179 29822 10205
rect 29870 10179 29884 10205
rect 29818 10178 29842 10179
rect 29870 10178 29894 10179
rect 29922 10178 29946 10206
rect 29974 10178 29998 10206
rect 30026 10205 30035 10206
rect 30034 10179 30035 10205
rect 30026 10178 30035 10179
rect 29573 10173 30035 10178
rect 31150 10094 31178 10822
rect 31374 10794 31402 11158
rect 31374 10094 31402 10766
rect 31934 10458 31962 11214
rect 31934 10425 31962 10430
rect 29414 10066 29498 10094
rect 29302 10010 29330 10015
rect 29414 10010 29442 10015
rect 29330 10009 29442 10010
rect 29330 9983 29415 10009
rect 29441 9983 29442 10009
rect 29330 9982 29442 9983
rect 29302 9944 29330 9982
rect 29078 9081 29106 9086
rect 29358 8833 29386 9982
rect 29414 9977 29442 9982
rect 29414 9618 29442 9623
rect 29414 9282 29442 9590
rect 29414 9225 29442 9254
rect 29414 9199 29415 9225
rect 29441 9199 29442 9225
rect 29414 9193 29442 9199
rect 29358 8807 29359 8833
rect 29385 8807 29386 8833
rect 29358 8777 29386 8807
rect 29358 8751 29359 8777
rect 29385 8751 29386 8777
rect 29358 8498 29386 8751
rect 29358 8465 29386 8470
rect 29022 8441 29050 8447
rect 29022 8415 29023 8441
rect 29049 8415 29050 8441
rect 29022 8050 29050 8415
rect 29022 7657 29050 8022
rect 29358 8050 29386 8055
rect 29470 8050 29498 10066
rect 31094 10066 31122 10071
rect 31150 10066 31234 10094
rect 30422 10009 30450 10015
rect 30422 9983 30423 10009
rect 30449 9983 30450 10009
rect 29573 9422 30035 9427
rect 29573 9421 29582 9422
rect 29573 9395 29574 9421
rect 29573 9394 29582 9395
rect 29610 9394 29634 9422
rect 29662 9394 29686 9422
rect 29714 9421 29738 9422
rect 29766 9421 29790 9422
rect 29724 9395 29738 9421
rect 29786 9395 29790 9421
rect 29714 9394 29738 9395
rect 29766 9394 29790 9395
rect 29818 9421 29842 9422
rect 29870 9421 29894 9422
rect 29818 9395 29822 9421
rect 29870 9395 29884 9421
rect 29818 9394 29842 9395
rect 29870 9394 29894 9395
rect 29922 9394 29946 9422
rect 29974 9394 29998 9422
rect 30026 9421 30035 9422
rect 30034 9395 30035 9421
rect 30026 9394 30035 9395
rect 29573 9389 30035 9394
rect 29694 9282 29722 9287
rect 29694 9235 29722 9254
rect 30422 9225 30450 9983
rect 31094 10009 31122 10038
rect 31094 9983 31095 10009
rect 31121 9983 31122 10009
rect 31038 9730 31066 9735
rect 30982 9617 31010 9623
rect 30982 9591 30983 9617
rect 31009 9591 31010 9617
rect 30422 9199 30423 9225
rect 30449 9199 30450 9225
rect 30422 9114 30450 9199
rect 30422 9081 30450 9086
rect 30478 9226 30506 9231
rect 29573 8638 30035 8643
rect 29573 8637 29582 8638
rect 29573 8611 29574 8637
rect 29573 8610 29582 8611
rect 29610 8610 29634 8638
rect 29662 8610 29686 8638
rect 29714 8637 29738 8638
rect 29766 8637 29790 8638
rect 29724 8611 29738 8637
rect 29786 8611 29790 8637
rect 29714 8610 29738 8611
rect 29766 8610 29790 8611
rect 29818 8637 29842 8638
rect 29870 8637 29894 8638
rect 29818 8611 29822 8637
rect 29870 8611 29884 8637
rect 29818 8610 29842 8611
rect 29870 8610 29894 8611
rect 29922 8610 29946 8638
rect 29974 8610 29998 8638
rect 30026 8637 30035 8638
rect 30034 8611 30035 8637
rect 30026 8610 30035 8611
rect 29573 8605 30035 8610
rect 29918 8498 29946 8503
rect 29918 8441 29946 8470
rect 29918 8415 29919 8441
rect 29945 8415 29946 8441
rect 29918 8409 29946 8415
rect 30478 8441 30506 9198
rect 30478 8415 30479 8441
rect 30505 8415 30506 8441
rect 29358 8049 29498 8050
rect 29358 8023 29359 8049
rect 29385 8023 29498 8049
rect 29358 8022 29498 8023
rect 29358 7994 29386 8022
rect 29022 7631 29023 7657
rect 29049 7631 29050 7657
rect 28742 6874 28770 6879
rect 28742 6827 28770 6846
rect 29022 6818 29050 7631
rect 29302 7993 29386 7994
rect 29302 7967 29359 7993
rect 29385 7967 29386 7993
rect 29302 7966 29386 7967
rect 29302 7657 29330 7966
rect 29358 7961 29386 7966
rect 29302 7631 29303 7657
rect 29329 7631 29330 7657
rect 29302 7625 29330 7631
rect 29470 7657 29498 8022
rect 29573 7854 30035 7859
rect 29573 7853 29582 7854
rect 29573 7827 29574 7853
rect 29573 7826 29582 7827
rect 29610 7826 29634 7854
rect 29662 7826 29686 7854
rect 29714 7853 29738 7854
rect 29766 7853 29790 7854
rect 29724 7827 29738 7853
rect 29786 7827 29790 7853
rect 29714 7826 29738 7827
rect 29766 7826 29790 7827
rect 29818 7853 29842 7854
rect 29870 7853 29894 7854
rect 29818 7827 29822 7853
rect 29870 7827 29884 7853
rect 29818 7826 29842 7827
rect 29870 7826 29894 7827
rect 29922 7826 29946 7854
rect 29974 7826 29998 7854
rect 30026 7853 30035 7854
rect 30034 7827 30035 7853
rect 30026 7826 30035 7827
rect 29573 7821 30035 7826
rect 29470 7631 29471 7657
rect 29497 7631 29498 7657
rect 29022 6785 29050 6790
rect 29190 7265 29218 7271
rect 29190 7239 29191 7265
rect 29217 7239 29218 7265
rect 29190 7209 29218 7239
rect 29190 7183 29191 7209
rect 29217 7183 29218 7209
rect 29190 6873 29218 7183
rect 29190 6847 29191 6873
rect 29217 6847 29218 6873
rect 28686 6762 28714 6767
rect 28686 6482 28714 6734
rect 29190 6762 29218 6847
rect 29190 6729 29218 6734
rect 29414 6873 29442 6879
rect 29414 6847 29415 6873
rect 29441 6847 29442 6873
rect 29414 6762 29442 6847
rect 29470 6874 29498 7631
rect 30478 7657 30506 8415
rect 30982 9114 31010 9591
rect 30982 8833 31010 9086
rect 31038 8890 31066 9702
rect 31094 9618 31122 9983
rect 31150 9618 31178 9623
rect 31122 9617 31178 9618
rect 31122 9591 31151 9617
rect 31177 9591 31178 9617
rect 31122 9590 31178 9591
rect 31094 9585 31122 9590
rect 31038 8857 31066 8862
rect 30982 8807 30983 8833
rect 31009 8807 31010 8833
rect 30982 8442 31010 8807
rect 30982 8409 31010 8414
rect 31150 8497 31178 9590
rect 31206 9282 31234 10066
rect 31262 10066 31402 10094
rect 31654 10401 31682 10407
rect 31654 10375 31655 10401
rect 31681 10375 31682 10401
rect 31654 10345 31682 10375
rect 31654 10319 31655 10345
rect 31681 10319 31682 10345
rect 31262 10019 31290 10038
rect 31374 9618 31402 9623
rect 31374 9571 31402 9590
rect 31374 9282 31402 9287
rect 31654 9282 31682 10319
rect 31990 10066 32018 11550
rect 32774 11578 32802 11583
rect 32774 11531 32802 11550
rect 32073 11382 32535 11387
rect 32073 11381 32082 11382
rect 32073 11355 32074 11381
rect 32073 11354 32082 11355
rect 32110 11354 32134 11382
rect 32162 11354 32186 11382
rect 32214 11381 32238 11382
rect 32266 11381 32290 11382
rect 32224 11355 32238 11381
rect 32286 11355 32290 11381
rect 32214 11354 32238 11355
rect 32266 11354 32290 11355
rect 32318 11381 32342 11382
rect 32370 11381 32394 11382
rect 32318 11355 32322 11381
rect 32370 11355 32384 11381
rect 32318 11354 32342 11355
rect 32370 11354 32394 11355
rect 32422 11354 32446 11382
rect 32474 11354 32498 11382
rect 32526 11381 32535 11382
rect 32534 11355 32535 11381
rect 32526 11354 32535 11355
rect 32073 11349 32535 11354
rect 32438 11186 32466 11191
rect 32438 11139 32466 11158
rect 32998 11186 33026 11191
rect 32998 10793 33026 11158
rect 33110 11185 33138 11887
rect 34573 11774 35035 11779
rect 34573 11773 34582 11774
rect 34573 11747 34574 11773
rect 34573 11746 34582 11747
rect 34610 11746 34634 11774
rect 34662 11746 34686 11774
rect 34714 11773 34738 11774
rect 34766 11773 34790 11774
rect 34724 11747 34738 11773
rect 34786 11747 34790 11773
rect 34714 11746 34738 11747
rect 34766 11746 34790 11747
rect 34818 11773 34842 11774
rect 34870 11773 34894 11774
rect 34818 11747 34822 11773
rect 34870 11747 34884 11773
rect 34818 11746 34842 11747
rect 34870 11746 34894 11747
rect 34922 11746 34946 11774
rect 34974 11746 34998 11774
rect 35026 11773 35035 11774
rect 35034 11747 35035 11773
rect 35026 11746 35035 11747
rect 34573 11741 35035 11746
rect 33110 11159 33111 11185
rect 33137 11159 33138 11185
rect 33110 11130 33138 11159
rect 33110 11064 33138 11102
rect 33894 11633 33922 11639
rect 33894 11607 33895 11633
rect 33921 11607 33922 11633
rect 33894 11577 33922 11607
rect 33894 11551 33895 11577
rect 33921 11551 33922 11577
rect 33894 11130 33922 11551
rect 35294 11522 35322 11527
rect 34958 11186 34986 11191
rect 34958 11139 34986 11158
rect 35238 11186 35266 11191
rect 35294 11186 35322 11494
rect 36974 11298 37002 19614
rect 37254 19530 37282 19614
rect 37408 19600 37464 20000
rect 37422 19530 37450 19600
rect 37254 19502 37450 19530
rect 37073 18438 37535 18443
rect 37073 18437 37082 18438
rect 37073 18411 37074 18437
rect 37073 18410 37082 18411
rect 37110 18410 37134 18438
rect 37162 18410 37186 18438
rect 37214 18437 37238 18438
rect 37266 18437 37290 18438
rect 37224 18411 37238 18437
rect 37286 18411 37290 18437
rect 37214 18410 37238 18411
rect 37266 18410 37290 18411
rect 37318 18437 37342 18438
rect 37370 18437 37394 18438
rect 37318 18411 37322 18437
rect 37370 18411 37384 18437
rect 37318 18410 37342 18411
rect 37370 18410 37394 18411
rect 37422 18410 37446 18438
rect 37474 18410 37498 18438
rect 37526 18437 37535 18438
rect 37534 18411 37535 18437
rect 37526 18410 37535 18411
rect 37073 18405 37535 18410
rect 37073 17654 37535 17659
rect 37073 17653 37082 17654
rect 37073 17627 37074 17653
rect 37073 17626 37082 17627
rect 37110 17626 37134 17654
rect 37162 17626 37186 17654
rect 37214 17653 37238 17654
rect 37266 17653 37290 17654
rect 37224 17627 37238 17653
rect 37286 17627 37290 17653
rect 37214 17626 37238 17627
rect 37266 17626 37290 17627
rect 37318 17653 37342 17654
rect 37370 17653 37394 17654
rect 37318 17627 37322 17653
rect 37370 17627 37384 17653
rect 37318 17626 37342 17627
rect 37370 17626 37394 17627
rect 37422 17626 37446 17654
rect 37474 17626 37498 17654
rect 37526 17653 37535 17654
rect 37534 17627 37535 17653
rect 37526 17626 37535 17627
rect 37073 17621 37535 17626
rect 37073 16870 37535 16875
rect 37073 16869 37082 16870
rect 37073 16843 37074 16869
rect 37073 16842 37082 16843
rect 37110 16842 37134 16870
rect 37162 16842 37186 16870
rect 37214 16869 37238 16870
rect 37266 16869 37290 16870
rect 37224 16843 37238 16869
rect 37286 16843 37290 16869
rect 37214 16842 37238 16843
rect 37266 16842 37290 16843
rect 37318 16869 37342 16870
rect 37370 16869 37394 16870
rect 37318 16843 37322 16869
rect 37370 16843 37384 16869
rect 37318 16842 37342 16843
rect 37370 16842 37394 16843
rect 37422 16842 37446 16870
rect 37474 16842 37498 16870
rect 37526 16869 37535 16870
rect 37534 16843 37535 16869
rect 37526 16842 37535 16843
rect 37073 16837 37535 16842
rect 37073 16086 37535 16091
rect 37073 16085 37082 16086
rect 37073 16059 37074 16085
rect 37073 16058 37082 16059
rect 37110 16058 37134 16086
rect 37162 16058 37186 16086
rect 37214 16085 37238 16086
rect 37266 16085 37290 16086
rect 37224 16059 37238 16085
rect 37286 16059 37290 16085
rect 37214 16058 37238 16059
rect 37266 16058 37290 16059
rect 37318 16085 37342 16086
rect 37370 16085 37394 16086
rect 37318 16059 37322 16085
rect 37370 16059 37384 16085
rect 37318 16058 37342 16059
rect 37370 16058 37394 16059
rect 37422 16058 37446 16086
rect 37474 16058 37498 16086
rect 37526 16085 37535 16086
rect 37534 16059 37535 16085
rect 37526 16058 37535 16059
rect 37073 16053 37535 16058
rect 37073 15302 37535 15307
rect 37073 15301 37082 15302
rect 37073 15275 37074 15301
rect 37073 15274 37082 15275
rect 37110 15274 37134 15302
rect 37162 15274 37186 15302
rect 37214 15301 37238 15302
rect 37266 15301 37290 15302
rect 37224 15275 37238 15301
rect 37286 15275 37290 15301
rect 37214 15274 37238 15275
rect 37266 15274 37290 15275
rect 37318 15301 37342 15302
rect 37370 15301 37394 15302
rect 37318 15275 37322 15301
rect 37370 15275 37384 15301
rect 37318 15274 37342 15275
rect 37370 15274 37394 15275
rect 37422 15274 37446 15302
rect 37474 15274 37498 15302
rect 37526 15301 37535 15302
rect 37534 15275 37535 15301
rect 37526 15274 37535 15275
rect 37073 15269 37535 15274
rect 37073 14518 37535 14523
rect 37073 14517 37082 14518
rect 37073 14491 37074 14517
rect 37073 14490 37082 14491
rect 37110 14490 37134 14518
rect 37162 14490 37186 14518
rect 37214 14517 37238 14518
rect 37266 14517 37290 14518
rect 37224 14491 37238 14517
rect 37286 14491 37290 14517
rect 37214 14490 37238 14491
rect 37266 14490 37290 14491
rect 37318 14517 37342 14518
rect 37370 14517 37394 14518
rect 37318 14491 37322 14517
rect 37370 14491 37384 14517
rect 37318 14490 37342 14491
rect 37370 14490 37394 14491
rect 37422 14490 37446 14518
rect 37474 14490 37498 14518
rect 37526 14517 37535 14518
rect 37534 14491 37535 14517
rect 37526 14490 37535 14491
rect 37073 14485 37535 14490
rect 37073 13734 37535 13739
rect 37073 13733 37082 13734
rect 37073 13707 37074 13733
rect 37073 13706 37082 13707
rect 37110 13706 37134 13734
rect 37162 13706 37186 13734
rect 37214 13733 37238 13734
rect 37266 13733 37290 13734
rect 37224 13707 37238 13733
rect 37286 13707 37290 13733
rect 37214 13706 37238 13707
rect 37266 13706 37290 13707
rect 37318 13733 37342 13734
rect 37370 13733 37394 13734
rect 37318 13707 37322 13733
rect 37370 13707 37384 13733
rect 37318 13706 37342 13707
rect 37370 13706 37394 13707
rect 37422 13706 37446 13734
rect 37474 13706 37498 13734
rect 37526 13733 37535 13734
rect 37534 13707 37535 13733
rect 37526 13706 37535 13707
rect 37073 13701 37535 13706
rect 37073 12950 37535 12955
rect 37073 12949 37082 12950
rect 37073 12923 37074 12949
rect 37073 12922 37082 12923
rect 37110 12922 37134 12950
rect 37162 12922 37186 12950
rect 37214 12949 37238 12950
rect 37266 12949 37290 12950
rect 37224 12923 37238 12949
rect 37286 12923 37290 12949
rect 37214 12922 37238 12923
rect 37266 12922 37290 12923
rect 37318 12949 37342 12950
rect 37370 12949 37394 12950
rect 37318 12923 37322 12949
rect 37370 12923 37384 12949
rect 37318 12922 37342 12923
rect 37370 12922 37394 12923
rect 37422 12922 37446 12950
rect 37474 12922 37498 12950
rect 37526 12949 37535 12950
rect 37534 12923 37535 12949
rect 37526 12922 37535 12923
rect 37073 12917 37535 12922
rect 37073 12166 37535 12171
rect 37073 12165 37082 12166
rect 37073 12139 37074 12165
rect 37073 12138 37082 12139
rect 37110 12138 37134 12166
rect 37162 12138 37186 12166
rect 37214 12165 37238 12166
rect 37266 12165 37290 12166
rect 37224 12139 37238 12165
rect 37286 12139 37290 12165
rect 37214 12138 37238 12139
rect 37266 12138 37290 12139
rect 37318 12165 37342 12166
rect 37370 12165 37394 12166
rect 37318 12139 37322 12165
rect 37370 12139 37384 12165
rect 37318 12138 37342 12139
rect 37370 12138 37394 12139
rect 37422 12138 37446 12166
rect 37474 12138 37498 12166
rect 37526 12165 37535 12166
rect 37534 12139 37535 12165
rect 37526 12138 37535 12139
rect 37073 12133 37535 12138
rect 37073 11382 37535 11387
rect 37073 11381 37082 11382
rect 37073 11355 37074 11381
rect 37073 11354 37082 11355
rect 37110 11354 37134 11382
rect 37162 11354 37186 11382
rect 37214 11381 37238 11382
rect 37266 11381 37290 11382
rect 37224 11355 37238 11381
rect 37286 11355 37290 11381
rect 37214 11354 37238 11355
rect 37266 11354 37290 11355
rect 37318 11381 37342 11382
rect 37370 11381 37394 11382
rect 37318 11355 37322 11381
rect 37370 11355 37384 11381
rect 37318 11354 37342 11355
rect 37370 11354 37394 11355
rect 37422 11354 37446 11382
rect 37474 11354 37498 11382
rect 37526 11381 37535 11382
rect 37534 11355 37535 11381
rect 37526 11354 37535 11355
rect 37073 11349 37535 11354
rect 36974 11270 37058 11298
rect 35238 11185 35322 11186
rect 35238 11159 35239 11185
rect 35265 11159 35322 11185
rect 35238 11158 35322 11159
rect 35238 11153 35266 11158
rect 32998 10767 32999 10793
rect 33025 10767 33026 10793
rect 32073 10598 32535 10603
rect 32073 10597 32082 10598
rect 32073 10571 32074 10597
rect 32073 10570 32082 10571
rect 32110 10570 32134 10598
rect 32162 10570 32186 10598
rect 32214 10597 32238 10598
rect 32266 10597 32290 10598
rect 32224 10571 32238 10597
rect 32286 10571 32290 10597
rect 32214 10570 32238 10571
rect 32266 10570 32290 10571
rect 32318 10597 32342 10598
rect 32370 10597 32394 10598
rect 32318 10571 32322 10597
rect 32370 10571 32384 10597
rect 32318 10570 32342 10571
rect 32370 10570 32394 10571
rect 32422 10570 32446 10598
rect 32474 10570 32498 10598
rect 32526 10597 32535 10598
rect 32534 10571 32535 10597
rect 32526 10570 32535 10571
rect 32073 10565 32535 10570
rect 32158 10458 32186 10463
rect 32158 10401 32186 10430
rect 32158 10375 32159 10401
rect 32185 10375 32186 10401
rect 32158 10369 32186 10375
rect 32606 10402 32634 10407
rect 31990 9730 32018 10038
rect 32073 9814 32535 9819
rect 32073 9813 32082 9814
rect 32073 9787 32074 9813
rect 32073 9786 32082 9787
rect 32110 9786 32134 9814
rect 32162 9786 32186 9814
rect 32214 9813 32238 9814
rect 32266 9813 32290 9814
rect 32224 9787 32238 9813
rect 32286 9787 32290 9813
rect 32214 9786 32238 9787
rect 32266 9786 32290 9787
rect 32318 9813 32342 9814
rect 32370 9813 32394 9814
rect 32318 9787 32322 9813
rect 32370 9787 32384 9813
rect 32318 9786 32342 9787
rect 32370 9786 32394 9787
rect 32422 9786 32446 9814
rect 32474 9786 32498 9814
rect 32526 9813 32535 9814
rect 32534 9787 32535 9813
rect 32526 9786 32535 9787
rect 32073 9781 32535 9786
rect 31990 9697 32018 9702
rect 31206 9281 31682 9282
rect 31206 9255 31375 9281
rect 31401 9255 31682 9281
rect 31206 9254 31682 9255
rect 32438 9618 32466 9623
rect 32606 9618 32634 10374
rect 32438 9617 32634 9618
rect 32438 9591 32439 9617
rect 32465 9591 32634 9617
rect 32438 9590 32634 9591
rect 32774 10009 32802 10015
rect 32774 9983 32775 10009
rect 32801 9983 32802 10009
rect 31150 8471 31151 8497
rect 31177 8471 31178 8497
rect 31150 8441 31178 8471
rect 31150 8415 31151 8441
rect 31177 8415 31178 8441
rect 30478 7631 30479 7657
rect 30505 7631 30506 7657
rect 30478 7546 30506 7631
rect 30982 8049 31010 8055
rect 30982 8023 30983 8049
rect 31009 8023 31010 8049
rect 30982 7546 31010 8023
rect 31150 8050 31178 8415
rect 31374 9225 31402 9254
rect 31374 9199 31375 9225
rect 31401 9199 31402 9225
rect 31374 8386 31402 9199
rect 32438 9226 32466 9590
rect 32438 9193 32466 9198
rect 32774 9170 32802 9983
rect 32774 9137 32802 9142
rect 32830 9618 32858 9623
rect 32073 9030 32535 9035
rect 32073 9029 32082 9030
rect 32073 9003 32074 9029
rect 32073 9002 32082 9003
rect 32110 9002 32134 9030
rect 32162 9002 32186 9030
rect 32214 9029 32238 9030
rect 32266 9029 32290 9030
rect 32224 9003 32238 9029
rect 32286 9003 32290 9029
rect 32214 9002 32238 9003
rect 32266 9002 32290 9003
rect 32318 9029 32342 9030
rect 32370 9029 32394 9030
rect 32318 9003 32322 9029
rect 32370 9003 32384 9029
rect 32318 9002 32342 9003
rect 32370 9002 32394 9003
rect 32422 9002 32446 9030
rect 32474 9002 32498 9030
rect 32526 9029 32535 9030
rect 32534 9003 32535 9029
rect 32526 9002 32535 9003
rect 32073 8997 32535 9002
rect 31374 8353 31402 8358
rect 31878 8833 31906 8839
rect 31878 8807 31879 8833
rect 31905 8807 31906 8833
rect 31878 8777 31906 8807
rect 31878 8751 31879 8777
rect 31905 8751 31906 8777
rect 31878 8386 31906 8751
rect 32158 8833 32186 8839
rect 32158 8807 32159 8833
rect 32185 8807 32186 8833
rect 31374 8050 31402 8055
rect 31150 8049 31402 8050
rect 31150 8023 31151 8049
rect 31177 8023 31375 8049
rect 31401 8023 31402 8049
rect 31150 8022 31402 8023
rect 31150 8017 31178 8022
rect 31374 7713 31402 8022
rect 31878 8050 31906 8358
rect 32046 8441 32074 8447
rect 32046 8415 32047 8441
rect 32073 8415 32074 8441
rect 32046 8330 32074 8415
rect 32158 8442 32186 8807
rect 32718 8834 32746 8839
rect 32830 8834 32858 9590
rect 32718 8833 32858 8834
rect 32718 8807 32719 8833
rect 32745 8807 32831 8833
rect 32857 8807 32858 8833
rect 32718 8806 32858 8807
rect 32718 8801 32746 8806
rect 32830 8801 32858 8806
rect 32942 9226 32970 9231
rect 32158 8409 32186 8414
rect 32214 8554 32242 8559
rect 32214 8442 32242 8526
rect 32326 8442 32354 8447
rect 32214 8441 32354 8442
rect 32214 8415 32215 8441
rect 32241 8415 32327 8441
rect 32353 8415 32354 8441
rect 32214 8414 32354 8415
rect 32214 8409 32242 8414
rect 32326 8409 32354 8414
rect 32886 8441 32914 8447
rect 32886 8415 32887 8441
rect 32913 8415 32914 8441
rect 31878 8017 31906 8022
rect 31934 8302 32074 8330
rect 31374 7687 31375 7713
rect 31401 7687 31402 7713
rect 31374 7657 31402 7687
rect 31374 7631 31375 7657
rect 31401 7631 31402 7657
rect 31374 7574 31402 7631
rect 31374 7546 31850 7574
rect 30478 7518 31010 7546
rect 30982 7265 31010 7518
rect 30982 7239 30983 7265
rect 31009 7239 31010 7265
rect 29573 7070 30035 7075
rect 29573 7069 29582 7070
rect 29573 7043 29574 7069
rect 29573 7042 29582 7043
rect 29610 7042 29634 7070
rect 29662 7042 29686 7070
rect 29714 7069 29738 7070
rect 29766 7069 29790 7070
rect 29724 7043 29738 7069
rect 29786 7043 29790 7069
rect 29714 7042 29738 7043
rect 29766 7042 29790 7043
rect 29818 7069 29842 7070
rect 29870 7069 29894 7070
rect 29818 7043 29822 7069
rect 29870 7043 29884 7069
rect 29818 7042 29842 7043
rect 29870 7042 29894 7043
rect 29922 7042 29946 7070
rect 29974 7042 29998 7070
rect 30026 7069 30035 7070
rect 30034 7043 30035 7069
rect 30026 7042 30035 7043
rect 29573 7037 30035 7042
rect 29470 6841 29498 6846
rect 30478 6873 30506 6879
rect 30478 6847 30479 6873
rect 30505 6847 30506 6873
rect 30478 6818 30506 6847
rect 30646 6874 30674 6879
rect 30646 6827 30674 6846
rect 30478 6785 30506 6790
rect 30926 6818 30954 6823
rect 29414 6729 29442 6734
rect 30310 6762 30338 6767
rect 28854 6482 28882 6487
rect 28686 6481 28882 6482
rect 28686 6455 28687 6481
rect 28713 6455 28855 6481
rect 28881 6455 28882 6481
rect 28686 6454 28882 6455
rect 28686 6449 28714 6454
rect 28854 6449 28882 6454
rect 30198 6482 30226 6487
rect 30310 6482 30338 6734
rect 30198 6481 30338 6482
rect 30198 6455 30199 6481
rect 30225 6455 30311 6481
rect 30337 6455 30338 6481
rect 30198 6454 30338 6455
rect 30030 6426 30058 6431
rect 30030 6425 30170 6426
rect 30030 6399 30031 6425
rect 30057 6399 30170 6425
rect 30030 6398 30170 6399
rect 30030 6393 30058 6398
rect 29573 6286 30035 6291
rect 29573 6285 29582 6286
rect 29573 6259 29574 6285
rect 29573 6258 29582 6259
rect 29610 6258 29634 6286
rect 29662 6258 29686 6286
rect 29714 6285 29738 6286
rect 29766 6285 29790 6286
rect 29724 6259 29738 6285
rect 29786 6259 29790 6285
rect 29714 6258 29738 6259
rect 29766 6258 29790 6259
rect 29818 6285 29842 6286
rect 29870 6285 29894 6286
rect 29818 6259 29822 6285
rect 29870 6259 29884 6285
rect 29818 6258 29842 6259
rect 29870 6258 29894 6259
rect 29922 6258 29946 6286
rect 29974 6258 29998 6286
rect 30026 6285 30035 6286
rect 30034 6259 30035 6285
rect 30026 6258 30035 6259
rect 29573 6253 30035 6258
rect 30086 6202 30114 6207
rect 29470 6146 29498 6151
rect 28742 6089 28770 6095
rect 28742 6063 28743 6089
rect 28769 6063 28770 6089
rect 28742 5866 28770 6063
rect 28742 5305 28770 5838
rect 28742 5279 28743 5305
rect 28769 5279 28770 5305
rect 28742 4521 28770 5279
rect 28742 4495 28743 4521
rect 28769 4495 28770 4521
rect 28742 4214 28770 4495
rect 29134 5697 29162 5703
rect 29134 5671 29135 5697
rect 29161 5671 29162 5697
rect 29134 5641 29162 5671
rect 29134 5615 29135 5641
rect 29161 5615 29162 5641
rect 29134 4913 29162 5615
rect 29470 5362 29498 6118
rect 29918 6146 29946 6151
rect 29918 6089 29946 6118
rect 29918 6063 29919 6089
rect 29945 6063 29946 6089
rect 29918 6057 29946 6063
rect 30086 5697 30114 6174
rect 30142 5810 30170 6398
rect 30142 5777 30170 5782
rect 30086 5671 30087 5697
rect 30113 5671 30114 5697
rect 29573 5502 30035 5507
rect 29573 5501 29582 5502
rect 29573 5475 29574 5501
rect 29573 5474 29582 5475
rect 29610 5474 29634 5502
rect 29662 5474 29686 5502
rect 29714 5501 29738 5502
rect 29766 5501 29790 5502
rect 29724 5475 29738 5501
rect 29786 5475 29790 5501
rect 29714 5474 29738 5475
rect 29766 5474 29790 5475
rect 29818 5501 29842 5502
rect 29870 5501 29894 5502
rect 29818 5475 29822 5501
rect 29870 5475 29884 5501
rect 29818 5474 29842 5475
rect 29870 5474 29894 5475
rect 29922 5474 29946 5502
rect 29974 5474 29998 5502
rect 30026 5501 30035 5502
rect 30034 5475 30035 5501
rect 30026 5474 30035 5475
rect 29573 5469 30035 5474
rect 29694 5362 29722 5367
rect 29470 5361 29722 5362
rect 29470 5335 29695 5361
rect 29721 5335 29722 5361
rect 29470 5334 29722 5335
rect 29470 5305 29498 5334
rect 29694 5329 29722 5334
rect 29470 5279 29471 5305
rect 29497 5279 29498 5305
rect 29470 5273 29498 5279
rect 29134 4887 29135 4913
rect 29161 4887 29162 4913
rect 29134 4857 29162 4887
rect 29134 4831 29135 4857
rect 29161 4831 29162 4857
rect 29134 4522 29162 4831
rect 30086 4913 30114 5671
rect 30142 5641 30170 5647
rect 30142 5615 30143 5641
rect 30169 5615 30170 5641
rect 30142 5306 30170 5615
rect 30142 5273 30170 5278
rect 30086 4887 30087 4913
rect 30113 4887 30114 4913
rect 29573 4718 30035 4723
rect 29573 4717 29582 4718
rect 29573 4691 29574 4717
rect 29573 4690 29582 4691
rect 29610 4690 29634 4718
rect 29662 4690 29686 4718
rect 29714 4717 29738 4718
rect 29766 4717 29790 4718
rect 29724 4691 29738 4717
rect 29786 4691 29790 4717
rect 29714 4690 29738 4691
rect 29766 4690 29790 4691
rect 29818 4717 29842 4718
rect 29870 4717 29894 4718
rect 29818 4691 29822 4717
rect 29870 4691 29884 4717
rect 29818 4690 29842 4691
rect 29870 4690 29894 4691
rect 29922 4690 29946 4718
rect 29974 4690 29998 4718
rect 30026 4717 30035 4718
rect 30034 4691 30035 4717
rect 30026 4690 30035 4691
rect 29573 4685 30035 4690
rect 29190 4522 29218 4527
rect 29414 4522 29442 4527
rect 29134 4521 29442 4522
rect 29134 4495 29191 4521
rect 29217 4495 29415 4521
rect 29441 4495 29442 4521
rect 29134 4494 29442 4495
rect 29190 4489 29218 4494
rect 28742 4186 29050 4214
rect 28630 3033 28658 3038
rect 29022 3737 29050 4186
rect 29022 3711 29023 3737
rect 29049 3711 29050 3737
rect 29022 2953 29050 3711
rect 29358 4129 29386 4494
rect 29414 4489 29442 4494
rect 29358 4103 29359 4129
rect 29385 4103 29386 4129
rect 29358 4073 29386 4103
rect 29358 4047 29359 4073
rect 29385 4047 29386 4073
rect 29358 3738 29386 4047
rect 30030 4073 30058 4079
rect 30030 4047 30031 4073
rect 30057 4047 30058 4073
rect 30030 4018 30058 4047
rect 30030 3985 30058 3990
rect 29573 3934 30035 3939
rect 29573 3933 29582 3934
rect 29573 3907 29574 3933
rect 29573 3906 29582 3907
rect 29610 3906 29634 3934
rect 29662 3906 29686 3934
rect 29714 3933 29738 3934
rect 29766 3933 29790 3934
rect 29724 3907 29738 3933
rect 29786 3907 29790 3933
rect 29714 3906 29738 3907
rect 29766 3906 29790 3907
rect 29818 3933 29842 3934
rect 29870 3933 29894 3934
rect 29818 3907 29822 3933
rect 29870 3907 29884 3933
rect 29818 3906 29842 3907
rect 29870 3906 29894 3907
rect 29922 3906 29946 3934
rect 29974 3906 29998 3934
rect 30026 3933 30035 3934
rect 30034 3907 30035 3933
rect 30026 3906 30035 3907
rect 29573 3901 30035 3906
rect 30030 3850 30058 3855
rect 29918 3793 29946 3799
rect 29918 3767 29919 3793
rect 29945 3767 29946 3793
rect 29470 3738 29498 3743
rect 29358 3710 29470 3738
rect 29358 3402 29386 3407
rect 29358 3346 29386 3374
rect 29470 3346 29498 3710
rect 29918 3738 29946 3767
rect 29918 3691 29946 3710
rect 29358 3345 29498 3346
rect 29358 3319 29359 3345
rect 29385 3319 29498 3345
rect 29358 3318 29498 3319
rect 29358 3289 29386 3318
rect 29358 3263 29359 3289
rect 29385 3263 29386 3289
rect 29358 3257 29386 3263
rect 29022 2927 29023 2953
rect 29049 2927 29050 2953
rect 28686 2674 28714 2679
rect 28462 2515 28490 2534
rect 28630 2562 28658 2567
rect 28294 2143 28295 2169
rect 28321 2143 28322 2169
rect 28294 2137 28322 2143
rect 27073 1974 27535 1979
rect 27073 1973 27082 1974
rect 27073 1947 27074 1973
rect 27073 1946 27082 1947
rect 27110 1946 27134 1974
rect 27162 1946 27186 1974
rect 27214 1973 27238 1974
rect 27266 1973 27290 1974
rect 27224 1947 27238 1973
rect 27286 1947 27290 1973
rect 27214 1946 27238 1947
rect 27266 1946 27290 1947
rect 27318 1973 27342 1974
rect 27370 1973 27394 1974
rect 27318 1947 27322 1973
rect 27370 1947 27384 1973
rect 27318 1946 27342 1947
rect 27370 1946 27394 1947
rect 27422 1946 27446 1974
rect 27474 1946 27498 1974
rect 27526 1973 27535 1974
rect 27534 1947 27535 1973
rect 27526 1946 27535 1947
rect 27073 1941 27535 1946
rect 27006 1862 27258 1890
rect 26894 1751 26895 1777
rect 26921 1751 26922 1777
rect 26894 1666 26922 1751
rect 27062 1777 27090 1783
rect 27062 1751 27063 1777
rect 27089 1751 27090 1777
rect 27062 1722 27090 1751
rect 27006 1694 27090 1722
rect 27006 1666 27034 1694
rect 26894 1638 27034 1666
rect 25606 462 25802 490
rect 25606 378 25634 462
rect 25774 400 25802 462
rect 27230 400 27258 1862
rect 28630 1777 28658 2534
rect 28630 1751 28631 1777
rect 28657 1751 28658 1777
rect 28630 1745 28658 1751
rect 28686 400 28714 2646
rect 29022 2562 29050 2927
rect 29302 2954 29330 2959
rect 29470 2954 29498 3318
rect 30030 3290 30058 3822
rect 30086 3794 30114 4887
rect 30198 4914 30226 6454
rect 30310 6449 30338 6454
rect 30926 6481 30954 6790
rect 30926 6455 30927 6481
rect 30953 6455 30954 6481
rect 30254 6089 30282 6095
rect 30254 6063 30255 6089
rect 30281 6063 30282 6089
rect 30254 5894 30282 6063
rect 30254 5866 30394 5894
rect 30310 5642 30338 5647
rect 30198 4214 30226 4886
rect 30086 3761 30114 3766
rect 30142 4186 30226 4214
rect 30254 5641 30338 5642
rect 30254 5615 30311 5641
rect 30337 5615 30338 5641
rect 30254 5614 30338 5615
rect 30254 5306 30282 5614
rect 30310 5609 30338 5614
rect 30142 3346 30170 4186
rect 30198 4130 30226 4135
rect 30254 4130 30282 5278
rect 30366 5305 30394 5866
rect 30366 5279 30367 5305
rect 30393 5279 30394 5305
rect 30310 4914 30338 4919
rect 30310 4867 30338 4886
rect 30366 4521 30394 5279
rect 30366 4495 30367 4521
rect 30393 4495 30394 4521
rect 30310 4130 30338 4135
rect 30198 4129 30338 4130
rect 30198 4103 30199 4129
rect 30225 4103 30311 4129
rect 30337 4103 30338 4129
rect 30198 4102 30338 4103
rect 30198 4097 30226 4102
rect 30310 4097 30338 4102
rect 30366 3737 30394 4495
rect 30366 3711 30367 3737
rect 30393 3711 30394 3737
rect 30198 3346 30226 3351
rect 30142 3345 30338 3346
rect 30142 3319 30199 3345
rect 30225 3319 30338 3345
rect 30142 3318 30338 3319
rect 30030 3243 30058 3262
rect 29573 3150 30035 3155
rect 29573 3149 29582 3150
rect 29573 3123 29574 3149
rect 29573 3122 29582 3123
rect 29610 3122 29634 3150
rect 29662 3122 29686 3150
rect 29714 3149 29738 3150
rect 29766 3149 29790 3150
rect 29724 3123 29738 3149
rect 29786 3123 29790 3149
rect 29714 3122 29738 3123
rect 29766 3122 29790 3123
rect 29818 3149 29842 3150
rect 29870 3149 29894 3150
rect 29818 3123 29822 3149
rect 29870 3123 29884 3149
rect 29818 3122 29842 3123
rect 29870 3122 29894 3123
rect 29922 3122 29946 3150
rect 29974 3122 29998 3150
rect 30026 3149 30035 3150
rect 30034 3123 30035 3149
rect 30026 3122 30035 3123
rect 29573 3117 30035 3122
rect 29302 2953 29498 2954
rect 29302 2927 29303 2953
rect 29329 2927 29471 2953
rect 29497 2927 29498 2953
rect 29302 2926 29498 2927
rect 29302 2921 29330 2926
rect 29022 2169 29050 2534
rect 29358 2561 29386 2926
rect 29470 2921 29498 2926
rect 29358 2535 29359 2561
rect 29385 2535 29386 2561
rect 29358 2505 29386 2535
rect 29358 2479 29359 2505
rect 29385 2479 29386 2505
rect 29358 2473 29386 2479
rect 30030 2562 30058 2567
rect 30198 2562 30226 3318
rect 30310 3289 30338 3318
rect 30310 3263 30311 3289
rect 30337 3263 30338 3289
rect 30310 3010 30338 3263
rect 30310 2977 30338 2982
rect 30030 2561 30226 2562
rect 30030 2535 30031 2561
rect 30057 2535 30199 2561
rect 30225 2535 30226 2561
rect 30030 2534 30226 2535
rect 30030 2506 30058 2534
rect 30198 2529 30226 2534
rect 30366 2953 30394 3711
rect 30366 2927 30367 2953
rect 30393 2927 30394 2953
rect 30366 2562 30394 2927
rect 30310 2506 30338 2511
rect 30030 2473 30058 2478
rect 30254 2505 30338 2506
rect 30254 2479 30311 2505
rect 30337 2479 30338 2505
rect 30254 2478 30338 2479
rect 29573 2366 30035 2371
rect 29573 2365 29582 2366
rect 29573 2339 29574 2365
rect 29573 2338 29582 2339
rect 29610 2338 29634 2366
rect 29662 2338 29686 2366
rect 29714 2365 29738 2366
rect 29766 2365 29790 2366
rect 29724 2339 29738 2365
rect 29786 2339 29790 2365
rect 29714 2338 29738 2339
rect 29766 2338 29790 2339
rect 29818 2365 29842 2366
rect 29870 2365 29894 2366
rect 29818 2339 29822 2365
rect 29870 2339 29884 2365
rect 29818 2338 29842 2339
rect 29870 2338 29894 2339
rect 29922 2338 29946 2366
rect 29974 2338 29998 2366
rect 30026 2365 30035 2366
rect 30034 2339 30035 2365
rect 30026 2338 30035 2339
rect 29573 2333 30035 2338
rect 29414 2226 29442 2231
rect 29022 2143 29023 2169
rect 29049 2143 29050 2169
rect 29022 2137 29050 2143
rect 29190 2170 29218 2175
rect 29414 2170 29442 2198
rect 29190 2169 29442 2170
rect 29190 2143 29191 2169
rect 29217 2143 29415 2169
rect 29441 2143 29442 2169
rect 29190 2142 29442 2143
rect 28798 1777 28826 1783
rect 28798 1751 28799 1777
rect 28825 1751 28826 1777
rect 28798 1666 28826 1751
rect 28798 1633 28826 1638
rect 29022 1778 29050 1783
rect 29190 1778 29218 2142
rect 29414 2137 29442 2142
rect 30254 2170 30282 2478
rect 30310 2473 30338 2478
rect 29022 1777 29218 1778
rect 29022 1751 29023 1777
rect 29049 1751 29218 1777
rect 29022 1750 29218 1751
rect 29022 1666 29050 1750
rect 30254 1722 30282 2142
rect 30366 2169 30394 2534
rect 30702 5697 30730 5703
rect 30702 5671 30703 5697
rect 30729 5671 30730 5697
rect 30702 4913 30730 5671
rect 30926 5698 30954 6455
rect 30982 6482 31010 7239
rect 31822 7265 31850 7546
rect 31822 7239 31823 7265
rect 31849 7239 31850 7265
rect 31822 7209 31850 7239
rect 31822 7183 31823 7209
rect 31849 7183 31850 7209
rect 31374 6873 31402 6879
rect 31374 6847 31375 6873
rect 31401 6847 31402 6873
rect 31374 6818 31402 6847
rect 31374 6785 31402 6790
rect 30982 6449 31010 6454
rect 30926 5665 30954 5670
rect 31374 6146 31402 6151
rect 31374 6089 31402 6118
rect 31374 6063 31375 6089
rect 31401 6063 31402 6089
rect 30702 4887 30703 4913
rect 30729 4887 30730 4913
rect 30702 4129 30730 4887
rect 31374 5361 31402 6063
rect 31822 5698 31850 7183
rect 31878 6818 31906 6823
rect 31878 6481 31906 6790
rect 31878 6455 31879 6481
rect 31905 6455 31906 6481
rect 31878 6425 31906 6455
rect 31878 6399 31879 6425
rect 31905 6399 31906 6425
rect 31878 6393 31906 6399
rect 31934 5810 31962 8302
rect 32073 8246 32535 8251
rect 32073 8245 32082 8246
rect 32073 8219 32074 8245
rect 32073 8218 32082 8219
rect 32110 8218 32134 8246
rect 32162 8218 32186 8246
rect 32214 8245 32238 8246
rect 32266 8245 32290 8246
rect 32224 8219 32238 8245
rect 32286 8219 32290 8245
rect 32214 8218 32238 8219
rect 32266 8218 32290 8219
rect 32318 8245 32342 8246
rect 32370 8245 32394 8246
rect 32318 8219 32322 8245
rect 32370 8219 32384 8245
rect 32318 8218 32342 8219
rect 32370 8218 32394 8219
rect 32422 8218 32446 8246
rect 32474 8218 32498 8246
rect 32526 8245 32535 8246
rect 32534 8219 32535 8245
rect 32526 8218 32535 8219
rect 32073 8213 32535 8218
rect 32438 8162 32466 8167
rect 32438 8049 32466 8134
rect 32438 8023 32439 8049
rect 32465 8023 32466 8049
rect 32102 7657 32130 7663
rect 32102 7631 32103 7657
rect 32129 7631 32130 7657
rect 32102 7546 32130 7631
rect 32158 7658 32186 7663
rect 32158 7611 32186 7630
rect 32326 7658 32354 7663
rect 32326 7611 32354 7630
rect 32438 7658 32466 8023
rect 32438 7625 32466 7630
rect 32886 7574 32914 8415
rect 32942 8442 32970 9198
rect 32998 8778 33026 10767
rect 33894 10849 33922 11102
rect 35294 11130 35322 11158
rect 35294 11097 35322 11102
rect 35854 11185 35882 11191
rect 35854 11159 35855 11185
rect 35881 11159 35882 11185
rect 35854 11130 35882 11159
rect 35854 11097 35882 11102
rect 36134 11186 36162 11191
rect 34573 10990 35035 10995
rect 34573 10989 34582 10990
rect 34573 10963 34574 10989
rect 34573 10962 34582 10963
rect 34610 10962 34634 10990
rect 34662 10962 34686 10990
rect 34714 10989 34738 10990
rect 34766 10989 34790 10990
rect 34724 10963 34738 10989
rect 34786 10963 34790 10989
rect 34714 10962 34738 10963
rect 34766 10962 34790 10963
rect 34818 10989 34842 10990
rect 34870 10989 34894 10990
rect 34818 10963 34822 10989
rect 34870 10963 34884 10989
rect 34818 10962 34842 10963
rect 34870 10962 34894 10963
rect 34922 10962 34946 10990
rect 34974 10962 34998 10990
rect 35026 10989 35035 10990
rect 35034 10963 35035 10989
rect 35026 10962 35035 10963
rect 34573 10957 35035 10962
rect 33894 10823 33895 10849
rect 33921 10823 33922 10849
rect 33894 10794 33922 10823
rect 35350 10849 35378 10855
rect 35350 10823 35351 10849
rect 35377 10823 35378 10849
rect 33894 10747 33922 10766
rect 34230 10793 34258 10799
rect 34230 10767 34231 10793
rect 34257 10767 34258 10793
rect 33110 10401 33138 10407
rect 33110 10375 33111 10401
rect 33137 10375 33138 10401
rect 33110 10345 33138 10375
rect 33110 10319 33111 10345
rect 33137 10319 33138 10345
rect 33110 9618 33138 10319
rect 34230 10094 34258 10767
rect 35350 10794 35378 10823
rect 35378 10766 35434 10794
rect 35350 10728 35378 10766
rect 34678 10402 34706 10407
rect 34510 10401 34706 10402
rect 34510 10375 34679 10401
rect 34705 10375 34706 10401
rect 34510 10374 34706 10375
rect 34510 10094 34538 10374
rect 34678 10369 34706 10374
rect 34573 10206 35035 10211
rect 34573 10205 34582 10206
rect 34573 10179 34574 10205
rect 34573 10178 34582 10179
rect 34610 10178 34634 10206
rect 34662 10178 34686 10206
rect 34714 10205 34738 10206
rect 34766 10205 34790 10206
rect 34724 10179 34738 10205
rect 34786 10179 34790 10205
rect 34714 10178 34738 10179
rect 34766 10178 34790 10179
rect 34818 10205 34842 10206
rect 34870 10205 34894 10206
rect 34818 10179 34822 10205
rect 34870 10179 34884 10205
rect 34818 10178 34842 10179
rect 34870 10178 34894 10179
rect 34922 10178 34946 10206
rect 34974 10178 34998 10206
rect 35026 10205 35035 10206
rect 35034 10179 35035 10205
rect 35026 10178 35035 10179
rect 34573 10173 35035 10178
rect 33110 9561 33138 9590
rect 33110 9535 33111 9561
rect 33137 9535 33138 9561
rect 33110 9226 33138 9535
rect 33838 10065 33866 10071
rect 33838 10039 33839 10065
rect 33865 10039 33866 10065
rect 33838 10009 33866 10039
rect 34230 10066 34538 10094
rect 35406 10094 35434 10766
rect 35630 10401 35658 10407
rect 35630 10375 35631 10401
rect 35657 10375 35658 10401
rect 35630 10345 35658 10375
rect 35630 10319 35631 10345
rect 35657 10319 35658 10345
rect 35630 10094 35658 10319
rect 34230 10033 34258 10038
rect 33838 9983 33839 10009
rect 33865 9983 33866 10009
rect 33390 9282 33418 9287
rect 33166 9226 33194 9231
rect 33390 9226 33418 9254
rect 33110 9225 33418 9226
rect 33110 9199 33167 9225
rect 33193 9199 33391 9225
rect 33417 9199 33418 9225
rect 33110 9198 33418 9199
rect 33166 9193 33194 9198
rect 33390 9193 33418 9198
rect 32998 8745 33026 8750
rect 32942 8409 32970 8414
rect 33334 8050 33362 8055
rect 33334 7993 33362 8022
rect 33726 8049 33754 8055
rect 33726 8023 33727 8049
rect 33753 8023 33754 8049
rect 33334 7967 33335 7993
rect 33361 7967 33362 7993
rect 33334 7714 33362 7967
rect 33614 7994 33642 7999
rect 33726 7994 33754 8023
rect 33614 7993 33754 7994
rect 33614 7967 33615 7993
rect 33641 7967 33754 7993
rect 33614 7966 33754 7967
rect 33614 7961 33642 7966
rect 33334 7681 33362 7686
rect 32102 7513 32130 7518
rect 32774 7546 32914 7574
rect 32606 7490 32634 7495
rect 32073 7462 32535 7467
rect 32073 7461 32082 7462
rect 32073 7435 32074 7461
rect 32073 7434 32082 7435
rect 32110 7434 32134 7462
rect 32162 7434 32186 7462
rect 32214 7461 32238 7462
rect 32266 7461 32290 7462
rect 32224 7435 32238 7461
rect 32286 7435 32290 7461
rect 32214 7434 32238 7435
rect 32266 7434 32290 7435
rect 32318 7461 32342 7462
rect 32370 7461 32394 7462
rect 32318 7435 32322 7461
rect 32370 7435 32384 7461
rect 32318 7434 32342 7435
rect 32370 7434 32394 7435
rect 32422 7434 32446 7462
rect 32474 7434 32498 7462
rect 32526 7461 32535 7462
rect 32534 7435 32535 7461
rect 32526 7434 32535 7435
rect 32073 7429 32535 7434
rect 32438 7266 32466 7271
rect 32046 6874 32074 6879
rect 31990 6873 32074 6874
rect 31990 6847 32047 6873
rect 32073 6847 32074 6873
rect 31990 6846 32074 6847
rect 31990 6202 32018 6846
rect 32046 6841 32074 6846
rect 32158 6874 32186 6879
rect 32326 6874 32354 6879
rect 32158 6873 32354 6874
rect 32158 6847 32159 6873
rect 32185 6847 32327 6873
rect 32353 6847 32354 6873
rect 32158 6846 32354 6847
rect 32158 6762 32186 6846
rect 32326 6841 32354 6846
rect 32158 6729 32186 6734
rect 32438 6762 32466 7238
rect 32438 6729 32466 6734
rect 32073 6678 32535 6683
rect 32073 6677 32082 6678
rect 32073 6651 32074 6677
rect 32073 6650 32082 6651
rect 32110 6650 32134 6678
rect 32162 6650 32186 6678
rect 32214 6677 32238 6678
rect 32266 6677 32290 6678
rect 32224 6651 32238 6677
rect 32286 6651 32290 6677
rect 32214 6650 32238 6651
rect 32266 6650 32290 6651
rect 32318 6677 32342 6678
rect 32370 6677 32394 6678
rect 32318 6651 32322 6677
rect 32370 6651 32384 6677
rect 32318 6650 32342 6651
rect 32370 6650 32394 6651
rect 32422 6650 32446 6678
rect 32474 6650 32498 6678
rect 32526 6677 32535 6678
rect 32534 6651 32535 6677
rect 32526 6650 32535 6651
rect 32073 6645 32535 6650
rect 32158 6482 32186 6487
rect 32158 6435 32186 6454
rect 31990 6169 32018 6174
rect 32046 6090 32074 6095
rect 31934 5777 31962 5782
rect 31990 6089 32074 6090
rect 31990 6063 32047 6089
rect 32073 6063 32074 6089
rect 31990 6062 32074 6063
rect 31878 5698 31906 5703
rect 31822 5697 31906 5698
rect 31822 5671 31879 5697
rect 31905 5671 31906 5697
rect 31822 5670 31906 5671
rect 31374 5335 31375 5361
rect 31401 5335 31402 5361
rect 31374 5305 31402 5335
rect 31374 5279 31375 5305
rect 31401 5279 31402 5305
rect 31374 4577 31402 5279
rect 31374 4551 31375 4577
rect 31401 4551 31402 4577
rect 31374 4522 31402 4551
rect 31878 5641 31906 5670
rect 31878 5615 31879 5641
rect 31905 5615 31906 5641
rect 31878 4913 31906 5615
rect 31878 4887 31879 4913
rect 31905 4887 31906 4913
rect 31878 4857 31906 4887
rect 31878 4831 31879 4857
rect 31905 4831 31906 4857
rect 31878 4522 31906 4831
rect 31374 4521 31906 4522
rect 31374 4495 31375 4521
rect 31401 4495 31906 4521
rect 31374 4494 31906 4495
rect 30702 4103 30703 4129
rect 30729 4103 30730 4129
rect 30702 3346 30730 4103
rect 31318 4130 31346 4135
rect 31318 3793 31346 4102
rect 31318 3767 31319 3793
rect 31345 3767 31346 3793
rect 31318 3738 31346 3767
rect 31318 3672 31346 3710
rect 30702 2562 30730 3318
rect 31374 3009 31402 4494
rect 31878 4129 31906 4494
rect 31878 4103 31879 4129
rect 31905 4103 31906 4129
rect 31878 4073 31906 4103
rect 31878 4047 31879 4073
rect 31905 4047 31906 4073
rect 31878 3402 31906 4047
rect 31878 3345 31906 3374
rect 31878 3319 31879 3345
rect 31905 3319 31906 3345
rect 31878 3289 31906 3319
rect 31878 3263 31879 3289
rect 31905 3263 31906 3289
rect 31878 3257 31906 3263
rect 31934 5306 31962 5311
rect 31374 2983 31375 3009
rect 31401 2983 31402 3009
rect 31374 2953 31402 2983
rect 31374 2927 31375 2953
rect 31401 2927 31402 2953
rect 30702 2515 30730 2534
rect 31262 2562 31290 2567
rect 31374 2562 31402 2927
rect 31262 2561 31402 2562
rect 31262 2535 31263 2561
rect 31289 2535 31375 2561
rect 31401 2535 31402 2561
rect 31262 2534 31402 2535
rect 30366 2143 30367 2169
rect 30393 2143 30394 2169
rect 30366 1777 30394 2143
rect 30366 1751 30367 1777
rect 30393 1751 30394 1777
rect 30366 1745 30394 1751
rect 31262 2226 31290 2534
rect 31374 2529 31402 2534
rect 31262 2169 31290 2198
rect 31262 2143 31263 2169
rect 31289 2143 31290 2169
rect 31262 1777 31290 2143
rect 31262 1751 31263 1777
rect 31289 1751 31290 1777
rect 29022 1633 29050 1638
rect 30142 1694 30282 1722
rect 31262 1721 31290 1751
rect 31262 1695 31263 1721
rect 31289 1695 31290 1721
rect 29573 1582 30035 1587
rect 29573 1581 29582 1582
rect 29573 1555 29574 1581
rect 29573 1554 29582 1555
rect 29610 1554 29634 1582
rect 29662 1554 29686 1582
rect 29714 1581 29738 1582
rect 29766 1581 29790 1582
rect 29724 1555 29738 1581
rect 29786 1555 29790 1581
rect 29714 1554 29738 1555
rect 29766 1554 29790 1555
rect 29818 1581 29842 1582
rect 29870 1581 29894 1582
rect 29818 1555 29822 1581
rect 29870 1555 29884 1581
rect 29818 1554 29842 1555
rect 29870 1554 29894 1555
rect 29922 1554 29946 1582
rect 29974 1554 29998 1582
rect 30026 1581 30035 1582
rect 30034 1555 30035 1581
rect 30026 1554 30035 1555
rect 29573 1549 30035 1554
rect 30142 400 30170 1694
rect 31262 1689 31290 1695
rect 31598 2450 31626 2455
rect 31598 1834 31626 2422
rect 31934 2226 31962 5278
rect 31990 5306 32018 6062
rect 32046 6057 32074 6062
rect 32158 6090 32186 6095
rect 32158 6043 32186 6062
rect 32326 6090 32354 6095
rect 32326 6043 32354 6062
rect 32073 5894 32535 5899
rect 32073 5893 32082 5894
rect 32073 5867 32074 5893
rect 32073 5866 32082 5867
rect 32110 5866 32134 5894
rect 32162 5866 32186 5894
rect 32214 5893 32238 5894
rect 32266 5893 32290 5894
rect 32224 5867 32238 5893
rect 32286 5867 32290 5893
rect 32214 5866 32238 5867
rect 32266 5866 32290 5867
rect 32318 5893 32342 5894
rect 32370 5893 32394 5894
rect 32318 5867 32322 5893
rect 32370 5867 32384 5893
rect 32318 5866 32342 5867
rect 32370 5866 32394 5867
rect 32422 5866 32446 5894
rect 32474 5866 32498 5894
rect 32526 5893 32535 5894
rect 32534 5867 32535 5893
rect 32526 5866 32535 5867
rect 32073 5861 32535 5866
rect 32158 5698 32186 5703
rect 32158 5651 32186 5670
rect 32046 5306 32074 5311
rect 31990 5305 32074 5306
rect 31990 5279 32047 5305
rect 32073 5279 32074 5305
rect 31990 5278 32074 5279
rect 31990 4522 32018 5278
rect 32046 5273 32074 5278
rect 32158 5306 32186 5311
rect 32158 5259 32186 5278
rect 32326 5306 32354 5311
rect 32326 5259 32354 5278
rect 32073 5110 32535 5115
rect 32073 5109 32082 5110
rect 32073 5083 32074 5109
rect 32073 5082 32082 5083
rect 32110 5082 32134 5110
rect 32162 5082 32186 5110
rect 32214 5109 32238 5110
rect 32266 5109 32290 5110
rect 32224 5083 32238 5109
rect 32286 5083 32290 5109
rect 32214 5082 32238 5083
rect 32266 5082 32290 5083
rect 32318 5109 32342 5110
rect 32370 5109 32394 5110
rect 32318 5083 32322 5109
rect 32370 5083 32384 5109
rect 32318 5082 32342 5083
rect 32370 5082 32394 5083
rect 32422 5082 32446 5110
rect 32474 5082 32498 5110
rect 32526 5109 32535 5110
rect 32534 5083 32535 5109
rect 32526 5082 32535 5083
rect 32073 5077 32535 5082
rect 32158 4914 32186 4919
rect 32158 4867 32186 4886
rect 32606 4690 32634 7462
rect 32774 7154 32802 7546
rect 32886 7513 32914 7518
rect 32942 7658 32970 7663
rect 32774 7121 32802 7126
rect 32886 7266 32914 7271
rect 32718 6482 32746 6487
rect 32718 6090 32746 6454
rect 32886 6370 32914 7238
rect 32886 6337 32914 6342
rect 32718 6089 32802 6090
rect 32718 6063 32719 6089
rect 32745 6063 32802 6089
rect 32718 6062 32802 6063
rect 32718 6057 32746 6062
rect 32606 4657 32634 4662
rect 32662 5698 32690 5703
rect 32662 4578 32690 5670
rect 32774 5306 32802 6062
rect 32774 5240 32802 5278
rect 32942 4970 32970 7630
rect 33726 7602 33754 7966
rect 33670 7490 33698 7495
rect 33334 7265 33362 7271
rect 33334 7239 33335 7265
rect 33361 7239 33362 7265
rect 33334 7209 33362 7239
rect 33334 7183 33335 7209
rect 33361 7183 33362 7209
rect 32998 6873 33026 6879
rect 32998 6847 32999 6873
rect 33025 6847 33026 6873
rect 32998 6762 33026 6847
rect 33334 6818 33362 7183
rect 33670 7265 33698 7462
rect 33670 7239 33671 7265
rect 33697 7239 33698 7265
rect 33670 7154 33698 7239
rect 33726 7265 33754 7574
rect 33726 7239 33727 7265
rect 33753 7239 33754 7265
rect 33726 7210 33754 7239
rect 33726 7177 33754 7182
rect 33838 7714 33866 9983
rect 34454 10009 34482 10066
rect 34454 9983 34455 10009
rect 34481 9983 34482 10009
rect 34454 9618 34482 9983
rect 35350 10065 35378 10071
rect 35406 10066 35658 10094
rect 35350 10039 35351 10065
rect 35377 10039 35378 10065
rect 35350 10009 35378 10039
rect 35350 9983 35351 10009
rect 35377 9983 35378 10009
rect 34454 9585 34482 9590
rect 34958 9618 34986 9623
rect 34958 9571 34986 9590
rect 35350 9562 35378 9983
rect 35350 9529 35378 9534
rect 34573 9422 35035 9427
rect 34573 9421 34582 9422
rect 34573 9395 34574 9421
rect 34573 9394 34582 9395
rect 34610 9394 34634 9422
rect 34662 9394 34686 9422
rect 34714 9421 34738 9422
rect 34766 9421 34790 9422
rect 34724 9395 34738 9421
rect 34786 9395 34790 9421
rect 34714 9394 34738 9395
rect 34766 9394 34790 9395
rect 34818 9421 34842 9422
rect 34870 9421 34894 9422
rect 34818 9395 34822 9421
rect 34870 9395 34884 9421
rect 34818 9394 34842 9395
rect 34870 9394 34894 9395
rect 34922 9394 34946 9422
rect 34974 9394 34998 9422
rect 35026 9421 35035 9422
rect 35034 9395 35035 9421
rect 35026 9394 35035 9395
rect 34573 9389 35035 9394
rect 34622 9282 34650 9287
rect 34174 9226 34202 9231
rect 34174 9179 34202 9198
rect 34622 9225 34650 9254
rect 34622 9199 34623 9225
rect 34649 9199 34650 9225
rect 34622 9193 34650 9199
rect 34846 9282 34874 9287
rect 34846 9225 34874 9254
rect 34846 9199 34847 9225
rect 34873 9199 34874 9225
rect 34846 9193 34874 9199
rect 35070 9282 35098 9287
rect 34958 8834 34986 8839
rect 34958 8787 34986 8806
rect 34573 8638 35035 8643
rect 34573 8637 34582 8638
rect 34573 8611 34574 8637
rect 34573 8610 34582 8611
rect 34610 8610 34634 8638
rect 34662 8610 34686 8638
rect 34714 8637 34738 8638
rect 34766 8637 34790 8638
rect 34724 8611 34738 8637
rect 34786 8611 34790 8637
rect 34714 8610 34738 8611
rect 34766 8610 34790 8611
rect 34818 8637 34842 8638
rect 34870 8637 34894 8638
rect 34818 8611 34822 8637
rect 34870 8611 34884 8637
rect 34818 8610 34842 8611
rect 34870 8610 34894 8611
rect 34922 8610 34946 8638
rect 34974 8610 34998 8638
rect 35026 8637 35035 8638
rect 35034 8611 35035 8637
rect 35026 8610 35035 8611
rect 34573 8605 35035 8610
rect 33894 8498 33922 8503
rect 33894 8442 33922 8470
rect 35070 8498 35098 9254
rect 35630 9226 35658 10066
rect 36078 10402 36106 10407
rect 35854 9617 35882 9623
rect 35854 9591 35855 9617
rect 35881 9591 35882 9617
rect 35854 9562 35882 9591
rect 35854 9515 35882 9534
rect 35630 9193 35658 9198
rect 35854 9226 35882 9231
rect 35238 9114 35266 9119
rect 35126 8498 35154 8503
rect 35070 8497 35154 8498
rect 35070 8471 35127 8497
rect 35153 8471 35154 8497
rect 35070 8470 35154 8471
rect 34398 8442 34426 8447
rect 33894 8441 33978 8442
rect 33894 8415 33895 8441
rect 33921 8415 33978 8441
rect 33894 8414 33978 8415
rect 33894 8409 33922 8414
rect 33838 7657 33866 7686
rect 33838 7631 33839 7657
rect 33865 7631 33866 7657
rect 33670 7121 33698 7126
rect 33334 6785 33362 6790
rect 33670 6929 33698 6935
rect 33670 6903 33671 6929
rect 33697 6903 33698 6929
rect 33670 6873 33698 6903
rect 33670 6847 33671 6873
rect 33697 6847 33698 6873
rect 32998 6729 33026 6734
rect 33670 6706 33698 6847
rect 33278 6481 33306 6487
rect 33278 6455 33279 6481
rect 33305 6455 33306 6481
rect 33278 6425 33306 6455
rect 33278 6399 33279 6425
rect 33305 6399 33306 6425
rect 33278 5866 33306 6399
rect 33614 6425 33642 6431
rect 33614 6399 33615 6425
rect 33641 6399 33642 6425
rect 33614 6202 33642 6399
rect 33614 6169 33642 6174
rect 33614 6089 33642 6095
rect 33614 6063 33615 6089
rect 33641 6063 33642 6089
rect 33278 5833 33306 5838
rect 33334 5922 33362 5927
rect 32942 4937 32970 4942
rect 33054 5810 33082 5815
rect 32662 4550 32802 4578
rect 32046 4522 32074 4527
rect 31990 4521 32074 4522
rect 31990 4495 32047 4521
rect 32073 4495 32074 4521
rect 31990 4494 32074 4495
rect 31990 3738 32018 4494
rect 32046 4489 32074 4494
rect 32214 4522 32242 4527
rect 32382 4522 32410 4527
rect 32214 4521 32410 4522
rect 32214 4495 32215 4521
rect 32241 4495 32383 4521
rect 32409 4495 32410 4521
rect 32214 4494 32410 4495
rect 32214 4489 32242 4494
rect 32382 4410 32410 4494
rect 32774 4521 32802 4550
rect 32774 4495 32775 4521
rect 32801 4495 32802 4521
rect 32382 4382 32634 4410
rect 32073 4326 32535 4331
rect 32073 4325 32082 4326
rect 32073 4299 32074 4325
rect 32073 4298 32082 4299
rect 32110 4298 32134 4326
rect 32162 4298 32186 4326
rect 32214 4325 32238 4326
rect 32266 4325 32290 4326
rect 32224 4299 32238 4325
rect 32286 4299 32290 4325
rect 32214 4298 32238 4299
rect 32266 4298 32290 4299
rect 32318 4325 32342 4326
rect 32370 4325 32394 4326
rect 32318 4299 32322 4325
rect 32370 4299 32384 4325
rect 32318 4298 32342 4299
rect 32370 4298 32394 4299
rect 32422 4298 32446 4326
rect 32474 4298 32498 4326
rect 32526 4325 32535 4326
rect 32534 4299 32535 4325
rect 32526 4298 32535 4299
rect 32073 4293 32535 4298
rect 32158 4129 32186 4135
rect 32158 4103 32159 4129
rect 32185 4103 32186 4129
rect 32158 4074 32186 4103
rect 32158 4041 32186 4046
rect 32046 3738 32074 3743
rect 31990 3737 32074 3738
rect 31990 3711 32047 3737
rect 32073 3711 32074 3737
rect 31990 3710 32074 3711
rect 31990 3290 32018 3710
rect 32046 3705 32074 3710
rect 32214 3738 32242 3743
rect 32382 3738 32410 3743
rect 32214 3737 32410 3738
rect 32214 3711 32215 3737
rect 32241 3711 32383 3737
rect 32409 3711 32410 3737
rect 32214 3710 32410 3711
rect 32214 3705 32242 3710
rect 32382 3682 32410 3710
rect 32606 3682 32634 4382
rect 32382 3654 32634 3682
rect 32073 3542 32535 3547
rect 32073 3541 32082 3542
rect 32073 3515 32074 3541
rect 32073 3514 32082 3515
rect 32110 3514 32134 3542
rect 32162 3514 32186 3542
rect 32214 3541 32238 3542
rect 32266 3541 32290 3542
rect 32224 3515 32238 3541
rect 32286 3515 32290 3541
rect 32214 3514 32238 3515
rect 32266 3514 32290 3515
rect 32318 3541 32342 3542
rect 32370 3541 32394 3542
rect 32318 3515 32322 3541
rect 32370 3515 32384 3541
rect 32318 3514 32342 3515
rect 32370 3514 32394 3515
rect 32422 3514 32446 3542
rect 32474 3514 32498 3542
rect 32526 3541 32535 3542
rect 32534 3515 32535 3541
rect 32526 3514 32535 3515
rect 32073 3509 32535 3514
rect 32158 3346 32186 3351
rect 32158 3299 32186 3318
rect 31990 3010 32018 3262
rect 32046 3010 32074 3015
rect 31990 2982 32046 3010
rect 32046 2963 32074 2982
rect 32214 2954 32242 2959
rect 32214 2907 32242 2926
rect 32382 2954 32410 2959
rect 32382 2907 32410 2926
rect 32606 2954 32634 3654
rect 32606 2921 32634 2926
rect 32774 3738 32802 4495
rect 32774 2953 32802 3710
rect 32774 2927 32775 2953
rect 32801 2927 32802 2953
rect 32073 2758 32535 2763
rect 32073 2757 32082 2758
rect 32073 2731 32074 2757
rect 32073 2730 32082 2731
rect 32110 2730 32134 2758
rect 32162 2730 32186 2758
rect 32214 2757 32238 2758
rect 32266 2757 32290 2758
rect 32224 2731 32238 2757
rect 32286 2731 32290 2757
rect 32214 2730 32238 2731
rect 32266 2730 32290 2731
rect 32318 2757 32342 2758
rect 32370 2757 32394 2758
rect 32318 2731 32322 2757
rect 32370 2731 32384 2757
rect 32318 2730 32342 2731
rect 32370 2730 32394 2731
rect 32422 2730 32446 2758
rect 32474 2730 32498 2758
rect 32526 2757 32535 2758
rect 32534 2731 32535 2757
rect 32526 2730 32535 2731
rect 32073 2725 32535 2730
rect 32438 2674 32466 2679
rect 32438 2562 32466 2646
rect 32774 2562 32802 2927
rect 32438 2561 32802 2562
rect 32438 2535 32439 2561
rect 32465 2535 32802 2561
rect 32438 2534 32802 2535
rect 32438 2529 32466 2534
rect 31822 2225 31962 2226
rect 31822 2199 31935 2225
rect 31961 2199 31962 2225
rect 31822 2198 31962 2199
rect 31654 2170 31682 2175
rect 31654 2123 31682 2142
rect 31822 2169 31850 2198
rect 31934 2193 31962 2198
rect 31822 2143 31823 2169
rect 31849 2143 31850 2169
rect 31822 2137 31850 2143
rect 32718 2169 32746 2534
rect 32718 2143 32719 2169
rect 32745 2143 32746 2169
rect 32073 1974 32535 1979
rect 32073 1973 32082 1974
rect 32073 1947 32074 1973
rect 32073 1946 32082 1947
rect 32110 1946 32134 1974
rect 32162 1946 32186 1974
rect 32214 1973 32238 1974
rect 32266 1973 32290 1974
rect 32224 1947 32238 1973
rect 32286 1947 32290 1973
rect 32214 1946 32238 1947
rect 32266 1946 32290 1947
rect 32318 1973 32342 1974
rect 32370 1973 32394 1974
rect 32318 1947 32322 1973
rect 32370 1947 32384 1973
rect 32318 1946 32342 1947
rect 32370 1946 32394 1947
rect 32422 1946 32446 1974
rect 32474 1946 32498 1974
rect 32526 1973 32535 1974
rect 32534 1947 32535 1973
rect 32526 1946 32535 1947
rect 32073 1941 32535 1946
rect 31598 400 31626 1806
rect 32550 1778 32578 1783
rect 32718 1778 32746 2143
rect 32550 1777 32746 1778
rect 32550 1751 32551 1777
rect 32577 1751 32746 1777
rect 32550 1750 32746 1751
rect 32550 1745 32578 1750
rect 33054 400 33082 5782
rect 33334 5697 33362 5894
rect 33334 5671 33335 5697
rect 33361 5671 33362 5697
rect 33334 5641 33362 5671
rect 33334 5615 33335 5641
rect 33361 5615 33362 5641
rect 33334 5609 33362 5615
rect 33614 5866 33642 6063
rect 33670 5922 33698 6678
rect 33670 5889 33698 5894
rect 33726 6426 33754 6431
rect 33334 5362 33362 5367
rect 33334 4913 33362 5334
rect 33614 5362 33642 5838
rect 33614 5329 33642 5334
rect 33670 5697 33698 5703
rect 33670 5671 33671 5697
rect 33697 5671 33698 5697
rect 33334 4887 33335 4913
rect 33361 4887 33362 4913
rect 33334 4857 33362 4887
rect 33334 4831 33335 4857
rect 33361 4831 33362 4857
rect 33334 4129 33362 4831
rect 33334 4103 33335 4129
rect 33361 4103 33362 4129
rect 33334 4073 33362 4103
rect 33334 4047 33335 4073
rect 33361 4047 33362 4073
rect 33334 3402 33362 4047
rect 33334 3345 33362 3374
rect 33334 3319 33335 3345
rect 33361 3319 33362 3345
rect 33334 3289 33362 3319
rect 33334 3263 33335 3289
rect 33361 3263 33362 3289
rect 33334 3257 33362 3263
rect 33670 4913 33698 5671
rect 33726 5642 33754 6398
rect 33782 6145 33810 6151
rect 33782 6119 33783 6145
rect 33809 6119 33810 6145
rect 33782 5866 33810 6119
rect 33782 5833 33810 5838
rect 33726 5595 33754 5614
rect 33838 5361 33866 7631
rect 33894 7993 33922 7999
rect 33894 7967 33895 7993
rect 33921 7967 33922 7993
rect 33894 7322 33922 7967
rect 33950 7574 33978 8414
rect 34398 8395 34426 8414
rect 34958 8442 34986 8447
rect 34958 8050 34986 8414
rect 35070 8441 35098 8470
rect 35126 8465 35154 8470
rect 35238 8498 35266 9086
rect 35854 8833 35882 9198
rect 35854 8807 35855 8833
rect 35881 8807 35882 8833
rect 35854 8777 35882 8807
rect 35854 8751 35855 8777
rect 35881 8751 35882 8777
rect 35854 8745 35882 8751
rect 35070 8415 35071 8441
rect 35097 8415 35098 8441
rect 35070 8409 35098 8415
rect 34958 8049 35098 8050
rect 34958 8023 34959 8049
rect 34985 8023 35098 8049
rect 34958 8022 35098 8023
rect 34958 8017 34986 8022
rect 34573 7854 35035 7859
rect 34573 7853 34582 7854
rect 34573 7827 34574 7853
rect 34573 7826 34582 7827
rect 34610 7826 34634 7854
rect 34662 7826 34686 7854
rect 34714 7853 34738 7854
rect 34766 7853 34790 7854
rect 34724 7827 34738 7853
rect 34786 7827 34790 7853
rect 34714 7826 34738 7827
rect 34766 7826 34790 7827
rect 34818 7853 34842 7854
rect 34870 7853 34894 7854
rect 34818 7827 34822 7853
rect 34870 7827 34884 7853
rect 34818 7826 34842 7827
rect 34870 7826 34894 7827
rect 34922 7826 34946 7854
rect 34974 7826 34998 7854
rect 35026 7853 35035 7854
rect 35034 7827 35035 7853
rect 35026 7826 35035 7827
rect 34573 7821 35035 7826
rect 34398 7657 34426 7663
rect 34398 7631 34399 7657
rect 34425 7631 34426 7657
rect 33950 7546 34034 7574
rect 33894 7289 33922 7294
rect 33894 7210 33922 7215
rect 33894 7163 33922 7182
rect 33950 6818 33978 6823
rect 33894 6426 33922 6431
rect 33894 6379 33922 6398
rect 33838 5335 33839 5361
rect 33865 5335 33866 5361
rect 33838 5305 33866 5335
rect 33838 5279 33839 5305
rect 33865 5279 33866 5305
rect 33838 5082 33866 5279
rect 33838 5049 33866 5054
rect 33894 5642 33922 5647
rect 33894 5250 33922 5614
rect 33670 4887 33671 4913
rect 33697 4887 33698 4913
rect 33670 4129 33698 4887
rect 33782 4914 33810 4919
rect 33894 4914 33922 5222
rect 33782 4913 33922 4914
rect 33782 4887 33783 4913
rect 33809 4887 33895 4913
rect 33921 4887 33922 4913
rect 33782 4886 33922 4887
rect 33782 4881 33810 4886
rect 33894 4881 33922 4886
rect 33838 4578 33866 4583
rect 33950 4578 33978 6790
rect 34006 6706 34034 7546
rect 34398 7546 34426 7631
rect 34398 6874 34426 7518
rect 34678 7266 34706 7271
rect 34678 7219 34706 7238
rect 34573 7070 35035 7075
rect 34573 7069 34582 7070
rect 34573 7043 34574 7069
rect 34573 7042 34582 7043
rect 34610 7042 34634 7070
rect 34662 7042 34686 7070
rect 34714 7069 34738 7070
rect 34766 7069 34790 7070
rect 34724 7043 34738 7069
rect 34786 7043 34790 7069
rect 34714 7042 34738 7043
rect 34766 7042 34790 7043
rect 34818 7069 34842 7070
rect 34870 7069 34894 7070
rect 34818 7043 34822 7069
rect 34870 7043 34884 7069
rect 34818 7042 34842 7043
rect 34870 7042 34894 7043
rect 34922 7042 34946 7070
rect 34974 7042 34998 7070
rect 35026 7069 35035 7070
rect 35034 7043 35035 7069
rect 35026 7042 35035 7043
rect 34573 7037 35035 7042
rect 34398 6808 34426 6846
rect 34678 6874 34706 6879
rect 34006 6673 34034 6678
rect 34398 6762 34426 6767
rect 34398 6089 34426 6734
rect 34678 6481 34706 6846
rect 35070 6762 35098 8022
rect 35238 7713 35266 8470
rect 35854 8049 35882 8055
rect 35854 8023 35855 8049
rect 35881 8023 35882 8049
rect 35854 7994 35882 8023
rect 35854 7993 35994 7994
rect 35854 7967 35855 7993
rect 35881 7967 35994 7993
rect 35854 7966 35994 7967
rect 35854 7961 35882 7966
rect 35238 7687 35239 7713
rect 35265 7687 35266 7713
rect 35238 7657 35266 7687
rect 35238 7631 35239 7657
rect 35265 7631 35266 7657
rect 35238 7625 35266 7631
rect 35630 7322 35658 7327
rect 35126 7265 35154 7271
rect 35126 7239 35127 7265
rect 35153 7239 35154 7265
rect 35126 6929 35154 7239
rect 35126 6903 35127 6929
rect 35153 6903 35154 6929
rect 35126 6873 35154 6903
rect 35126 6847 35127 6873
rect 35153 6847 35154 6873
rect 35126 6818 35154 6847
rect 35126 6785 35154 6790
rect 35350 7265 35378 7271
rect 35350 7239 35351 7265
rect 35377 7239 35378 7265
rect 35350 6818 35378 7239
rect 35070 6729 35098 6734
rect 34678 6455 34679 6481
rect 34705 6455 34706 6481
rect 34678 6449 34706 6455
rect 35238 6482 35266 6487
rect 35350 6482 35378 6790
rect 35238 6481 35378 6482
rect 35238 6455 35239 6481
rect 35265 6455 35351 6481
rect 35377 6455 35378 6481
rect 35238 6454 35378 6455
rect 35238 6449 35266 6454
rect 35350 6449 35378 6454
rect 35518 7154 35546 7159
rect 34573 6286 35035 6291
rect 34573 6285 34582 6286
rect 34573 6259 34574 6285
rect 34573 6258 34582 6259
rect 34610 6258 34634 6286
rect 34662 6258 34686 6286
rect 34714 6285 34738 6286
rect 34766 6285 34790 6286
rect 34724 6259 34738 6285
rect 34786 6259 34790 6285
rect 34714 6258 34738 6259
rect 34766 6258 34790 6259
rect 34818 6285 34842 6286
rect 34870 6285 34894 6286
rect 34818 6259 34822 6285
rect 34870 6259 34884 6285
rect 34818 6258 34842 6259
rect 34870 6258 34894 6259
rect 34922 6258 34946 6286
rect 34974 6258 34998 6286
rect 35026 6285 35035 6286
rect 35034 6259 35035 6285
rect 35026 6258 35035 6259
rect 34573 6253 35035 6258
rect 34398 6063 34399 6089
rect 34425 6063 34426 6089
rect 34398 5698 34426 6063
rect 35126 6145 35154 6151
rect 35126 6119 35127 6145
rect 35153 6119 35154 6145
rect 35126 6089 35154 6119
rect 35126 6063 35127 6089
rect 35153 6063 35154 6089
rect 35126 5922 35154 6063
rect 34958 5698 34986 5703
rect 35126 5698 35154 5894
rect 35518 6090 35546 7126
rect 35630 6930 35658 7294
rect 35742 7210 35770 7215
rect 35742 6930 35770 7182
rect 35910 6930 35938 6935
rect 35630 6929 35714 6930
rect 35630 6903 35631 6929
rect 35657 6903 35714 6929
rect 35630 6902 35714 6903
rect 35630 6897 35658 6902
rect 35630 6090 35658 6095
rect 35518 6089 35658 6090
rect 35518 6063 35631 6089
rect 35657 6063 35658 6089
rect 35518 6062 35658 6063
rect 35350 5698 35378 5703
rect 34398 5697 35098 5698
rect 34398 5671 34959 5697
rect 34985 5671 35098 5697
rect 34398 5670 35098 5671
rect 34958 5665 34986 5670
rect 34573 5502 35035 5507
rect 34573 5501 34582 5502
rect 34573 5475 34574 5501
rect 34573 5474 34582 5475
rect 34610 5474 34634 5502
rect 34662 5474 34686 5502
rect 34714 5501 34738 5502
rect 34766 5501 34790 5502
rect 34724 5475 34738 5501
rect 34786 5475 34790 5501
rect 34714 5474 34738 5475
rect 34766 5474 34790 5475
rect 34818 5501 34842 5502
rect 34870 5501 34894 5502
rect 34818 5475 34822 5501
rect 34870 5475 34884 5501
rect 34818 5474 34842 5475
rect 34870 5474 34894 5475
rect 34922 5474 34946 5502
rect 34974 5474 34998 5502
rect 35026 5501 35035 5502
rect 35034 5475 35035 5501
rect 35026 5474 35035 5475
rect 34573 5469 35035 5474
rect 33838 4577 33978 4578
rect 33838 4551 33839 4577
rect 33865 4551 33978 4577
rect 33838 4550 33978 4551
rect 34174 5306 34202 5311
rect 34174 4914 34202 5278
rect 33838 4521 33866 4550
rect 33838 4495 33839 4521
rect 33865 4495 33866 4521
rect 33670 4103 33671 4129
rect 33697 4103 33698 4129
rect 33670 3345 33698 4103
rect 33670 3319 33671 3345
rect 33697 3319 33698 3345
rect 33670 3010 33698 3319
rect 33334 2898 33362 2903
rect 33334 2618 33362 2870
rect 33334 2561 33362 2590
rect 33334 2535 33335 2561
rect 33361 2535 33362 2561
rect 33334 2505 33362 2535
rect 33670 2562 33698 2982
rect 33670 2515 33698 2534
rect 33782 4129 33810 4135
rect 33782 4103 33783 4129
rect 33809 4103 33810 4129
rect 33782 3346 33810 4103
rect 33838 3794 33866 4495
rect 34174 4522 34202 4886
rect 34510 5082 34538 5087
rect 34510 4522 34538 5054
rect 34678 4914 34706 4919
rect 34678 4867 34706 4886
rect 34573 4718 35035 4723
rect 34573 4717 34582 4718
rect 34573 4691 34574 4717
rect 34573 4690 34582 4691
rect 34610 4690 34634 4718
rect 34662 4690 34686 4718
rect 34714 4717 34738 4718
rect 34766 4717 34790 4718
rect 34724 4691 34738 4717
rect 34786 4691 34790 4717
rect 34714 4690 34738 4691
rect 34766 4690 34790 4691
rect 34818 4717 34842 4718
rect 34870 4717 34894 4718
rect 34818 4691 34822 4717
rect 34870 4691 34884 4717
rect 34818 4690 34842 4691
rect 34870 4690 34894 4691
rect 34922 4690 34946 4718
rect 34974 4690 34998 4718
rect 35026 4717 35035 4718
rect 35034 4691 35035 4717
rect 35026 4690 35035 4691
rect 34573 4685 35035 4690
rect 34622 4606 34874 4634
rect 34622 4522 34650 4606
rect 34510 4521 34650 4522
rect 34510 4495 34623 4521
rect 34649 4495 34650 4521
rect 34510 4494 34650 4495
rect 34174 4456 34202 4494
rect 34622 4489 34650 4494
rect 34678 4522 34706 4527
rect 33950 4129 33978 4135
rect 34678 4130 34706 4494
rect 33950 4103 33951 4129
rect 33977 4103 33978 4129
rect 33894 3794 33922 3799
rect 33838 3793 33922 3794
rect 33838 3767 33895 3793
rect 33921 3767 33922 3793
rect 33838 3766 33922 3767
rect 33782 2954 33810 3318
rect 33782 2562 33810 2926
rect 33894 3737 33922 3766
rect 33894 3711 33895 3737
rect 33921 3711 33922 3737
rect 33894 3290 33922 3711
rect 33950 3346 33978 4103
rect 34510 4129 34706 4130
rect 34510 4103 34679 4129
rect 34705 4103 34706 4129
rect 34510 4102 34706 4103
rect 34174 3738 34202 3743
rect 34174 3691 34202 3710
rect 34510 3346 34538 4102
rect 34678 4097 34706 4102
rect 34846 4521 34874 4606
rect 34846 4495 34847 4521
rect 34873 4495 34874 4521
rect 34846 4130 34874 4495
rect 35070 4410 35098 5670
rect 35070 4377 35098 4382
rect 35126 5697 35378 5698
rect 35126 5671 35127 5697
rect 35153 5671 35351 5697
rect 35377 5671 35378 5697
rect 35126 5670 35378 5671
rect 34846 4097 34874 4102
rect 34573 3934 35035 3939
rect 34573 3933 34582 3934
rect 34573 3907 34574 3933
rect 34573 3906 34582 3907
rect 34610 3906 34634 3934
rect 34662 3906 34686 3934
rect 34714 3933 34738 3934
rect 34766 3933 34790 3934
rect 34724 3907 34738 3933
rect 34786 3907 34790 3933
rect 34714 3906 34738 3907
rect 34766 3906 34790 3907
rect 34818 3933 34842 3934
rect 34870 3933 34894 3934
rect 34818 3907 34822 3933
rect 34870 3907 34884 3933
rect 34818 3906 34842 3907
rect 34870 3906 34894 3907
rect 34922 3906 34946 3934
rect 34974 3906 34998 3934
rect 35026 3933 35035 3934
rect 35034 3907 35035 3933
rect 35026 3906 35035 3907
rect 34573 3901 35035 3906
rect 35126 3793 35154 5670
rect 35350 5665 35378 5670
rect 35238 5361 35266 5367
rect 35238 5335 35239 5361
rect 35265 5335 35266 5361
rect 35238 5306 35266 5335
rect 35238 5259 35266 5278
rect 35126 3767 35127 3793
rect 35153 3767 35154 3793
rect 35070 3738 35098 3743
rect 35126 3738 35154 3767
rect 35070 3737 35154 3738
rect 35070 3711 35071 3737
rect 35097 3711 35154 3737
rect 35070 3710 35154 3711
rect 35182 4130 35210 4135
rect 34678 3346 34706 3351
rect 33950 3299 33978 3318
rect 34454 3345 34706 3346
rect 34454 3319 34679 3345
rect 34705 3319 34706 3345
rect 34454 3318 34706 3319
rect 33894 3009 33922 3262
rect 33894 2983 33895 3009
rect 33921 2983 33922 3009
rect 33894 2953 33922 2983
rect 33894 2927 33895 2953
rect 33921 2927 33922 2953
rect 33894 2898 33922 2927
rect 33894 2865 33922 2870
rect 34454 2953 34482 3318
rect 34678 3313 34706 3318
rect 34573 3150 35035 3155
rect 34573 3149 34582 3150
rect 34573 3123 34574 3149
rect 34573 3122 34582 3123
rect 34610 3122 34634 3150
rect 34662 3122 34686 3150
rect 34714 3149 34738 3150
rect 34766 3149 34790 3150
rect 34724 3123 34738 3149
rect 34786 3123 34790 3149
rect 34714 3122 34738 3123
rect 34766 3122 34790 3123
rect 34818 3149 34842 3150
rect 34870 3149 34894 3150
rect 34818 3123 34822 3149
rect 34870 3123 34884 3149
rect 34818 3122 34842 3123
rect 34870 3122 34894 3123
rect 34922 3122 34946 3150
rect 34974 3122 34998 3150
rect 35026 3149 35035 3150
rect 35034 3123 35035 3149
rect 35026 3122 35035 3123
rect 34573 3117 35035 3122
rect 34454 2927 34455 2953
rect 34481 2927 34482 2953
rect 33894 2562 33922 2567
rect 34454 2562 34482 2927
rect 34678 2618 34706 2623
rect 34678 2562 34706 2590
rect 33782 2561 33922 2562
rect 33782 2535 33783 2561
rect 33809 2535 33895 2561
rect 33921 2535 33922 2561
rect 33782 2534 33922 2535
rect 33782 2529 33810 2534
rect 33894 2529 33922 2534
rect 34398 2561 34706 2562
rect 34398 2535 34679 2561
rect 34705 2535 34706 2561
rect 34398 2534 34706 2535
rect 33334 2479 33335 2505
rect 33361 2479 33362 2505
rect 33334 2473 33362 2479
rect 33278 2170 33306 2175
rect 33446 2170 33474 2175
rect 33278 2169 33474 2170
rect 33278 2143 33279 2169
rect 33305 2143 33447 2169
rect 33473 2143 33474 2169
rect 33278 2142 33474 2143
rect 33278 2137 33306 2142
rect 33446 1777 33474 2142
rect 33446 1751 33447 1777
rect 33473 1751 33474 1777
rect 33446 1722 33474 1751
rect 34398 2169 34426 2534
rect 34678 2529 34706 2534
rect 34398 2143 34399 2169
rect 34425 2143 34426 2169
rect 34398 1777 34426 2143
rect 34398 1751 34399 1777
rect 34425 1751 34426 1777
rect 34398 1745 34426 1751
rect 34510 2450 34538 2455
rect 33446 1689 33474 1694
rect 34510 400 34538 2422
rect 34573 2366 35035 2371
rect 34573 2365 34582 2366
rect 34573 2339 34574 2365
rect 34573 2338 34582 2339
rect 34610 2338 34634 2366
rect 34662 2338 34686 2366
rect 34714 2365 34738 2366
rect 34766 2365 34790 2366
rect 34724 2339 34738 2365
rect 34786 2339 34790 2365
rect 34714 2338 34738 2339
rect 34766 2338 34790 2339
rect 34818 2365 34842 2366
rect 34870 2365 34894 2366
rect 34818 2339 34822 2365
rect 34870 2339 34884 2365
rect 34818 2338 34842 2339
rect 34870 2338 34894 2339
rect 34922 2338 34946 2366
rect 34974 2338 34998 2366
rect 35026 2365 35035 2366
rect 35034 2339 35035 2365
rect 35026 2338 35035 2339
rect 34573 2333 35035 2338
rect 35070 1722 35098 3710
rect 35070 1689 35098 1694
rect 35182 3346 35210 4102
rect 35350 4130 35378 4135
rect 35350 4083 35378 4102
rect 35294 3402 35322 3407
rect 35294 3346 35322 3374
rect 35182 3345 35322 3346
rect 35182 3319 35183 3345
rect 35209 3319 35322 3345
rect 35182 3318 35322 3319
rect 35182 3009 35210 3318
rect 35182 2983 35183 3009
rect 35209 2983 35210 3009
rect 35182 2953 35210 2983
rect 35182 2927 35183 2953
rect 35209 2927 35210 2953
rect 35182 2562 35210 2927
rect 35350 2562 35378 2567
rect 35182 2561 35378 2562
rect 35182 2535 35183 2561
rect 35209 2535 35351 2561
rect 35377 2535 35378 2561
rect 35182 2534 35378 2535
rect 35182 2225 35210 2534
rect 35350 2529 35378 2534
rect 35518 2506 35546 6062
rect 35630 6057 35658 6062
rect 35630 5978 35658 5983
rect 35630 5305 35658 5950
rect 35630 5279 35631 5305
rect 35657 5279 35658 5305
rect 35630 4522 35658 5279
rect 35686 4914 35714 6902
rect 35742 6929 35938 6930
rect 35742 6903 35743 6929
rect 35769 6903 35911 6929
rect 35937 6903 35938 6929
rect 35742 6902 35938 6903
rect 35742 6897 35770 6902
rect 35910 6897 35938 6902
rect 35686 4881 35714 4886
rect 35742 6090 35770 6095
rect 35910 6090 35938 6095
rect 35742 6089 35938 6090
rect 35742 6063 35743 6089
rect 35769 6063 35911 6089
rect 35937 6063 35938 6089
rect 35742 6062 35938 6063
rect 35742 5305 35770 6062
rect 35910 6057 35938 6062
rect 35966 5698 35994 7966
rect 36078 7266 36106 10374
rect 36134 10401 36162 11158
rect 36134 10375 36135 10401
rect 36161 10375 36162 10401
rect 36134 9617 36162 10375
rect 36190 11185 36218 11191
rect 36190 11159 36191 11185
rect 36217 11159 36218 11185
rect 36190 9954 36218 11159
rect 36694 11186 36722 11191
rect 36806 11186 36834 11191
rect 36694 11185 36834 11186
rect 36694 11159 36695 11185
rect 36721 11159 36807 11185
rect 36833 11159 36834 11185
rect 36694 11158 36834 11159
rect 36694 11130 36722 11158
rect 36806 11153 36834 11158
rect 36694 10402 36722 11102
rect 37030 10682 37058 11270
rect 36974 10654 37058 10682
rect 36974 10514 37002 10654
rect 37073 10598 37535 10603
rect 37073 10597 37082 10598
rect 37073 10571 37074 10597
rect 37073 10570 37082 10571
rect 37110 10570 37134 10598
rect 37162 10570 37186 10598
rect 37214 10597 37238 10598
rect 37266 10597 37290 10598
rect 37224 10571 37238 10597
rect 37286 10571 37290 10597
rect 37214 10570 37238 10571
rect 37266 10570 37290 10571
rect 37318 10597 37342 10598
rect 37370 10597 37394 10598
rect 37318 10571 37322 10597
rect 37370 10571 37384 10597
rect 37318 10570 37342 10571
rect 37370 10570 37394 10571
rect 37422 10570 37446 10598
rect 37474 10570 37498 10598
rect 37526 10597 37535 10598
rect 37534 10571 37535 10597
rect 37526 10570 37535 10571
rect 37073 10565 37535 10570
rect 36974 10486 37058 10514
rect 36862 10402 36890 10407
rect 36694 10401 36890 10402
rect 36694 10375 36695 10401
rect 36721 10375 36863 10401
rect 36889 10375 36890 10401
rect 36694 10374 36890 10375
rect 36694 10369 36722 10374
rect 36190 9921 36218 9926
rect 36694 10009 36722 10015
rect 36694 9983 36695 10009
rect 36721 9983 36722 10009
rect 36694 9954 36722 9983
rect 36694 9921 36722 9926
rect 36134 9591 36135 9617
rect 36161 9591 36162 9617
rect 36134 9170 36162 9591
rect 36134 8106 36162 9142
rect 36358 9618 36386 9623
rect 36358 8946 36386 9590
rect 36862 9562 36890 10374
rect 37030 9954 37058 10486
rect 36694 9225 36722 9231
rect 36694 9199 36695 9225
rect 36721 9199 36722 9225
rect 36694 9170 36722 9199
rect 36694 9137 36722 9142
rect 36358 8918 36722 8946
rect 36358 8833 36386 8918
rect 36358 8807 36359 8833
rect 36385 8807 36386 8833
rect 36358 8801 36386 8807
rect 36414 8834 36442 8839
rect 36134 8073 36162 8078
rect 36414 8050 36442 8806
rect 36694 8441 36722 8918
rect 36862 8778 36890 9534
rect 36918 9926 37058 9954
rect 37646 10065 37674 10071
rect 37646 10039 37647 10065
rect 37673 10039 37674 10065
rect 37646 10009 37674 10039
rect 37646 9983 37647 10009
rect 37673 9983 37674 10009
rect 36918 9114 36946 9926
rect 37073 9814 37535 9819
rect 37073 9813 37082 9814
rect 37073 9787 37074 9813
rect 37073 9786 37082 9787
rect 37110 9786 37134 9814
rect 37162 9786 37186 9814
rect 37214 9813 37238 9814
rect 37266 9813 37290 9814
rect 37224 9787 37238 9813
rect 37286 9787 37290 9813
rect 37214 9786 37238 9787
rect 37266 9786 37290 9787
rect 37318 9813 37342 9814
rect 37370 9813 37394 9814
rect 37318 9787 37322 9813
rect 37370 9787 37384 9813
rect 37318 9786 37342 9787
rect 37370 9786 37394 9787
rect 37422 9786 37446 9814
rect 37474 9786 37498 9814
rect 37526 9813 37535 9814
rect 37534 9787 37535 9813
rect 37526 9786 37535 9787
rect 37073 9781 37535 9786
rect 37310 9617 37338 9623
rect 37310 9591 37311 9617
rect 37337 9591 37338 9617
rect 37310 9561 37338 9591
rect 37310 9535 37311 9561
rect 37337 9535 37338 9561
rect 37310 9226 37338 9535
rect 37646 9281 37674 9983
rect 37646 9255 37647 9281
rect 37673 9255 37674 9281
rect 37310 9193 37338 9198
rect 37590 9226 37618 9231
rect 37646 9226 37674 9255
rect 37618 9198 37674 9226
rect 36918 9081 36946 9086
rect 37073 9030 37535 9035
rect 37073 9029 37082 9030
rect 37073 9003 37074 9029
rect 37073 9002 37082 9003
rect 37110 9002 37134 9030
rect 37162 9002 37186 9030
rect 37214 9029 37238 9030
rect 37266 9029 37290 9030
rect 37224 9003 37238 9029
rect 37286 9003 37290 9029
rect 37214 9002 37238 9003
rect 37266 9002 37290 9003
rect 37318 9029 37342 9030
rect 37370 9029 37394 9030
rect 37318 9003 37322 9029
rect 37370 9003 37384 9029
rect 37318 9002 37342 9003
rect 37370 9002 37394 9003
rect 37422 9002 37446 9030
rect 37474 9002 37498 9030
rect 37526 9029 37535 9030
rect 37534 9003 37535 9029
rect 37526 9002 37535 9003
rect 37073 8997 37535 9002
rect 36862 8745 36890 8750
rect 37310 8833 37338 8839
rect 37310 8807 37311 8833
rect 37337 8807 37338 8833
rect 37310 8778 37338 8807
rect 37310 8731 37338 8750
rect 36694 8415 36695 8441
rect 36721 8415 36722 8441
rect 36694 8409 36722 8415
rect 37073 8246 37535 8251
rect 37073 8245 37082 8246
rect 37073 8219 37074 8245
rect 37073 8218 37082 8219
rect 37110 8218 37134 8246
rect 37162 8218 37186 8246
rect 37214 8245 37238 8246
rect 37266 8245 37290 8246
rect 37224 8219 37238 8245
rect 37286 8219 37290 8245
rect 37214 8218 37238 8219
rect 37266 8218 37290 8219
rect 37318 8245 37342 8246
rect 37370 8245 37394 8246
rect 37318 8219 37322 8245
rect 37370 8219 37384 8245
rect 37318 8218 37342 8219
rect 37370 8218 37394 8219
rect 37422 8218 37446 8246
rect 37474 8218 37498 8246
rect 37526 8245 37535 8246
rect 37534 8219 37535 8245
rect 37526 8218 37535 8219
rect 37073 8213 37535 8218
rect 36414 8049 36722 8050
rect 36414 8023 36415 8049
rect 36441 8023 36722 8049
rect 36414 8022 36722 8023
rect 36414 8017 36442 8022
rect 36694 7657 36722 8022
rect 37310 8049 37338 8055
rect 37310 8023 37311 8049
rect 37337 8023 37338 8049
rect 37310 7994 37338 8023
rect 37590 7994 37618 9198
rect 37646 8778 37674 8783
rect 37646 8497 37674 8750
rect 37646 8471 37647 8497
rect 37673 8471 37674 8497
rect 37646 8441 37674 8471
rect 37646 8415 37647 8441
rect 37673 8415 37674 8441
rect 37646 8409 37674 8415
rect 37310 7993 37674 7994
rect 37310 7967 37311 7993
rect 37337 7967 37674 7993
rect 37310 7966 37674 7967
rect 37310 7961 37338 7966
rect 36694 7631 36695 7657
rect 36721 7631 36722 7657
rect 36694 7625 36722 7631
rect 37646 7713 37674 7966
rect 37646 7687 37647 7713
rect 37673 7687 37674 7713
rect 37646 7657 37674 7687
rect 37646 7631 37647 7657
rect 37673 7631 37674 7657
rect 37646 7625 37674 7631
rect 37073 7462 37535 7467
rect 37073 7461 37082 7462
rect 37073 7435 37074 7461
rect 37073 7434 37082 7435
rect 37110 7434 37134 7462
rect 37162 7434 37186 7462
rect 37214 7461 37238 7462
rect 37266 7461 37290 7462
rect 37224 7435 37238 7461
rect 37286 7435 37290 7461
rect 37214 7434 37238 7435
rect 37266 7434 37290 7435
rect 37318 7461 37342 7462
rect 37370 7461 37394 7462
rect 37318 7435 37322 7461
rect 37370 7435 37384 7461
rect 37318 7434 37342 7435
rect 37370 7434 37394 7435
rect 37422 7434 37446 7462
rect 37474 7434 37498 7462
rect 37526 7461 37535 7462
rect 37534 7435 37535 7461
rect 37526 7434 37535 7435
rect 37073 7429 37535 7434
rect 36078 7233 36106 7238
rect 36414 7266 36442 7271
rect 36414 7219 36442 7238
rect 36694 7266 36722 7271
rect 36694 6873 36722 7238
rect 37310 7265 37338 7271
rect 37310 7239 37311 7265
rect 37337 7239 37338 7265
rect 37310 7210 37338 7239
rect 37310 7209 37674 7210
rect 37310 7183 37311 7209
rect 37337 7183 37674 7209
rect 37310 7182 37674 7183
rect 37310 7177 37338 7182
rect 36694 6847 36695 6873
rect 36721 6847 36722 6873
rect 36694 6841 36722 6847
rect 37646 6929 37674 7182
rect 37646 6903 37647 6929
rect 37673 6903 37674 6929
rect 37646 6873 37674 6903
rect 37646 6847 37647 6873
rect 37673 6847 37674 6873
rect 36134 6762 36162 6767
rect 36134 6481 36162 6734
rect 36134 6455 36135 6481
rect 36161 6455 36162 6481
rect 36134 6449 36162 6455
rect 36694 6762 36722 6767
rect 36694 6089 36722 6734
rect 37073 6678 37535 6683
rect 37073 6677 37082 6678
rect 37073 6651 37074 6677
rect 37073 6650 37082 6651
rect 37110 6650 37134 6678
rect 37162 6650 37186 6678
rect 37214 6677 37238 6678
rect 37266 6677 37290 6678
rect 37224 6651 37238 6677
rect 37286 6651 37290 6677
rect 37214 6650 37238 6651
rect 37266 6650 37290 6651
rect 37318 6677 37342 6678
rect 37370 6677 37394 6678
rect 37318 6651 37322 6677
rect 37370 6651 37384 6677
rect 37318 6650 37342 6651
rect 37370 6650 37394 6651
rect 37422 6650 37446 6678
rect 37474 6650 37498 6678
rect 37526 6677 37535 6678
rect 37534 6651 37535 6677
rect 37526 6650 37535 6651
rect 37073 6645 37535 6650
rect 37310 6482 37338 6487
rect 37646 6482 37674 6847
rect 37310 6481 37674 6482
rect 37310 6455 37311 6481
rect 37337 6455 37674 6481
rect 37310 6454 37674 6455
rect 37310 6425 37338 6454
rect 37310 6399 37311 6425
rect 37337 6399 37338 6425
rect 37310 6393 37338 6399
rect 36694 6063 36695 6089
rect 36721 6063 36722 6089
rect 36694 6057 36722 6063
rect 37646 6145 37674 6454
rect 37646 6119 37647 6145
rect 37673 6119 37674 6145
rect 37646 6089 37674 6119
rect 37646 6063 37647 6089
rect 37673 6063 37674 6089
rect 37073 5894 37535 5899
rect 37073 5893 37082 5894
rect 37073 5867 37074 5893
rect 37073 5866 37082 5867
rect 37110 5866 37134 5894
rect 37162 5866 37186 5894
rect 37214 5893 37238 5894
rect 37266 5893 37290 5894
rect 37224 5867 37238 5893
rect 37286 5867 37290 5893
rect 37214 5866 37238 5867
rect 37266 5866 37290 5867
rect 37318 5893 37342 5894
rect 37370 5893 37394 5894
rect 37318 5867 37322 5893
rect 37370 5867 37384 5893
rect 37318 5866 37342 5867
rect 37370 5866 37394 5867
rect 37422 5866 37446 5894
rect 37474 5866 37498 5894
rect 37526 5893 37535 5894
rect 37534 5867 37535 5893
rect 37526 5866 37535 5867
rect 37073 5861 37535 5866
rect 35742 5279 35743 5305
rect 35769 5279 35770 5305
rect 35742 5250 35770 5279
rect 35686 4522 35714 4527
rect 35630 4521 35714 4522
rect 35630 4495 35687 4521
rect 35713 4495 35714 4521
rect 35630 4494 35714 4495
rect 35686 4466 35714 4494
rect 35686 4433 35714 4438
rect 35742 3794 35770 5222
rect 35910 5305 35938 5311
rect 35910 5279 35911 5305
rect 35937 5279 35938 5305
rect 35910 5250 35938 5279
rect 35910 5217 35938 5222
rect 35966 5306 35994 5670
rect 35966 5026 35994 5278
rect 35854 4998 35994 5026
rect 36134 5697 36162 5703
rect 36134 5671 36135 5697
rect 36161 5671 36162 5697
rect 35854 4913 35882 4998
rect 36134 4970 36162 5671
rect 37142 5698 37170 5703
rect 37142 5641 37170 5670
rect 37142 5615 37143 5641
rect 37169 5615 37170 5641
rect 35854 4887 35855 4913
rect 35881 4887 35882 4913
rect 35854 4857 35882 4887
rect 35854 4831 35855 4857
rect 35881 4831 35882 4857
rect 35854 4825 35882 4831
rect 36078 4914 36106 4919
rect 35910 4578 35938 4583
rect 35854 4577 35938 4578
rect 35854 4551 35911 4577
rect 35937 4551 35938 4577
rect 35854 4550 35938 4551
rect 35798 4522 35826 4527
rect 35854 4522 35882 4550
rect 35910 4545 35938 4550
rect 35798 4521 35882 4522
rect 35798 4495 35799 4521
rect 35825 4495 35882 4521
rect 35798 4494 35882 4495
rect 35798 4489 35826 4494
rect 35518 2473 35546 2478
rect 35686 3737 35714 3743
rect 35686 3711 35687 3737
rect 35713 3711 35714 3737
rect 35686 2953 35714 3711
rect 35742 3626 35770 3766
rect 35742 3598 35826 3626
rect 35742 3402 35770 3407
rect 35742 3345 35770 3374
rect 35742 3319 35743 3345
rect 35769 3319 35770 3345
rect 35742 3313 35770 3319
rect 35742 3010 35770 3015
rect 35742 2963 35770 2982
rect 35686 2927 35687 2953
rect 35713 2927 35714 2953
rect 35686 2562 35714 2927
rect 35182 2199 35183 2225
rect 35209 2199 35210 2225
rect 35182 2169 35210 2199
rect 35182 2143 35183 2169
rect 35209 2143 35210 2169
rect 35182 1777 35210 2143
rect 35182 1751 35183 1777
rect 35209 1751 35210 1777
rect 35182 1721 35210 1751
rect 35686 2169 35714 2534
rect 35686 2143 35687 2169
rect 35713 2143 35714 2169
rect 35686 1778 35714 2143
rect 35798 2226 35826 3598
rect 35854 3346 35882 4494
rect 35910 3794 35938 3799
rect 35910 3747 35938 3766
rect 35854 3010 35882 3318
rect 35910 3010 35938 3015
rect 35854 2982 35910 3010
rect 35910 2963 35938 2982
rect 35910 2226 35938 2231
rect 35798 2225 35938 2226
rect 35798 2199 35911 2225
rect 35937 2199 35938 2225
rect 35798 2198 35938 2199
rect 35798 2169 35826 2198
rect 35910 2193 35938 2198
rect 35798 2143 35799 2169
rect 35825 2143 35826 2169
rect 35798 2137 35826 2143
rect 35686 1745 35714 1750
rect 35182 1695 35183 1721
rect 35209 1695 35210 1721
rect 35182 1689 35210 1695
rect 36078 1694 36106 4886
rect 36134 4913 36162 4942
rect 36134 4887 36135 4913
rect 36161 4887 36162 4913
rect 36134 4881 36162 4887
rect 36694 5305 36722 5311
rect 36694 5279 36695 5305
rect 36721 5279 36722 5305
rect 36694 4970 36722 5279
rect 37142 5306 37170 5615
rect 37590 5641 37618 5647
rect 37590 5615 37591 5641
rect 37617 5615 37618 5641
rect 37366 5306 37394 5311
rect 37142 5305 37394 5306
rect 37142 5279 37143 5305
rect 37169 5279 37367 5305
rect 37393 5279 37394 5305
rect 37142 5278 37394 5279
rect 37142 5194 37170 5278
rect 37366 5273 37394 5278
rect 36974 5166 37170 5194
rect 36974 5026 37002 5166
rect 37073 5110 37535 5115
rect 37073 5109 37082 5110
rect 37073 5083 37074 5109
rect 37073 5082 37082 5083
rect 37110 5082 37134 5110
rect 37162 5082 37186 5110
rect 37214 5109 37238 5110
rect 37266 5109 37290 5110
rect 37224 5083 37238 5109
rect 37286 5083 37290 5109
rect 37214 5082 37238 5083
rect 37266 5082 37290 5083
rect 37318 5109 37342 5110
rect 37370 5109 37394 5110
rect 37318 5083 37322 5109
rect 37370 5083 37384 5109
rect 37318 5082 37342 5083
rect 37370 5082 37394 5083
rect 37422 5082 37446 5110
rect 37474 5082 37498 5110
rect 37526 5109 37535 5110
rect 37534 5083 37535 5109
rect 37526 5082 37535 5083
rect 37073 5077 37535 5082
rect 36974 4998 37058 5026
rect 36694 4521 36722 4942
rect 36694 4495 36695 4521
rect 36721 4495 36722 4521
rect 36694 4489 36722 4495
rect 36862 4970 36890 4975
rect 36134 4129 36162 4135
rect 36134 4103 36135 4129
rect 36161 4103 36162 4129
rect 36134 3345 36162 4103
rect 36134 3319 36135 3345
rect 36161 3319 36162 3345
rect 36134 2954 36162 3319
rect 36694 3402 36722 3407
rect 36694 3346 36722 3374
rect 36862 3346 36890 4942
rect 37030 4802 37058 4998
rect 37310 4970 37338 4975
rect 37310 4913 37338 4942
rect 37310 4887 37311 4913
rect 37337 4887 37338 4913
rect 37310 4857 37338 4887
rect 37590 4914 37618 5615
rect 37590 4867 37618 4886
rect 37646 4970 37674 6063
rect 37702 5642 37730 5647
rect 37870 5642 37898 5647
rect 37702 5641 37898 5642
rect 37702 5615 37703 5641
rect 37729 5615 37871 5641
rect 37897 5615 37898 5641
rect 37702 5614 37898 5615
rect 37702 5250 37730 5614
rect 37870 5609 37898 5614
rect 37702 5217 37730 5222
rect 38150 5305 38178 5311
rect 38150 5279 38151 5305
rect 38177 5279 38178 5305
rect 37310 4831 37311 4857
rect 37337 4831 37338 4857
rect 37310 4825 37338 4831
rect 36974 4774 37058 4802
rect 36974 4130 37002 4774
rect 37646 4577 37674 4942
rect 37758 4914 37786 4919
rect 37870 4914 37898 4919
rect 37758 4913 37898 4914
rect 37758 4887 37759 4913
rect 37785 4887 37871 4913
rect 37897 4887 37898 4913
rect 37758 4886 37898 4887
rect 37758 4881 37786 4886
rect 37646 4551 37647 4577
rect 37673 4551 37674 4577
rect 37646 4521 37674 4551
rect 37870 4578 37898 4886
rect 38150 4914 38178 5279
rect 38262 5305 38290 5311
rect 38262 5279 38263 5305
rect 38289 5279 38290 5305
rect 38262 5250 38290 5279
rect 38262 5217 38290 5222
rect 38430 5305 38458 5311
rect 38430 5279 38431 5305
rect 38457 5279 38458 5305
rect 38430 5250 38458 5279
rect 38430 5217 38458 5222
rect 38598 5250 38626 5255
rect 38598 5026 38626 5222
rect 38598 4998 38682 5026
rect 37898 4550 37954 4578
rect 37870 4545 37898 4550
rect 37646 4495 37647 4521
rect 37673 4495 37674 4521
rect 37646 4489 37674 4495
rect 37590 4466 37618 4471
rect 37073 4326 37535 4331
rect 37073 4325 37082 4326
rect 37073 4299 37074 4325
rect 37073 4298 37082 4299
rect 37110 4298 37134 4326
rect 37162 4298 37186 4326
rect 37214 4325 37238 4326
rect 37266 4325 37290 4326
rect 37224 4299 37238 4325
rect 37286 4299 37290 4325
rect 37214 4298 37238 4299
rect 37266 4298 37290 4299
rect 37318 4325 37342 4326
rect 37370 4325 37394 4326
rect 37318 4299 37322 4325
rect 37370 4299 37384 4325
rect 37318 4298 37342 4299
rect 37370 4298 37394 4299
rect 37422 4298 37446 4326
rect 37474 4298 37498 4326
rect 37526 4325 37535 4326
rect 37534 4299 37535 4325
rect 37526 4298 37535 4299
rect 37073 4293 37535 4298
rect 37086 4130 37114 4135
rect 36974 4129 37114 4130
rect 36974 4103 37087 4129
rect 37113 4103 37114 4129
rect 36974 4102 37114 4103
rect 37086 4073 37114 4102
rect 37086 4047 37087 4073
rect 37113 4047 37114 4073
rect 37086 4041 37114 4047
rect 37590 4129 37618 4438
rect 37590 4103 37591 4129
rect 37617 4103 37618 4129
rect 36918 3794 36946 3799
rect 36918 3793 37002 3794
rect 36918 3767 36919 3793
rect 36945 3767 37002 3793
rect 36918 3766 37002 3767
rect 36918 3761 36946 3766
rect 36974 3737 37002 3766
rect 36974 3711 36975 3737
rect 37001 3711 37002 3737
rect 36974 3458 37002 3711
rect 37073 3542 37535 3547
rect 37073 3541 37082 3542
rect 37073 3515 37074 3541
rect 37073 3514 37082 3515
rect 37110 3514 37134 3542
rect 37162 3514 37186 3542
rect 37214 3541 37238 3542
rect 37266 3541 37290 3542
rect 37224 3515 37238 3541
rect 37286 3515 37290 3541
rect 37214 3514 37238 3515
rect 37266 3514 37290 3515
rect 37318 3541 37342 3542
rect 37370 3541 37394 3542
rect 37318 3515 37322 3541
rect 37370 3515 37384 3541
rect 37318 3514 37342 3515
rect 37370 3514 37394 3515
rect 37422 3514 37446 3542
rect 37474 3514 37498 3542
rect 37526 3541 37535 3542
rect 37534 3515 37535 3541
rect 37526 3514 37535 3515
rect 37073 3509 37535 3514
rect 36974 3430 37058 3458
rect 36694 3345 36890 3346
rect 36694 3319 36695 3345
rect 36721 3319 36863 3345
rect 36889 3319 36890 3345
rect 36694 3318 36890 3319
rect 36694 3313 36722 3318
rect 36134 2618 36162 2926
rect 36694 2954 36722 2959
rect 36694 2907 36722 2926
rect 36862 2954 36890 3318
rect 37030 3290 37058 3430
rect 37030 3010 37058 3262
rect 36134 2561 36162 2590
rect 36134 2535 36135 2561
rect 36161 2535 36162 2561
rect 36134 2529 36162 2535
rect 36694 2562 36722 2567
rect 36862 2562 36890 2926
rect 36974 2982 37058 3010
rect 37590 3346 37618 4103
rect 37646 4410 37674 4415
rect 37646 3737 37674 4382
rect 37702 4130 37730 4135
rect 37702 4083 37730 4102
rect 37870 4130 37898 4135
rect 37870 4083 37898 4102
rect 37646 3711 37647 3737
rect 37673 3711 37674 3737
rect 37646 3705 37674 3711
rect 36974 2674 37002 2982
rect 37142 2954 37170 2959
rect 37142 2907 37170 2926
rect 37366 2954 37394 2959
rect 37366 2907 37394 2926
rect 37073 2758 37535 2763
rect 37073 2757 37082 2758
rect 37073 2731 37074 2757
rect 37073 2730 37082 2731
rect 37110 2730 37134 2758
rect 37162 2730 37186 2758
rect 37214 2757 37238 2758
rect 37266 2757 37290 2758
rect 37224 2731 37238 2757
rect 37286 2731 37290 2757
rect 37214 2730 37238 2731
rect 37266 2730 37290 2731
rect 37318 2757 37342 2758
rect 37370 2757 37394 2758
rect 37318 2731 37322 2757
rect 37370 2731 37384 2757
rect 37318 2730 37342 2731
rect 37370 2730 37394 2731
rect 37422 2730 37446 2758
rect 37474 2730 37498 2758
rect 37526 2757 37535 2758
rect 37534 2731 37535 2757
rect 37526 2730 37535 2731
rect 37073 2725 37535 2730
rect 36974 2646 37226 2674
rect 36694 2561 36890 2562
rect 36694 2535 36695 2561
rect 36721 2535 36863 2561
rect 36889 2535 36890 2561
rect 36694 2534 36890 2535
rect 36694 2529 36722 2534
rect 36862 2529 36890 2534
rect 37198 2170 37226 2646
rect 37590 2561 37618 3318
rect 37926 3345 37954 4550
rect 38150 4577 38178 4886
rect 38654 4914 38682 4998
rect 38766 4914 38794 4919
rect 38654 4913 38794 4914
rect 38654 4887 38655 4913
rect 38681 4887 38767 4913
rect 38793 4887 38794 4913
rect 38654 4886 38794 4887
rect 38654 4881 38682 4886
rect 38150 4551 38151 4577
rect 38177 4551 38178 4577
rect 38150 4545 38178 4551
rect 38262 4578 38290 4583
rect 38262 4531 38290 4550
rect 38430 4578 38458 4583
rect 38430 4531 38458 4550
rect 38710 4578 38738 4886
rect 38766 4881 38794 4886
rect 38878 4914 38906 4919
rect 38906 4886 38962 4914
rect 38878 4867 38906 4886
rect 38710 4577 38850 4578
rect 38710 4551 38711 4577
rect 38737 4551 38850 4577
rect 38710 4550 38850 4551
rect 38710 4545 38738 4550
rect 38262 4130 38290 4135
rect 38262 3794 38290 4102
rect 38654 4130 38682 4135
rect 38766 4130 38794 4550
rect 38822 4521 38850 4550
rect 38822 4495 38823 4521
rect 38849 4495 38850 4521
rect 38822 4489 38850 4495
rect 38934 4521 38962 4886
rect 38934 4495 38935 4521
rect 38961 4495 38962 4521
rect 38934 4489 38962 4495
rect 38682 4129 38794 4130
rect 38682 4103 38767 4129
rect 38793 4103 38794 4129
rect 38682 4102 38794 4103
rect 38654 4064 38682 4102
rect 38430 3794 38458 3799
rect 38262 3793 38458 3794
rect 38262 3767 38263 3793
rect 38289 3767 38431 3793
rect 38457 3767 38458 3793
rect 38262 3766 38458 3767
rect 38262 3761 38290 3766
rect 38430 3761 38458 3766
rect 38710 3794 38738 4102
rect 38766 4097 38794 4102
rect 38934 4074 38962 4079
rect 38934 4073 39018 4074
rect 38934 4047 38935 4073
rect 38961 4047 39018 4073
rect 38934 4046 39018 4047
rect 38934 4041 38962 4046
rect 38710 3793 38850 3794
rect 38710 3767 38711 3793
rect 38737 3767 38850 3793
rect 38710 3766 38850 3767
rect 38710 3761 38738 3766
rect 37926 3319 37927 3345
rect 37953 3319 37954 3345
rect 37590 2535 37591 2561
rect 37617 2535 37618 2561
rect 37590 2529 37618 2535
rect 37702 3290 37730 3295
rect 37702 3010 37730 3262
rect 37926 3290 37954 3319
rect 37926 3257 37954 3262
rect 38150 3737 38178 3743
rect 38150 3711 38151 3737
rect 38177 3711 38178 3737
rect 38150 3346 38178 3711
rect 37702 2562 37730 2982
rect 38150 3009 38178 3318
rect 38654 3346 38682 3351
rect 38766 3346 38794 3766
rect 38822 3737 38850 3766
rect 38822 3711 38823 3737
rect 38849 3711 38850 3737
rect 38822 3705 38850 3711
rect 38990 3738 39018 4046
rect 38990 3737 39074 3738
rect 38990 3711 38991 3737
rect 39017 3711 39074 3737
rect 38990 3710 39074 3711
rect 38990 3705 39018 3710
rect 38654 3345 38794 3346
rect 38654 3319 38655 3345
rect 38681 3319 38767 3345
rect 38793 3319 38794 3345
rect 38654 3318 38794 3319
rect 38654 3313 38682 3318
rect 38150 2983 38151 3009
rect 38177 2983 38178 3009
rect 37870 2562 37898 2567
rect 37702 2561 37898 2562
rect 37702 2535 37703 2561
rect 37729 2535 37871 2561
rect 37897 2535 37898 2561
rect 37702 2534 37898 2535
rect 37702 2529 37730 2534
rect 37870 2529 37898 2534
rect 38150 2562 38178 2983
rect 38150 2529 38178 2534
rect 38262 3290 38290 3295
rect 38262 3010 38290 3262
rect 38430 3010 38458 3015
rect 38262 3009 38458 3010
rect 38262 2983 38263 3009
rect 38289 2983 38431 3009
rect 38457 2983 38458 3009
rect 38262 2982 38458 2983
rect 37310 2170 37338 2175
rect 37198 2169 37338 2170
rect 37198 2143 37199 2169
rect 37225 2143 37311 2169
rect 37337 2143 37338 2169
rect 37198 2142 37338 2143
rect 37198 2137 37226 2142
rect 37310 2137 37338 2142
rect 37590 2169 37618 2175
rect 37590 2143 37591 2169
rect 37617 2143 37618 2169
rect 37073 1974 37535 1979
rect 37073 1973 37082 1974
rect 37073 1947 37074 1973
rect 37073 1946 37082 1947
rect 37110 1946 37134 1974
rect 37162 1946 37186 1974
rect 37214 1973 37238 1974
rect 37266 1973 37290 1974
rect 37224 1947 37238 1973
rect 37286 1947 37290 1973
rect 37214 1946 37238 1947
rect 37266 1946 37290 1947
rect 37318 1973 37342 1974
rect 37370 1973 37394 1974
rect 37318 1947 37322 1973
rect 37370 1947 37384 1973
rect 37318 1946 37342 1947
rect 37370 1946 37394 1947
rect 37422 1946 37446 1974
rect 37474 1946 37498 1974
rect 37526 1973 37535 1974
rect 37534 1947 37535 1973
rect 37526 1946 37535 1947
rect 37073 1941 37535 1946
rect 36190 1890 36218 1895
rect 36190 1777 36218 1862
rect 37590 1890 37618 2143
rect 37590 1857 37618 1862
rect 38150 2169 38178 2175
rect 38150 2143 38151 2169
rect 38177 2143 38178 2169
rect 38150 1834 38178 2143
rect 36190 1751 36191 1777
rect 36217 1751 36218 1777
rect 36190 1745 36218 1751
rect 37142 1777 37170 1783
rect 37142 1751 37143 1777
rect 37169 1751 37170 1777
rect 35966 1666 36106 1694
rect 37142 1722 37170 1751
rect 37142 1689 37170 1694
rect 37422 1778 37450 1783
rect 34573 1582 35035 1587
rect 34573 1581 34582 1582
rect 34573 1555 34574 1581
rect 34573 1554 34582 1555
rect 34610 1554 34634 1582
rect 34662 1554 34686 1582
rect 34714 1581 34738 1582
rect 34766 1581 34790 1582
rect 34724 1555 34738 1581
rect 34786 1555 34790 1581
rect 34714 1554 34738 1555
rect 34766 1554 34790 1555
rect 34818 1581 34842 1582
rect 34870 1581 34894 1582
rect 34818 1555 34822 1581
rect 34870 1555 34884 1581
rect 34818 1554 34842 1555
rect 34870 1554 34894 1555
rect 34922 1554 34946 1582
rect 34974 1554 34998 1582
rect 35026 1581 35035 1582
rect 35034 1555 35035 1581
rect 35026 1554 35035 1555
rect 34573 1549 35035 1554
rect 35966 400 35994 1666
rect 37422 400 37450 1750
rect 38150 1777 38178 1806
rect 38150 1751 38151 1777
rect 38177 1751 38178 1777
rect 38150 1745 38178 1751
rect 38262 1778 38290 2982
rect 38430 2618 38458 2982
rect 38710 3010 38738 3318
rect 38766 3313 38794 3318
rect 38878 3345 38906 3351
rect 38878 3319 38879 3345
rect 38905 3319 38906 3345
rect 38710 3009 38850 3010
rect 38710 2983 38711 3009
rect 38737 2983 38850 3009
rect 38710 2982 38850 2983
rect 38710 2977 38738 2982
rect 38430 2585 38458 2590
rect 38766 2561 38794 2982
rect 38822 2953 38850 2982
rect 38822 2927 38823 2953
rect 38849 2927 38850 2953
rect 38822 2921 38850 2927
rect 38878 2954 38906 3319
rect 38934 2954 38962 2959
rect 38878 2953 38962 2954
rect 38878 2927 38935 2953
rect 38961 2927 38962 2953
rect 38878 2926 38962 2927
rect 38766 2535 38767 2561
rect 38793 2535 38794 2561
rect 38654 2506 38682 2511
rect 38766 2506 38794 2535
rect 38654 2505 38794 2506
rect 38654 2479 38655 2505
rect 38681 2479 38794 2505
rect 38654 2478 38794 2479
rect 38822 2618 38850 2623
rect 38654 2394 38682 2478
rect 38486 2366 38682 2394
rect 38318 2170 38346 2175
rect 38486 2170 38514 2366
rect 38822 2282 38850 2590
rect 38878 2562 38906 2926
rect 38934 2921 38962 2926
rect 38906 2534 38962 2562
rect 38878 2515 38906 2534
rect 38710 2254 38906 2282
rect 38710 2225 38738 2254
rect 38710 2199 38711 2225
rect 38737 2199 38738 2225
rect 38710 2193 38738 2199
rect 38878 2225 38906 2254
rect 38878 2199 38879 2225
rect 38905 2199 38906 2225
rect 38878 2193 38906 2199
rect 38318 2169 38514 2170
rect 38318 2143 38319 2169
rect 38345 2143 38487 2169
rect 38513 2143 38514 2169
rect 38318 2142 38514 2143
rect 38318 2137 38346 2142
rect 38430 1778 38458 1783
rect 38262 1777 38458 1778
rect 38262 1751 38263 1777
rect 38289 1751 38431 1777
rect 38457 1751 38458 1777
rect 38262 1750 38458 1751
rect 38486 1778 38514 2142
rect 38934 1946 38962 2534
rect 38990 2506 39018 2511
rect 39046 2506 39074 3710
rect 39018 2478 39074 2506
rect 38990 2225 39018 2478
rect 38990 2199 38991 2225
rect 39017 2199 39018 2225
rect 38990 2193 39018 2199
rect 38934 1918 39018 1946
rect 38934 1834 38962 1839
rect 38654 1778 38682 1783
rect 38486 1750 38654 1778
rect 38262 1745 38290 1750
rect 38430 1745 38458 1750
rect 38654 1712 38682 1750
rect 38822 1778 38850 1797
rect 38822 1745 38850 1750
rect 38934 1777 38962 1806
rect 38934 1751 38935 1777
rect 38961 1751 38962 1777
rect 38934 1745 38962 1751
rect 38990 1694 39018 1918
rect 38878 1666 39018 1694
rect 38878 400 38906 1666
rect 25438 350 25634 378
rect 25760 0 25816 400
rect 27216 0 27272 400
rect 28672 0 28728 400
rect 30128 0 30184 400
rect 31584 0 31640 400
rect 33040 0 33096 400
rect 34496 0 34552 400
rect 35952 0 36008 400
rect 37408 0 37464 400
rect 38864 0 38920 400
<< via2 >>
rect 2082 18437 2110 18438
rect 2082 18411 2100 18437
rect 2100 18411 2110 18437
rect 2082 18410 2110 18411
rect 2134 18437 2162 18438
rect 2134 18411 2136 18437
rect 2136 18411 2162 18437
rect 2134 18410 2162 18411
rect 2186 18437 2214 18438
rect 2238 18437 2266 18438
rect 2186 18411 2198 18437
rect 2198 18411 2214 18437
rect 2238 18411 2260 18437
rect 2260 18411 2266 18437
rect 2186 18410 2214 18411
rect 2238 18410 2266 18411
rect 2290 18410 2318 18438
rect 2342 18437 2370 18438
rect 2394 18437 2422 18438
rect 2342 18411 2348 18437
rect 2348 18411 2370 18437
rect 2394 18411 2410 18437
rect 2410 18411 2422 18437
rect 2342 18410 2370 18411
rect 2394 18410 2422 18411
rect 2446 18437 2474 18438
rect 2446 18411 2472 18437
rect 2472 18411 2474 18437
rect 2446 18410 2474 18411
rect 2498 18437 2526 18438
rect 2498 18411 2508 18437
rect 2508 18411 2526 18437
rect 2498 18410 2526 18411
rect 2082 17653 2110 17654
rect 2082 17627 2100 17653
rect 2100 17627 2110 17653
rect 2082 17626 2110 17627
rect 2134 17653 2162 17654
rect 2134 17627 2136 17653
rect 2136 17627 2162 17653
rect 2134 17626 2162 17627
rect 2186 17653 2214 17654
rect 2238 17653 2266 17654
rect 2186 17627 2198 17653
rect 2198 17627 2214 17653
rect 2238 17627 2260 17653
rect 2260 17627 2266 17653
rect 2186 17626 2214 17627
rect 2238 17626 2266 17627
rect 2290 17626 2318 17654
rect 2342 17653 2370 17654
rect 2394 17653 2422 17654
rect 2342 17627 2348 17653
rect 2348 17627 2370 17653
rect 2394 17627 2410 17653
rect 2410 17627 2422 17653
rect 2342 17626 2370 17627
rect 2394 17626 2422 17627
rect 2446 17653 2474 17654
rect 2446 17627 2472 17653
rect 2472 17627 2474 17653
rect 2446 17626 2474 17627
rect 2498 17653 2526 17654
rect 2498 17627 2508 17653
rect 2508 17627 2526 17653
rect 2498 17626 2526 17627
rect 2082 16869 2110 16870
rect 2082 16843 2100 16869
rect 2100 16843 2110 16869
rect 2082 16842 2110 16843
rect 2134 16869 2162 16870
rect 2134 16843 2136 16869
rect 2136 16843 2162 16869
rect 2134 16842 2162 16843
rect 2186 16869 2214 16870
rect 2238 16869 2266 16870
rect 2186 16843 2198 16869
rect 2198 16843 2214 16869
rect 2238 16843 2260 16869
rect 2260 16843 2266 16869
rect 2186 16842 2214 16843
rect 2238 16842 2266 16843
rect 2290 16842 2318 16870
rect 2342 16869 2370 16870
rect 2394 16869 2422 16870
rect 2342 16843 2348 16869
rect 2348 16843 2370 16869
rect 2394 16843 2410 16869
rect 2410 16843 2422 16869
rect 2342 16842 2370 16843
rect 2394 16842 2422 16843
rect 2446 16869 2474 16870
rect 2446 16843 2472 16869
rect 2472 16843 2474 16869
rect 2446 16842 2474 16843
rect 2498 16869 2526 16870
rect 2498 16843 2508 16869
rect 2508 16843 2526 16869
rect 2498 16842 2526 16843
rect 2082 16085 2110 16086
rect 2082 16059 2100 16085
rect 2100 16059 2110 16085
rect 2082 16058 2110 16059
rect 2134 16085 2162 16086
rect 2134 16059 2136 16085
rect 2136 16059 2162 16085
rect 2134 16058 2162 16059
rect 2186 16085 2214 16086
rect 2238 16085 2266 16086
rect 2186 16059 2198 16085
rect 2198 16059 2214 16085
rect 2238 16059 2260 16085
rect 2260 16059 2266 16085
rect 2186 16058 2214 16059
rect 2238 16058 2266 16059
rect 2290 16058 2318 16086
rect 2342 16085 2370 16086
rect 2394 16085 2422 16086
rect 2342 16059 2348 16085
rect 2348 16059 2370 16085
rect 2394 16059 2410 16085
rect 2410 16059 2422 16085
rect 2342 16058 2370 16059
rect 2394 16058 2422 16059
rect 2446 16085 2474 16086
rect 2446 16059 2472 16085
rect 2472 16059 2474 16085
rect 2446 16058 2474 16059
rect 2498 16085 2526 16086
rect 2498 16059 2508 16085
rect 2508 16059 2526 16085
rect 2498 16058 2526 16059
rect 2082 15301 2110 15302
rect 2082 15275 2100 15301
rect 2100 15275 2110 15301
rect 2082 15274 2110 15275
rect 2134 15301 2162 15302
rect 2134 15275 2136 15301
rect 2136 15275 2162 15301
rect 2134 15274 2162 15275
rect 2186 15301 2214 15302
rect 2238 15301 2266 15302
rect 2186 15275 2198 15301
rect 2198 15275 2214 15301
rect 2238 15275 2260 15301
rect 2260 15275 2266 15301
rect 2186 15274 2214 15275
rect 2238 15274 2266 15275
rect 2290 15274 2318 15302
rect 2342 15301 2370 15302
rect 2394 15301 2422 15302
rect 2342 15275 2348 15301
rect 2348 15275 2370 15301
rect 2394 15275 2410 15301
rect 2410 15275 2422 15301
rect 2342 15274 2370 15275
rect 2394 15274 2422 15275
rect 2446 15301 2474 15302
rect 2446 15275 2472 15301
rect 2472 15275 2474 15301
rect 2446 15274 2474 15275
rect 2498 15301 2526 15302
rect 2498 15275 2508 15301
rect 2508 15275 2526 15301
rect 2498 15274 2526 15275
rect 1974 14686 2002 14714
rect 1582 9198 1610 9226
rect 2478 14713 2506 14714
rect 2478 14687 2479 14713
rect 2479 14687 2505 14713
rect 2505 14687 2506 14713
rect 2478 14686 2506 14687
rect 2082 14517 2110 14518
rect 2082 14491 2100 14517
rect 2100 14491 2110 14517
rect 2082 14490 2110 14491
rect 2134 14517 2162 14518
rect 2134 14491 2136 14517
rect 2136 14491 2162 14517
rect 2134 14490 2162 14491
rect 2186 14517 2214 14518
rect 2238 14517 2266 14518
rect 2186 14491 2198 14517
rect 2198 14491 2214 14517
rect 2238 14491 2260 14517
rect 2260 14491 2266 14517
rect 2186 14490 2214 14491
rect 2238 14490 2266 14491
rect 2290 14490 2318 14518
rect 2342 14517 2370 14518
rect 2394 14517 2422 14518
rect 2342 14491 2348 14517
rect 2348 14491 2370 14517
rect 2394 14491 2410 14517
rect 2410 14491 2422 14517
rect 2342 14490 2370 14491
rect 2394 14490 2422 14491
rect 2446 14517 2474 14518
rect 2446 14491 2472 14517
rect 2472 14491 2474 14517
rect 2446 14490 2474 14491
rect 2498 14517 2526 14518
rect 2498 14491 2508 14517
rect 2508 14491 2526 14517
rect 2498 14490 2526 14491
rect 4582 18045 4610 18046
rect 4582 18019 4600 18045
rect 4600 18019 4610 18045
rect 4582 18018 4610 18019
rect 4634 18045 4662 18046
rect 4634 18019 4636 18045
rect 4636 18019 4662 18045
rect 4634 18018 4662 18019
rect 4686 18045 4714 18046
rect 4738 18045 4766 18046
rect 4686 18019 4698 18045
rect 4698 18019 4714 18045
rect 4738 18019 4760 18045
rect 4760 18019 4766 18045
rect 4686 18018 4714 18019
rect 4738 18018 4766 18019
rect 4790 18018 4818 18046
rect 4842 18045 4870 18046
rect 4894 18045 4922 18046
rect 4842 18019 4848 18045
rect 4848 18019 4870 18045
rect 4894 18019 4910 18045
rect 4910 18019 4922 18045
rect 4842 18018 4870 18019
rect 4894 18018 4922 18019
rect 4946 18045 4974 18046
rect 4946 18019 4972 18045
rect 4972 18019 4974 18045
rect 4946 18018 4974 18019
rect 4998 18045 5026 18046
rect 4998 18019 5008 18045
rect 5008 18019 5026 18045
rect 4998 18018 5026 18019
rect 4582 17261 4610 17262
rect 4582 17235 4600 17261
rect 4600 17235 4610 17261
rect 4582 17234 4610 17235
rect 4634 17261 4662 17262
rect 4634 17235 4636 17261
rect 4636 17235 4662 17261
rect 4634 17234 4662 17235
rect 4686 17261 4714 17262
rect 4738 17261 4766 17262
rect 4686 17235 4698 17261
rect 4698 17235 4714 17261
rect 4738 17235 4760 17261
rect 4760 17235 4766 17261
rect 4686 17234 4714 17235
rect 4738 17234 4766 17235
rect 4790 17234 4818 17262
rect 4842 17261 4870 17262
rect 4894 17261 4922 17262
rect 4842 17235 4848 17261
rect 4848 17235 4870 17261
rect 4894 17235 4910 17261
rect 4910 17235 4922 17261
rect 4842 17234 4870 17235
rect 4894 17234 4922 17235
rect 4946 17261 4974 17262
rect 4946 17235 4972 17261
rect 4972 17235 4974 17261
rect 4946 17234 4974 17235
rect 4998 17261 5026 17262
rect 4998 17235 5008 17261
rect 5008 17235 5026 17261
rect 4998 17234 5026 17235
rect 4582 16477 4610 16478
rect 4582 16451 4600 16477
rect 4600 16451 4610 16477
rect 4582 16450 4610 16451
rect 4634 16477 4662 16478
rect 4634 16451 4636 16477
rect 4636 16451 4662 16477
rect 4634 16450 4662 16451
rect 4686 16477 4714 16478
rect 4738 16477 4766 16478
rect 4686 16451 4698 16477
rect 4698 16451 4714 16477
rect 4738 16451 4760 16477
rect 4760 16451 4766 16477
rect 4686 16450 4714 16451
rect 4738 16450 4766 16451
rect 4790 16450 4818 16478
rect 4842 16477 4870 16478
rect 4894 16477 4922 16478
rect 4842 16451 4848 16477
rect 4848 16451 4870 16477
rect 4894 16451 4910 16477
rect 4910 16451 4922 16477
rect 4842 16450 4870 16451
rect 4894 16450 4922 16451
rect 4946 16477 4974 16478
rect 4946 16451 4972 16477
rect 4972 16451 4974 16477
rect 4946 16450 4974 16451
rect 4998 16477 5026 16478
rect 4998 16451 5008 16477
rect 5008 16451 5026 16477
rect 4998 16450 5026 16451
rect 4582 15693 4610 15694
rect 4582 15667 4600 15693
rect 4600 15667 4610 15693
rect 4582 15666 4610 15667
rect 4634 15693 4662 15694
rect 4634 15667 4636 15693
rect 4636 15667 4662 15693
rect 4634 15666 4662 15667
rect 4686 15693 4714 15694
rect 4738 15693 4766 15694
rect 4686 15667 4698 15693
rect 4698 15667 4714 15693
rect 4738 15667 4760 15693
rect 4760 15667 4766 15693
rect 4686 15666 4714 15667
rect 4738 15666 4766 15667
rect 4790 15666 4818 15694
rect 4842 15693 4870 15694
rect 4894 15693 4922 15694
rect 4842 15667 4848 15693
rect 4848 15667 4870 15693
rect 4894 15667 4910 15693
rect 4910 15667 4922 15693
rect 4842 15666 4870 15667
rect 4894 15666 4922 15667
rect 4946 15693 4974 15694
rect 4946 15667 4972 15693
rect 4972 15667 4974 15693
rect 4946 15666 4974 15667
rect 4998 15693 5026 15694
rect 4998 15667 5008 15693
rect 5008 15667 5026 15693
rect 4998 15666 5026 15667
rect 2646 14686 2674 14714
rect 2082 13733 2110 13734
rect 2082 13707 2100 13733
rect 2100 13707 2110 13733
rect 2082 13706 2110 13707
rect 2134 13733 2162 13734
rect 2134 13707 2136 13733
rect 2136 13707 2162 13733
rect 2134 13706 2162 13707
rect 2186 13733 2214 13734
rect 2238 13733 2266 13734
rect 2186 13707 2198 13733
rect 2198 13707 2214 13733
rect 2238 13707 2260 13733
rect 2260 13707 2266 13733
rect 2186 13706 2214 13707
rect 2238 13706 2266 13707
rect 2290 13706 2318 13734
rect 2342 13733 2370 13734
rect 2394 13733 2422 13734
rect 2342 13707 2348 13733
rect 2348 13707 2370 13733
rect 2394 13707 2410 13733
rect 2410 13707 2422 13733
rect 2342 13706 2370 13707
rect 2394 13706 2422 13707
rect 2446 13733 2474 13734
rect 2446 13707 2472 13733
rect 2472 13707 2474 13733
rect 2446 13706 2474 13707
rect 2498 13733 2526 13734
rect 2498 13707 2508 13733
rect 2508 13707 2526 13733
rect 2498 13706 2526 13707
rect 2758 14294 2786 14322
rect 3318 14294 3346 14322
rect 3822 15105 3850 15106
rect 3822 15079 3823 15105
rect 3823 15079 3849 15105
rect 3849 15079 3850 15105
rect 3822 15078 3850 15079
rect 5558 15105 5586 15106
rect 5558 15079 5559 15105
rect 5559 15079 5585 15105
rect 5585 15079 5586 15105
rect 5558 15078 5586 15079
rect 4582 14909 4610 14910
rect 4582 14883 4600 14909
rect 4600 14883 4610 14909
rect 4582 14882 4610 14883
rect 4634 14909 4662 14910
rect 4634 14883 4636 14909
rect 4636 14883 4662 14909
rect 4634 14882 4662 14883
rect 4686 14909 4714 14910
rect 4738 14909 4766 14910
rect 4686 14883 4698 14909
rect 4698 14883 4714 14909
rect 4738 14883 4760 14909
rect 4760 14883 4766 14909
rect 4686 14882 4714 14883
rect 4738 14882 4766 14883
rect 4790 14882 4818 14910
rect 4842 14909 4870 14910
rect 4894 14909 4922 14910
rect 4842 14883 4848 14909
rect 4848 14883 4870 14909
rect 4894 14883 4910 14909
rect 4910 14883 4922 14909
rect 4842 14882 4870 14883
rect 4894 14882 4922 14883
rect 4946 14909 4974 14910
rect 4946 14883 4972 14909
rect 4972 14883 4974 14909
rect 4946 14882 4974 14883
rect 4998 14909 5026 14910
rect 4998 14883 5008 14909
rect 5008 14883 5026 14909
rect 4998 14882 5026 14883
rect 3822 14321 3850 14322
rect 3822 14295 3823 14321
rect 3823 14295 3849 14321
rect 3849 14295 3850 14321
rect 3822 14294 3850 14295
rect 5558 14686 5586 14714
rect 4582 14125 4610 14126
rect 4582 14099 4600 14125
rect 4600 14099 4610 14125
rect 4582 14098 4610 14099
rect 4634 14125 4662 14126
rect 4634 14099 4636 14125
rect 4636 14099 4662 14125
rect 4634 14098 4662 14099
rect 4686 14125 4714 14126
rect 4738 14125 4766 14126
rect 4686 14099 4698 14125
rect 4698 14099 4714 14125
rect 4738 14099 4760 14125
rect 4760 14099 4766 14125
rect 4686 14098 4714 14099
rect 4738 14098 4766 14099
rect 4790 14098 4818 14126
rect 4842 14125 4870 14126
rect 4894 14125 4922 14126
rect 4842 14099 4848 14125
rect 4848 14099 4870 14125
rect 4894 14099 4910 14125
rect 4910 14099 4922 14125
rect 4842 14098 4870 14099
rect 4894 14098 4922 14099
rect 4946 14125 4974 14126
rect 4946 14099 4972 14125
rect 4972 14099 4974 14125
rect 4946 14098 4974 14099
rect 4998 14125 5026 14126
rect 4998 14099 5008 14125
rect 5008 14099 5026 14125
rect 4998 14098 5026 14099
rect 1974 13118 2002 13146
rect 2366 13145 2394 13146
rect 2366 13119 2367 13145
rect 2367 13119 2393 13145
rect 2393 13119 2394 13145
rect 2366 13118 2394 13119
rect 2082 12949 2110 12950
rect 2082 12923 2100 12949
rect 2100 12923 2110 12949
rect 2082 12922 2110 12923
rect 2134 12949 2162 12950
rect 2134 12923 2136 12949
rect 2136 12923 2162 12949
rect 2134 12922 2162 12923
rect 2186 12949 2214 12950
rect 2238 12949 2266 12950
rect 2186 12923 2198 12949
rect 2198 12923 2214 12949
rect 2238 12923 2260 12949
rect 2260 12923 2266 12949
rect 2186 12922 2214 12923
rect 2238 12922 2266 12923
rect 2290 12922 2318 12950
rect 2342 12949 2370 12950
rect 2394 12949 2422 12950
rect 2342 12923 2348 12949
rect 2348 12923 2370 12949
rect 2394 12923 2410 12949
rect 2410 12923 2422 12949
rect 2342 12922 2370 12923
rect 2394 12922 2422 12923
rect 2446 12949 2474 12950
rect 2446 12923 2472 12949
rect 2472 12923 2474 12949
rect 2446 12922 2474 12923
rect 2498 12949 2526 12950
rect 2498 12923 2508 12949
rect 2508 12923 2526 12949
rect 2498 12922 2526 12923
rect 2478 12753 2506 12754
rect 2478 12727 2479 12753
rect 2479 12727 2505 12753
rect 2505 12727 2506 12753
rect 2478 12726 2506 12727
rect 1750 8833 1778 8834
rect 1750 8807 1751 8833
rect 1751 8807 1777 8833
rect 1777 8807 1778 8833
rect 1750 8806 1778 8807
rect 2082 12165 2110 12166
rect 2082 12139 2100 12165
rect 2100 12139 2110 12165
rect 2082 12138 2110 12139
rect 2134 12165 2162 12166
rect 2134 12139 2136 12165
rect 2136 12139 2162 12165
rect 2134 12138 2162 12139
rect 2186 12165 2214 12166
rect 2238 12165 2266 12166
rect 2186 12139 2198 12165
rect 2198 12139 2214 12165
rect 2238 12139 2260 12165
rect 2260 12139 2266 12165
rect 2186 12138 2214 12139
rect 2238 12138 2266 12139
rect 2290 12138 2318 12166
rect 2342 12165 2370 12166
rect 2394 12165 2422 12166
rect 2342 12139 2348 12165
rect 2348 12139 2370 12165
rect 2394 12139 2410 12165
rect 2410 12139 2422 12165
rect 2342 12138 2370 12139
rect 2394 12138 2422 12139
rect 2446 12165 2474 12166
rect 2446 12139 2472 12165
rect 2472 12139 2474 12165
rect 2446 12138 2474 12139
rect 2498 12165 2526 12166
rect 2498 12139 2508 12165
rect 2508 12139 2526 12165
rect 2498 12138 2526 12139
rect 2758 12726 2786 12754
rect 2082 11381 2110 11382
rect 2082 11355 2100 11381
rect 2100 11355 2110 11381
rect 2082 11354 2110 11355
rect 2134 11381 2162 11382
rect 2134 11355 2136 11381
rect 2136 11355 2162 11381
rect 2134 11354 2162 11355
rect 2186 11381 2214 11382
rect 2238 11381 2266 11382
rect 2186 11355 2198 11381
rect 2198 11355 2214 11381
rect 2238 11355 2260 11381
rect 2260 11355 2266 11381
rect 2186 11354 2214 11355
rect 2238 11354 2266 11355
rect 2290 11354 2318 11382
rect 2342 11381 2370 11382
rect 2394 11381 2422 11382
rect 2342 11355 2348 11381
rect 2348 11355 2370 11381
rect 2394 11355 2410 11381
rect 2410 11355 2422 11381
rect 2342 11354 2370 11355
rect 2394 11354 2422 11355
rect 2446 11381 2474 11382
rect 2446 11355 2472 11381
rect 2472 11355 2474 11381
rect 2446 11354 2474 11355
rect 2498 11381 2526 11382
rect 2498 11355 2508 11381
rect 2508 11355 2526 11381
rect 2498 11354 2526 11355
rect 2082 10597 2110 10598
rect 2082 10571 2100 10597
rect 2100 10571 2110 10597
rect 2082 10570 2110 10571
rect 2134 10597 2162 10598
rect 2134 10571 2136 10597
rect 2136 10571 2162 10597
rect 2134 10570 2162 10571
rect 2186 10597 2214 10598
rect 2238 10597 2266 10598
rect 2186 10571 2198 10597
rect 2198 10571 2214 10597
rect 2238 10571 2260 10597
rect 2260 10571 2266 10597
rect 2186 10570 2214 10571
rect 2238 10570 2266 10571
rect 2290 10570 2318 10598
rect 2342 10597 2370 10598
rect 2394 10597 2422 10598
rect 2342 10571 2348 10597
rect 2348 10571 2370 10597
rect 2394 10571 2410 10597
rect 2410 10571 2422 10597
rect 2342 10570 2370 10571
rect 2394 10570 2422 10571
rect 2446 10597 2474 10598
rect 2446 10571 2472 10597
rect 2472 10571 2474 10597
rect 2446 10570 2474 10571
rect 2498 10597 2526 10598
rect 2498 10571 2508 10597
rect 2508 10571 2526 10597
rect 2498 10570 2526 10571
rect 2082 9813 2110 9814
rect 2082 9787 2100 9813
rect 2100 9787 2110 9813
rect 2082 9786 2110 9787
rect 2134 9813 2162 9814
rect 2134 9787 2136 9813
rect 2136 9787 2162 9813
rect 2134 9786 2162 9787
rect 2186 9813 2214 9814
rect 2238 9813 2266 9814
rect 2186 9787 2198 9813
rect 2198 9787 2214 9813
rect 2238 9787 2260 9813
rect 2260 9787 2266 9813
rect 2186 9786 2214 9787
rect 2238 9786 2266 9787
rect 2290 9786 2318 9814
rect 2342 9813 2370 9814
rect 2394 9813 2422 9814
rect 2342 9787 2348 9813
rect 2348 9787 2370 9813
rect 2394 9787 2410 9813
rect 2410 9787 2422 9813
rect 2342 9786 2370 9787
rect 2394 9786 2422 9787
rect 2446 9813 2474 9814
rect 2446 9787 2472 9813
rect 2472 9787 2474 9813
rect 2446 9786 2474 9787
rect 2498 9813 2526 9814
rect 2498 9787 2508 9813
rect 2508 9787 2526 9813
rect 2498 9786 2526 9787
rect 1918 9225 1946 9226
rect 1918 9199 1919 9225
rect 1919 9199 1945 9225
rect 1945 9199 1946 9225
rect 1918 9198 1946 9199
rect 2478 9198 2506 9226
rect 3038 9225 3066 9226
rect 3038 9199 3039 9225
rect 3039 9199 3065 9225
rect 3065 9199 3066 9225
rect 3038 9198 3066 9199
rect 2082 9029 2110 9030
rect 2082 9003 2100 9029
rect 2100 9003 2110 9029
rect 2082 9002 2110 9003
rect 2134 9029 2162 9030
rect 2134 9003 2136 9029
rect 2136 9003 2162 9029
rect 2134 9002 2162 9003
rect 2186 9029 2214 9030
rect 2238 9029 2266 9030
rect 2186 9003 2198 9029
rect 2198 9003 2214 9029
rect 2238 9003 2260 9029
rect 2260 9003 2266 9029
rect 2186 9002 2214 9003
rect 2238 9002 2266 9003
rect 2290 9002 2318 9030
rect 2342 9029 2370 9030
rect 2394 9029 2422 9030
rect 2342 9003 2348 9029
rect 2348 9003 2370 9029
rect 2394 9003 2410 9029
rect 2410 9003 2422 9029
rect 2342 9002 2370 9003
rect 2394 9002 2422 9003
rect 2446 9029 2474 9030
rect 2446 9003 2472 9029
rect 2472 9003 2474 9029
rect 2446 9002 2474 9003
rect 2498 9029 2526 9030
rect 2498 9003 2508 9029
rect 2508 9003 2526 9029
rect 2498 9002 2526 9003
rect 1918 8414 1946 8442
rect 1974 8833 2002 8834
rect 1974 8807 1975 8833
rect 1975 8807 2001 8833
rect 2001 8807 2002 8833
rect 1974 8806 2002 8807
rect 1022 7966 1050 7994
rect 2310 8806 2338 8834
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 2534 8470 2562 8498
rect 2082 8245 2110 8246
rect 2082 8219 2100 8245
rect 2100 8219 2110 8245
rect 2082 8218 2110 8219
rect 2134 8245 2162 8246
rect 2134 8219 2136 8245
rect 2136 8219 2162 8245
rect 2134 8218 2162 8219
rect 2186 8245 2214 8246
rect 2238 8245 2266 8246
rect 2186 8219 2198 8245
rect 2198 8219 2214 8245
rect 2238 8219 2260 8245
rect 2260 8219 2266 8245
rect 2186 8218 2214 8219
rect 2238 8218 2266 8219
rect 2290 8218 2318 8246
rect 2342 8245 2370 8246
rect 2394 8245 2422 8246
rect 2342 8219 2348 8245
rect 2348 8219 2370 8245
rect 2394 8219 2410 8245
rect 2410 8219 2422 8245
rect 2342 8218 2370 8219
rect 2394 8218 2422 8219
rect 2446 8245 2474 8246
rect 2446 8219 2472 8245
rect 2472 8219 2474 8245
rect 2446 8218 2474 8219
rect 2498 8245 2526 8246
rect 2498 8219 2508 8245
rect 2508 8219 2526 8245
rect 2498 8218 2526 8219
rect 2926 8078 2954 8106
rect 1806 7265 1834 7266
rect 1806 7239 1807 7265
rect 1807 7239 1833 7265
rect 1833 7239 1834 7265
rect 1806 7238 1834 7239
rect 2590 7630 2618 7658
rect 2082 7461 2110 7462
rect 2082 7435 2100 7461
rect 2100 7435 2110 7461
rect 2082 7434 2110 7435
rect 2134 7461 2162 7462
rect 2134 7435 2136 7461
rect 2136 7435 2162 7461
rect 2134 7434 2162 7435
rect 2186 7461 2214 7462
rect 2238 7461 2266 7462
rect 2186 7435 2198 7461
rect 2198 7435 2214 7461
rect 2238 7435 2260 7461
rect 2260 7435 2266 7461
rect 2186 7434 2214 7435
rect 2238 7434 2266 7435
rect 2290 7434 2318 7462
rect 2342 7461 2370 7462
rect 2394 7461 2422 7462
rect 2342 7435 2348 7461
rect 2348 7435 2370 7461
rect 2394 7435 2410 7461
rect 2410 7435 2422 7461
rect 2342 7434 2370 7435
rect 2394 7434 2422 7435
rect 2446 7461 2474 7462
rect 2446 7435 2472 7461
rect 2472 7435 2474 7461
rect 2446 7434 2474 7435
rect 2498 7461 2526 7462
rect 2498 7435 2508 7461
rect 2508 7435 2526 7461
rect 2498 7434 2526 7435
rect 2030 7265 2058 7266
rect 2030 7239 2031 7265
rect 2031 7239 2057 7265
rect 2057 7239 2058 7265
rect 2030 7238 2058 7239
rect 2366 7238 2394 7266
rect 2082 6677 2110 6678
rect 2082 6651 2100 6677
rect 2100 6651 2110 6677
rect 2082 6650 2110 6651
rect 2134 6677 2162 6678
rect 2134 6651 2136 6677
rect 2136 6651 2162 6677
rect 2134 6650 2162 6651
rect 2186 6677 2214 6678
rect 2238 6677 2266 6678
rect 2186 6651 2198 6677
rect 2198 6651 2214 6677
rect 2238 6651 2260 6677
rect 2260 6651 2266 6677
rect 2186 6650 2214 6651
rect 2238 6650 2266 6651
rect 2290 6650 2318 6678
rect 2342 6677 2370 6678
rect 2394 6677 2422 6678
rect 2342 6651 2348 6677
rect 2348 6651 2370 6677
rect 2394 6651 2410 6677
rect 2410 6651 2422 6677
rect 2342 6650 2370 6651
rect 2394 6650 2422 6651
rect 2446 6677 2474 6678
rect 2446 6651 2472 6677
rect 2472 6651 2474 6677
rect 2446 6650 2474 6651
rect 2498 6677 2526 6678
rect 2498 6651 2508 6677
rect 2508 6651 2526 6677
rect 2498 6650 2526 6651
rect 2590 6062 2618 6090
rect 2082 5893 2110 5894
rect 2082 5867 2100 5893
rect 2100 5867 2110 5893
rect 2082 5866 2110 5867
rect 2134 5893 2162 5894
rect 2134 5867 2136 5893
rect 2136 5867 2162 5893
rect 2134 5866 2162 5867
rect 2186 5893 2214 5894
rect 2238 5893 2266 5894
rect 2186 5867 2198 5893
rect 2198 5867 2214 5893
rect 2238 5867 2260 5893
rect 2260 5867 2266 5893
rect 2186 5866 2214 5867
rect 2238 5866 2266 5867
rect 2290 5866 2318 5894
rect 2342 5893 2370 5894
rect 2394 5893 2422 5894
rect 2342 5867 2348 5893
rect 2348 5867 2370 5893
rect 2394 5867 2410 5893
rect 2410 5867 2422 5893
rect 2342 5866 2370 5867
rect 2394 5866 2422 5867
rect 2446 5893 2474 5894
rect 2446 5867 2472 5893
rect 2472 5867 2474 5893
rect 2446 5866 2474 5867
rect 2498 5893 2526 5894
rect 2498 5867 2508 5893
rect 2508 5867 2526 5893
rect 2498 5866 2526 5867
rect 2082 5109 2110 5110
rect 2082 5083 2100 5109
rect 2100 5083 2110 5109
rect 2082 5082 2110 5083
rect 2134 5109 2162 5110
rect 2134 5083 2136 5109
rect 2136 5083 2162 5109
rect 2134 5082 2162 5083
rect 2186 5109 2214 5110
rect 2238 5109 2266 5110
rect 2186 5083 2198 5109
rect 2198 5083 2214 5109
rect 2238 5083 2260 5109
rect 2260 5083 2266 5109
rect 2186 5082 2214 5083
rect 2238 5082 2266 5083
rect 2290 5082 2318 5110
rect 2342 5109 2370 5110
rect 2394 5109 2422 5110
rect 2342 5083 2348 5109
rect 2348 5083 2370 5109
rect 2394 5083 2410 5109
rect 2410 5083 2422 5109
rect 2342 5082 2370 5083
rect 2394 5082 2422 5083
rect 2446 5109 2474 5110
rect 2446 5083 2472 5109
rect 2472 5083 2474 5109
rect 2446 5082 2474 5083
rect 2498 5109 2526 5110
rect 2498 5083 2508 5109
rect 2508 5083 2526 5109
rect 2498 5082 2526 5083
rect 2082 4325 2110 4326
rect 2082 4299 2100 4325
rect 2100 4299 2110 4325
rect 2082 4298 2110 4299
rect 2134 4325 2162 4326
rect 2134 4299 2136 4325
rect 2136 4299 2162 4325
rect 2134 4298 2162 4299
rect 2186 4325 2214 4326
rect 2238 4325 2266 4326
rect 2186 4299 2198 4325
rect 2198 4299 2214 4325
rect 2238 4299 2260 4325
rect 2260 4299 2266 4325
rect 2186 4298 2214 4299
rect 2238 4298 2266 4299
rect 2290 4298 2318 4326
rect 2342 4325 2370 4326
rect 2394 4325 2422 4326
rect 2342 4299 2348 4325
rect 2348 4299 2370 4325
rect 2394 4299 2410 4325
rect 2410 4299 2422 4325
rect 2342 4298 2370 4299
rect 2394 4298 2422 4299
rect 2446 4325 2474 4326
rect 2446 4299 2472 4325
rect 2472 4299 2474 4325
rect 2446 4298 2474 4299
rect 2498 4325 2526 4326
rect 2498 4299 2508 4325
rect 2508 4299 2526 4325
rect 2498 4298 2526 4299
rect 2590 4158 2618 4186
rect 2082 3541 2110 3542
rect 2082 3515 2100 3541
rect 2100 3515 2110 3541
rect 2082 3514 2110 3515
rect 2134 3541 2162 3542
rect 2134 3515 2136 3541
rect 2136 3515 2162 3541
rect 2134 3514 2162 3515
rect 2186 3541 2214 3542
rect 2238 3541 2266 3542
rect 2186 3515 2198 3541
rect 2198 3515 2214 3541
rect 2238 3515 2260 3541
rect 2260 3515 2266 3541
rect 2186 3514 2214 3515
rect 2238 3514 2266 3515
rect 2290 3514 2318 3542
rect 2342 3541 2370 3542
rect 2394 3541 2422 3542
rect 2342 3515 2348 3541
rect 2348 3515 2370 3541
rect 2394 3515 2410 3541
rect 2410 3515 2422 3541
rect 2342 3514 2370 3515
rect 2394 3514 2422 3515
rect 2446 3541 2474 3542
rect 2446 3515 2472 3541
rect 2472 3515 2474 3541
rect 2446 3514 2474 3515
rect 2498 3541 2526 3542
rect 2498 3515 2508 3541
rect 2508 3515 2526 3541
rect 2498 3514 2526 3515
rect 2478 3345 2506 3346
rect 2478 3319 2479 3345
rect 2479 3319 2505 3345
rect 2505 3319 2506 3345
rect 2478 3318 2506 3319
rect 2082 2757 2110 2758
rect 2082 2731 2100 2757
rect 2100 2731 2110 2757
rect 2082 2730 2110 2731
rect 2134 2757 2162 2758
rect 2134 2731 2136 2757
rect 2136 2731 2162 2757
rect 2134 2730 2162 2731
rect 2186 2757 2214 2758
rect 2238 2757 2266 2758
rect 2186 2731 2198 2757
rect 2198 2731 2214 2757
rect 2238 2731 2260 2757
rect 2260 2731 2266 2757
rect 2186 2730 2214 2731
rect 2238 2730 2266 2731
rect 2290 2730 2318 2758
rect 2342 2757 2370 2758
rect 2394 2757 2422 2758
rect 2342 2731 2348 2757
rect 2348 2731 2370 2757
rect 2394 2731 2410 2757
rect 2410 2731 2422 2757
rect 2342 2730 2370 2731
rect 2394 2730 2422 2731
rect 2446 2757 2474 2758
rect 2446 2731 2472 2757
rect 2472 2731 2474 2757
rect 2446 2730 2474 2731
rect 2498 2757 2526 2758
rect 2498 2731 2508 2757
rect 2508 2731 2526 2757
rect 2498 2730 2526 2731
rect 1638 2478 1666 2506
rect 2478 2561 2506 2562
rect 2478 2535 2479 2561
rect 2479 2535 2505 2561
rect 2505 2535 2506 2561
rect 2478 2534 2506 2535
rect 2030 2198 2058 2226
rect 2478 2198 2506 2226
rect 2082 1973 2110 1974
rect 2082 1947 2100 1973
rect 2100 1947 2110 1973
rect 2082 1946 2110 1947
rect 2134 1973 2162 1974
rect 2134 1947 2136 1973
rect 2136 1947 2162 1973
rect 2134 1946 2162 1947
rect 2186 1973 2214 1974
rect 2238 1973 2266 1974
rect 2186 1947 2198 1973
rect 2198 1947 2214 1973
rect 2238 1947 2260 1973
rect 2260 1947 2266 1973
rect 2186 1946 2214 1947
rect 2238 1946 2266 1947
rect 2290 1946 2318 1974
rect 2342 1973 2370 1974
rect 2394 1973 2422 1974
rect 2342 1947 2348 1973
rect 2348 1947 2370 1973
rect 2394 1947 2410 1973
rect 2410 1947 2422 1973
rect 2342 1946 2370 1947
rect 2394 1946 2422 1947
rect 2446 1973 2474 1974
rect 2446 1947 2472 1973
rect 2472 1947 2474 1973
rect 2446 1946 2474 1947
rect 2498 1973 2526 1974
rect 2498 1947 2508 1973
rect 2508 1947 2526 1973
rect 2498 1946 2526 1947
rect 2478 1638 2506 1666
rect 3038 7657 3066 7658
rect 3038 7631 3039 7657
rect 3039 7631 3065 7657
rect 3065 7631 3066 7657
rect 3038 7630 3066 7631
rect 4582 13341 4610 13342
rect 4582 13315 4600 13341
rect 4600 13315 4610 13341
rect 4582 13314 4610 13315
rect 4634 13341 4662 13342
rect 4634 13315 4636 13341
rect 4636 13315 4662 13341
rect 4634 13314 4662 13315
rect 4686 13341 4714 13342
rect 4738 13341 4766 13342
rect 4686 13315 4698 13341
rect 4698 13315 4714 13341
rect 4738 13315 4760 13341
rect 4760 13315 4766 13341
rect 4686 13314 4714 13315
rect 4738 13314 4766 13315
rect 4790 13314 4818 13342
rect 4842 13341 4870 13342
rect 4894 13341 4922 13342
rect 4842 13315 4848 13341
rect 4848 13315 4870 13341
rect 4894 13315 4910 13341
rect 4910 13315 4922 13341
rect 4842 13314 4870 13315
rect 4894 13314 4922 13315
rect 4946 13341 4974 13342
rect 4946 13315 4972 13341
rect 4972 13315 4974 13341
rect 4946 13314 4974 13315
rect 4998 13341 5026 13342
rect 4998 13315 5008 13341
rect 5008 13315 5026 13341
rect 4998 13314 5026 13315
rect 6118 15078 6146 15106
rect 6118 14798 6146 14826
rect 6118 14713 6146 14714
rect 6118 14687 6119 14713
rect 6119 14687 6145 14713
rect 6145 14687 6146 14713
rect 6118 14686 6146 14687
rect 5894 13510 5922 13538
rect 5558 12753 5586 12754
rect 5558 12727 5559 12753
rect 5559 12727 5585 12753
rect 5585 12727 5586 12753
rect 5558 12726 5586 12727
rect 4582 12557 4610 12558
rect 4582 12531 4600 12557
rect 4600 12531 4610 12557
rect 4582 12530 4610 12531
rect 4634 12557 4662 12558
rect 4634 12531 4636 12557
rect 4636 12531 4662 12557
rect 4634 12530 4662 12531
rect 4686 12557 4714 12558
rect 4738 12557 4766 12558
rect 4686 12531 4698 12557
rect 4698 12531 4714 12557
rect 4738 12531 4760 12557
rect 4760 12531 4766 12557
rect 4686 12530 4714 12531
rect 4738 12530 4766 12531
rect 4790 12530 4818 12558
rect 4842 12557 4870 12558
rect 4894 12557 4922 12558
rect 4842 12531 4848 12557
rect 4848 12531 4870 12557
rect 4894 12531 4910 12557
rect 4910 12531 4922 12557
rect 4842 12530 4870 12531
rect 4894 12530 4922 12531
rect 4946 12557 4974 12558
rect 4946 12531 4972 12557
rect 4972 12531 4974 12557
rect 4946 12530 4974 12531
rect 4998 12557 5026 12558
rect 4998 12531 5008 12557
rect 5008 12531 5026 12557
rect 4998 12530 5026 12531
rect 6118 12726 6146 12754
rect 6118 12361 6146 12362
rect 6118 12335 6119 12361
rect 6119 12335 6145 12361
rect 6145 12335 6146 12361
rect 6118 12334 6146 12335
rect 6454 13537 6482 13538
rect 6454 13511 6455 13537
rect 6455 13511 6481 13537
rect 6481 13511 6482 13537
rect 6454 13510 6482 13511
rect 6454 12697 6482 12698
rect 6454 12671 6455 12697
rect 6455 12671 6481 12697
rect 6481 12671 6482 12697
rect 6454 12670 6482 12671
rect 4582 11773 4610 11774
rect 4582 11747 4600 11773
rect 4600 11747 4610 11773
rect 4582 11746 4610 11747
rect 4634 11773 4662 11774
rect 4634 11747 4636 11773
rect 4636 11747 4662 11773
rect 4634 11746 4662 11747
rect 4686 11773 4714 11774
rect 4738 11773 4766 11774
rect 4686 11747 4698 11773
rect 4698 11747 4714 11773
rect 4738 11747 4760 11773
rect 4760 11747 4766 11773
rect 4686 11746 4714 11747
rect 4738 11746 4766 11747
rect 4790 11746 4818 11774
rect 4842 11773 4870 11774
rect 4894 11773 4922 11774
rect 4842 11747 4848 11773
rect 4848 11747 4870 11773
rect 4894 11747 4910 11773
rect 4910 11747 4922 11773
rect 4842 11746 4870 11747
rect 4894 11746 4922 11747
rect 4946 11773 4974 11774
rect 4946 11747 4972 11773
rect 4972 11747 4974 11773
rect 4946 11746 4974 11747
rect 4998 11773 5026 11774
rect 4998 11747 5008 11773
rect 5008 11747 5026 11773
rect 4998 11746 5026 11747
rect 4582 10989 4610 10990
rect 4582 10963 4600 10989
rect 4600 10963 4610 10989
rect 4582 10962 4610 10963
rect 4634 10989 4662 10990
rect 4634 10963 4636 10989
rect 4636 10963 4662 10989
rect 4634 10962 4662 10963
rect 4686 10989 4714 10990
rect 4738 10989 4766 10990
rect 4686 10963 4698 10989
rect 4698 10963 4714 10989
rect 4738 10963 4760 10989
rect 4760 10963 4766 10989
rect 4686 10962 4714 10963
rect 4738 10962 4766 10963
rect 4790 10962 4818 10990
rect 4842 10989 4870 10990
rect 4894 10989 4922 10990
rect 4842 10963 4848 10989
rect 4848 10963 4870 10989
rect 4894 10963 4910 10989
rect 4910 10963 4922 10989
rect 4842 10962 4870 10963
rect 4894 10962 4922 10963
rect 4946 10989 4974 10990
rect 4946 10963 4972 10989
rect 4972 10963 4974 10989
rect 4946 10962 4974 10963
rect 4998 10989 5026 10990
rect 4998 10963 5008 10989
rect 5008 10963 5026 10989
rect 4998 10962 5026 10963
rect 4582 10205 4610 10206
rect 4582 10179 4600 10205
rect 4600 10179 4610 10205
rect 4582 10178 4610 10179
rect 4634 10205 4662 10206
rect 4634 10179 4636 10205
rect 4636 10179 4662 10205
rect 4634 10178 4662 10179
rect 4686 10205 4714 10206
rect 4738 10205 4766 10206
rect 4686 10179 4698 10205
rect 4698 10179 4714 10205
rect 4738 10179 4760 10205
rect 4760 10179 4766 10205
rect 4686 10178 4714 10179
rect 4738 10178 4766 10179
rect 4790 10178 4818 10206
rect 4842 10205 4870 10206
rect 4894 10205 4922 10206
rect 4842 10179 4848 10205
rect 4848 10179 4870 10205
rect 4894 10179 4910 10205
rect 4910 10179 4922 10205
rect 4842 10178 4870 10179
rect 4894 10178 4922 10179
rect 4946 10205 4974 10206
rect 4946 10179 4972 10205
rect 4972 10179 4974 10205
rect 4946 10178 4974 10179
rect 4998 10205 5026 10206
rect 4998 10179 5008 10205
rect 5008 10179 5026 10205
rect 4998 10178 5026 10179
rect 3598 8441 3626 8442
rect 3598 8415 3599 8441
rect 3599 8415 3625 8441
rect 3625 8415 3626 8441
rect 3598 8414 3626 8415
rect 3598 6790 3626 6818
rect 3710 8862 3738 8890
rect 3038 6089 3066 6090
rect 3038 6063 3039 6089
rect 3039 6063 3065 6089
rect 3065 6063 3066 6089
rect 3038 6062 3066 6063
rect 3598 6089 3626 6090
rect 3598 6063 3599 6089
rect 3599 6063 3625 6089
rect 3625 6063 3626 6089
rect 3598 6062 3626 6063
rect 3038 4158 3066 4186
rect 3542 4214 3570 4242
rect 3038 3318 3066 3346
rect 3038 2534 3066 2562
rect 3038 2169 3066 2170
rect 3038 2143 3039 2169
rect 3039 2143 3065 2169
rect 3065 2143 3066 2169
rect 3038 2142 3066 2143
rect 3486 2169 3514 2170
rect 3486 2143 3487 2169
rect 3487 2143 3513 2169
rect 3513 2143 3514 2169
rect 3486 2142 3514 2143
rect 3486 1806 3514 1834
rect 2926 1694 2954 1722
rect 2534 1470 2562 1498
rect 4998 9561 5026 9562
rect 4998 9535 4999 9561
rect 4999 9535 5025 9561
rect 5025 9535 5026 9561
rect 4998 9534 5026 9535
rect 4582 9421 4610 9422
rect 4582 9395 4600 9421
rect 4600 9395 4610 9421
rect 4582 9394 4610 9395
rect 4634 9421 4662 9422
rect 4634 9395 4636 9421
rect 4636 9395 4662 9421
rect 4634 9394 4662 9395
rect 4686 9421 4714 9422
rect 4738 9421 4766 9422
rect 4686 9395 4698 9421
rect 4698 9395 4714 9421
rect 4738 9395 4760 9421
rect 4760 9395 4766 9421
rect 4686 9394 4714 9395
rect 4738 9394 4766 9395
rect 4790 9394 4818 9422
rect 4842 9421 4870 9422
rect 4894 9421 4922 9422
rect 4842 9395 4848 9421
rect 4848 9395 4870 9421
rect 4894 9395 4910 9421
rect 4910 9395 4922 9421
rect 4842 9394 4870 9395
rect 4894 9394 4922 9395
rect 4946 9421 4974 9422
rect 4946 9395 4972 9421
rect 4972 9395 4974 9421
rect 4946 9394 4974 9395
rect 4998 9421 5026 9422
rect 4998 9395 5008 9421
rect 5008 9395 5026 9421
rect 4998 9394 5026 9395
rect 4494 9198 4522 9226
rect 4494 8833 4522 8834
rect 4494 8807 4495 8833
rect 4495 8807 4521 8833
rect 4521 8807 4522 8833
rect 4494 8806 4522 8807
rect 4582 8637 4610 8638
rect 4582 8611 4600 8637
rect 4600 8611 4610 8637
rect 4582 8610 4610 8611
rect 4634 8637 4662 8638
rect 4634 8611 4636 8637
rect 4636 8611 4662 8637
rect 4634 8610 4662 8611
rect 4686 8637 4714 8638
rect 4738 8637 4766 8638
rect 4686 8611 4698 8637
rect 4698 8611 4714 8637
rect 4738 8611 4760 8637
rect 4760 8611 4766 8637
rect 4686 8610 4714 8611
rect 4738 8610 4766 8611
rect 4790 8610 4818 8638
rect 4842 8637 4870 8638
rect 4894 8637 4922 8638
rect 4842 8611 4848 8637
rect 4848 8611 4870 8637
rect 4894 8611 4910 8637
rect 4910 8611 4922 8637
rect 4842 8610 4870 8611
rect 4894 8610 4922 8611
rect 4946 8637 4974 8638
rect 4946 8611 4972 8637
rect 4972 8611 4974 8637
rect 4946 8610 4974 8611
rect 4998 8637 5026 8638
rect 4998 8611 5008 8637
rect 5008 8611 5026 8637
rect 4998 8610 5026 8611
rect 4214 8470 4242 8498
rect 4582 7853 4610 7854
rect 4582 7827 4600 7853
rect 4600 7827 4610 7853
rect 4582 7826 4610 7827
rect 4634 7853 4662 7854
rect 4634 7827 4636 7853
rect 4636 7827 4662 7853
rect 4634 7826 4662 7827
rect 4686 7853 4714 7854
rect 4738 7853 4766 7854
rect 4686 7827 4698 7853
rect 4698 7827 4714 7853
rect 4738 7827 4760 7853
rect 4760 7827 4766 7853
rect 4686 7826 4714 7827
rect 4738 7826 4766 7827
rect 4790 7826 4818 7854
rect 4842 7853 4870 7854
rect 4894 7853 4922 7854
rect 4842 7827 4848 7853
rect 4848 7827 4870 7853
rect 4894 7827 4910 7853
rect 4910 7827 4922 7853
rect 4842 7826 4870 7827
rect 4894 7826 4922 7827
rect 4946 7853 4974 7854
rect 4946 7827 4972 7853
rect 4972 7827 4974 7853
rect 4946 7826 4974 7827
rect 4998 7853 5026 7854
rect 4998 7827 5008 7853
rect 5008 7827 5026 7853
rect 4998 7826 5026 7827
rect 5894 9926 5922 9954
rect 6454 9561 6482 9562
rect 6454 9535 6455 9561
rect 6455 9535 6481 9561
rect 6481 9535 6482 9561
rect 6454 9534 6482 9535
rect 5950 8833 5978 8834
rect 5950 8807 5951 8833
rect 5951 8807 5977 8833
rect 5977 8807 5978 8833
rect 5950 8806 5978 8807
rect 6230 8806 6258 8834
rect 7082 18437 7110 18438
rect 7082 18411 7100 18437
rect 7100 18411 7110 18437
rect 7082 18410 7110 18411
rect 7134 18437 7162 18438
rect 7134 18411 7136 18437
rect 7136 18411 7162 18437
rect 7134 18410 7162 18411
rect 7186 18437 7214 18438
rect 7238 18437 7266 18438
rect 7186 18411 7198 18437
rect 7198 18411 7214 18437
rect 7238 18411 7260 18437
rect 7260 18411 7266 18437
rect 7186 18410 7214 18411
rect 7238 18410 7266 18411
rect 7290 18410 7318 18438
rect 7342 18437 7370 18438
rect 7394 18437 7422 18438
rect 7342 18411 7348 18437
rect 7348 18411 7370 18437
rect 7394 18411 7410 18437
rect 7410 18411 7422 18437
rect 7342 18410 7370 18411
rect 7394 18410 7422 18411
rect 7446 18437 7474 18438
rect 7446 18411 7472 18437
rect 7472 18411 7474 18437
rect 7446 18410 7474 18411
rect 7498 18437 7526 18438
rect 7498 18411 7508 18437
rect 7508 18411 7526 18437
rect 7498 18410 7526 18411
rect 12082 18437 12110 18438
rect 12082 18411 12100 18437
rect 12100 18411 12110 18437
rect 12082 18410 12110 18411
rect 12134 18437 12162 18438
rect 12134 18411 12136 18437
rect 12136 18411 12162 18437
rect 12134 18410 12162 18411
rect 12186 18437 12214 18438
rect 12238 18437 12266 18438
rect 12186 18411 12198 18437
rect 12198 18411 12214 18437
rect 12238 18411 12260 18437
rect 12260 18411 12266 18437
rect 12186 18410 12214 18411
rect 12238 18410 12266 18411
rect 12290 18410 12318 18438
rect 12342 18437 12370 18438
rect 12394 18437 12422 18438
rect 12342 18411 12348 18437
rect 12348 18411 12370 18437
rect 12394 18411 12410 18437
rect 12410 18411 12422 18437
rect 12342 18410 12370 18411
rect 12394 18410 12422 18411
rect 12446 18437 12474 18438
rect 12446 18411 12472 18437
rect 12472 18411 12474 18437
rect 12446 18410 12474 18411
rect 12498 18437 12526 18438
rect 12498 18411 12508 18437
rect 12508 18411 12526 18437
rect 12498 18410 12526 18411
rect 17082 18437 17110 18438
rect 17082 18411 17100 18437
rect 17100 18411 17110 18437
rect 17082 18410 17110 18411
rect 17134 18437 17162 18438
rect 17134 18411 17136 18437
rect 17136 18411 17162 18437
rect 17134 18410 17162 18411
rect 17186 18437 17214 18438
rect 17238 18437 17266 18438
rect 17186 18411 17198 18437
rect 17198 18411 17214 18437
rect 17238 18411 17260 18437
rect 17260 18411 17266 18437
rect 17186 18410 17214 18411
rect 17238 18410 17266 18411
rect 17290 18410 17318 18438
rect 17342 18437 17370 18438
rect 17394 18437 17422 18438
rect 17342 18411 17348 18437
rect 17348 18411 17370 18437
rect 17394 18411 17410 18437
rect 17410 18411 17422 18437
rect 17342 18410 17370 18411
rect 17394 18410 17422 18411
rect 17446 18437 17474 18438
rect 17446 18411 17472 18437
rect 17472 18411 17474 18437
rect 17446 18410 17474 18411
rect 17498 18437 17526 18438
rect 17498 18411 17508 18437
rect 17508 18411 17526 18437
rect 17498 18410 17526 18411
rect 9582 18045 9610 18046
rect 9582 18019 9600 18045
rect 9600 18019 9610 18045
rect 9582 18018 9610 18019
rect 9634 18045 9662 18046
rect 9634 18019 9636 18045
rect 9636 18019 9662 18045
rect 9634 18018 9662 18019
rect 9686 18045 9714 18046
rect 9738 18045 9766 18046
rect 9686 18019 9698 18045
rect 9698 18019 9714 18045
rect 9738 18019 9760 18045
rect 9760 18019 9766 18045
rect 9686 18018 9714 18019
rect 9738 18018 9766 18019
rect 9790 18018 9818 18046
rect 9842 18045 9870 18046
rect 9894 18045 9922 18046
rect 9842 18019 9848 18045
rect 9848 18019 9870 18045
rect 9894 18019 9910 18045
rect 9910 18019 9922 18045
rect 9842 18018 9870 18019
rect 9894 18018 9922 18019
rect 9946 18045 9974 18046
rect 9946 18019 9972 18045
rect 9972 18019 9974 18045
rect 9946 18018 9974 18019
rect 9998 18045 10026 18046
rect 9998 18019 10008 18045
rect 10008 18019 10026 18045
rect 9998 18018 10026 18019
rect 9254 17822 9282 17850
rect 7082 17653 7110 17654
rect 7082 17627 7100 17653
rect 7100 17627 7110 17653
rect 7082 17626 7110 17627
rect 7134 17653 7162 17654
rect 7134 17627 7136 17653
rect 7136 17627 7162 17653
rect 7134 17626 7162 17627
rect 7186 17653 7214 17654
rect 7238 17653 7266 17654
rect 7186 17627 7198 17653
rect 7198 17627 7214 17653
rect 7238 17627 7260 17653
rect 7260 17627 7266 17653
rect 7186 17626 7214 17627
rect 7238 17626 7266 17627
rect 7290 17626 7318 17654
rect 7342 17653 7370 17654
rect 7394 17653 7422 17654
rect 7342 17627 7348 17653
rect 7348 17627 7370 17653
rect 7394 17627 7410 17653
rect 7410 17627 7422 17653
rect 7342 17626 7370 17627
rect 7394 17626 7422 17627
rect 7446 17653 7474 17654
rect 7446 17627 7472 17653
rect 7472 17627 7474 17653
rect 7446 17626 7474 17627
rect 7498 17653 7526 17654
rect 7498 17627 7508 17653
rect 7508 17627 7526 17653
rect 7498 17626 7526 17627
rect 9814 17849 9842 17850
rect 9814 17823 9815 17849
rect 9815 17823 9841 17849
rect 9841 17823 9842 17849
rect 9814 17822 9842 17823
rect 7082 16869 7110 16870
rect 7082 16843 7100 16869
rect 7100 16843 7110 16869
rect 7082 16842 7110 16843
rect 7134 16869 7162 16870
rect 7134 16843 7136 16869
rect 7136 16843 7162 16869
rect 7134 16842 7162 16843
rect 7186 16869 7214 16870
rect 7238 16869 7266 16870
rect 7186 16843 7198 16869
rect 7198 16843 7214 16869
rect 7238 16843 7260 16869
rect 7260 16843 7266 16869
rect 7186 16842 7214 16843
rect 7238 16842 7266 16843
rect 7290 16842 7318 16870
rect 7342 16869 7370 16870
rect 7394 16869 7422 16870
rect 7342 16843 7348 16869
rect 7348 16843 7370 16869
rect 7394 16843 7410 16869
rect 7410 16843 7422 16869
rect 7342 16842 7370 16843
rect 7394 16842 7422 16843
rect 7446 16869 7474 16870
rect 7446 16843 7472 16869
rect 7472 16843 7474 16869
rect 7446 16842 7474 16843
rect 7498 16869 7526 16870
rect 7498 16843 7508 16869
rect 7508 16843 7526 16869
rect 7498 16842 7526 16843
rect 7798 16673 7826 16674
rect 7798 16647 7799 16673
rect 7799 16647 7825 16673
rect 7825 16647 7826 16673
rect 7798 16646 7826 16647
rect 7082 16085 7110 16086
rect 7082 16059 7100 16085
rect 7100 16059 7110 16085
rect 7082 16058 7110 16059
rect 7134 16085 7162 16086
rect 7134 16059 7136 16085
rect 7136 16059 7162 16085
rect 7134 16058 7162 16059
rect 7186 16085 7214 16086
rect 7238 16085 7266 16086
rect 7186 16059 7198 16085
rect 7198 16059 7214 16085
rect 7238 16059 7260 16085
rect 7260 16059 7266 16085
rect 7186 16058 7214 16059
rect 7238 16058 7266 16059
rect 7290 16058 7318 16086
rect 7342 16085 7370 16086
rect 7394 16085 7422 16086
rect 7342 16059 7348 16085
rect 7348 16059 7370 16085
rect 7394 16059 7410 16085
rect 7410 16059 7422 16085
rect 7342 16058 7370 16059
rect 7394 16058 7422 16059
rect 7446 16085 7474 16086
rect 7446 16059 7472 16085
rect 7472 16059 7474 16085
rect 7446 16058 7474 16059
rect 7498 16085 7526 16086
rect 7498 16059 7508 16085
rect 7508 16059 7526 16085
rect 7498 16058 7526 16059
rect 6790 8806 6818 8834
rect 6902 14798 6930 14826
rect 6902 14630 6930 14658
rect 5894 7966 5922 7994
rect 6230 7630 6258 7658
rect 4582 7069 4610 7070
rect 4582 7043 4600 7069
rect 4600 7043 4610 7069
rect 4582 7042 4610 7043
rect 4634 7069 4662 7070
rect 4634 7043 4636 7069
rect 4636 7043 4662 7069
rect 4634 7042 4662 7043
rect 4686 7069 4714 7070
rect 4738 7069 4766 7070
rect 4686 7043 4698 7069
rect 4698 7043 4714 7069
rect 4738 7043 4760 7069
rect 4760 7043 4766 7069
rect 4686 7042 4714 7043
rect 4738 7042 4766 7043
rect 4790 7042 4818 7070
rect 4842 7069 4870 7070
rect 4894 7069 4922 7070
rect 4842 7043 4848 7069
rect 4848 7043 4870 7069
rect 4894 7043 4910 7069
rect 4910 7043 4922 7069
rect 4842 7042 4870 7043
rect 4894 7042 4922 7043
rect 4946 7069 4974 7070
rect 4946 7043 4972 7069
rect 4972 7043 4974 7069
rect 4946 7042 4974 7043
rect 4998 7069 5026 7070
rect 4998 7043 5008 7069
rect 5008 7043 5026 7069
rect 4998 7042 5026 7043
rect 4102 6790 4130 6818
rect 5278 6790 5306 6818
rect 4582 6285 4610 6286
rect 4582 6259 4600 6285
rect 4600 6259 4610 6285
rect 4582 6258 4610 6259
rect 4634 6285 4662 6286
rect 4634 6259 4636 6285
rect 4636 6259 4662 6285
rect 4634 6258 4662 6259
rect 4686 6285 4714 6286
rect 4738 6285 4766 6286
rect 4686 6259 4698 6285
rect 4698 6259 4714 6285
rect 4738 6259 4760 6285
rect 4760 6259 4766 6285
rect 4686 6258 4714 6259
rect 4738 6258 4766 6259
rect 4790 6258 4818 6286
rect 4842 6285 4870 6286
rect 4894 6285 4922 6286
rect 4842 6259 4848 6285
rect 4848 6259 4870 6285
rect 4894 6259 4910 6285
rect 4910 6259 4922 6285
rect 4842 6258 4870 6259
rect 4894 6258 4922 6259
rect 4946 6285 4974 6286
rect 4946 6259 4972 6285
rect 4972 6259 4974 6285
rect 4946 6258 4974 6259
rect 4998 6285 5026 6286
rect 4998 6259 5008 6285
rect 5008 6259 5026 6285
rect 4998 6258 5026 6259
rect 3710 4214 3738 4242
rect 4102 6062 4130 6090
rect 4998 5697 5026 5698
rect 4998 5671 4999 5697
rect 4999 5671 5025 5697
rect 5025 5671 5026 5697
rect 4998 5670 5026 5671
rect 4582 5501 4610 5502
rect 4582 5475 4600 5501
rect 4600 5475 4610 5501
rect 4582 5474 4610 5475
rect 4634 5501 4662 5502
rect 4634 5475 4636 5501
rect 4636 5475 4662 5501
rect 4634 5474 4662 5475
rect 4686 5501 4714 5502
rect 4738 5501 4766 5502
rect 4686 5475 4698 5501
rect 4698 5475 4714 5501
rect 4738 5475 4760 5501
rect 4760 5475 4766 5501
rect 4686 5474 4714 5475
rect 4738 5474 4766 5475
rect 4790 5474 4818 5502
rect 4842 5501 4870 5502
rect 4894 5501 4922 5502
rect 4842 5475 4848 5501
rect 4848 5475 4870 5501
rect 4894 5475 4910 5501
rect 4910 5475 4922 5501
rect 4842 5474 4870 5475
rect 4894 5474 4922 5475
rect 4946 5501 4974 5502
rect 4946 5475 4972 5501
rect 4972 5475 4974 5501
rect 4946 5474 4974 5475
rect 4998 5501 5026 5502
rect 4998 5475 5008 5501
rect 5008 5475 5026 5501
rect 4998 5474 5026 5475
rect 4494 5054 4522 5082
rect 4998 5054 5026 5082
rect 3598 4102 3626 4130
rect 5838 5697 5866 5698
rect 5838 5671 5839 5697
rect 5839 5671 5865 5697
rect 5865 5671 5866 5697
rect 5838 5670 5866 5671
rect 5950 5054 5978 5082
rect 4582 4717 4610 4718
rect 4582 4691 4600 4717
rect 4600 4691 4610 4717
rect 4582 4690 4610 4691
rect 4634 4717 4662 4718
rect 4634 4691 4636 4717
rect 4636 4691 4662 4717
rect 4634 4690 4662 4691
rect 4686 4717 4714 4718
rect 4738 4717 4766 4718
rect 4686 4691 4698 4717
rect 4698 4691 4714 4717
rect 4738 4691 4760 4717
rect 4760 4691 4766 4717
rect 4686 4690 4714 4691
rect 4738 4690 4766 4691
rect 4790 4690 4818 4718
rect 4842 4717 4870 4718
rect 4894 4717 4922 4718
rect 4842 4691 4848 4717
rect 4848 4691 4870 4717
rect 4894 4691 4910 4717
rect 4910 4691 4922 4717
rect 4842 4690 4870 4691
rect 4894 4690 4922 4691
rect 4946 4717 4974 4718
rect 4946 4691 4972 4717
rect 4972 4691 4974 4717
rect 4946 4690 4974 4691
rect 4998 4717 5026 4718
rect 4998 4691 5008 4717
rect 5008 4691 5026 4717
rect 4998 4690 5026 4691
rect 4494 4521 4522 4522
rect 4494 4495 4495 4521
rect 4495 4495 4521 4521
rect 4521 4495 4522 4521
rect 4494 4494 4522 4495
rect 4774 4494 4802 4522
rect 4102 4129 4130 4130
rect 4102 4103 4103 4129
rect 4103 4103 4129 4129
rect 4129 4103 4130 4129
rect 4102 4102 4130 4103
rect 5278 4129 5306 4130
rect 5278 4103 5279 4129
rect 5279 4103 5305 4129
rect 5305 4103 5306 4129
rect 5278 4102 5306 4103
rect 4582 3933 4610 3934
rect 4582 3907 4600 3933
rect 4600 3907 4610 3933
rect 4582 3906 4610 3907
rect 4634 3933 4662 3934
rect 4634 3907 4636 3933
rect 4636 3907 4662 3933
rect 4634 3906 4662 3907
rect 4686 3933 4714 3934
rect 4738 3933 4766 3934
rect 4686 3907 4698 3933
rect 4698 3907 4714 3933
rect 4738 3907 4760 3933
rect 4760 3907 4766 3933
rect 4686 3906 4714 3907
rect 4738 3906 4766 3907
rect 4790 3906 4818 3934
rect 4842 3933 4870 3934
rect 4894 3933 4922 3934
rect 4842 3907 4848 3933
rect 4848 3907 4870 3933
rect 4894 3907 4910 3933
rect 4910 3907 4922 3933
rect 4842 3906 4870 3907
rect 4894 3906 4922 3907
rect 4946 3933 4974 3934
rect 4946 3907 4972 3933
rect 4972 3907 4974 3933
rect 4946 3906 4974 3907
rect 4998 3933 5026 3934
rect 4998 3907 5008 3933
rect 5008 3907 5026 3933
rect 4998 3906 5026 3907
rect 6454 6062 6482 6090
rect 6118 5305 6146 5306
rect 6118 5279 6119 5305
rect 6119 5279 6145 5305
rect 6145 5279 6146 5305
rect 6118 5278 6146 5279
rect 6454 4913 6482 4914
rect 6454 4887 6455 4913
rect 6455 4887 6481 4913
rect 6481 4887 6482 4913
rect 6454 4886 6482 4887
rect 6790 4886 6818 4914
rect 6790 4521 6818 4522
rect 6790 4495 6791 4521
rect 6791 4495 6817 4521
rect 6817 4495 6818 4521
rect 6790 4494 6818 4495
rect 7082 15301 7110 15302
rect 7082 15275 7100 15301
rect 7100 15275 7110 15301
rect 7082 15274 7110 15275
rect 7134 15301 7162 15302
rect 7134 15275 7136 15301
rect 7136 15275 7162 15301
rect 7134 15274 7162 15275
rect 7186 15301 7214 15302
rect 7238 15301 7266 15302
rect 7186 15275 7198 15301
rect 7198 15275 7214 15301
rect 7238 15275 7260 15301
rect 7260 15275 7266 15301
rect 7186 15274 7214 15275
rect 7238 15274 7266 15275
rect 7290 15274 7318 15302
rect 7342 15301 7370 15302
rect 7394 15301 7422 15302
rect 7342 15275 7348 15301
rect 7348 15275 7370 15301
rect 7394 15275 7410 15301
rect 7410 15275 7422 15301
rect 7342 15274 7370 15275
rect 7394 15274 7422 15275
rect 7446 15301 7474 15302
rect 7446 15275 7472 15301
rect 7472 15275 7474 15301
rect 7446 15274 7474 15275
rect 7498 15301 7526 15302
rect 7498 15275 7508 15301
rect 7508 15275 7526 15301
rect 7498 15274 7526 15275
rect 7082 14517 7110 14518
rect 7082 14491 7100 14517
rect 7100 14491 7110 14517
rect 7082 14490 7110 14491
rect 7134 14517 7162 14518
rect 7134 14491 7136 14517
rect 7136 14491 7162 14517
rect 7134 14490 7162 14491
rect 7186 14517 7214 14518
rect 7238 14517 7266 14518
rect 7186 14491 7198 14517
rect 7198 14491 7214 14517
rect 7238 14491 7260 14517
rect 7260 14491 7266 14517
rect 7186 14490 7214 14491
rect 7238 14490 7266 14491
rect 7290 14490 7318 14518
rect 7342 14517 7370 14518
rect 7394 14517 7422 14518
rect 7342 14491 7348 14517
rect 7348 14491 7370 14517
rect 7394 14491 7410 14517
rect 7410 14491 7422 14517
rect 7342 14490 7370 14491
rect 7394 14490 7422 14491
rect 7446 14517 7474 14518
rect 7446 14491 7472 14517
rect 7472 14491 7474 14517
rect 7446 14490 7474 14491
rect 7498 14517 7526 14518
rect 7498 14491 7508 14517
rect 7508 14491 7526 14517
rect 7498 14490 7526 14491
rect 11102 17822 11130 17850
rect 9582 17261 9610 17262
rect 9582 17235 9600 17261
rect 9600 17235 9610 17261
rect 9582 17234 9610 17235
rect 9634 17261 9662 17262
rect 9634 17235 9636 17261
rect 9636 17235 9662 17261
rect 9634 17234 9662 17235
rect 9686 17261 9714 17262
rect 9738 17261 9766 17262
rect 9686 17235 9698 17261
rect 9698 17235 9714 17261
rect 9738 17235 9760 17261
rect 9760 17235 9766 17261
rect 9686 17234 9714 17235
rect 9738 17234 9766 17235
rect 9790 17234 9818 17262
rect 9842 17261 9870 17262
rect 9894 17261 9922 17262
rect 9842 17235 9848 17261
rect 9848 17235 9870 17261
rect 9894 17235 9910 17261
rect 9910 17235 9922 17261
rect 9842 17234 9870 17235
rect 9894 17234 9922 17235
rect 9946 17261 9974 17262
rect 9946 17235 9972 17261
rect 9972 17235 9974 17261
rect 9946 17234 9974 17235
rect 9998 17261 10026 17262
rect 9998 17235 10008 17261
rect 10008 17235 10026 17261
rect 9998 17234 10026 17235
rect 9254 16646 9282 16674
rect 7798 14686 7826 14714
rect 7082 13733 7110 13734
rect 7082 13707 7100 13733
rect 7100 13707 7110 13733
rect 7082 13706 7110 13707
rect 7134 13733 7162 13734
rect 7134 13707 7136 13733
rect 7136 13707 7162 13733
rect 7134 13706 7162 13707
rect 7186 13733 7214 13734
rect 7238 13733 7266 13734
rect 7186 13707 7198 13733
rect 7198 13707 7214 13733
rect 7238 13707 7260 13733
rect 7260 13707 7266 13733
rect 7186 13706 7214 13707
rect 7238 13706 7266 13707
rect 7290 13706 7318 13734
rect 7342 13733 7370 13734
rect 7394 13733 7422 13734
rect 7342 13707 7348 13733
rect 7348 13707 7370 13733
rect 7394 13707 7410 13733
rect 7410 13707 7422 13733
rect 7342 13706 7370 13707
rect 7394 13706 7422 13707
rect 7446 13733 7474 13734
rect 7446 13707 7472 13733
rect 7472 13707 7474 13733
rect 7446 13706 7474 13707
rect 7498 13733 7526 13734
rect 7498 13707 7508 13733
rect 7508 13707 7526 13733
rect 7498 13706 7526 13707
rect 7082 12949 7110 12950
rect 7082 12923 7100 12949
rect 7100 12923 7110 12949
rect 7082 12922 7110 12923
rect 7134 12949 7162 12950
rect 7134 12923 7136 12949
rect 7136 12923 7162 12949
rect 7134 12922 7162 12923
rect 7186 12949 7214 12950
rect 7238 12949 7266 12950
rect 7186 12923 7198 12949
rect 7198 12923 7214 12949
rect 7238 12923 7260 12949
rect 7260 12923 7266 12949
rect 7186 12922 7214 12923
rect 7238 12922 7266 12923
rect 7290 12922 7318 12950
rect 7342 12949 7370 12950
rect 7394 12949 7422 12950
rect 7342 12923 7348 12949
rect 7348 12923 7370 12949
rect 7394 12923 7410 12949
rect 7410 12923 7422 12949
rect 7342 12922 7370 12923
rect 7394 12922 7422 12923
rect 7446 12949 7474 12950
rect 7446 12923 7472 12949
rect 7472 12923 7474 12949
rect 7446 12922 7474 12923
rect 7498 12949 7526 12950
rect 7498 12923 7508 12949
rect 7508 12923 7526 12949
rect 7498 12922 7526 12923
rect 7014 12670 7042 12698
rect 7014 12417 7042 12418
rect 7014 12391 7015 12417
rect 7015 12391 7041 12417
rect 7041 12391 7042 12417
rect 7014 12390 7042 12391
rect 7574 12361 7602 12362
rect 7574 12335 7575 12361
rect 7575 12335 7601 12361
rect 7601 12335 7602 12361
rect 7574 12334 7602 12335
rect 7082 12165 7110 12166
rect 7082 12139 7100 12165
rect 7100 12139 7110 12165
rect 7082 12138 7110 12139
rect 7134 12165 7162 12166
rect 7134 12139 7136 12165
rect 7136 12139 7162 12165
rect 7134 12138 7162 12139
rect 7186 12165 7214 12166
rect 7238 12165 7266 12166
rect 7186 12139 7198 12165
rect 7198 12139 7214 12165
rect 7238 12139 7260 12165
rect 7260 12139 7266 12165
rect 7186 12138 7214 12139
rect 7238 12138 7266 12139
rect 7290 12138 7318 12166
rect 7342 12165 7370 12166
rect 7394 12165 7422 12166
rect 7342 12139 7348 12165
rect 7348 12139 7370 12165
rect 7394 12139 7410 12165
rect 7410 12139 7422 12165
rect 7342 12138 7370 12139
rect 7394 12138 7422 12139
rect 7446 12165 7474 12166
rect 7446 12139 7472 12165
rect 7472 12139 7474 12165
rect 7446 12138 7474 12139
rect 7498 12165 7526 12166
rect 7498 12139 7508 12165
rect 7508 12139 7526 12165
rect 7498 12138 7526 12139
rect 7574 11774 7602 11802
rect 8470 14713 8498 14714
rect 8470 14687 8471 14713
rect 8471 14687 8497 14713
rect 8497 14687 8498 14713
rect 8470 14686 8498 14687
rect 8974 14686 9002 14714
rect 8974 14321 9002 14322
rect 8974 14295 8975 14321
rect 8975 14295 9001 14321
rect 9001 14295 9002 14321
rect 8974 14294 9002 14295
rect 9582 16477 9610 16478
rect 9582 16451 9600 16477
rect 9600 16451 9610 16477
rect 9582 16450 9610 16451
rect 9634 16477 9662 16478
rect 9634 16451 9636 16477
rect 9636 16451 9662 16477
rect 9634 16450 9662 16451
rect 9686 16477 9714 16478
rect 9738 16477 9766 16478
rect 9686 16451 9698 16477
rect 9698 16451 9714 16477
rect 9738 16451 9760 16477
rect 9760 16451 9766 16477
rect 9686 16450 9714 16451
rect 9738 16450 9766 16451
rect 9790 16450 9818 16478
rect 9842 16477 9870 16478
rect 9894 16477 9922 16478
rect 9842 16451 9848 16477
rect 9848 16451 9870 16477
rect 9894 16451 9910 16477
rect 9910 16451 9922 16477
rect 9842 16450 9870 16451
rect 9894 16450 9922 16451
rect 9946 16477 9974 16478
rect 9946 16451 9972 16477
rect 9972 16451 9974 16477
rect 9946 16450 9974 16451
rect 9998 16477 10026 16478
rect 9998 16451 10008 16477
rect 10008 16451 10026 16477
rect 9998 16450 10026 16451
rect 10094 16281 10122 16282
rect 10094 16255 10095 16281
rect 10095 16255 10121 16281
rect 10121 16255 10122 16281
rect 10094 16254 10122 16255
rect 10430 15833 10458 15834
rect 10430 15807 10431 15833
rect 10431 15807 10457 15833
rect 10457 15807 10458 15833
rect 10430 15806 10458 15807
rect 9582 15693 9610 15694
rect 9582 15667 9600 15693
rect 9600 15667 9610 15693
rect 9582 15666 9610 15667
rect 9634 15693 9662 15694
rect 9634 15667 9636 15693
rect 9636 15667 9662 15693
rect 9634 15666 9662 15667
rect 9686 15693 9714 15694
rect 9738 15693 9766 15694
rect 9686 15667 9698 15693
rect 9698 15667 9714 15693
rect 9738 15667 9760 15693
rect 9760 15667 9766 15693
rect 9686 15666 9714 15667
rect 9738 15666 9766 15667
rect 9790 15666 9818 15694
rect 9842 15693 9870 15694
rect 9894 15693 9922 15694
rect 9842 15667 9848 15693
rect 9848 15667 9870 15693
rect 9894 15667 9910 15693
rect 9910 15667 9922 15693
rect 9842 15666 9870 15667
rect 9894 15666 9922 15667
rect 9946 15693 9974 15694
rect 9946 15667 9972 15693
rect 9972 15667 9974 15693
rect 9946 15666 9974 15667
rect 9998 15693 10026 15694
rect 9998 15667 10008 15693
rect 10008 15667 10026 15693
rect 9998 15666 10026 15667
rect 10038 15497 10066 15498
rect 10038 15471 10039 15497
rect 10039 15471 10065 15497
rect 10065 15471 10066 15497
rect 10038 15470 10066 15471
rect 10990 16281 11018 16282
rect 10990 16255 10991 16281
rect 10991 16255 11017 16281
rect 11017 16255 11018 16281
rect 10990 16254 11018 16255
rect 10990 15806 11018 15834
rect 11270 15497 11298 15498
rect 11270 15471 11271 15497
rect 11271 15471 11297 15497
rect 11297 15471 11298 15497
rect 11270 15470 11298 15471
rect 9582 14909 9610 14910
rect 9582 14883 9600 14909
rect 9600 14883 9610 14909
rect 9582 14882 9610 14883
rect 9634 14909 9662 14910
rect 9634 14883 9636 14909
rect 9636 14883 9662 14909
rect 9634 14882 9662 14883
rect 9686 14909 9714 14910
rect 9738 14909 9766 14910
rect 9686 14883 9698 14909
rect 9698 14883 9714 14909
rect 9738 14883 9760 14909
rect 9760 14883 9766 14909
rect 9686 14882 9714 14883
rect 9738 14882 9766 14883
rect 9790 14882 9818 14910
rect 9842 14909 9870 14910
rect 9894 14909 9922 14910
rect 9842 14883 9848 14909
rect 9848 14883 9870 14909
rect 9894 14883 9910 14909
rect 9910 14883 9922 14909
rect 9842 14882 9870 14883
rect 9894 14882 9922 14883
rect 9946 14909 9974 14910
rect 9946 14883 9972 14909
rect 9972 14883 9974 14909
rect 9946 14882 9974 14883
rect 9998 14909 10026 14910
rect 9998 14883 10008 14909
rect 10008 14883 10026 14909
rect 9998 14882 10026 14883
rect 8862 13846 8890 13874
rect 8358 12417 8386 12418
rect 8358 12391 8359 12417
rect 8359 12391 8385 12417
rect 8385 12391 8386 12417
rect 8358 12390 8386 12391
rect 8078 11774 8106 11802
rect 7082 11381 7110 11382
rect 7082 11355 7100 11381
rect 7100 11355 7110 11381
rect 7082 11354 7110 11355
rect 7134 11381 7162 11382
rect 7134 11355 7136 11381
rect 7136 11355 7162 11381
rect 7134 11354 7162 11355
rect 7186 11381 7214 11382
rect 7238 11381 7266 11382
rect 7186 11355 7198 11381
rect 7198 11355 7214 11381
rect 7238 11355 7260 11381
rect 7260 11355 7266 11381
rect 7186 11354 7214 11355
rect 7238 11354 7266 11355
rect 7290 11354 7318 11382
rect 7342 11381 7370 11382
rect 7394 11381 7422 11382
rect 7342 11355 7348 11381
rect 7348 11355 7370 11381
rect 7394 11355 7410 11381
rect 7410 11355 7422 11381
rect 7342 11354 7370 11355
rect 7394 11354 7422 11355
rect 7446 11381 7474 11382
rect 7446 11355 7472 11381
rect 7472 11355 7474 11381
rect 7446 11354 7474 11355
rect 7498 11381 7526 11382
rect 7498 11355 7508 11381
rect 7508 11355 7526 11381
rect 7498 11354 7526 11355
rect 8470 11102 8498 11130
rect 7082 10597 7110 10598
rect 7082 10571 7100 10597
rect 7100 10571 7110 10597
rect 7082 10570 7110 10571
rect 7134 10597 7162 10598
rect 7134 10571 7136 10597
rect 7136 10571 7162 10597
rect 7134 10570 7162 10571
rect 7186 10597 7214 10598
rect 7238 10597 7266 10598
rect 7186 10571 7198 10597
rect 7198 10571 7214 10597
rect 7238 10571 7260 10597
rect 7260 10571 7266 10597
rect 7186 10570 7214 10571
rect 7238 10570 7266 10571
rect 7290 10570 7318 10598
rect 7342 10597 7370 10598
rect 7394 10597 7422 10598
rect 7342 10571 7348 10597
rect 7348 10571 7370 10597
rect 7394 10571 7410 10597
rect 7410 10571 7422 10597
rect 7342 10570 7370 10571
rect 7394 10570 7422 10571
rect 7446 10597 7474 10598
rect 7446 10571 7472 10597
rect 7472 10571 7474 10597
rect 7446 10570 7474 10571
rect 7498 10597 7526 10598
rect 7498 10571 7508 10597
rect 7508 10571 7526 10597
rect 7498 10570 7526 10571
rect 7082 9813 7110 9814
rect 7082 9787 7100 9813
rect 7100 9787 7110 9813
rect 7082 9786 7110 9787
rect 7134 9813 7162 9814
rect 7134 9787 7136 9813
rect 7136 9787 7162 9813
rect 7134 9786 7162 9787
rect 7186 9813 7214 9814
rect 7238 9813 7266 9814
rect 7186 9787 7198 9813
rect 7198 9787 7214 9813
rect 7238 9787 7260 9813
rect 7260 9787 7266 9813
rect 7186 9786 7214 9787
rect 7238 9786 7266 9787
rect 7290 9786 7318 9814
rect 7342 9813 7370 9814
rect 7394 9813 7422 9814
rect 7342 9787 7348 9813
rect 7348 9787 7370 9813
rect 7394 9787 7410 9813
rect 7410 9787 7422 9813
rect 7342 9786 7370 9787
rect 7394 9786 7422 9787
rect 7446 9813 7474 9814
rect 7446 9787 7472 9813
rect 7472 9787 7474 9813
rect 7446 9786 7474 9787
rect 7498 9813 7526 9814
rect 7498 9787 7508 9813
rect 7508 9787 7526 9813
rect 7498 9786 7526 9787
rect 7014 9534 7042 9562
rect 7082 9029 7110 9030
rect 7082 9003 7100 9029
rect 7100 9003 7110 9029
rect 7082 9002 7110 9003
rect 7134 9029 7162 9030
rect 7134 9003 7136 9029
rect 7136 9003 7162 9029
rect 7134 9002 7162 9003
rect 7186 9029 7214 9030
rect 7238 9029 7266 9030
rect 7186 9003 7198 9029
rect 7198 9003 7214 9029
rect 7238 9003 7260 9029
rect 7260 9003 7266 9029
rect 7186 9002 7214 9003
rect 7238 9002 7266 9003
rect 7290 9002 7318 9030
rect 7342 9029 7370 9030
rect 7394 9029 7422 9030
rect 7342 9003 7348 9029
rect 7348 9003 7370 9029
rect 7394 9003 7410 9029
rect 7410 9003 7422 9029
rect 7342 9002 7370 9003
rect 7394 9002 7422 9003
rect 7446 9029 7474 9030
rect 7446 9003 7472 9029
rect 7472 9003 7474 9029
rect 7446 9002 7474 9003
rect 7498 9029 7526 9030
rect 7498 9003 7508 9029
rect 7508 9003 7526 9029
rect 7498 9002 7526 9003
rect 7082 8245 7110 8246
rect 7082 8219 7100 8245
rect 7100 8219 7110 8245
rect 7082 8218 7110 8219
rect 7134 8245 7162 8246
rect 7134 8219 7136 8245
rect 7136 8219 7162 8245
rect 7134 8218 7162 8219
rect 7186 8245 7214 8246
rect 7238 8245 7266 8246
rect 7186 8219 7198 8245
rect 7198 8219 7214 8245
rect 7238 8219 7260 8245
rect 7260 8219 7266 8245
rect 7186 8218 7214 8219
rect 7238 8218 7266 8219
rect 7290 8218 7318 8246
rect 7342 8245 7370 8246
rect 7394 8245 7422 8246
rect 7342 8219 7348 8245
rect 7348 8219 7370 8245
rect 7394 8219 7410 8245
rect 7410 8219 7422 8245
rect 7342 8218 7370 8219
rect 7394 8218 7422 8219
rect 7446 8245 7474 8246
rect 7446 8219 7472 8245
rect 7472 8219 7474 8245
rect 7446 8218 7474 8219
rect 7498 8245 7526 8246
rect 7498 8219 7508 8245
rect 7508 8219 7526 8245
rect 7498 8218 7526 8219
rect 7014 7630 7042 7658
rect 8358 8497 8386 8498
rect 8358 8471 8359 8497
rect 8359 8471 8385 8497
rect 8385 8471 8386 8497
rect 8358 8470 8386 8471
rect 7082 7461 7110 7462
rect 7082 7435 7100 7461
rect 7100 7435 7110 7461
rect 7082 7434 7110 7435
rect 7134 7461 7162 7462
rect 7134 7435 7136 7461
rect 7136 7435 7162 7461
rect 7134 7434 7162 7435
rect 7186 7461 7214 7462
rect 7238 7461 7266 7462
rect 7186 7435 7198 7461
rect 7198 7435 7214 7461
rect 7238 7435 7260 7461
rect 7260 7435 7266 7461
rect 7186 7434 7214 7435
rect 7238 7434 7266 7435
rect 7290 7434 7318 7462
rect 7342 7461 7370 7462
rect 7394 7461 7422 7462
rect 7342 7435 7348 7461
rect 7348 7435 7370 7461
rect 7394 7435 7410 7461
rect 7410 7435 7422 7461
rect 7342 7434 7370 7435
rect 7394 7434 7422 7435
rect 7446 7461 7474 7462
rect 7446 7435 7472 7461
rect 7472 7435 7474 7461
rect 7446 7434 7474 7435
rect 7498 7461 7526 7462
rect 7498 7435 7508 7461
rect 7508 7435 7526 7461
rect 7498 7434 7526 7435
rect 7742 7657 7770 7658
rect 7742 7631 7743 7657
rect 7743 7631 7769 7657
rect 7769 7631 7770 7657
rect 7742 7630 7770 7631
rect 7966 7657 7994 7658
rect 7966 7631 7967 7657
rect 7967 7631 7993 7657
rect 7993 7631 7994 7657
rect 7966 7630 7994 7631
rect 8470 7630 8498 7658
rect 7082 6677 7110 6678
rect 7082 6651 7100 6677
rect 7100 6651 7110 6677
rect 7082 6650 7110 6651
rect 7134 6677 7162 6678
rect 7134 6651 7136 6677
rect 7136 6651 7162 6677
rect 7134 6650 7162 6651
rect 7186 6677 7214 6678
rect 7238 6677 7266 6678
rect 7186 6651 7198 6677
rect 7198 6651 7214 6677
rect 7238 6651 7260 6677
rect 7260 6651 7266 6677
rect 7186 6650 7214 6651
rect 7238 6650 7266 6651
rect 7290 6650 7318 6678
rect 7342 6677 7370 6678
rect 7394 6677 7422 6678
rect 7342 6651 7348 6677
rect 7348 6651 7370 6677
rect 7394 6651 7410 6677
rect 7410 6651 7422 6677
rect 7342 6650 7370 6651
rect 7394 6650 7422 6651
rect 7446 6677 7474 6678
rect 7446 6651 7472 6677
rect 7472 6651 7474 6677
rect 7446 6650 7474 6651
rect 7498 6677 7526 6678
rect 7498 6651 7508 6677
rect 7508 6651 7526 6677
rect 7498 6650 7526 6651
rect 7014 6089 7042 6090
rect 7014 6063 7015 6089
rect 7015 6063 7041 6089
rect 7041 6063 7042 6089
rect 7014 6062 7042 6063
rect 7082 5893 7110 5894
rect 7082 5867 7100 5893
rect 7100 5867 7110 5893
rect 7082 5866 7110 5867
rect 7134 5893 7162 5894
rect 7134 5867 7136 5893
rect 7136 5867 7162 5893
rect 7134 5866 7162 5867
rect 7186 5893 7214 5894
rect 7238 5893 7266 5894
rect 7186 5867 7198 5893
rect 7198 5867 7214 5893
rect 7238 5867 7260 5893
rect 7260 5867 7266 5893
rect 7186 5866 7214 5867
rect 7238 5866 7266 5867
rect 7290 5866 7318 5894
rect 7342 5893 7370 5894
rect 7394 5893 7422 5894
rect 7342 5867 7348 5893
rect 7348 5867 7370 5893
rect 7394 5867 7410 5893
rect 7410 5867 7422 5893
rect 7342 5866 7370 5867
rect 7394 5866 7422 5867
rect 7446 5893 7474 5894
rect 7446 5867 7472 5893
rect 7472 5867 7474 5893
rect 7446 5866 7474 5867
rect 7498 5893 7526 5894
rect 7498 5867 7508 5893
rect 7508 5867 7526 5893
rect 7498 5866 7526 5867
rect 7574 5838 7602 5866
rect 8358 6062 8386 6090
rect 8078 5838 8106 5866
rect 7294 5305 7322 5306
rect 7294 5279 7295 5305
rect 7295 5279 7321 5305
rect 7321 5279 7322 5305
rect 7294 5278 7322 5279
rect 8078 5278 8106 5306
rect 7082 5109 7110 5110
rect 7082 5083 7100 5109
rect 7100 5083 7110 5109
rect 7082 5082 7110 5083
rect 7134 5109 7162 5110
rect 7134 5083 7136 5109
rect 7136 5083 7162 5109
rect 7134 5082 7162 5083
rect 7186 5109 7214 5110
rect 7238 5109 7266 5110
rect 7186 5083 7198 5109
rect 7198 5083 7214 5109
rect 7238 5083 7260 5109
rect 7260 5083 7266 5109
rect 7186 5082 7214 5083
rect 7238 5082 7266 5083
rect 7290 5082 7318 5110
rect 7342 5109 7370 5110
rect 7394 5109 7422 5110
rect 7342 5083 7348 5109
rect 7348 5083 7370 5109
rect 7394 5083 7410 5109
rect 7410 5083 7422 5109
rect 7342 5082 7370 5083
rect 7394 5082 7422 5083
rect 7446 5109 7474 5110
rect 7446 5083 7472 5109
rect 7472 5083 7474 5109
rect 7446 5082 7474 5083
rect 7498 5109 7526 5110
rect 7498 5083 7508 5109
rect 7508 5083 7526 5109
rect 7498 5082 7526 5083
rect 7014 4494 7042 4522
rect 7082 4325 7110 4326
rect 7082 4299 7100 4325
rect 7100 4299 7110 4325
rect 7082 4298 7110 4299
rect 7134 4325 7162 4326
rect 7134 4299 7136 4325
rect 7136 4299 7162 4325
rect 7134 4298 7162 4299
rect 7186 4325 7214 4326
rect 7238 4325 7266 4326
rect 7186 4299 7198 4325
rect 7198 4299 7214 4325
rect 7238 4299 7260 4325
rect 7260 4299 7266 4325
rect 7186 4298 7214 4299
rect 7238 4298 7266 4299
rect 7290 4298 7318 4326
rect 7342 4325 7370 4326
rect 7394 4325 7422 4326
rect 7342 4299 7348 4325
rect 7348 4299 7370 4325
rect 7394 4299 7410 4325
rect 7410 4299 7422 4325
rect 7342 4298 7370 4299
rect 7394 4298 7422 4299
rect 7446 4325 7474 4326
rect 7446 4299 7472 4325
rect 7472 4299 7474 4325
rect 7446 4298 7474 4299
rect 7498 4325 7526 4326
rect 7498 4299 7508 4325
rect 7508 4299 7526 4325
rect 7498 4298 7526 4299
rect 5950 4102 5978 4130
rect 6454 4129 6482 4130
rect 6454 4103 6455 4129
rect 6455 4103 6481 4129
rect 6481 4103 6482 4129
rect 6454 4102 6482 4103
rect 5278 3710 5306 3738
rect 5838 3737 5866 3738
rect 5838 3711 5839 3737
rect 5839 3711 5865 3737
rect 5865 3711 5866 3737
rect 5838 3710 5866 3711
rect 4582 3149 4610 3150
rect 4582 3123 4600 3149
rect 4600 3123 4610 3149
rect 4582 3122 4610 3123
rect 4634 3149 4662 3150
rect 4634 3123 4636 3149
rect 4636 3123 4662 3149
rect 4634 3122 4662 3123
rect 4686 3149 4714 3150
rect 4738 3149 4766 3150
rect 4686 3123 4698 3149
rect 4698 3123 4714 3149
rect 4738 3123 4760 3149
rect 4760 3123 4766 3149
rect 4686 3122 4714 3123
rect 4738 3122 4766 3123
rect 4790 3122 4818 3150
rect 4842 3149 4870 3150
rect 4894 3149 4922 3150
rect 4842 3123 4848 3149
rect 4848 3123 4870 3149
rect 4894 3123 4910 3149
rect 4910 3123 4922 3149
rect 4842 3122 4870 3123
rect 4894 3122 4922 3123
rect 4946 3149 4974 3150
rect 4946 3123 4972 3149
rect 4972 3123 4974 3149
rect 4946 3122 4974 3123
rect 4998 3149 5026 3150
rect 4998 3123 5008 3149
rect 5008 3123 5026 3149
rect 4998 3122 5026 3123
rect 4494 2478 4522 2506
rect 5390 3430 5418 3458
rect 4998 2505 5026 2506
rect 4998 2479 4999 2505
rect 4999 2479 5025 2505
rect 5025 2479 5026 2505
rect 4998 2478 5026 2479
rect 4582 2365 4610 2366
rect 4582 2339 4600 2365
rect 4600 2339 4610 2365
rect 4582 2338 4610 2339
rect 4634 2365 4662 2366
rect 4634 2339 4636 2365
rect 4636 2339 4662 2365
rect 4634 2338 4662 2339
rect 4686 2365 4714 2366
rect 4738 2365 4766 2366
rect 4686 2339 4698 2365
rect 4698 2339 4714 2365
rect 4738 2339 4760 2365
rect 4760 2339 4766 2365
rect 4686 2338 4714 2339
rect 4738 2338 4766 2339
rect 4790 2338 4818 2366
rect 4842 2365 4870 2366
rect 4894 2365 4922 2366
rect 4842 2339 4848 2365
rect 4848 2339 4870 2365
rect 4894 2339 4910 2365
rect 4910 2339 4922 2365
rect 4842 2338 4870 2339
rect 4894 2338 4922 2339
rect 4946 2365 4974 2366
rect 4946 2339 4972 2365
rect 4972 2339 4974 2365
rect 4946 2338 4974 2339
rect 4998 2365 5026 2366
rect 4998 2339 5008 2365
rect 5008 2339 5026 2365
rect 4998 2338 5026 2339
rect 3822 1806 3850 1834
rect 4438 2225 4466 2226
rect 4438 2199 4439 2225
rect 4439 2199 4465 2225
rect 4465 2199 4466 2225
rect 4438 2198 4466 2199
rect 4438 1721 4466 1722
rect 4438 1695 4439 1721
rect 4439 1695 4465 1721
rect 4465 1695 4466 1721
rect 4438 1694 4466 1695
rect 4582 1581 4610 1582
rect 4582 1555 4600 1581
rect 4600 1555 4610 1581
rect 4582 1554 4610 1555
rect 4634 1581 4662 1582
rect 4634 1555 4636 1581
rect 4636 1555 4662 1581
rect 4634 1554 4662 1555
rect 4686 1581 4714 1582
rect 4738 1581 4766 1582
rect 4686 1555 4698 1581
rect 4698 1555 4714 1581
rect 4738 1555 4760 1581
rect 4760 1555 4766 1581
rect 4686 1554 4714 1555
rect 4738 1554 4766 1555
rect 4790 1554 4818 1582
rect 4842 1581 4870 1582
rect 4894 1581 4922 1582
rect 4842 1555 4848 1581
rect 4848 1555 4870 1581
rect 4894 1555 4910 1581
rect 4910 1555 4922 1581
rect 4842 1554 4870 1555
rect 4894 1554 4922 1555
rect 4946 1581 4974 1582
rect 4946 1555 4972 1581
rect 4972 1555 4974 1581
rect 4946 1554 4974 1555
rect 4998 1581 5026 1582
rect 4998 1555 5008 1581
rect 5008 1555 5026 1581
rect 4998 1554 5026 1555
rect 6454 3710 6482 3738
rect 6454 3289 6482 3290
rect 6454 3263 6455 3289
rect 6455 3263 6481 3289
rect 6481 3263 6482 3289
rect 6454 3262 6482 3263
rect 5894 2169 5922 2170
rect 5894 2143 5895 2169
rect 5895 2143 5921 2169
rect 5921 2143 5922 2169
rect 5894 2142 5922 2143
rect 6342 2478 6370 2506
rect 5502 1806 5530 1834
rect 6510 1750 6538 1778
rect 6398 1414 6426 1442
rect 7014 4158 7042 4186
rect 6958 3737 6986 3738
rect 6958 3711 6959 3737
rect 6959 3711 6985 3737
rect 6985 3711 6986 3737
rect 6958 3710 6986 3711
rect 8470 4521 8498 4522
rect 8470 4495 8471 4521
rect 8471 4495 8497 4521
rect 8497 4495 8498 4521
rect 8470 4494 8498 4495
rect 8470 4158 8498 4186
rect 7082 3541 7110 3542
rect 7082 3515 7100 3541
rect 7100 3515 7110 3541
rect 7082 3514 7110 3515
rect 7134 3541 7162 3542
rect 7134 3515 7136 3541
rect 7136 3515 7162 3541
rect 7134 3514 7162 3515
rect 7186 3541 7214 3542
rect 7238 3541 7266 3542
rect 7186 3515 7198 3541
rect 7198 3515 7214 3541
rect 7238 3515 7260 3541
rect 7260 3515 7266 3541
rect 7186 3514 7214 3515
rect 7238 3514 7266 3515
rect 7290 3514 7318 3542
rect 7342 3541 7370 3542
rect 7394 3541 7422 3542
rect 7342 3515 7348 3541
rect 7348 3515 7370 3541
rect 7394 3515 7410 3541
rect 7410 3515 7422 3541
rect 7342 3514 7370 3515
rect 7394 3514 7422 3515
rect 7446 3541 7474 3542
rect 7446 3515 7472 3541
rect 7472 3515 7474 3541
rect 7446 3514 7474 3515
rect 7498 3541 7526 3542
rect 7498 3515 7508 3541
rect 7508 3515 7526 3541
rect 7498 3514 7526 3515
rect 8078 3374 8106 3402
rect 8358 3737 8386 3738
rect 8358 3711 8359 3737
rect 8359 3711 8385 3737
rect 8385 3711 8386 3737
rect 8358 3710 8386 3711
rect 7014 3262 7042 3290
rect 10374 14321 10402 14322
rect 10374 14295 10375 14321
rect 10375 14295 10401 14321
rect 10401 14295 10402 14321
rect 10374 14294 10402 14295
rect 9582 14125 9610 14126
rect 9582 14099 9600 14125
rect 9600 14099 9610 14125
rect 9582 14098 9610 14099
rect 9634 14125 9662 14126
rect 9634 14099 9636 14125
rect 9636 14099 9662 14125
rect 9634 14098 9662 14099
rect 9686 14125 9714 14126
rect 9738 14125 9766 14126
rect 9686 14099 9698 14125
rect 9698 14099 9714 14125
rect 9738 14099 9760 14125
rect 9760 14099 9766 14125
rect 9686 14098 9714 14099
rect 9738 14098 9766 14099
rect 9790 14098 9818 14126
rect 9842 14125 9870 14126
rect 9894 14125 9922 14126
rect 9842 14099 9848 14125
rect 9848 14099 9870 14125
rect 9894 14099 9910 14125
rect 9910 14099 9922 14125
rect 9842 14098 9870 14099
rect 9894 14098 9922 14099
rect 9946 14125 9974 14126
rect 9946 14099 9972 14125
rect 9972 14099 9974 14125
rect 9946 14098 9974 14099
rect 9998 14125 10026 14126
rect 9998 14099 10008 14125
rect 10008 14099 10026 14125
rect 9998 14098 10026 14099
rect 9582 13341 9610 13342
rect 9582 13315 9600 13341
rect 9600 13315 9610 13341
rect 9582 13314 9610 13315
rect 9634 13341 9662 13342
rect 9634 13315 9636 13341
rect 9636 13315 9662 13341
rect 9634 13314 9662 13315
rect 9686 13341 9714 13342
rect 9738 13341 9766 13342
rect 9686 13315 9698 13341
rect 9698 13315 9714 13341
rect 9738 13315 9760 13341
rect 9760 13315 9766 13341
rect 9686 13314 9714 13315
rect 9738 13314 9766 13315
rect 9790 13314 9818 13342
rect 9842 13341 9870 13342
rect 9894 13341 9922 13342
rect 9842 13315 9848 13341
rect 9848 13315 9870 13341
rect 9894 13315 9910 13341
rect 9910 13315 9922 13341
rect 9842 13314 9870 13315
rect 9894 13314 9922 13315
rect 9946 13341 9974 13342
rect 9946 13315 9972 13341
rect 9972 13315 9974 13341
rect 9946 13314 9974 13315
rect 9998 13341 10026 13342
rect 9998 13315 10008 13341
rect 10008 13315 10026 13341
rect 9998 13314 10026 13315
rect 9582 12557 9610 12558
rect 9582 12531 9600 12557
rect 9600 12531 9610 12557
rect 9582 12530 9610 12531
rect 9634 12557 9662 12558
rect 9634 12531 9636 12557
rect 9636 12531 9662 12557
rect 9634 12530 9662 12531
rect 9686 12557 9714 12558
rect 9738 12557 9766 12558
rect 9686 12531 9698 12557
rect 9698 12531 9714 12557
rect 9738 12531 9760 12557
rect 9760 12531 9766 12557
rect 9686 12530 9714 12531
rect 9738 12530 9766 12531
rect 9790 12530 9818 12558
rect 9842 12557 9870 12558
rect 9894 12557 9922 12558
rect 9842 12531 9848 12557
rect 9848 12531 9870 12557
rect 9894 12531 9910 12557
rect 9910 12531 9922 12557
rect 9842 12530 9870 12531
rect 9894 12530 9922 12531
rect 9946 12557 9974 12558
rect 9946 12531 9972 12557
rect 9972 12531 9974 12557
rect 9946 12530 9974 12531
rect 9998 12557 10026 12558
rect 9998 12531 10008 12557
rect 10008 12531 10026 12557
rect 9998 12530 10026 12531
rect 9534 12334 9562 12362
rect 10430 13537 10458 13538
rect 10430 13511 10431 13537
rect 10431 13511 10457 13537
rect 10457 13511 10458 13537
rect 10430 13510 10458 13511
rect 10766 13510 10794 13538
rect 10094 12361 10122 12362
rect 10094 12335 10095 12361
rect 10095 12335 10121 12361
rect 10121 12335 10122 12361
rect 10094 12334 10122 12335
rect 8974 11969 9002 11970
rect 8974 11943 8975 11969
rect 8975 11943 9001 11969
rect 9001 11943 9002 11969
rect 8974 11942 9002 11943
rect 9702 11969 9730 11970
rect 9702 11943 9703 11969
rect 9703 11943 9729 11969
rect 9729 11943 9730 11969
rect 9702 11942 9730 11943
rect 11270 12361 11298 12362
rect 11270 12335 11271 12361
rect 11271 12335 11297 12361
rect 11297 12335 11298 12361
rect 11270 12334 11298 12335
rect 10374 11969 10402 11970
rect 10374 11943 10375 11969
rect 10375 11943 10401 11969
rect 10401 11943 10402 11969
rect 10374 11942 10402 11943
rect 9478 11774 9506 11802
rect 9582 11773 9610 11774
rect 9582 11747 9600 11773
rect 9600 11747 9610 11773
rect 9582 11746 9610 11747
rect 9634 11773 9662 11774
rect 9634 11747 9636 11773
rect 9636 11747 9662 11773
rect 9634 11746 9662 11747
rect 9686 11773 9714 11774
rect 9738 11773 9766 11774
rect 9686 11747 9698 11773
rect 9698 11747 9714 11773
rect 9738 11747 9760 11773
rect 9760 11747 9766 11773
rect 9686 11746 9714 11747
rect 9738 11746 9766 11747
rect 9790 11746 9818 11774
rect 9842 11773 9870 11774
rect 9894 11773 9922 11774
rect 9842 11747 9848 11773
rect 9848 11747 9870 11773
rect 9894 11747 9910 11773
rect 9910 11747 9922 11773
rect 9842 11746 9870 11747
rect 9894 11746 9922 11747
rect 9946 11773 9974 11774
rect 9946 11747 9972 11773
rect 9972 11747 9974 11773
rect 9946 11746 9974 11747
rect 9998 11773 10026 11774
rect 9998 11747 10008 11773
rect 10008 11747 10026 11773
rect 9998 11746 10026 11747
rect 8974 11129 9002 11130
rect 8974 11103 8975 11129
rect 8975 11103 9001 11129
rect 9001 11103 9002 11129
rect 8974 11102 9002 11103
rect 13398 18214 13426 18242
rect 12082 17653 12110 17654
rect 12082 17627 12100 17653
rect 12100 17627 12110 17653
rect 12082 17626 12110 17627
rect 12134 17653 12162 17654
rect 12134 17627 12136 17653
rect 12136 17627 12162 17653
rect 12134 17626 12162 17627
rect 12186 17653 12214 17654
rect 12238 17653 12266 17654
rect 12186 17627 12198 17653
rect 12198 17627 12214 17653
rect 12238 17627 12260 17653
rect 12260 17627 12266 17653
rect 12186 17626 12214 17627
rect 12238 17626 12266 17627
rect 12290 17626 12318 17654
rect 12342 17653 12370 17654
rect 12394 17653 12422 17654
rect 12342 17627 12348 17653
rect 12348 17627 12370 17653
rect 12394 17627 12410 17653
rect 12410 17627 12422 17653
rect 12342 17626 12370 17627
rect 12394 17626 12422 17627
rect 12446 17653 12474 17654
rect 12446 17627 12472 17653
rect 12472 17627 12474 17653
rect 12446 17626 12474 17627
rect 12498 17653 12526 17654
rect 12498 17627 12508 17653
rect 12508 17627 12526 17653
rect 12498 17626 12526 17627
rect 12614 17318 12642 17346
rect 14630 18241 14658 18242
rect 14630 18215 14631 18241
rect 14631 18215 14657 18241
rect 14657 18215 14658 18241
rect 14630 18214 14658 18215
rect 15078 18214 15106 18242
rect 14582 18045 14610 18046
rect 14582 18019 14600 18045
rect 14600 18019 14610 18045
rect 14582 18018 14610 18019
rect 14634 18045 14662 18046
rect 14634 18019 14636 18045
rect 14636 18019 14662 18045
rect 14634 18018 14662 18019
rect 14686 18045 14714 18046
rect 14738 18045 14766 18046
rect 14686 18019 14698 18045
rect 14698 18019 14714 18045
rect 14738 18019 14760 18045
rect 14760 18019 14766 18045
rect 14686 18018 14714 18019
rect 14738 18018 14766 18019
rect 14790 18018 14818 18046
rect 14842 18045 14870 18046
rect 14894 18045 14922 18046
rect 14842 18019 14848 18045
rect 14848 18019 14870 18045
rect 14894 18019 14910 18045
rect 14910 18019 14922 18045
rect 14842 18018 14870 18019
rect 14894 18018 14922 18019
rect 14946 18045 14974 18046
rect 14946 18019 14972 18045
rect 14972 18019 14974 18045
rect 14946 18018 14974 18019
rect 14998 18045 15026 18046
rect 14998 18019 15008 18045
rect 15008 18019 15026 18045
rect 14998 18018 15026 18019
rect 14238 17822 14266 17850
rect 14574 17849 14602 17850
rect 14574 17823 14575 17849
rect 14575 17823 14601 17849
rect 14601 17823 14602 17849
rect 14574 17822 14602 17823
rect 12082 16869 12110 16870
rect 12082 16843 12100 16869
rect 12100 16843 12110 16869
rect 12082 16842 12110 16843
rect 12134 16869 12162 16870
rect 12134 16843 12136 16869
rect 12136 16843 12162 16869
rect 12134 16842 12162 16843
rect 12186 16869 12214 16870
rect 12238 16869 12266 16870
rect 12186 16843 12198 16869
rect 12198 16843 12214 16869
rect 12238 16843 12260 16869
rect 12260 16843 12266 16869
rect 12186 16842 12214 16843
rect 12238 16842 12266 16843
rect 12290 16842 12318 16870
rect 12342 16869 12370 16870
rect 12394 16869 12422 16870
rect 12342 16843 12348 16869
rect 12348 16843 12370 16869
rect 12394 16843 12410 16869
rect 12410 16843 12422 16869
rect 12342 16842 12370 16843
rect 12394 16842 12422 16843
rect 12446 16869 12474 16870
rect 12446 16843 12472 16869
rect 12472 16843 12474 16869
rect 12446 16842 12474 16843
rect 12498 16869 12526 16870
rect 12498 16843 12508 16869
rect 12508 16843 12526 16869
rect 12498 16842 12526 16843
rect 11830 16646 11858 16674
rect 12222 16673 12250 16674
rect 12222 16647 12223 16673
rect 12223 16647 12249 16673
rect 12249 16647 12250 16673
rect 12222 16646 12250 16647
rect 12446 16673 12474 16674
rect 12446 16647 12447 16673
rect 12447 16647 12473 16673
rect 12473 16647 12474 16673
rect 12446 16646 12474 16647
rect 11830 16281 11858 16282
rect 11830 16255 11831 16281
rect 11831 16255 11857 16281
rect 11857 16255 11858 16281
rect 11830 16254 11858 16255
rect 11942 16281 11970 16282
rect 11942 16255 11943 16281
rect 11943 16255 11969 16281
rect 11969 16255 11970 16281
rect 11942 16254 11970 16255
rect 12082 16085 12110 16086
rect 12082 16059 12100 16085
rect 12100 16059 12110 16085
rect 12082 16058 12110 16059
rect 12134 16085 12162 16086
rect 12134 16059 12136 16085
rect 12136 16059 12162 16085
rect 12134 16058 12162 16059
rect 12186 16085 12214 16086
rect 12238 16085 12266 16086
rect 12186 16059 12198 16085
rect 12198 16059 12214 16085
rect 12238 16059 12260 16085
rect 12260 16059 12266 16085
rect 12186 16058 12214 16059
rect 12238 16058 12266 16059
rect 12290 16058 12318 16086
rect 12342 16085 12370 16086
rect 12394 16085 12422 16086
rect 12342 16059 12348 16085
rect 12348 16059 12370 16085
rect 12394 16059 12410 16085
rect 12410 16059 12422 16085
rect 12342 16058 12370 16059
rect 12394 16058 12422 16059
rect 12446 16085 12474 16086
rect 12446 16059 12472 16085
rect 12472 16059 12474 16085
rect 12446 16058 12474 16059
rect 12498 16085 12526 16086
rect 12498 16059 12508 16085
rect 12508 16059 12526 16085
rect 12498 16058 12526 16059
rect 11830 15974 11858 16002
rect 12222 15974 12250 16002
rect 12446 15974 12474 16002
rect 13286 15918 13314 15946
rect 12082 15301 12110 15302
rect 12082 15275 12100 15301
rect 12100 15275 12110 15301
rect 12082 15274 12110 15275
rect 12134 15301 12162 15302
rect 12134 15275 12136 15301
rect 12136 15275 12162 15301
rect 12134 15274 12162 15275
rect 12186 15301 12214 15302
rect 12238 15301 12266 15302
rect 12186 15275 12198 15301
rect 12198 15275 12214 15301
rect 12238 15275 12260 15301
rect 12260 15275 12266 15301
rect 12186 15274 12214 15275
rect 12238 15274 12266 15275
rect 12290 15274 12318 15302
rect 12342 15301 12370 15302
rect 12394 15301 12422 15302
rect 12342 15275 12348 15301
rect 12348 15275 12370 15301
rect 12394 15275 12410 15301
rect 12410 15275 12422 15301
rect 12342 15274 12370 15275
rect 12394 15274 12422 15275
rect 12446 15301 12474 15302
rect 12446 15275 12472 15301
rect 12472 15275 12474 15301
rect 12446 15274 12474 15275
rect 12498 15301 12526 15302
rect 12498 15275 12508 15301
rect 12508 15275 12526 15301
rect 12498 15274 12526 15275
rect 12082 14517 12110 14518
rect 12082 14491 12100 14517
rect 12100 14491 12110 14517
rect 12082 14490 12110 14491
rect 12134 14517 12162 14518
rect 12134 14491 12136 14517
rect 12136 14491 12162 14517
rect 12134 14490 12162 14491
rect 12186 14517 12214 14518
rect 12238 14517 12266 14518
rect 12186 14491 12198 14517
rect 12198 14491 12214 14517
rect 12238 14491 12260 14517
rect 12260 14491 12266 14517
rect 12186 14490 12214 14491
rect 12238 14490 12266 14491
rect 12290 14490 12318 14518
rect 12342 14517 12370 14518
rect 12394 14517 12422 14518
rect 12342 14491 12348 14517
rect 12348 14491 12370 14517
rect 12394 14491 12410 14517
rect 12410 14491 12422 14517
rect 12342 14490 12370 14491
rect 12394 14490 12422 14491
rect 12446 14517 12474 14518
rect 12446 14491 12472 14517
rect 12472 14491 12474 14517
rect 12446 14490 12474 14491
rect 12498 14517 12526 14518
rect 12498 14491 12508 14517
rect 12508 14491 12526 14517
rect 12498 14490 12526 14491
rect 15806 17822 15834 17850
rect 14582 17261 14610 17262
rect 14582 17235 14600 17261
rect 14600 17235 14610 17261
rect 14582 17234 14610 17235
rect 14634 17261 14662 17262
rect 14634 17235 14636 17261
rect 14636 17235 14662 17261
rect 14634 17234 14662 17235
rect 14686 17261 14714 17262
rect 14738 17261 14766 17262
rect 14686 17235 14698 17261
rect 14698 17235 14714 17261
rect 14738 17235 14760 17261
rect 14760 17235 14766 17261
rect 14686 17234 14714 17235
rect 14738 17234 14766 17235
rect 14790 17234 14818 17262
rect 14842 17261 14870 17262
rect 14894 17261 14922 17262
rect 14842 17235 14848 17261
rect 14848 17235 14870 17261
rect 14894 17235 14910 17261
rect 14910 17235 14922 17261
rect 14842 17234 14870 17235
rect 14894 17234 14922 17235
rect 14946 17261 14974 17262
rect 14946 17235 14972 17261
rect 14972 17235 14974 17261
rect 14946 17234 14974 17235
rect 14998 17261 15026 17262
rect 14998 17235 15008 17261
rect 15008 17235 15026 17261
rect 14998 17234 15026 17235
rect 14238 16673 14266 16674
rect 14238 16647 14239 16673
rect 14239 16647 14265 16673
rect 14265 16647 14266 16673
rect 14238 16646 14266 16647
rect 13734 15918 13762 15946
rect 17082 17653 17110 17654
rect 17082 17627 17100 17653
rect 17100 17627 17110 17653
rect 17082 17626 17110 17627
rect 17134 17653 17162 17654
rect 17134 17627 17136 17653
rect 17136 17627 17162 17653
rect 17134 17626 17162 17627
rect 17186 17653 17214 17654
rect 17238 17653 17266 17654
rect 17186 17627 17198 17653
rect 17198 17627 17214 17653
rect 17238 17627 17260 17653
rect 17260 17627 17266 17653
rect 17186 17626 17214 17627
rect 17238 17626 17266 17627
rect 17290 17626 17318 17654
rect 17342 17653 17370 17654
rect 17394 17653 17422 17654
rect 17342 17627 17348 17653
rect 17348 17627 17370 17653
rect 17394 17627 17410 17653
rect 17410 17627 17422 17653
rect 17342 17626 17370 17627
rect 17394 17626 17422 17627
rect 17446 17653 17474 17654
rect 17446 17627 17472 17653
rect 17472 17627 17474 17653
rect 17446 17626 17474 17627
rect 17498 17653 17526 17654
rect 17498 17627 17508 17653
rect 17508 17627 17526 17653
rect 17498 17626 17526 17627
rect 14582 16477 14610 16478
rect 14582 16451 14600 16477
rect 14600 16451 14610 16477
rect 14582 16450 14610 16451
rect 14634 16477 14662 16478
rect 14634 16451 14636 16477
rect 14636 16451 14662 16477
rect 14634 16450 14662 16451
rect 14686 16477 14714 16478
rect 14738 16477 14766 16478
rect 14686 16451 14698 16477
rect 14698 16451 14714 16477
rect 14738 16451 14760 16477
rect 14760 16451 14766 16477
rect 14686 16450 14714 16451
rect 14738 16450 14766 16451
rect 14790 16450 14818 16478
rect 14842 16477 14870 16478
rect 14894 16477 14922 16478
rect 14842 16451 14848 16477
rect 14848 16451 14870 16477
rect 14894 16451 14910 16477
rect 14910 16451 14922 16477
rect 14842 16450 14870 16451
rect 14894 16450 14922 16451
rect 14946 16477 14974 16478
rect 14946 16451 14972 16477
rect 14972 16451 14974 16477
rect 14946 16450 14974 16451
rect 14998 16477 15026 16478
rect 14998 16451 15008 16477
rect 15008 16451 15026 16477
rect 14998 16450 15026 16451
rect 15974 16142 16002 16170
rect 16758 16673 16786 16674
rect 16758 16647 16759 16673
rect 16759 16647 16785 16673
rect 16785 16647 16786 16673
rect 16758 16646 16786 16647
rect 16254 16254 16282 16282
rect 14582 15693 14610 15694
rect 14582 15667 14600 15693
rect 14600 15667 14610 15693
rect 14582 15666 14610 15667
rect 14634 15693 14662 15694
rect 14634 15667 14636 15693
rect 14636 15667 14662 15693
rect 14634 15666 14662 15667
rect 14686 15693 14714 15694
rect 14738 15693 14766 15694
rect 14686 15667 14698 15693
rect 14698 15667 14714 15693
rect 14738 15667 14760 15693
rect 14760 15667 14766 15693
rect 14686 15666 14714 15667
rect 14738 15666 14766 15667
rect 14790 15666 14818 15694
rect 14842 15693 14870 15694
rect 14894 15693 14922 15694
rect 14842 15667 14848 15693
rect 14848 15667 14870 15693
rect 14894 15667 14910 15693
rect 14910 15667 14922 15693
rect 14842 15666 14870 15667
rect 14894 15666 14922 15667
rect 14946 15693 14974 15694
rect 14946 15667 14972 15693
rect 14972 15667 14974 15693
rect 14946 15666 14974 15667
rect 14998 15693 15026 15694
rect 14998 15667 15008 15693
rect 15008 15667 15026 15693
rect 14998 15666 15026 15667
rect 16310 16142 16338 16170
rect 17082 16869 17110 16870
rect 17082 16843 17100 16869
rect 17100 16843 17110 16869
rect 17082 16842 17110 16843
rect 17134 16869 17162 16870
rect 17134 16843 17136 16869
rect 17136 16843 17162 16869
rect 17134 16842 17162 16843
rect 17186 16869 17214 16870
rect 17238 16869 17266 16870
rect 17186 16843 17198 16869
rect 17198 16843 17214 16869
rect 17238 16843 17260 16869
rect 17260 16843 17266 16869
rect 17186 16842 17214 16843
rect 17238 16842 17266 16843
rect 17290 16842 17318 16870
rect 17342 16869 17370 16870
rect 17394 16869 17422 16870
rect 17342 16843 17348 16869
rect 17348 16843 17370 16869
rect 17394 16843 17410 16869
rect 17410 16843 17422 16869
rect 17342 16842 17370 16843
rect 17394 16842 17422 16843
rect 17446 16869 17474 16870
rect 17446 16843 17472 16869
rect 17472 16843 17474 16869
rect 17446 16842 17474 16843
rect 17498 16869 17526 16870
rect 17498 16843 17508 16869
rect 17508 16843 17526 16869
rect 17498 16842 17526 16843
rect 16926 16673 16954 16674
rect 16926 16647 16927 16673
rect 16927 16647 16953 16673
rect 16953 16647 16954 16673
rect 16926 16646 16954 16647
rect 16814 16281 16842 16282
rect 16814 16255 16815 16281
rect 16815 16255 16841 16281
rect 16841 16255 16842 16281
rect 16814 16254 16842 16255
rect 16814 16142 16842 16170
rect 11998 13902 12026 13930
rect 12446 13929 12474 13930
rect 12446 13903 12447 13929
rect 12447 13903 12473 13929
rect 12473 13903 12474 13929
rect 12446 13902 12474 13903
rect 12082 13733 12110 13734
rect 12082 13707 12100 13733
rect 12100 13707 12110 13733
rect 12082 13706 12110 13707
rect 12134 13733 12162 13734
rect 12134 13707 12136 13733
rect 12136 13707 12162 13733
rect 12134 13706 12162 13707
rect 12186 13733 12214 13734
rect 12238 13733 12266 13734
rect 12186 13707 12198 13733
rect 12198 13707 12214 13733
rect 12238 13707 12260 13733
rect 12260 13707 12266 13733
rect 12186 13706 12214 13707
rect 12238 13706 12266 13707
rect 12290 13706 12318 13734
rect 12342 13733 12370 13734
rect 12394 13733 12422 13734
rect 12342 13707 12348 13733
rect 12348 13707 12370 13733
rect 12394 13707 12410 13733
rect 12410 13707 12422 13733
rect 12342 13706 12370 13707
rect 12394 13706 12422 13707
rect 12446 13733 12474 13734
rect 12446 13707 12472 13733
rect 12472 13707 12474 13733
rect 12446 13706 12474 13707
rect 12498 13733 12526 13734
rect 12498 13707 12508 13733
rect 12508 13707 12526 13733
rect 12498 13706 12526 13707
rect 12222 13510 12250 13538
rect 12950 13537 12978 13538
rect 12950 13511 12951 13537
rect 12951 13511 12977 13537
rect 12977 13511 12978 13537
rect 12950 13510 12978 13511
rect 14582 14909 14610 14910
rect 14582 14883 14600 14909
rect 14600 14883 14610 14909
rect 14582 14882 14610 14883
rect 14634 14909 14662 14910
rect 14634 14883 14636 14909
rect 14636 14883 14662 14909
rect 14634 14882 14662 14883
rect 14686 14909 14714 14910
rect 14738 14909 14766 14910
rect 14686 14883 14698 14909
rect 14698 14883 14714 14909
rect 14738 14883 14760 14909
rect 14760 14883 14766 14909
rect 14686 14882 14714 14883
rect 14738 14882 14766 14883
rect 14790 14882 14818 14910
rect 14842 14909 14870 14910
rect 14894 14909 14922 14910
rect 14842 14883 14848 14909
rect 14848 14883 14870 14909
rect 14894 14883 14910 14909
rect 14910 14883 14922 14909
rect 14842 14882 14870 14883
rect 14894 14882 14922 14883
rect 14946 14909 14974 14910
rect 14946 14883 14972 14909
rect 14972 14883 14974 14909
rect 14946 14882 14974 14883
rect 14998 14909 15026 14910
rect 14998 14883 15008 14909
rect 15008 14883 15026 14909
rect 14998 14882 15026 14883
rect 15190 14294 15218 14322
rect 14582 14125 14610 14126
rect 14582 14099 14600 14125
rect 14600 14099 14610 14125
rect 14582 14098 14610 14099
rect 14634 14125 14662 14126
rect 14634 14099 14636 14125
rect 14636 14099 14662 14125
rect 14634 14098 14662 14099
rect 14686 14125 14714 14126
rect 14738 14125 14766 14126
rect 14686 14099 14698 14125
rect 14698 14099 14714 14125
rect 14738 14099 14760 14125
rect 14760 14099 14766 14125
rect 14686 14098 14714 14099
rect 14738 14098 14766 14099
rect 14790 14098 14818 14126
rect 14842 14125 14870 14126
rect 14894 14125 14922 14126
rect 14842 14099 14848 14125
rect 14848 14099 14870 14125
rect 14894 14099 14910 14125
rect 14910 14099 14922 14125
rect 14842 14098 14870 14099
rect 14894 14098 14922 14099
rect 14946 14125 14974 14126
rect 14946 14099 14972 14125
rect 14972 14099 14974 14125
rect 14946 14098 14974 14099
rect 14998 14125 15026 14126
rect 14998 14099 15008 14125
rect 15008 14099 15026 14125
rect 14998 14098 15026 14099
rect 13678 13510 13706 13538
rect 13230 13398 13258 13426
rect 14462 13902 14490 13930
rect 13734 13398 13762 13426
rect 13790 13454 13818 13482
rect 14126 13454 14154 13482
rect 14910 13929 14938 13930
rect 14910 13903 14911 13929
rect 14911 13903 14937 13929
rect 14937 13903 14938 13929
rect 14910 13902 14938 13903
rect 17082 16085 17110 16086
rect 17082 16059 17100 16085
rect 17100 16059 17110 16085
rect 17082 16058 17110 16059
rect 17134 16085 17162 16086
rect 17134 16059 17136 16085
rect 17136 16059 17162 16085
rect 17134 16058 17162 16059
rect 17186 16085 17214 16086
rect 17238 16085 17266 16086
rect 17186 16059 17198 16085
rect 17198 16059 17214 16085
rect 17238 16059 17260 16085
rect 17260 16059 17266 16085
rect 17186 16058 17214 16059
rect 17238 16058 17266 16059
rect 17290 16058 17318 16086
rect 17342 16085 17370 16086
rect 17394 16085 17422 16086
rect 17342 16059 17348 16085
rect 17348 16059 17370 16085
rect 17394 16059 17410 16085
rect 17410 16059 17422 16085
rect 17342 16058 17370 16059
rect 17394 16058 17422 16059
rect 17446 16085 17474 16086
rect 17446 16059 17472 16085
rect 17472 16059 17474 16085
rect 17446 16058 17474 16059
rect 17498 16085 17526 16086
rect 17498 16059 17508 16085
rect 17508 16059 17526 16085
rect 17498 16058 17526 16059
rect 16254 14321 16282 14322
rect 16254 14295 16255 14321
rect 16255 14295 16281 14321
rect 16281 14295 16282 14321
rect 16254 14294 16282 14295
rect 16310 15134 16338 15162
rect 15974 14265 16002 14266
rect 15974 14239 15975 14265
rect 15975 14239 16001 14265
rect 16001 14239 16002 14265
rect 15974 14238 16002 14239
rect 15974 13902 16002 13930
rect 14406 13510 14434 13538
rect 11774 12753 11802 12754
rect 11774 12727 11775 12753
rect 11775 12727 11801 12753
rect 11801 12727 11802 12753
rect 11774 12726 11802 12727
rect 11270 11942 11298 11970
rect 12082 12949 12110 12950
rect 12082 12923 12100 12949
rect 12100 12923 12110 12949
rect 12082 12922 12110 12923
rect 12134 12949 12162 12950
rect 12134 12923 12136 12949
rect 12136 12923 12162 12949
rect 12134 12922 12162 12923
rect 12186 12949 12214 12950
rect 12238 12949 12266 12950
rect 12186 12923 12198 12949
rect 12198 12923 12214 12949
rect 12238 12923 12260 12949
rect 12260 12923 12266 12949
rect 12186 12922 12214 12923
rect 12238 12922 12266 12923
rect 12290 12922 12318 12950
rect 12342 12949 12370 12950
rect 12394 12949 12422 12950
rect 12342 12923 12348 12949
rect 12348 12923 12370 12949
rect 12394 12923 12410 12949
rect 12410 12923 12422 12949
rect 12342 12922 12370 12923
rect 12394 12922 12422 12923
rect 12446 12949 12474 12950
rect 12446 12923 12472 12949
rect 12472 12923 12474 12949
rect 12446 12922 12474 12923
rect 12498 12949 12526 12950
rect 12498 12923 12508 12949
rect 12508 12923 12526 12949
rect 12498 12922 12526 12923
rect 14582 13341 14610 13342
rect 14582 13315 14600 13341
rect 14600 13315 14610 13341
rect 14582 13314 14610 13315
rect 14634 13341 14662 13342
rect 14634 13315 14636 13341
rect 14636 13315 14662 13341
rect 14634 13314 14662 13315
rect 14686 13341 14714 13342
rect 14738 13341 14766 13342
rect 14686 13315 14698 13341
rect 14698 13315 14714 13341
rect 14738 13315 14760 13341
rect 14760 13315 14766 13341
rect 14686 13314 14714 13315
rect 14738 13314 14766 13315
rect 14790 13314 14818 13342
rect 14842 13341 14870 13342
rect 14894 13341 14922 13342
rect 14842 13315 14848 13341
rect 14848 13315 14870 13341
rect 14894 13315 14910 13341
rect 14910 13315 14922 13341
rect 14842 13314 14870 13315
rect 14894 13314 14922 13315
rect 14946 13341 14974 13342
rect 14946 13315 14972 13341
rect 14972 13315 14974 13341
rect 14946 13314 14974 13315
rect 14998 13341 15026 13342
rect 14998 13315 15008 13341
rect 15008 13315 15026 13341
rect 14998 13314 15026 13315
rect 15134 13145 15162 13146
rect 15134 13119 15135 13145
rect 15135 13119 15161 13145
rect 15161 13119 15162 13145
rect 15134 13118 15162 13119
rect 13230 12753 13258 12754
rect 13230 12727 13231 12753
rect 13231 12727 13257 12753
rect 13257 12727 13258 12753
rect 13230 12726 13258 12727
rect 16366 14238 16394 14266
rect 17082 15301 17110 15302
rect 17082 15275 17100 15301
rect 17100 15275 17110 15301
rect 17082 15274 17110 15275
rect 17134 15301 17162 15302
rect 17134 15275 17136 15301
rect 17136 15275 17162 15301
rect 17134 15274 17162 15275
rect 17186 15301 17214 15302
rect 17238 15301 17266 15302
rect 17186 15275 17198 15301
rect 17198 15275 17214 15301
rect 17238 15275 17260 15301
rect 17260 15275 17266 15301
rect 17186 15274 17214 15275
rect 17238 15274 17266 15275
rect 17290 15274 17318 15302
rect 17342 15301 17370 15302
rect 17394 15301 17422 15302
rect 17342 15275 17348 15301
rect 17348 15275 17370 15301
rect 17394 15275 17410 15301
rect 17410 15275 17422 15301
rect 17342 15274 17370 15275
rect 17394 15274 17422 15275
rect 17446 15301 17474 15302
rect 17446 15275 17472 15301
rect 17472 15275 17474 15301
rect 17446 15274 17474 15275
rect 17498 15301 17526 15302
rect 17498 15275 17508 15301
rect 17508 15275 17526 15301
rect 17498 15274 17526 15275
rect 16926 15134 16954 15162
rect 16814 14294 16842 14322
rect 17082 14517 17110 14518
rect 17082 14491 17100 14517
rect 17100 14491 17110 14517
rect 17082 14490 17110 14491
rect 17134 14517 17162 14518
rect 17134 14491 17136 14517
rect 17136 14491 17162 14517
rect 17134 14490 17162 14491
rect 17186 14517 17214 14518
rect 17238 14517 17266 14518
rect 17186 14491 17198 14517
rect 17198 14491 17214 14517
rect 17238 14491 17260 14517
rect 17260 14491 17266 14517
rect 17186 14490 17214 14491
rect 17238 14490 17266 14491
rect 17290 14490 17318 14518
rect 17342 14517 17370 14518
rect 17394 14517 17422 14518
rect 17342 14491 17348 14517
rect 17348 14491 17370 14517
rect 17394 14491 17410 14517
rect 17410 14491 17422 14517
rect 17342 14490 17370 14491
rect 17394 14490 17422 14491
rect 17446 14517 17474 14518
rect 17446 14491 17472 14517
rect 17472 14491 17474 14517
rect 17446 14490 17474 14491
rect 17498 14517 17526 14518
rect 17498 14491 17508 14517
rect 17508 14491 17526 14517
rect 17498 14490 17526 14491
rect 16982 14238 17010 14266
rect 17430 14265 17458 14266
rect 17430 14239 17431 14265
rect 17431 14239 17457 14265
rect 17457 14239 17458 14265
rect 17430 14238 17458 14239
rect 17082 13733 17110 13734
rect 17082 13707 17100 13733
rect 17100 13707 17110 13733
rect 17082 13706 17110 13707
rect 17134 13733 17162 13734
rect 17134 13707 17136 13733
rect 17136 13707 17162 13733
rect 17134 13706 17162 13707
rect 17186 13733 17214 13734
rect 17238 13733 17266 13734
rect 17186 13707 17198 13733
rect 17198 13707 17214 13733
rect 17238 13707 17260 13733
rect 17260 13707 17266 13733
rect 17186 13706 17214 13707
rect 17238 13706 17266 13707
rect 17290 13706 17318 13734
rect 17342 13733 17370 13734
rect 17394 13733 17422 13734
rect 17342 13707 17348 13733
rect 17348 13707 17370 13733
rect 17394 13707 17410 13733
rect 17410 13707 17422 13733
rect 17342 13706 17370 13707
rect 17394 13706 17422 13707
rect 17446 13733 17474 13734
rect 17446 13707 17472 13733
rect 17472 13707 17474 13733
rect 17446 13706 17474 13707
rect 17498 13733 17526 13734
rect 17498 13707 17508 13733
rect 17508 13707 17526 13733
rect 17498 13706 17526 13707
rect 16814 13426 16842 13454
rect 15470 13118 15498 13146
rect 15750 13118 15778 13146
rect 14582 12557 14610 12558
rect 14582 12531 14600 12557
rect 14600 12531 14610 12557
rect 14582 12530 14610 12531
rect 14634 12557 14662 12558
rect 14634 12531 14636 12557
rect 14636 12531 14662 12557
rect 14634 12530 14662 12531
rect 14686 12557 14714 12558
rect 14738 12557 14766 12558
rect 14686 12531 14698 12557
rect 14698 12531 14714 12557
rect 14738 12531 14760 12557
rect 14760 12531 14766 12557
rect 14686 12530 14714 12531
rect 14738 12530 14766 12531
rect 14790 12530 14818 12558
rect 14842 12557 14870 12558
rect 14894 12557 14922 12558
rect 14842 12531 14848 12557
rect 14848 12531 14870 12557
rect 14894 12531 14910 12557
rect 14910 12531 14922 12557
rect 14842 12530 14870 12531
rect 14894 12530 14922 12531
rect 14946 12557 14974 12558
rect 14946 12531 14972 12557
rect 14972 12531 14974 12557
rect 14946 12530 14974 12531
rect 14998 12557 15026 12558
rect 14998 12531 15008 12557
rect 15008 12531 15026 12557
rect 14998 12530 15026 12531
rect 11718 11942 11746 11970
rect 12082 12165 12110 12166
rect 12082 12139 12100 12165
rect 12100 12139 12110 12165
rect 12082 12138 12110 12139
rect 12134 12165 12162 12166
rect 12134 12139 12136 12165
rect 12136 12139 12162 12165
rect 12134 12138 12162 12139
rect 12186 12165 12214 12166
rect 12238 12165 12266 12166
rect 12186 12139 12198 12165
rect 12198 12139 12214 12165
rect 12238 12139 12260 12165
rect 12260 12139 12266 12165
rect 12186 12138 12214 12139
rect 12238 12138 12266 12139
rect 12290 12138 12318 12166
rect 12342 12165 12370 12166
rect 12394 12165 12422 12166
rect 12342 12139 12348 12165
rect 12348 12139 12370 12165
rect 12394 12139 12410 12165
rect 12410 12139 12422 12165
rect 12342 12138 12370 12139
rect 12394 12138 12422 12139
rect 12446 12165 12474 12166
rect 12446 12139 12472 12165
rect 12472 12139 12474 12165
rect 12446 12138 12474 12139
rect 12498 12165 12526 12166
rect 12498 12139 12508 12165
rect 12508 12139 12526 12165
rect 12498 12138 12526 12139
rect 10374 11129 10402 11130
rect 10374 11103 10375 11129
rect 10375 11103 10401 11129
rect 10401 11103 10402 11129
rect 10374 11102 10402 11103
rect 9582 10989 9610 10990
rect 9582 10963 9600 10989
rect 9600 10963 9610 10989
rect 9582 10962 9610 10963
rect 9634 10989 9662 10990
rect 9634 10963 9636 10989
rect 9636 10963 9662 10989
rect 9634 10962 9662 10963
rect 9686 10989 9714 10990
rect 9738 10989 9766 10990
rect 9686 10963 9698 10989
rect 9698 10963 9714 10989
rect 9738 10963 9760 10989
rect 9760 10963 9766 10989
rect 9686 10962 9714 10963
rect 9738 10962 9766 10963
rect 9790 10962 9818 10990
rect 9842 10989 9870 10990
rect 9894 10989 9922 10990
rect 9842 10963 9848 10989
rect 9848 10963 9870 10989
rect 9894 10963 9910 10989
rect 9910 10963 9922 10989
rect 9842 10962 9870 10963
rect 9894 10962 9922 10963
rect 9946 10989 9974 10990
rect 9946 10963 9972 10989
rect 9972 10963 9974 10989
rect 9946 10962 9974 10963
rect 9998 10989 10026 10990
rect 9998 10963 10008 10989
rect 10008 10963 10026 10989
rect 9998 10962 10026 10963
rect 9582 10205 9610 10206
rect 9582 10179 9600 10205
rect 9600 10179 9610 10205
rect 9582 10178 9610 10179
rect 9634 10205 9662 10206
rect 9634 10179 9636 10205
rect 9636 10179 9662 10205
rect 9634 10178 9662 10179
rect 9686 10205 9714 10206
rect 9738 10205 9766 10206
rect 9686 10179 9698 10205
rect 9698 10179 9714 10205
rect 9738 10179 9760 10205
rect 9760 10179 9766 10205
rect 9686 10178 9714 10179
rect 9738 10178 9766 10179
rect 9790 10178 9818 10206
rect 9842 10205 9870 10206
rect 9894 10205 9922 10206
rect 9842 10179 9848 10205
rect 9848 10179 9870 10205
rect 9894 10179 9910 10205
rect 9910 10179 9922 10205
rect 9842 10178 9870 10179
rect 9894 10178 9922 10179
rect 9946 10205 9974 10206
rect 9946 10179 9972 10205
rect 9972 10179 9974 10205
rect 9946 10178 9974 10179
rect 9998 10205 10026 10206
rect 9998 10179 10008 10205
rect 10008 10179 10026 10205
rect 9998 10178 10026 10179
rect 12082 11381 12110 11382
rect 12082 11355 12100 11381
rect 12100 11355 12110 11381
rect 12082 11354 12110 11355
rect 12134 11381 12162 11382
rect 12134 11355 12136 11381
rect 12136 11355 12162 11381
rect 12134 11354 12162 11355
rect 12186 11381 12214 11382
rect 12238 11381 12266 11382
rect 12186 11355 12198 11381
rect 12198 11355 12214 11381
rect 12238 11355 12260 11381
rect 12260 11355 12266 11381
rect 12186 11354 12214 11355
rect 12238 11354 12266 11355
rect 12290 11354 12318 11382
rect 12342 11381 12370 11382
rect 12394 11381 12422 11382
rect 12342 11355 12348 11381
rect 12348 11355 12370 11381
rect 12394 11355 12410 11381
rect 12410 11355 12422 11381
rect 12342 11354 12370 11355
rect 12394 11354 12422 11355
rect 12446 11381 12474 11382
rect 12446 11355 12472 11381
rect 12472 11355 12474 11381
rect 12446 11354 12474 11355
rect 12498 11381 12526 11382
rect 12498 11355 12508 11381
rect 12508 11355 12526 11381
rect 12498 11354 12526 11355
rect 16030 12390 16058 12418
rect 16422 12417 16450 12418
rect 16422 12391 16423 12417
rect 16423 12391 16449 12417
rect 16449 12391 16450 12417
rect 16422 12390 16450 12391
rect 13230 11158 13258 11186
rect 13510 11185 13538 11186
rect 13510 11159 13511 11185
rect 13511 11159 13537 11185
rect 13537 11159 13538 11185
rect 13510 11158 13538 11159
rect 12082 10597 12110 10598
rect 12082 10571 12100 10597
rect 12100 10571 12110 10597
rect 12082 10570 12110 10571
rect 12134 10597 12162 10598
rect 12134 10571 12136 10597
rect 12136 10571 12162 10597
rect 12134 10570 12162 10571
rect 12186 10597 12214 10598
rect 12238 10597 12266 10598
rect 12186 10571 12198 10597
rect 12198 10571 12214 10597
rect 12238 10571 12260 10597
rect 12260 10571 12266 10597
rect 12186 10570 12214 10571
rect 12238 10570 12266 10571
rect 12290 10570 12318 10598
rect 12342 10597 12370 10598
rect 12394 10597 12422 10598
rect 12342 10571 12348 10597
rect 12348 10571 12370 10597
rect 12394 10571 12410 10597
rect 12410 10571 12422 10597
rect 12342 10570 12370 10571
rect 12394 10570 12422 10571
rect 12446 10597 12474 10598
rect 12446 10571 12472 10597
rect 12472 10571 12474 10597
rect 12446 10570 12474 10571
rect 12498 10597 12526 10598
rect 12498 10571 12508 10597
rect 12508 10571 12526 10597
rect 12498 10570 12526 10571
rect 9582 9421 9610 9422
rect 9582 9395 9600 9421
rect 9600 9395 9610 9421
rect 9582 9394 9610 9395
rect 9634 9421 9662 9422
rect 9634 9395 9636 9421
rect 9636 9395 9662 9421
rect 9634 9394 9662 9395
rect 9686 9421 9714 9422
rect 9738 9421 9766 9422
rect 9686 9395 9698 9421
rect 9698 9395 9714 9421
rect 9738 9395 9760 9421
rect 9760 9395 9766 9421
rect 9686 9394 9714 9395
rect 9738 9394 9766 9395
rect 9790 9394 9818 9422
rect 9842 9421 9870 9422
rect 9894 9421 9922 9422
rect 9842 9395 9848 9421
rect 9848 9395 9870 9421
rect 9894 9395 9910 9421
rect 9910 9395 9922 9421
rect 9842 9394 9870 9395
rect 9894 9394 9922 9395
rect 9946 9421 9974 9422
rect 9946 9395 9972 9421
rect 9972 9395 9974 9421
rect 9946 9394 9974 9395
rect 9998 9421 10026 9422
rect 9998 9395 10008 9421
rect 10008 9395 10026 9421
rect 9998 9394 10026 9395
rect 9478 9198 9506 9226
rect 9254 8414 9282 8442
rect 9254 7630 9282 7658
rect 8862 3430 8890 3458
rect 8974 4494 9002 4522
rect 9422 4102 9450 4130
rect 8974 3345 9002 3346
rect 8974 3319 8975 3345
rect 8975 3319 9001 3345
rect 9001 3319 9002 3345
rect 8974 3318 9002 3319
rect 7082 2757 7110 2758
rect 7082 2731 7100 2757
rect 7100 2731 7110 2757
rect 7082 2730 7110 2731
rect 7134 2757 7162 2758
rect 7134 2731 7136 2757
rect 7136 2731 7162 2757
rect 7134 2730 7162 2731
rect 7186 2757 7214 2758
rect 7238 2757 7266 2758
rect 7186 2731 7198 2757
rect 7198 2731 7214 2757
rect 7238 2731 7260 2757
rect 7260 2731 7266 2757
rect 7186 2730 7214 2731
rect 7238 2730 7266 2731
rect 7290 2730 7318 2758
rect 7342 2757 7370 2758
rect 7394 2757 7422 2758
rect 7342 2731 7348 2757
rect 7348 2731 7370 2757
rect 7394 2731 7410 2757
rect 7410 2731 7422 2757
rect 7342 2730 7370 2731
rect 7394 2730 7422 2731
rect 7446 2757 7474 2758
rect 7446 2731 7472 2757
rect 7472 2731 7474 2757
rect 7446 2730 7474 2731
rect 7498 2757 7526 2758
rect 7498 2731 7508 2757
rect 7508 2731 7526 2757
rect 7498 2730 7526 2731
rect 7294 2169 7322 2170
rect 7294 2143 7295 2169
rect 7295 2143 7321 2169
rect 7321 2143 7322 2169
rect 7294 2142 7322 2143
rect 7574 2142 7602 2170
rect 7082 1973 7110 1974
rect 7082 1947 7100 1973
rect 7100 1947 7110 1973
rect 7082 1946 7110 1947
rect 7134 1973 7162 1974
rect 7134 1947 7136 1973
rect 7136 1947 7162 1973
rect 7134 1946 7162 1947
rect 7186 1973 7214 1974
rect 7238 1973 7266 1974
rect 7186 1947 7198 1973
rect 7198 1947 7214 1973
rect 7238 1947 7260 1973
rect 7260 1947 7266 1973
rect 7186 1946 7214 1947
rect 7238 1946 7266 1947
rect 7290 1946 7318 1974
rect 7342 1973 7370 1974
rect 7394 1973 7422 1974
rect 7342 1947 7348 1973
rect 7348 1947 7370 1973
rect 7394 1947 7410 1973
rect 7410 1947 7422 1973
rect 7342 1946 7370 1947
rect 7394 1946 7422 1947
rect 7446 1973 7474 1974
rect 7446 1947 7472 1973
rect 7472 1947 7474 1973
rect 7446 1946 7474 1947
rect 7498 1973 7526 1974
rect 7498 1947 7508 1973
rect 7508 1947 7526 1973
rect 7498 1946 7526 1947
rect 7798 2142 7826 2170
rect 8470 2478 8498 2506
rect 8974 2505 9002 2506
rect 8974 2479 8975 2505
rect 8975 2479 9001 2505
rect 9001 2479 9002 2505
rect 8974 2478 9002 2479
rect 7574 1862 7602 1890
rect 8302 1862 8330 1890
rect 8134 1777 8162 1778
rect 8134 1751 8135 1777
rect 8135 1751 8161 1777
rect 8161 1751 8162 1777
rect 8134 1750 8162 1751
rect 9422 1862 9450 1890
rect 9814 9225 9842 9226
rect 9814 9199 9815 9225
rect 9815 9199 9841 9225
rect 9841 9199 9842 9225
rect 9814 9198 9842 9199
rect 9582 8637 9610 8638
rect 9582 8611 9600 8637
rect 9600 8611 9610 8637
rect 9582 8610 9610 8611
rect 9634 8637 9662 8638
rect 9634 8611 9636 8637
rect 9636 8611 9662 8637
rect 9634 8610 9662 8611
rect 9686 8637 9714 8638
rect 9738 8637 9766 8638
rect 9686 8611 9698 8637
rect 9698 8611 9714 8637
rect 9738 8611 9760 8637
rect 9760 8611 9766 8637
rect 9686 8610 9714 8611
rect 9738 8610 9766 8611
rect 9790 8610 9818 8638
rect 9842 8637 9870 8638
rect 9894 8637 9922 8638
rect 9842 8611 9848 8637
rect 9848 8611 9870 8637
rect 9894 8611 9910 8637
rect 9910 8611 9922 8637
rect 9842 8610 9870 8611
rect 9894 8610 9922 8611
rect 9946 8637 9974 8638
rect 9946 8611 9972 8637
rect 9972 8611 9974 8637
rect 9946 8610 9974 8611
rect 9998 8637 10026 8638
rect 9998 8611 10008 8637
rect 10008 8611 10026 8637
rect 9998 8610 10026 8611
rect 10262 8470 10290 8498
rect 9814 8441 9842 8442
rect 9814 8415 9815 8441
rect 9815 8415 9841 8441
rect 9841 8415 9842 8441
rect 9814 8414 9842 8415
rect 9582 7853 9610 7854
rect 9582 7827 9600 7853
rect 9600 7827 9610 7853
rect 9582 7826 9610 7827
rect 9634 7853 9662 7854
rect 9634 7827 9636 7853
rect 9636 7827 9662 7853
rect 9634 7826 9662 7827
rect 9686 7853 9714 7854
rect 9738 7853 9766 7854
rect 9686 7827 9698 7853
rect 9698 7827 9714 7853
rect 9738 7827 9760 7853
rect 9760 7827 9766 7853
rect 9686 7826 9714 7827
rect 9738 7826 9766 7827
rect 9790 7826 9818 7854
rect 9842 7853 9870 7854
rect 9894 7853 9922 7854
rect 9842 7827 9848 7853
rect 9848 7827 9870 7853
rect 9894 7827 9910 7853
rect 9910 7827 9922 7853
rect 9842 7826 9870 7827
rect 9894 7826 9922 7827
rect 9946 7853 9974 7854
rect 9946 7827 9972 7853
rect 9972 7827 9974 7853
rect 9946 7826 9974 7827
rect 9998 7853 10026 7854
rect 9998 7827 10008 7853
rect 10008 7827 10026 7853
rect 9998 7826 10026 7827
rect 9814 7657 9842 7658
rect 9814 7631 9815 7657
rect 9815 7631 9841 7657
rect 9841 7631 9842 7657
rect 9814 7630 9842 7631
rect 10206 7518 10234 7546
rect 9582 7069 9610 7070
rect 9582 7043 9600 7069
rect 9600 7043 9610 7069
rect 9582 7042 9610 7043
rect 9634 7069 9662 7070
rect 9634 7043 9636 7069
rect 9636 7043 9662 7069
rect 9634 7042 9662 7043
rect 9686 7069 9714 7070
rect 9738 7069 9766 7070
rect 9686 7043 9698 7069
rect 9698 7043 9714 7069
rect 9738 7043 9760 7069
rect 9760 7043 9766 7069
rect 9686 7042 9714 7043
rect 9738 7042 9766 7043
rect 9790 7042 9818 7070
rect 9842 7069 9870 7070
rect 9894 7069 9922 7070
rect 9842 7043 9848 7069
rect 9848 7043 9870 7069
rect 9894 7043 9910 7069
rect 9910 7043 9922 7069
rect 9842 7042 9870 7043
rect 9894 7042 9922 7043
rect 9946 7069 9974 7070
rect 9946 7043 9972 7069
rect 9972 7043 9974 7069
rect 9946 7042 9974 7043
rect 9998 7069 10026 7070
rect 9998 7043 10008 7069
rect 10008 7043 10026 7069
rect 9998 7042 10026 7043
rect 10206 6454 10234 6482
rect 10878 7574 10906 7602
rect 11886 9646 11914 9674
rect 12446 10009 12474 10010
rect 12446 9983 12447 10009
rect 12447 9983 12473 10009
rect 12473 9983 12474 10009
rect 12446 9982 12474 9983
rect 11550 8441 11578 8442
rect 11550 8415 11551 8441
rect 11551 8415 11577 8441
rect 11577 8415 11578 8441
rect 11550 8414 11578 8415
rect 12950 9982 12978 10010
rect 12082 9813 12110 9814
rect 12082 9787 12100 9813
rect 12100 9787 12110 9813
rect 12082 9786 12110 9787
rect 12134 9813 12162 9814
rect 12134 9787 12136 9813
rect 12136 9787 12162 9813
rect 12134 9786 12162 9787
rect 12186 9813 12214 9814
rect 12238 9813 12266 9814
rect 12186 9787 12198 9813
rect 12198 9787 12214 9813
rect 12238 9787 12260 9813
rect 12260 9787 12266 9813
rect 12186 9786 12214 9787
rect 12238 9786 12266 9787
rect 12290 9786 12318 9814
rect 12342 9813 12370 9814
rect 12394 9813 12422 9814
rect 12342 9787 12348 9813
rect 12348 9787 12370 9813
rect 12394 9787 12410 9813
rect 12410 9787 12422 9813
rect 12342 9786 12370 9787
rect 12394 9786 12422 9787
rect 12446 9813 12474 9814
rect 12446 9787 12472 9813
rect 12472 9787 12474 9813
rect 12446 9786 12474 9787
rect 12498 9813 12526 9814
rect 12498 9787 12508 9813
rect 12508 9787 12526 9813
rect 12498 9786 12526 9787
rect 12054 9646 12082 9674
rect 12950 9561 12978 9562
rect 12950 9535 12951 9561
rect 12951 9535 12977 9561
rect 12977 9535 12978 9561
rect 12950 9534 12978 9535
rect 13510 9646 13538 9674
rect 12082 9029 12110 9030
rect 12082 9003 12100 9029
rect 12100 9003 12110 9029
rect 12082 9002 12110 9003
rect 12134 9029 12162 9030
rect 12134 9003 12136 9029
rect 12136 9003 12162 9029
rect 12134 9002 12162 9003
rect 12186 9029 12214 9030
rect 12238 9029 12266 9030
rect 12186 9003 12198 9029
rect 12198 9003 12214 9029
rect 12238 9003 12260 9029
rect 12260 9003 12266 9029
rect 12186 9002 12214 9003
rect 12238 9002 12266 9003
rect 12290 9002 12318 9030
rect 12342 9029 12370 9030
rect 12394 9029 12422 9030
rect 12342 9003 12348 9029
rect 12348 9003 12370 9029
rect 12394 9003 12410 9029
rect 12410 9003 12422 9029
rect 12342 9002 12370 9003
rect 12394 9002 12422 9003
rect 12446 9029 12474 9030
rect 12446 9003 12472 9029
rect 12472 9003 12474 9029
rect 12446 9002 12474 9003
rect 12498 9029 12526 9030
rect 12498 9003 12508 9029
rect 12508 9003 12526 9029
rect 12498 9002 12526 9003
rect 11942 8358 11970 8386
rect 11998 8414 12026 8442
rect 13510 8833 13538 8834
rect 13510 8807 13511 8833
rect 13511 8807 13537 8833
rect 13537 8807 13538 8833
rect 13510 8806 13538 8807
rect 14582 11773 14610 11774
rect 14582 11747 14600 11773
rect 14600 11747 14610 11773
rect 14582 11746 14610 11747
rect 14634 11773 14662 11774
rect 14634 11747 14636 11773
rect 14636 11747 14662 11773
rect 14634 11746 14662 11747
rect 14686 11773 14714 11774
rect 14738 11773 14766 11774
rect 14686 11747 14698 11773
rect 14698 11747 14714 11773
rect 14738 11747 14760 11773
rect 14760 11747 14766 11773
rect 14686 11746 14714 11747
rect 14738 11746 14766 11747
rect 14790 11746 14818 11774
rect 14842 11773 14870 11774
rect 14894 11773 14922 11774
rect 14842 11747 14848 11773
rect 14848 11747 14870 11773
rect 14894 11747 14910 11773
rect 14910 11747 14922 11773
rect 14842 11746 14870 11747
rect 14894 11746 14922 11747
rect 14946 11773 14974 11774
rect 14946 11747 14972 11773
rect 14972 11747 14974 11773
rect 14946 11746 14974 11747
rect 14998 11773 15026 11774
rect 14998 11747 15008 11773
rect 15008 11747 15026 11773
rect 14998 11746 15026 11747
rect 15862 11969 15890 11970
rect 15862 11943 15863 11969
rect 15863 11943 15889 11969
rect 15889 11943 15890 11969
rect 15862 11942 15890 11943
rect 15078 11606 15106 11634
rect 14582 10989 14610 10990
rect 14582 10963 14600 10989
rect 14600 10963 14610 10989
rect 14582 10962 14610 10963
rect 14634 10989 14662 10990
rect 14634 10963 14636 10989
rect 14636 10963 14662 10989
rect 14634 10962 14662 10963
rect 14686 10989 14714 10990
rect 14738 10989 14766 10990
rect 14686 10963 14698 10989
rect 14698 10963 14714 10989
rect 14738 10963 14760 10989
rect 14760 10963 14766 10989
rect 14686 10962 14714 10963
rect 14738 10962 14766 10963
rect 14790 10962 14818 10990
rect 14842 10989 14870 10990
rect 14894 10989 14922 10990
rect 14842 10963 14848 10989
rect 14848 10963 14870 10989
rect 14894 10963 14910 10989
rect 14910 10963 14922 10989
rect 14842 10962 14870 10963
rect 14894 10962 14922 10963
rect 14946 10989 14974 10990
rect 14946 10963 14972 10989
rect 14972 10963 14974 10989
rect 14946 10962 14974 10963
rect 14998 10989 15026 10990
rect 14998 10963 15008 10989
rect 15008 10963 15026 10989
rect 14998 10962 15026 10963
rect 16198 11633 16226 11634
rect 16198 11607 16199 11633
rect 16199 11607 16225 11633
rect 16225 11607 16226 11633
rect 16198 11606 16226 11607
rect 16758 11606 16786 11634
rect 14582 10205 14610 10206
rect 14582 10179 14600 10205
rect 14600 10179 14610 10205
rect 14582 10178 14610 10179
rect 14634 10205 14662 10206
rect 14634 10179 14636 10205
rect 14636 10179 14662 10205
rect 14634 10178 14662 10179
rect 14686 10205 14714 10206
rect 14738 10205 14766 10206
rect 14686 10179 14698 10205
rect 14698 10179 14714 10205
rect 14738 10179 14760 10205
rect 14760 10179 14766 10205
rect 14686 10178 14714 10179
rect 14738 10178 14766 10179
rect 14790 10178 14818 10206
rect 14842 10205 14870 10206
rect 14894 10205 14922 10206
rect 14842 10179 14848 10205
rect 14848 10179 14870 10205
rect 14894 10179 14910 10205
rect 14910 10179 14922 10205
rect 14842 10178 14870 10179
rect 14894 10178 14922 10179
rect 14946 10205 14974 10206
rect 14946 10179 14972 10205
rect 14972 10179 14974 10205
rect 14946 10178 14974 10179
rect 14998 10205 15026 10206
rect 14998 10179 15008 10205
rect 15008 10179 15026 10205
rect 14998 10178 15026 10179
rect 16366 10401 16394 10402
rect 16366 10375 16367 10401
rect 16367 10375 16393 10401
rect 16393 10375 16394 10401
rect 16366 10374 16394 10375
rect 14406 9561 14434 9562
rect 14406 9535 14407 9561
rect 14407 9535 14433 9561
rect 14433 9535 14434 9561
rect 14406 9534 14434 9535
rect 14582 9421 14610 9422
rect 14582 9395 14600 9421
rect 14600 9395 14610 9421
rect 14582 9394 14610 9395
rect 14634 9421 14662 9422
rect 14634 9395 14636 9421
rect 14636 9395 14662 9421
rect 14634 9394 14662 9395
rect 14686 9421 14714 9422
rect 14738 9421 14766 9422
rect 14686 9395 14698 9421
rect 14698 9395 14714 9421
rect 14738 9395 14760 9421
rect 14760 9395 14766 9421
rect 14686 9394 14714 9395
rect 14738 9394 14766 9395
rect 14790 9394 14818 9422
rect 14842 9421 14870 9422
rect 14894 9421 14922 9422
rect 14842 9395 14848 9421
rect 14848 9395 14870 9421
rect 14894 9395 14910 9421
rect 14910 9395 14922 9421
rect 14842 9394 14870 9395
rect 14894 9394 14922 9395
rect 14946 9421 14974 9422
rect 14946 9395 14972 9421
rect 14972 9395 14974 9421
rect 14946 9394 14974 9395
rect 14998 9421 15026 9422
rect 14998 9395 15008 9421
rect 15008 9395 15026 9421
rect 14998 9394 15026 9395
rect 14070 8806 14098 8834
rect 12222 8358 12250 8386
rect 12082 8245 12110 8246
rect 12082 8219 12100 8245
rect 12100 8219 12110 8245
rect 12082 8218 12110 8219
rect 12134 8245 12162 8246
rect 12134 8219 12136 8245
rect 12136 8219 12162 8245
rect 12134 8218 12162 8219
rect 12186 8245 12214 8246
rect 12238 8245 12266 8246
rect 12186 8219 12198 8245
rect 12198 8219 12214 8245
rect 12238 8219 12260 8245
rect 12260 8219 12266 8245
rect 12186 8218 12214 8219
rect 12238 8218 12266 8219
rect 12290 8218 12318 8246
rect 12342 8245 12370 8246
rect 12394 8245 12422 8246
rect 12342 8219 12348 8245
rect 12348 8219 12370 8245
rect 12394 8219 12410 8245
rect 12410 8219 12422 8245
rect 12342 8218 12370 8219
rect 12394 8218 12422 8219
rect 12446 8245 12474 8246
rect 12446 8219 12472 8245
rect 12472 8219 12474 8245
rect 12446 8218 12474 8219
rect 12498 8245 12526 8246
rect 12498 8219 12508 8245
rect 12508 8219 12526 8245
rect 12498 8218 12526 8219
rect 12054 8049 12082 8050
rect 12054 8023 12055 8049
rect 12055 8023 12081 8049
rect 12081 8023 12082 8049
rect 12054 8022 12082 8023
rect 11774 7574 11802 7602
rect 11942 7574 11970 7602
rect 12446 7966 12474 7994
rect 13398 8049 13426 8050
rect 13398 8023 13399 8049
rect 13399 8023 13425 8049
rect 13425 8023 13426 8049
rect 13398 8022 13426 8023
rect 12222 7574 12250 7602
rect 9582 6285 9610 6286
rect 9582 6259 9600 6285
rect 9600 6259 9610 6285
rect 9582 6258 9610 6259
rect 9634 6285 9662 6286
rect 9634 6259 9636 6285
rect 9636 6259 9662 6285
rect 9634 6258 9662 6259
rect 9686 6285 9714 6286
rect 9738 6285 9766 6286
rect 9686 6259 9698 6285
rect 9698 6259 9714 6285
rect 9738 6259 9760 6285
rect 9760 6259 9766 6285
rect 9686 6258 9714 6259
rect 9738 6258 9766 6259
rect 9790 6258 9818 6286
rect 9842 6285 9870 6286
rect 9894 6285 9922 6286
rect 9842 6259 9848 6285
rect 9848 6259 9870 6285
rect 9894 6259 9910 6285
rect 9910 6259 9922 6285
rect 9842 6258 9870 6259
rect 9894 6258 9922 6259
rect 9946 6285 9974 6286
rect 9946 6259 9972 6285
rect 9972 6259 9974 6285
rect 9946 6258 9974 6259
rect 9998 6285 10026 6286
rect 9998 6259 10008 6285
rect 10008 6259 10026 6285
rect 9998 6258 10026 6259
rect 12082 7461 12110 7462
rect 12082 7435 12100 7461
rect 12100 7435 12110 7461
rect 12082 7434 12110 7435
rect 12134 7461 12162 7462
rect 12134 7435 12136 7461
rect 12136 7435 12162 7461
rect 12134 7434 12162 7435
rect 12186 7461 12214 7462
rect 12238 7461 12266 7462
rect 12186 7435 12198 7461
rect 12198 7435 12214 7461
rect 12238 7435 12260 7461
rect 12260 7435 12266 7461
rect 12186 7434 12214 7435
rect 12238 7434 12266 7435
rect 12290 7434 12318 7462
rect 12342 7461 12370 7462
rect 12394 7461 12422 7462
rect 12342 7435 12348 7461
rect 12348 7435 12370 7461
rect 12394 7435 12410 7461
rect 12410 7435 12422 7461
rect 12342 7434 12370 7435
rect 12394 7434 12422 7435
rect 12446 7461 12474 7462
rect 12446 7435 12472 7461
rect 12472 7435 12474 7461
rect 12446 7434 12474 7435
rect 12498 7461 12526 7462
rect 12498 7435 12508 7461
rect 12508 7435 12526 7461
rect 12498 7434 12526 7435
rect 9582 5501 9610 5502
rect 9582 5475 9600 5501
rect 9600 5475 9610 5501
rect 9582 5474 9610 5475
rect 9634 5501 9662 5502
rect 9634 5475 9636 5501
rect 9636 5475 9662 5501
rect 9634 5474 9662 5475
rect 9686 5501 9714 5502
rect 9738 5501 9766 5502
rect 9686 5475 9698 5501
rect 9698 5475 9714 5501
rect 9738 5475 9760 5501
rect 9760 5475 9766 5501
rect 9686 5474 9714 5475
rect 9738 5474 9766 5475
rect 9790 5474 9818 5502
rect 9842 5501 9870 5502
rect 9894 5501 9922 5502
rect 9842 5475 9848 5501
rect 9848 5475 9870 5501
rect 9894 5475 9910 5501
rect 9910 5475 9922 5501
rect 9842 5474 9870 5475
rect 9894 5474 9922 5475
rect 9946 5501 9974 5502
rect 9946 5475 9972 5501
rect 9972 5475 9974 5501
rect 9946 5474 9974 5475
rect 9998 5501 10026 5502
rect 9998 5475 10008 5501
rect 10008 5475 10026 5501
rect 9998 5474 10026 5475
rect 9582 4717 9610 4718
rect 9582 4691 9600 4717
rect 9600 4691 9610 4717
rect 9582 4690 9610 4691
rect 9634 4717 9662 4718
rect 9634 4691 9636 4717
rect 9636 4691 9662 4717
rect 9634 4690 9662 4691
rect 9686 4717 9714 4718
rect 9738 4717 9766 4718
rect 9686 4691 9698 4717
rect 9698 4691 9714 4717
rect 9738 4691 9760 4717
rect 9760 4691 9766 4717
rect 9686 4690 9714 4691
rect 9738 4690 9766 4691
rect 9790 4690 9818 4718
rect 9842 4717 9870 4718
rect 9894 4717 9922 4718
rect 9842 4691 9848 4717
rect 9848 4691 9870 4717
rect 9894 4691 9910 4717
rect 9910 4691 9922 4717
rect 9842 4690 9870 4691
rect 9894 4690 9922 4691
rect 9946 4717 9974 4718
rect 9946 4691 9972 4717
rect 9972 4691 9974 4717
rect 9946 4690 9974 4691
rect 9998 4717 10026 4718
rect 9998 4691 10008 4717
rect 10008 4691 10026 4717
rect 9998 4690 10026 4691
rect 9534 4129 9562 4130
rect 9534 4103 9535 4129
rect 9535 4103 9561 4129
rect 9561 4103 9562 4129
rect 9534 4102 9562 4103
rect 10038 4102 10066 4130
rect 9582 3933 9610 3934
rect 9582 3907 9600 3933
rect 9600 3907 9610 3933
rect 9582 3906 9610 3907
rect 9634 3933 9662 3934
rect 9634 3907 9636 3933
rect 9636 3907 9662 3933
rect 9634 3906 9662 3907
rect 9686 3933 9714 3934
rect 9738 3933 9766 3934
rect 9686 3907 9698 3933
rect 9698 3907 9714 3933
rect 9738 3907 9760 3933
rect 9760 3907 9766 3933
rect 9686 3906 9714 3907
rect 9738 3906 9766 3907
rect 9790 3906 9818 3934
rect 9842 3933 9870 3934
rect 9894 3933 9922 3934
rect 9842 3907 9848 3933
rect 9848 3907 9870 3933
rect 9894 3907 9910 3933
rect 9910 3907 9922 3933
rect 9842 3906 9870 3907
rect 9894 3906 9922 3907
rect 9946 3933 9974 3934
rect 9946 3907 9972 3933
rect 9972 3907 9974 3933
rect 9946 3906 9974 3907
rect 9998 3933 10026 3934
rect 9998 3907 10008 3933
rect 10008 3907 10026 3933
rect 9998 3906 10026 3907
rect 9534 3374 9562 3402
rect 10038 3374 10066 3402
rect 10262 3737 10290 3738
rect 10262 3711 10263 3737
rect 10263 3711 10289 3737
rect 10289 3711 10290 3737
rect 10262 3710 10290 3711
rect 9582 3149 9610 3150
rect 9582 3123 9600 3149
rect 9600 3123 9610 3149
rect 9582 3122 9610 3123
rect 9634 3149 9662 3150
rect 9634 3123 9636 3149
rect 9636 3123 9662 3149
rect 9634 3122 9662 3123
rect 9686 3149 9714 3150
rect 9738 3149 9766 3150
rect 9686 3123 9698 3149
rect 9698 3123 9714 3149
rect 9738 3123 9760 3149
rect 9760 3123 9766 3149
rect 9686 3122 9714 3123
rect 9738 3122 9766 3123
rect 9790 3122 9818 3150
rect 9842 3149 9870 3150
rect 9894 3149 9922 3150
rect 9842 3123 9848 3149
rect 9848 3123 9870 3149
rect 9894 3123 9910 3149
rect 9910 3123 9922 3149
rect 9842 3122 9870 3123
rect 9894 3122 9922 3123
rect 9946 3149 9974 3150
rect 9946 3123 9972 3149
rect 9972 3123 9974 3149
rect 9946 3122 9974 3123
rect 9998 3149 10026 3150
rect 9998 3123 10008 3149
rect 10008 3123 10026 3149
rect 9998 3122 10026 3123
rect 10318 6481 10346 6482
rect 10318 6455 10319 6481
rect 10319 6455 10345 6481
rect 10345 6455 10346 6481
rect 10318 6454 10346 6455
rect 11774 6873 11802 6874
rect 11774 6847 11775 6873
rect 11775 6847 11801 6873
rect 11801 6847 11802 6873
rect 11774 6846 11802 6847
rect 14582 8637 14610 8638
rect 14582 8611 14600 8637
rect 14600 8611 14610 8637
rect 14582 8610 14610 8611
rect 14634 8637 14662 8638
rect 14634 8611 14636 8637
rect 14636 8611 14662 8637
rect 14634 8610 14662 8611
rect 14686 8637 14714 8638
rect 14738 8637 14766 8638
rect 14686 8611 14698 8637
rect 14698 8611 14714 8637
rect 14738 8611 14760 8637
rect 14760 8611 14766 8637
rect 14686 8610 14714 8611
rect 14738 8610 14766 8611
rect 14790 8610 14818 8638
rect 14842 8637 14870 8638
rect 14894 8637 14922 8638
rect 14842 8611 14848 8637
rect 14848 8611 14870 8637
rect 14894 8611 14910 8637
rect 14910 8611 14922 8637
rect 14842 8610 14870 8611
rect 14894 8610 14922 8611
rect 14946 8637 14974 8638
rect 14946 8611 14972 8637
rect 14972 8611 14974 8637
rect 14946 8610 14974 8611
rect 14998 8637 15026 8638
rect 14998 8611 15008 8637
rect 15008 8611 15026 8637
rect 14998 8610 15026 8611
rect 14406 8414 14434 8442
rect 14966 8441 14994 8442
rect 14966 8415 14967 8441
rect 14967 8415 14993 8441
rect 14993 8415 14994 8441
rect 14966 8414 14994 8415
rect 15526 9142 15554 9170
rect 14182 7993 14210 7994
rect 14182 7967 14183 7993
rect 14183 7967 14209 7993
rect 14209 7967 14210 7993
rect 14182 7966 14210 7967
rect 14582 7853 14610 7854
rect 14582 7827 14600 7853
rect 14600 7827 14610 7853
rect 14582 7826 14610 7827
rect 14634 7853 14662 7854
rect 14634 7827 14636 7853
rect 14636 7827 14662 7853
rect 14634 7826 14662 7827
rect 14686 7853 14714 7854
rect 14738 7853 14766 7854
rect 14686 7827 14698 7853
rect 14698 7827 14714 7853
rect 14738 7827 14760 7853
rect 14760 7827 14766 7853
rect 14686 7826 14714 7827
rect 14738 7826 14766 7827
rect 14790 7826 14818 7854
rect 14842 7853 14870 7854
rect 14894 7853 14922 7854
rect 14842 7827 14848 7853
rect 14848 7827 14870 7853
rect 14894 7827 14910 7853
rect 14910 7827 14922 7853
rect 14842 7826 14870 7827
rect 14894 7826 14922 7827
rect 14946 7853 14974 7854
rect 14946 7827 14972 7853
rect 14972 7827 14974 7853
rect 14946 7826 14974 7827
rect 14998 7853 15026 7854
rect 14998 7827 15008 7853
rect 15008 7827 15026 7853
rect 14998 7826 15026 7827
rect 14070 7657 14098 7658
rect 14070 7631 14071 7657
rect 14071 7631 14097 7657
rect 14097 7631 14098 7657
rect 14070 7630 14098 7631
rect 11998 6873 12026 6874
rect 11998 6847 11999 6873
rect 11999 6847 12025 6873
rect 12025 6847 12026 6873
rect 11998 6846 12026 6847
rect 12222 6846 12250 6874
rect 14294 6873 14322 6874
rect 14294 6847 14295 6873
rect 14295 6847 14321 6873
rect 14321 6847 14322 6873
rect 14294 6846 14322 6847
rect 12082 6677 12110 6678
rect 12082 6651 12100 6677
rect 12100 6651 12110 6677
rect 12082 6650 12110 6651
rect 12134 6677 12162 6678
rect 12134 6651 12136 6677
rect 12136 6651 12162 6677
rect 12134 6650 12162 6651
rect 12186 6677 12214 6678
rect 12238 6677 12266 6678
rect 12186 6651 12198 6677
rect 12198 6651 12214 6677
rect 12238 6651 12260 6677
rect 12260 6651 12266 6677
rect 12186 6650 12214 6651
rect 12238 6650 12266 6651
rect 12290 6650 12318 6678
rect 12342 6677 12370 6678
rect 12394 6677 12422 6678
rect 12342 6651 12348 6677
rect 12348 6651 12370 6677
rect 12394 6651 12410 6677
rect 12410 6651 12422 6677
rect 12342 6650 12370 6651
rect 12394 6650 12422 6651
rect 12446 6677 12474 6678
rect 12446 6651 12472 6677
rect 12472 6651 12474 6677
rect 12446 6650 12474 6651
rect 12498 6677 12526 6678
rect 12498 6651 12508 6677
rect 12508 6651 12526 6677
rect 12498 6650 12526 6651
rect 11998 6454 12026 6482
rect 12334 6481 12362 6482
rect 12334 6455 12335 6481
rect 12335 6455 12361 6481
rect 12361 6455 12362 6481
rect 12334 6454 12362 6455
rect 12446 6089 12474 6090
rect 12446 6063 12447 6089
rect 12447 6063 12473 6089
rect 12473 6063 12474 6089
rect 12446 6062 12474 6063
rect 12950 6062 12978 6090
rect 10486 3737 10514 3738
rect 10486 3711 10487 3737
rect 10487 3711 10513 3737
rect 10513 3711 10514 3737
rect 10486 3710 10514 3711
rect 10318 3318 10346 3346
rect 10262 2505 10290 2506
rect 10262 2479 10263 2505
rect 10263 2479 10289 2505
rect 10289 2479 10290 2505
rect 10262 2478 10290 2479
rect 9582 2365 9610 2366
rect 9582 2339 9600 2365
rect 9600 2339 9610 2365
rect 9582 2338 9610 2339
rect 9634 2365 9662 2366
rect 9634 2339 9636 2365
rect 9636 2339 9662 2365
rect 9634 2338 9662 2339
rect 9686 2365 9714 2366
rect 9738 2365 9766 2366
rect 9686 2339 9698 2365
rect 9698 2339 9714 2365
rect 9738 2339 9760 2365
rect 9760 2339 9766 2365
rect 9686 2338 9714 2339
rect 9738 2338 9766 2339
rect 9790 2338 9818 2366
rect 9842 2365 9870 2366
rect 9894 2365 9922 2366
rect 9842 2339 9848 2365
rect 9848 2339 9870 2365
rect 9894 2339 9910 2365
rect 9910 2339 9922 2365
rect 9842 2338 9870 2339
rect 9894 2338 9922 2339
rect 9946 2365 9974 2366
rect 9946 2339 9972 2365
rect 9972 2339 9974 2365
rect 9946 2338 9974 2339
rect 9998 2365 10026 2366
rect 9998 2339 10008 2365
rect 10008 2339 10026 2365
rect 9998 2338 10026 2339
rect 10038 2169 10066 2170
rect 10038 2143 10039 2169
rect 10039 2143 10065 2169
rect 10065 2143 10066 2169
rect 10038 2142 10066 2143
rect 12082 5893 12110 5894
rect 12082 5867 12100 5893
rect 12100 5867 12110 5893
rect 12082 5866 12110 5867
rect 12134 5893 12162 5894
rect 12134 5867 12136 5893
rect 12136 5867 12162 5893
rect 12134 5866 12162 5867
rect 12186 5893 12214 5894
rect 12238 5893 12266 5894
rect 12186 5867 12198 5893
rect 12198 5867 12214 5893
rect 12238 5867 12260 5893
rect 12260 5867 12266 5893
rect 12186 5866 12214 5867
rect 12238 5866 12266 5867
rect 12290 5866 12318 5894
rect 12342 5893 12370 5894
rect 12394 5893 12422 5894
rect 12342 5867 12348 5893
rect 12348 5867 12370 5893
rect 12394 5867 12410 5893
rect 12410 5867 12422 5893
rect 12342 5866 12370 5867
rect 12394 5866 12422 5867
rect 12446 5893 12474 5894
rect 12446 5867 12472 5893
rect 12472 5867 12474 5893
rect 12446 5866 12474 5867
rect 12498 5893 12526 5894
rect 12498 5867 12508 5893
rect 12508 5867 12526 5893
rect 12498 5866 12526 5867
rect 12446 5305 12474 5306
rect 12446 5279 12447 5305
rect 12447 5279 12473 5305
rect 12473 5279 12474 5305
rect 12446 5278 12474 5279
rect 12950 5278 12978 5306
rect 12082 5109 12110 5110
rect 12082 5083 12100 5109
rect 12100 5083 12110 5109
rect 12082 5082 12110 5083
rect 12134 5109 12162 5110
rect 12134 5083 12136 5109
rect 12136 5083 12162 5109
rect 12134 5082 12162 5083
rect 12186 5109 12214 5110
rect 12238 5109 12266 5110
rect 12186 5083 12198 5109
rect 12198 5083 12214 5109
rect 12238 5083 12260 5109
rect 12260 5083 12266 5109
rect 12186 5082 12214 5083
rect 12238 5082 12266 5083
rect 12290 5082 12318 5110
rect 12342 5109 12370 5110
rect 12394 5109 12422 5110
rect 12342 5083 12348 5109
rect 12348 5083 12370 5109
rect 12394 5083 12410 5109
rect 12410 5083 12422 5109
rect 12342 5082 12370 5083
rect 12394 5082 12422 5083
rect 12446 5109 12474 5110
rect 12446 5083 12472 5109
rect 12472 5083 12474 5109
rect 12446 5082 12474 5083
rect 12498 5109 12526 5110
rect 12498 5083 12508 5109
rect 12508 5083 12526 5109
rect 12498 5082 12526 5083
rect 12950 4857 12978 4858
rect 12950 4831 12951 4857
rect 12951 4831 12977 4857
rect 12977 4831 12978 4857
rect 12950 4830 12978 4831
rect 12670 4606 12698 4634
rect 12446 4521 12474 4522
rect 12446 4495 12447 4521
rect 12447 4495 12473 4521
rect 12473 4495 12474 4521
rect 12446 4494 12474 4495
rect 12082 4325 12110 4326
rect 12082 4299 12100 4325
rect 12100 4299 12110 4325
rect 12082 4298 12110 4299
rect 12134 4325 12162 4326
rect 12134 4299 12136 4325
rect 12136 4299 12162 4325
rect 12134 4298 12162 4299
rect 12186 4325 12214 4326
rect 12238 4325 12266 4326
rect 12186 4299 12198 4325
rect 12198 4299 12214 4325
rect 12238 4299 12260 4325
rect 12260 4299 12266 4325
rect 12186 4298 12214 4299
rect 12238 4298 12266 4299
rect 12290 4298 12318 4326
rect 12342 4325 12370 4326
rect 12394 4325 12422 4326
rect 12342 4299 12348 4325
rect 12348 4299 12370 4325
rect 12394 4299 12410 4325
rect 12410 4299 12422 4325
rect 12342 4298 12370 4299
rect 12394 4298 12422 4299
rect 12446 4325 12474 4326
rect 12446 4299 12472 4325
rect 12472 4299 12474 4325
rect 12446 4298 12474 4299
rect 12498 4325 12526 4326
rect 12498 4299 12508 4325
rect 12508 4299 12526 4325
rect 12498 4298 12526 4299
rect 12446 3737 12474 3738
rect 12446 3711 12447 3737
rect 12447 3711 12473 3737
rect 12473 3711 12474 3737
rect 12446 3710 12474 3711
rect 12082 3541 12110 3542
rect 12082 3515 12100 3541
rect 12100 3515 12110 3541
rect 12082 3514 12110 3515
rect 12134 3541 12162 3542
rect 12134 3515 12136 3541
rect 12136 3515 12162 3541
rect 12134 3514 12162 3515
rect 12186 3541 12214 3542
rect 12238 3541 12266 3542
rect 12186 3515 12198 3541
rect 12198 3515 12214 3541
rect 12238 3515 12260 3541
rect 12260 3515 12266 3541
rect 12186 3514 12214 3515
rect 12238 3514 12266 3515
rect 12290 3514 12318 3542
rect 12342 3541 12370 3542
rect 12394 3541 12422 3542
rect 12342 3515 12348 3541
rect 12348 3515 12370 3541
rect 12394 3515 12410 3541
rect 12410 3515 12422 3541
rect 12342 3514 12370 3515
rect 12394 3514 12422 3515
rect 12446 3541 12474 3542
rect 12446 3515 12472 3541
rect 12472 3515 12474 3541
rect 12446 3514 12474 3515
rect 12498 3541 12526 3542
rect 12498 3515 12508 3541
rect 12508 3515 12526 3541
rect 12498 3514 12526 3515
rect 12054 3374 12082 3402
rect 12446 3009 12474 3010
rect 12446 2983 12447 3009
rect 12447 2983 12473 3009
rect 12473 2983 12474 3009
rect 12446 2982 12474 2983
rect 12082 2757 12110 2758
rect 12082 2731 12100 2757
rect 12100 2731 12110 2757
rect 12082 2730 12110 2731
rect 12134 2757 12162 2758
rect 12134 2731 12136 2757
rect 12136 2731 12162 2757
rect 12134 2730 12162 2731
rect 12186 2757 12214 2758
rect 12238 2757 12266 2758
rect 12186 2731 12198 2757
rect 12198 2731 12214 2757
rect 12238 2731 12260 2757
rect 12260 2731 12266 2757
rect 12186 2730 12214 2731
rect 12238 2730 12266 2731
rect 12290 2730 12318 2758
rect 12342 2757 12370 2758
rect 12394 2757 12422 2758
rect 12342 2731 12348 2757
rect 12348 2731 12370 2757
rect 12394 2731 12410 2757
rect 12410 2731 12422 2757
rect 12342 2730 12370 2731
rect 12394 2730 12422 2731
rect 12446 2757 12474 2758
rect 12446 2731 12472 2757
rect 12472 2731 12474 2757
rect 12446 2730 12474 2731
rect 12498 2757 12526 2758
rect 12498 2731 12508 2757
rect 12508 2731 12526 2757
rect 12498 2730 12526 2731
rect 11214 2142 11242 2170
rect 11998 2198 12026 2226
rect 12446 2225 12474 2226
rect 12446 2199 12447 2225
rect 12447 2199 12473 2225
rect 12473 2199 12474 2225
rect 12446 2198 12474 2199
rect 12082 1973 12110 1974
rect 12082 1947 12100 1973
rect 12100 1947 12110 1973
rect 12082 1946 12110 1947
rect 12134 1973 12162 1974
rect 12134 1947 12136 1973
rect 12136 1947 12162 1973
rect 12134 1946 12162 1947
rect 12186 1973 12214 1974
rect 12238 1973 12266 1974
rect 12186 1947 12198 1973
rect 12198 1947 12214 1973
rect 12238 1947 12260 1973
rect 12260 1947 12266 1973
rect 12186 1946 12214 1947
rect 12238 1946 12266 1947
rect 12290 1946 12318 1974
rect 12342 1973 12370 1974
rect 12394 1973 12422 1974
rect 12342 1947 12348 1973
rect 12348 1947 12370 1973
rect 12394 1947 12410 1973
rect 12410 1947 12422 1973
rect 12342 1946 12370 1947
rect 12394 1946 12422 1947
rect 12446 1973 12474 1974
rect 12446 1947 12472 1973
rect 12472 1947 12474 1973
rect 12446 1946 12474 1947
rect 12498 1973 12526 1974
rect 12498 1947 12508 1973
rect 12508 1947 12526 1973
rect 12498 1946 12526 1947
rect 9582 1581 9610 1582
rect 9582 1555 9600 1581
rect 9600 1555 9610 1581
rect 9582 1554 9610 1555
rect 9634 1581 9662 1582
rect 9634 1555 9636 1581
rect 9636 1555 9662 1581
rect 9634 1554 9662 1555
rect 9686 1581 9714 1582
rect 9738 1581 9766 1582
rect 9686 1555 9698 1581
rect 9698 1555 9714 1581
rect 9738 1555 9760 1581
rect 9760 1555 9766 1581
rect 9686 1554 9714 1555
rect 9738 1554 9766 1555
rect 9790 1554 9818 1582
rect 9842 1581 9870 1582
rect 9894 1581 9922 1582
rect 9842 1555 9848 1581
rect 9848 1555 9870 1581
rect 9894 1555 9910 1581
rect 9910 1555 9922 1581
rect 9842 1554 9870 1555
rect 9894 1554 9922 1555
rect 9946 1581 9974 1582
rect 9946 1555 9972 1581
rect 9972 1555 9974 1581
rect 9946 1554 9974 1555
rect 9998 1581 10026 1582
rect 9998 1555 10008 1581
rect 10008 1555 10026 1581
rect 9998 1554 10026 1555
rect 12726 4494 12754 4522
rect 12950 3710 12978 3738
rect 13342 6062 13370 6090
rect 14582 7069 14610 7070
rect 14582 7043 14600 7069
rect 14600 7043 14610 7069
rect 14582 7042 14610 7043
rect 14634 7069 14662 7070
rect 14634 7043 14636 7069
rect 14636 7043 14662 7069
rect 14634 7042 14662 7043
rect 14686 7069 14714 7070
rect 14738 7069 14766 7070
rect 14686 7043 14698 7069
rect 14698 7043 14714 7069
rect 14738 7043 14760 7069
rect 14760 7043 14766 7069
rect 14686 7042 14714 7043
rect 14738 7042 14766 7043
rect 14790 7042 14818 7070
rect 14842 7069 14870 7070
rect 14894 7069 14922 7070
rect 14842 7043 14848 7069
rect 14848 7043 14870 7069
rect 14894 7043 14910 7069
rect 14910 7043 14922 7069
rect 14842 7042 14870 7043
rect 14894 7042 14922 7043
rect 14946 7069 14974 7070
rect 14946 7043 14972 7069
rect 14972 7043 14974 7069
rect 14946 7042 14974 7043
rect 14998 7069 15026 7070
rect 14998 7043 15008 7069
rect 15008 7043 15026 7069
rect 14998 7042 15026 7043
rect 14406 6873 14434 6874
rect 14406 6847 14407 6873
rect 14407 6847 14433 6873
rect 14433 6847 14434 6873
rect 14406 6846 14434 6847
rect 15078 6846 15106 6874
rect 15190 7630 15218 7658
rect 14582 6285 14610 6286
rect 14582 6259 14600 6285
rect 14600 6259 14610 6285
rect 14582 6258 14610 6259
rect 14634 6285 14662 6286
rect 14634 6259 14636 6285
rect 14636 6259 14662 6285
rect 14634 6258 14662 6259
rect 14686 6285 14714 6286
rect 14738 6285 14766 6286
rect 14686 6259 14698 6285
rect 14698 6259 14714 6285
rect 14738 6259 14760 6285
rect 14760 6259 14766 6285
rect 14686 6258 14714 6259
rect 14738 6258 14766 6259
rect 14790 6258 14818 6286
rect 14842 6285 14870 6286
rect 14894 6285 14922 6286
rect 14842 6259 14848 6285
rect 14848 6259 14870 6285
rect 14894 6259 14910 6285
rect 14910 6259 14922 6285
rect 14842 6258 14870 6259
rect 14894 6258 14922 6259
rect 14946 6285 14974 6286
rect 14946 6259 14972 6285
rect 14972 6259 14974 6285
rect 14946 6258 14974 6259
rect 14998 6285 15026 6286
rect 14998 6259 15008 6285
rect 15008 6259 15026 6285
rect 14998 6258 15026 6259
rect 14462 6118 14490 6146
rect 13510 6062 13538 6090
rect 13958 6089 13986 6090
rect 13958 6063 13959 6089
rect 13959 6063 13985 6089
rect 13985 6063 13986 6089
rect 13958 6062 13986 6063
rect 14854 6145 14882 6146
rect 14854 6119 14855 6145
rect 14855 6119 14881 6145
rect 14881 6119 14882 6145
rect 14854 6118 14882 6119
rect 15190 6089 15218 6090
rect 15190 6063 15191 6089
rect 15191 6063 15217 6089
rect 15217 6063 15218 6089
rect 15190 6062 15218 6063
rect 14582 5501 14610 5502
rect 14582 5475 14600 5501
rect 14600 5475 14610 5501
rect 14582 5474 14610 5475
rect 14634 5501 14662 5502
rect 14634 5475 14636 5501
rect 14636 5475 14662 5501
rect 14634 5474 14662 5475
rect 14686 5501 14714 5502
rect 14738 5501 14766 5502
rect 14686 5475 14698 5501
rect 14698 5475 14714 5501
rect 14738 5475 14760 5501
rect 14760 5475 14766 5501
rect 14686 5474 14714 5475
rect 14738 5474 14766 5475
rect 14790 5474 14818 5502
rect 14842 5501 14870 5502
rect 14894 5501 14922 5502
rect 14842 5475 14848 5501
rect 14848 5475 14870 5501
rect 14894 5475 14910 5501
rect 14910 5475 14922 5501
rect 14842 5474 14870 5475
rect 14894 5474 14922 5475
rect 14946 5501 14974 5502
rect 14946 5475 14972 5501
rect 14972 5475 14974 5501
rect 14946 5474 14974 5475
rect 14998 5501 15026 5502
rect 14998 5475 15008 5501
rect 15008 5475 15026 5501
rect 14998 5474 15026 5475
rect 13342 3710 13370 3738
rect 12726 3345 12754 3346
rect 12726 3319 12727 3345
rect 12727 3319 12753 3345
rect 12753 3319 12754 3345
rect 12726 3318 12754 3319
rect 12726 2982 12754 3010
rect 12726 2198 12754 2226
rect 14182 5278 14210 5306
rect 14462 5305 14490 5306
rect 14462 5279 14463 5305
rect 14463 5279 14489 5305
rect 14489 5279 14490 5305
rect 14462 5278 14490 5279
rect 14182 4857 14210 4858
rect 14182 4831 14183 4857
rect 14183 4831 14209 4857
rect 14209 4831 14210 4857
rect 14182 4830 14210 4831
rect 14582 4717 14610 4718
rect 14582 4691 14600 4717
rect 14600 4691 14610 4717
rect 14582 4690 14610 4691
rect 14634 4717 14662 4718
rect 14634 4691 14636 4717
rect 14636 4691 14662 4717
rect 14634 4690 14662 4691
rect 14686 4717 14714 4718
rect 14738 4717 14766 4718
rect 14686 4691 14698 4717
rect 14698 4691 14714 4717
rect 14738 4691 14760 4717
rect 14760 4691 14766 4717
rect 14686 4690 14714 4691
rect 14738 4690 14766 4691
rect 14790 4690 14818 4718
rect 14842 4717 14870 4718
rect 14894 4717 14922 4718
rect 14842 4691 14848 4717
rect 14848 4691 14870 4717
rect 14894 4691 14910 4717
rect 14910 4691 14922 4717
rect 14842 4690 14870 4691
rect 14894 4690 14922 4691
rect 14946 4717 14974 4718
rect 14946 4691 14972 4717
rect 14972 4691 14974 4717
rect 14946 4690 14974 4691
rect 14998 4717 15026 4718
rect 14998 4691 15008 4717
rect 15008 4691 15026 4717
rect 14998 4690 15026 4691
rect 15694 8441 15722 8442
rect 15694 8415 15695 8441
rect 15695 8415 15721 8441
rect 15721 8415 15722 8441
rect 15694 8414 15722 8415
rect 15918 8441 15946 8442
rect 15918 8415 15919 8441
rect 15919 8415 15945 8441
rect 15945 8415 15946 8441
rect 15918 8414 15946 8415
rect 16198 6873 16226 6874
rect 16198 6847 16199 6873
rect 16199 6847 16225 6873
rect 16225 6847 16226 6873
rect 16198 6846 16226 6847
rect 16758 7630 16786 7658
rect 22082 18437 22110 18438
rect 22082 18411 22100 18437
rect 22100 18411 22110 18437
rect 22082 18410 22110 18411
rect 22134 18437 22162 18438
rect 22134 18411 22136 18437
rect 22136 18411 22162 18437
rect 22134 18410 22162 18411
rect 22186 18437 22214 18438
rect 22238 18437 22266 18438
rect 22186 18411 22198 18437
rect 22198 18411 22214 18437
rect 22238 18411 22260 18437
rect 22260 18411 22266 18437
rect 22186 18410 22214 18411
rect 22238 18410 22266 18411
rect 22290 18410 22318 18438
rect 22342 18437 22370 18438
rect 22394 18437 22422 18438
rect 22342 18411 22348 18437
rect 22348 18411 22370 18437
rect 22394 18411 22410 18437
rect 22410 18411 22422 18437
rect 22342 18410 22370 18411
rect 22394 18410 22422 18411
rect 22446 18437 22474 18438
rect 22446 18411 22472 18437
rect 22472 18411 22474 18437
rect 22446 18410 22474 18411
rect 22498 18437 22526 18438
rect 22498 18411 22508 18437
rect 22508 18411 22526 18437
rect 22498 18410 22526 18411
rect 19582 18045 19610 18046
rect 19582 18019 19600 18045
rect 19600 18019 19610 18045
rect 19582 18018 19610 18019
rect 19634 18045 19662 18046
rect 19634 18019 19636 18045
rect 19636 18019 19662 18045
rect 19634 18018 19662 18019
rect 19686 18045 19714 18046
rect 19738 18045 19766 18046
rect 19686 18019 19698 18045
rect 19698 18019 19714 18045
rect 19738 18019 19760 18045
rect 19760 18019 19766 18045
rect 19686 18018 19714 18019
rect 19738 18018 19766 18019
rect 19790 18018 19818 18046
rect 19842 18045 19870 18046
rect 19894 18045 19922 18046
rect 19842 18019 19848 18045
rect 19848 18019 19870 18045
rect 19894 18019 19910 18045
rect 19910 18019 19922 18045
rect 19842 18018 19870 18019
rect 19894 18018 19922 18019
rect 19946 18045 19974 18046
rect 19946 18019 19972 18045
rect 19972 18019 19974 18045
rect 19946 18018 19974 18019
rect 19998 18045 20026 18046
rect 19998 18019 20008 18045
rect 20008 18019 20026 18045
rect 19998 18018 20026 18019
rect 22082 17653 22110 17654
rect 22082 17627 22100 17653
rect 22100 17627 22110 17653
rect 22082 17626 22110 17627
rect 22134 17653 22162 17654
rect 22134 17627 22136 17653
rect 22136 17627 22162 17653
rect 22134 17626 22162 17627
rect 22186 17653 22214 17654
rect 22238 17653 22266 17654
rect 22186 17627 22198 17653
rect 22198 17627 22214 17653
rect 22238 17627 22260 17653
rect 22260 17627 22266 17653
rect 22186 17626 22214 17627
rect 22238 17626 22266 17627
rect 22290 17626 22318 17654
rect 22342 17653 22370 17654
rect 22394 17653 22422 17654
rect 22342 17627 22348 17653
rect 22348 17627 22370 17653
rect 22394 17627 22410 17653
rect 22410 17627 22422 17653
rect 22342 17626 22370 17627
rect 22394 17626 22422 17627
rect 22446 17653 22474 17654
rect 22446 17627 22472 17653
rect 22472 17627 22474 17653
rect 22446 17626 22474 17627
rect 22498 17653 22526 17654
rect 22498 17627 22508 17653
rect 22508 17627 22526 17653
rect 22498 17626 22526 17627
rect 18494 17318 18522 17346
rect 17598 13454 17626 13482
rect 19582 17261 19610 17262
rect 19582 17235 19600 17261
rect 19600 17235 19610 17261
rect 19582 17234 19610 17235
rect 19634 17261 19662 17262
rect 19634 17235 19636 17261
rect 19636 17235 19662 17261
rect 19634 17234 19662 17235
rect 19686 17261 19714 17262
rect 19738 17261 19766 17262
rect 19686 17235 19698 17261
rect 19698 17235 19714 17261
rect 19738 17235 19760 17261
rect 19760 17235 19766 17261
rect 19686 17234 19714 17235
rect 19738 17234 19766 17235
rect 19790 17234 19818 17262
rect 19842 17261 19870 17262
rect 19894 17261 19922 17262
rect 19842 17235 19848 17261
rect 19848 17235 19870 17261
rect 19894 17235 19910 17261
rect 19910 17235 19922 17261
rect 19842 17234 19870 17235
rect 19894 17234 19922 17235
rect 19946 17261 19974 17262
rect 19946 17235 19972 17261
rect 19972 17235 19974 17261
rect 19946 17234 19974 17235
rect 19998 17261 20026 17262
rect 19998 17235 20008 17261
rect 20008 17235 20026 17261
rect 19998 17234 20026 17235
rect 22082 16869 22110 16870
rect 22082 16843 22100 16869
rect 22100 16843 22110 16869
rect 22082 16842 22110 16843
rect 22134 16869 22162 16870
rect 22134 16843 22136 16869
rect 22136 16843 22162 16869
rect 22134 16842 22162 16843
rect 22186 16869 22214 16870
rect 22238 16869 22266 16870
rect 22186 16843 22198 16869
rect 22198 16843 22214 16869
rect 22238 16843 22260 16869
rect 22260 16843 22266 16869
rect 22186 16842 22214 16843
rect 22238 16842 22266 16843
rect 22290 16842 22318 16870
rect 22342 16869 22370 16870
rect 22394 16869 22422 16870
rect 22342 16843 22348 16869
rect 22348 16843 22370 16869
rect 22394 16843 22410 16869
rect 22410 16843 22422 16869
rect 22342 16842 22370 16843
rect 22394 16842 22422 16843
rect 22446 16869 22474 16870
rect 22446 16843 22472 16869
rect 22472 16843 22474 16869
rect 22446 16842 22474 16843
rect 22498 16869 22526 16870
rect 22498 16843 22508 16869
rect 22508 16843 22526 16869
rect 22498 16842 22526 16843
rect 19582 16477 19610 16478
rect 19582 16451 19600 16477
rect 19600 16451 19610 16477
rect 19582 16450 19610 16451
rect 19634 16477 19662 16478
rect 19634 16451 19636 16477
rect 19636 16451 19662 16477
rect 19634 16450 19662 16451
rect 19686 16477 19714 16478
rect 19738 16477 19766 16478
rect 19686 16451 19698 16477
rect 19698 16451 19714 16477
rect 19738 16451 19760 16477
rect 19760 16451 19766 16477
rect 19686 16450 19714 16451
rect 19738 16450 19766 16451
rect 19790 16450 19818 16478
rect 19842 16477 19870 16478
rect 19894 16477 19922 16478
rect 19842 16451 19848 16477
rect 19848 16451 19870 16477
rect 19894 16451 19910 16477
rect 19910 16451 19922 16477
rect 19842 16450 19870 16451
rect 19894 16450 19922 16451
rect 19946 16477 19974 16478
rect 19946 16451 19972 16477
rect 19972 16451 19974 16477
rect 19946 16450 19974 16451
rect 19998 16477 20026 16478
rect 19998 16451 20008 16477
rect 20008 16451 20026 16477
rect 19998 16450 20026 16451
rect 18494 16366 18522 16394
rect 17878 15974 17906 16002
rect 17082 12949 17110 12950
rect 17082 12923 17100 12949
rect 17100 12923 17110 12949
rect 17082 12922 17110 12923
rect 17134 12949 17162 12950
rect 17134 12923 17136 12949
rect 17136 12923 17162 12949
rect 17134 12922 17162 12923
rect 17186 12949 17214 12950
rect 17238 12949 17266 12950
rect 17186 12923 17198 12949
rect 17198 12923 17214 12949
rect 17238 12923 17260 12949
rect 17260 12923 17266 12949
rect 17186 12922 17214 12923
rect 17238 12922 17266 12923
rect 17290 12922 17318 12950
rect 17342 12949 17370 12950
rect 17394 12949 17422 12950
rect 17342 12923 17348 12949
rect 17348 12923 17370 12949
rect 17394 12923 17410 12949
rect 17410 12923 17422 12949
rect 17342 12922 17370 12923
rect 17394 12922 17422 12923
rect 17446 12949 17474 12950
rect 17446 12923 17472 12949
rect 17472 12923 17474 12949
rect 17446 12922 17474 12923
rect 17498 12949 17526 12950
rect 17498 12923 17508 12949
rect 17508 12923 17526 12949
rect 17498 12922 17526 12923
rect 18270 15862 18298 15890
rect 17934 14238 17962 14266
rect 27082 18437 27110 18438
rect 27082 18411 27100 18437
rect 27100 18411 27110 18437
rect 27082 18410 27110 18411
rect 27134 18437 27162 18438
rect 27134 18411 27136 18437
rect 27136 18411 27162 18437
rect 27134 18410 27162 18411
rect 27186 18437 27214 18438
rect 27238 18437 27266 18438
rect 27186 18411 27198 18437
rect 27198 18411 27214 18437
rect 27238 18411 27260 18437
rect 27260 18411 27266 18437
rect 27186 18410 27214 18411
rect 27238 18410 27266 18411
rect 27290 18410 27318 18438
rect 27342 18437 27370 18438
rect 27394 18437 27422 18438
rect 27342 18411 27348 18437
rect 27348 18411 27370 18437
rect 27394 18411 27410 18437
rect 27410 18411 27422 18437
rect 27342 18410 27370 18411
rect 27394 18410 27422 18411
rect 27446 18437 27474 18438
rect 27446 18411 27472 18437
rect 27472 18411 27474 18437
rect 27446 18410 27474 18411
rect 27498 18437 27526 18438
rect 27498 18411 27508 18437
rect 27508 18411 27526 18437
rect 27498 18410 27526 18411
rect 24582 18045 24610 18046
rect 24582 18019 24600 18045
rect 24600 18019 24610 18045
rect 24582 18018 24610 18019
rect 24634 18045 24662 18046
rect 24634 18019 24636 18045
rect 24636 18019 24662 18045
rect 24634 18018 24662 18019
rect 24686 18045 24714 18046
rect 24738 18045 24766 18046
rect 24686 18019 24698 18045
rect 24698 18019 24714 18045
rect 24738 18019 24760 18045
rect 24760 18019 24766 18045
rect 24686 18018 24714 18019
rect 24738 18018 24766 18019
rect 24790 18018 24818 18046
rect 24842 18045 24870 18046
rect 24894 18045 24922 18046
rect 24842 18019 24848 18045
rect 24848 18019 24870 18045
rect 24894 18019 24910 18045
rect 24910 18019 24922 18045
rect 24842 18018 24870 18019
rect 24894 18018 24922 18019
rect 24946 18045 24974 18046
rect 24946 18019 24972 18045
rect 24972 18019 24974 18045
rect 24946 18018 24974 18019
rect 24998 18045 25026 18046
rect 24998 18019 25008 18045
rect 25008 18019 25026 18045
rect 24998 18018 25026 18019
rect 27082 17653 27110 17654
rect 27082 17627 27100 17653
rect 27100 17627 27110 17653
rect 27082 17626 27110 17627
rect 27134 17653 27162 17654
rect 27134 17627 27136 17653
rect 27136 17627 27162 17653
rect 27134 17626 27162 17627
rect 27186 17653 27214 17654
rect 27238 17653 27266 17654
rect 27186 17627 27198 17653
rect 27198 17627 27214 17653
rect 27238 17627 27260 17653
rect 27260 17627 27266 17653
rect 27186 17626 27214 17627
rect 27238 17626 27266 17627
rect 27290 17626 27318 17654
rect 27342 17653 27370 17654
rect 27394 17653 27422 17654
rect 27342 17627 27348 17653
rect 27348 17627 27370 17653
rect 27394 17627 27410 17653
rect 27410 17627 27422 17653
rect 27342 17626 27370 17627
rect 27394 17626 27422 17627
rect 27446 17653 27474 17654
rect 27446 17627 27472 17653
rect 27472 17627 27474 17653
rect 27446 17626 27474 17627
rect 27498 17653 27526 17654
rect 27498 17627 27508 17653
rect 27508 17627 27526 17653
rect 27498 17626 27526 17627
rect 24582 17261 24610 17262
rect 24582 17235 24600 17261
rect 24600 17235 24610 17261
rect 24582 17234 24610 17235
rect 24634 17261 24662 17262
rect 24634 17235 24636 17261
rect 24636 17235 24662 17261
rect 24634 17234 24662 17235
rect 24686 17261 24714 17262
rect 24738 17261 24766 17262
rect 24686 17235 24698 17261
rect 24698 17235 24714 17261
rect 24738 17235 24760 17261
rect 24760 17235 24766 17261
rect 24686 17234 24714 17235
rect 24738 17234 24766 17235
rect 24790 17234 24818 17262
rect 24842 17261 24870 17262
rect 24894 17261 24922 17262
rect 24842 17235 24848 17261
rect 24848 17235 24870 17261
rect 24894 17235 24910 17261
rect 24910 17235 24922 17261
rect 24842 17234 24870 17235
rect 24894 17234 24922 17235
rect 24946 17261 24974 17262
rect 24946 17235 24972 17261
rect 24972 17235 24974 17261
rect 24946 17234 24974 17235
rect 24998 17261 25026 17262
rect 24998 17235 25008 17261
rect 25008 17235 25026 17261
rect 24998 17234 25026 17235
rect 27082 16869 27110 16870
rect 27082 16843 27100 16869
rect 27100 16843 27110 16869
rect 27082 16842 27110 16843
rect 27134 16869 27162 16870
rect 27134 16843 27136 16869
rect 27136 16843 27162 16869
rect 27134 16842 27162 16843
rect 27186 16869 27214 16870
rect 27238 16869 27266 16870
rect 27186 16843 27198 16869
rect 27198 16843 27214 16869
rect 27238 16843 27260 16869
rect 27260 16843 27266 16869
rect 27186 16842 27214 16843
rect 27238 16842 27266 16843
rect 27290 16842 27318 16870
rect 27342 16869 27370 16870
rect 27394 16869 27422 16870
rect 27342 16843 27348 16869
rect 27348 16843 27370 16869
rect 27394 16843 27410 16869
rect 27410 16843 27422 16869
rect 27342 16842 27370 16843
rect 27394 16842 27422 16843
rect 27446 16869 27474 16870
rect 27446 16843 27472 16869
rect 27472 16843 27474 16869
rect 27446 16842 27474 16843
rect 27498 16869 27526 16870
rect 27498 16843 27508 16869
rect 27508 16843 27526 16869
rect 27498 16842 27526 16843
rect 24582 16477 24610 16478
rect 24582 16451 24600 16477
rect 24600 16451 24610 16477
rect 24582 16450 24610 16451
rect 24634 16477 24662 16478
rect 24634 16451 24636 16477
rect 24636 16451 24662 16477
rect 24634 16450 24662 16451
rect 24686 16477 24714 16478
rect 24738 16477 24766 16478
rect 24686 16451 24698 16477
rect 24698 16451 24714 16477
rect 24738 16451 24760 16477
rect 24760 16451 24766 16477
rect 24686 16450 24714 16451
rect 24738 16450 24766 16451
rect 24790 16450 24818 16478
rect 24842 16477 24870 16478
rect 24894 16477 24922 16478
rect 24842 16451 24848 16477
rect 24848 16451 24870 16477
rect 24894 16451 24910 16477
rect 24910 16451 24922 16477
rect 24842 16450 24870 16451
rect 24894 16450 24922 16451
rect 24946 16477 24974 16478
rect 24946 16451 24972 16477
rect 24972 16451 24974 16477
rect 24946 16450 24974 16451
rect 24998 16477 25026 16478
rect 24998 16451 25008 16477
rect 25008 16451 25026 16477
rect 24998 16450 25026 16451
rect 22582 16254 22610 16282
rect 24094 16366 24122 16394
rect 22082 16085 22110 16086
rect 22082 16059 22100 16085
rect 22100 16059 22110 16085
rect 22082 16058 22110 16059
rect 22134 16085 22162 16086
rect 22134 16059 22136 16085
rect 22136 16059 22162 16085
rect 22134 16058 22162 16059
rect 22186 16085 22214 16086
rect 22238 16085 22266 16086
rect 22186 16059 22198 16085
rect 22198 16059 22214 16085
rect 22238 16059 22260 16085
rect 22260 16059 22266 16085
rect 22186 16058 22214 16059
rect 22238 16058 22266 16059
rect 22290 16058 22318 16086
rect 22342 16085 22370 16086
rect 22394 16085 22422 16086
rect 22342 16059 22348 16085
rect 22348 16059 22370 16085
rect 22394 16059 22410 16085
rect 22410 16059 22422 16085
rect 22342 16058 22370 16059
rect 22394 16058 22422 16059
rect 22446 16085 22474 16086
rect 22446 16059 22472 16085
rect 22472 16059 22474 16085
rect 22446 16058 22474 16059
rect 22498 16085 22526 16086
rect 22498 16059 22508 16085
rect 22508 16059 22526 16085
rect 22498 16058 22526 16059
rect 18718 15974 18746 16002
rect 19222 15974 19250 16002
rect 18774 15889 18802 15890
rect 18774 15863 18775 15889
rect 18775 15863 18801 15889
rect 18801 15863 18802 15889
rect 18774 15862 18802 15863
rect 18270 14294 18298 14322
rect 19582 15693 19610 15694
rect 19582 15667 19600 15693
rect 19600 15667 19610 15693
rect 19582 15666 19610 15667
rect 19634 15693 19662 15694
rect 19634 15667 19636 15693
rect 19636 15667 19662 15693
rect 19634 15666 19662 15667
rect 19686 15693 19714 15694
rect 19738 15693 19766 15694
rect 19686 15667 19698 15693
rect 19698 15667 19714 15693
rect 19738 15667 19760 15693
rect 19760 15667 19766 15693
rect 19686 15666 19714 15667
rect 19738 15666 19766 15667
rect 19790 15666 19818 15694
rect 19842 15693 19870 15694
rect 19894 15693 19922 15694
rect 19842 15667 19848 15693
rect 19848 15667 19870 15693
rect 19894 15667 19910 15693
rect 19910 15667 19922 15693
rect 19842 15666 19870 15667
rect 19894 15666 19922 15667
rect 19946 15693 19974 15694
rect 19946 15667 19972 15693
rect 19972 15667 19974 15693
rect 19946 15666 19974 15667
rect 19998 15693 20026 15694
rect 19998 15667 20008 15693
rect 20008 15667 20026 15693
rect 19998 15666 20026 15667
rect 19582 14909 19610 14910
rect 19582 14883 19600 14909
rect 19600 14883 19610 14909
rect 19582 14882 19610 14883
rect 19634 14909 19662 14910
rect 19634 14883 19636 14909
rect 19636 14883 19662 14909
rect 19634 14882 19662 14883
rect 19686 14909 19714 14910
rect 19738 14909 19766 14910
rect 19686 14883 19698 14909
rect 19698 14883 19714 14909
rect 19738 14883 19760 14909
rect 19760 14883 19766 14909
rect 19686 14882 19714 14883
rect 19738 14882 19766 14883
rect 19790 14882 19818 14910
rect 19842 14909 19870 14910
rect 19894 14909 19922 14910
rect 19842 14883 19848 14909
rect 19848 14883 19870 14909
rect 19894 14883 19910 14909
rect 19910 14883 19922 14909
rect 19842 14882 19870 14883
rect 19894 14882 19922 14883
rect 19946 14909 19974 14910
rect 19946 14883 19972 14909
rect 19972 14883 19974 14909
rect 19946 14882 19974 14883
rect 19998 14909 20026 14910
rect 19998 14883 20008 14909
rect 20008 14883 20026 14909
rect 19998 14882 20026 14883
rect 19446 14321 19474 14322
rect 19446 14295 19447 14321
rect 19447 14295 19473 14321
rect 19473 14295 19474 14321
rect 19446 14294 19474 14295
rect 20790 14630 20818 14658
rect 22082 15301 22110 15302
rect 22082 15275 22100 15301
rect 22100 15275 22110 15301
rect 22082 15274 22110 15275
rect 22134 15301 22162 15302
rect 22134 15275 22136 15301
rect 22136 15275 22162 15301
rect 22134 15274 22162 15275
rect 22186 15301 22214 15302
rect 22238 15301 22266 15302
rect 22186 15275 22198 15301
rect 22198 15275 22214 15301
rect 22238 15275 22260 15301
rect 22260 15275 22266 15301
rect 22186 15274 22214 15275
rect 22238 15274 22266 15275
rect 22290 15274 22318 15302
rect 22342 15301 22370 15302
rect 22394 15301 22422 15302
rect 22342 15275 22348 15301
rect 22348 15275 22370 15301
rect 22394 15275 22410 15301
rect 22410 15275 22422 15301
rect 22342 15274 22370 15275
rect 22394 15274 22422 15275
rect 22446 15301 22474 15302
rect 22446 15275 22472 15301
rect 22472 15275 22474 15301
rect 22446 15274 22474 15275
rect 22498 15301 22526 15302
rect 22498 15275 22508 15301
rect 22508 15275 22526 15301
rect 22498 15274 22526 15275
rect 19582 14125 19610 14126
rect 19582 14099 19600 14125
rect 19600 14099 19610 14125
rect 19582 14098 19610 14099
rect 19634 14125 19662 14126
rect 19634 14099 19636 14125
rect 19636 14099 19662 14125
rect 19634 14098 19662 14099
rect 19686 14125 19714 14126
rect 19738 14125 19766 14126
rect 19686 14099 19698 14125
rect 19698 14099 19714 14125
rect 19738 14099 19760 14125
rect 19760 14099 19766 14125
rect 19686 14098 19714 14099
rect 19738 14098 19766 14099
rect 19790 14098 19818 14126
rect 19842 14125 19870 14126
rect 19894 14125 19922 14126
rect 19842 14099 19848 14125
rect 19848 14099 19870 14125
rect 19894 14099 19910 14125
rect 19910 14099 19922 14125
rect 19842 14098 19870 14099
rect 19894 14098 19922 14099
rect 19946 14125 19974 14126
rect 19946 14099 19972 14125
rect 19972 14099 19974 14125
rect 19946 14098 19974 14099
rect 19998 14125 20026 14126
rect 19998 14099 20008 14125
rect 20008 14099 20026 14125
rect 19998 14098 20026 14099
rect 20678 14321 20706 14322
rect 20678 14295 20679 14321
rect 20679 14295 20705 14321
rect 20705 14295 20706 14321
rect 20678 14294 20706 14295
rect 22582 14630 22610 14658
rect 22082 14517 22110 14518
rect 22082 14491 22100 14517
rect 22100 14491 22110 14517
rect 22082 14490 22110 14491
rect 22134 14517 22162 14518
rect 22134 14491 22136 14517
rect 22136 14491 22162 14517
rect 22134 14490 22162 14491
rect 22186 14517 22214 14518
rect 22238 14517 22266 14518
rect 22186 14491 22198 14517
rect 22198 14491 22214 14517
rect 22238 14491 22260 14517
rect 22260 14491 22266 14517
rect 22186 14490 22214 14491
rect 22238 14490 22266 14491
rect 22290 14490 22318 14518
rect 22342 14517 22370 14518
rect 22394 14517 22422 14518
rect 22342 14491 22348 14517
rect 22348 14491 22370 14517
rect 22394 14491 22410 14517
rect 22410 14491 22422 14517
rect 22342 14490 22370 14491
rect 22394 14490 22422 14491
rect 22446 14517 22474 14518
rect 22446 14491 22472 14517
rect 22472 14491 22474 14517
rect 22446 14490 22474 14491
rect 22498 14517 22526 14518
rect 22498 14491 22508 14517
rect 22508 14491 22526 14517
rect 22498 14490 22526 14491
rect 21014 14321 21042 14322
rect 21014 14295 21015 14321
rect 21015 14295 21041 14321
rect 21041 14295 21042 14321
rect 21014 14294 21042 14295
rect 17990 13145 18018 13146
rect 17990 13119 17991 13145
rect 17991 13119 18017 13145
rect 18017 13119 18018 13145
rect 17990 13118 18018 13119
rect 18550 13398 18578 13426
rect 19054 13398 19082 13426
rect 19582 13341 19610 13342
rect 19582 13315 19600 13341
rect 19600 13315 19610 13341
rect 19582 13314 19610 13315
rect 19634 13341 19662 13342
rect 19634 13315 19636 13341
rect 19636 13315 19662 13341
rect 19634 13314 19662 13315
rect 19686 13341 19714 13342
rect 19738 13341 19766 13342
rect 19686 13315 19698 13341
rect 19698 13315 19714 13341
rect 19738 13315 19760 13341
rect 19760 13315 19766 13341
rect 19686 13314 19714 13315
rect 19738 13314 19766 13315
rect 19790 13314 19818 13342
rect 19842 13341 19870 13342
rect 19894 13341 19922 13342
rect 19842 13315 19848 13341
rect 19848 13315 19870 13341
rect 19894 13315 19910 13341
rect 19910 13315 19922 13341
rect 19842 13314 19870 13315
rect 19894 13314 19922 13315
rect 19946 13341 19974 13342
rect 19946 13315 19972 13341
rect 19972 13315 19974 13341
rect 19946 13314 19974 13315
rect 19998 13341 20026 13342
rect 19998 13315 20008 13341
rect 20008 13315 20026 13341
rect 19998 13314 20026 13315
rect 17082 12165 17110 12166
rect 17082 12139 17100 12165
rect 17100 12139 17110 12165
rect 17082 12138 17110 12139
rect 17134 12165 17162 12166
rect 17134 12139 17136 12165
rect 17136 12139 17162 12165
rect 17134 12138 17162 12139
rect 17186 12165 17214 12166
rect 17238 12165 17266 12166
rect 17186 12139 17198 12165
rect 17198 12139 17214 12165
rect 17238 12139 17260 12165
rect 17260 12139 17266 12165
rect 17186 12138 17214 12139
rect 17238 12138 17266 12139
rect 17290 12138 17318 12166
rect 17342 12165 17370 12166
rect 17394 12165 17422 12166
rect 17342 12139 17348 12165
rect 17348 12139 17370 12165
rect 17394 12139 17410 12165
rect 17410 12139 17422 12165
rect 17342 12138 17370 12139
rect 17394 12138 17422 12139
rect 17446 12165 17474 12166
rect 17446 12139 17472 12165
rect 17472 12139 17474 12165
rect 17446 12138 17474 12139
rect 17498 12165 17526 12166
rect 17498 12139 17508 12165
rect 17508 12139 17526 12165
rect 17498 12138 17526 12139
rect 16926 11942 16954 11970
rect 19446 13145 19474 13146
rect 19446 13119 19447 13145
rect 19447 13119 19473 13145
rect 19473 13119 19474 13145
rect 19446 13118 19474 13119
rect 18774 12614 18802 12642
rect 19446 12670 19474 12698
rect 19950 12697 19978 12698
rect 19950 12671 19951 12697
rect 19951 12671 19977 12697
rect 19977 12671 19978 12697
rect 19950 12670 19978 12671
rect 19582 12557 19610 12558
rect 19582 12531 19600 12557
rect 19600 12531 19610 12557
rect 19582 12530 19610 12531
rect 19634 12557 19662 12558
rect 19634 12531 19636 12557
rect 19636 12531 19662 12557
rect 19634 12530 19662 12531
rect 19686 12557 19714 12558
rect 19738 12557 19766 12558
rect 19686 12531 19698 12557
rect 19698 12531 19714 12557
rect 19738 12531 19760 12557
rect 19760 12531 19766 12557
rect 19686 12530 19714 12531
rect 19738 12530 19766 12531
rect 19790 12530 19818 12558
rect 19842 12557 19870 12558
rect 19894 12557 19922 12558
rect 19842 12531 19848 12557
rect 19848 12531 19870 12557
rect 19894 12531 19910 12557
rect 19910 12531 19922 12557
rect 19842 12530 19870 12531
rect 19894 12530 19922 12531
rect 19946 12557 19974 12558
rect 19946 12531 19972 12557
rect 19972 12531 19974 12557
rect 19946 12530 19974 12531
rect 19998 12557 20026 12558
rect 19998 12531 20008 12557
rect 20008 12531 20026 12557
rect 19998 12530 20026 12531
rect 19950 11969 19978 11970
rect 19950 11943 19951 11969
rect 19951 11943 19977 11969
rect 19977 11943 19978 11969
rect 19950 11942 19978 11943
rect 20118 11942 20146 11970
rect 20510 12614 20538 12642
rect 19582 11773 19610 11774
rect 19582 11747 19600 11773
rect 19600 11747 19610 11773
rect 19582 11746 19610 11747
rect 19634 11773 19662 11774
rect 19634 11747 19636 11773
rect 19636 11747 19662 11773
rect 19634 11746 19662 11747
rect 19686 11773 19714 11774
rect 19738 11773 19766 11774
rect 19686 11747 19698 11773
rect 19698 11747 19714 11773
rect 19738 11747 19760 11773
rect 19760 11747 19766 11773
rect 19686 11746 19714 11747
rect 19738 11746 19766 11747
rect 19790 11746 19818 11774
rect 19842 11773 19870 11774
rect 19894 11773 19922 11774
rect 19842 11747 19848 11773
rect 19848 11747 19870 11773
rect 19894 11747 19910 11773
rect 19910 11747 19922 11773
rect 19842 11746 19870 11747
rect 19894 11746 19922 11747
rect 19946 11773 19974 11774
rect 19946 11747 19972 11773
rect 19972 11747 19974 11773
rect 19946 11746 19974 11747
rect 19998 11773 20026 11774
rect 19998 11747 20008 11773
rect 20008 11747 20026 11773
rect 19998 11746 20026 11747
rect 17082 11381 17110 11382
rect 17082 11355 17100 11381
rect 17100 11355 17110 11381
rect 17082 11354 17110 11355
rect 17134 11381 17162 11382
rect 17134 11355 17136 11381
rect 17136 11355 17162 11381
rect 17134 11354 17162 11355
rect 17186 11381 17214 11382
rect 17238 11381 17266 11382
rect 17186 11355 17198 11381
rect 17198 11355 17214 11381
rect 17238 11355 17260 11381
rect 17260 11355 17266 11381
rect 17186 11354 17214 11355
rect 17238 11354 17266 11355
rect 17290 11354 17318 11382
rect 17342 11381 17370 11382
rect 17394 11381 17422 11382
rect 17342 11355 17348 11381
rect 17348 11355 17370 11381
rect 17394 11355 17410 11381
rect 17410 11355 17422 11381
rect 17342 11354 17370 11355
rect 17394 11354 17422 11355
rect 17446 11381 17474 11382
rect 17446 11355 17472 11381
rect 17472 11355 17474 11381
rect 17446 11354 17474 11355
rect 17498 11381 17526 11382
rect 17498 11355 17508 11381
rect 17508 11355 17526 11381
rect 17498 11354 17526 11355
rect 17654 10710 17682 10738
rect 17082 10597 17110 10598
rect 17082 10571 17100 10597
rect 17100 10571 17110 10597
rect 17082 10570 17110 10571
rect 17134 10597 17162 10598
rect 17134 10571 17136 10597
rect 17136 10571 17162 10597
rect 17134 10570 17162 10571
rect 17186 10597 17214 10598
rect 17238 10597 17266 10598
rect 17186 10571 17198 10597
rect 17198 10571 17214 10597
rect 17238 10571 17260 10597
rect 17260 10571 17266 10597
rect 17186 10570 17214 10571
rect 17238 10570 17266 10571
rect 17290 10570 17318 10598
rect 17342 10597 17370 10598
rect 17394 10597 17422 10598
rect 17342 10571 17348 10597
rect 17348 10571 17370 10597
rect 17394 10571 17410 10597
rect 17410 10571 17422 10597
rect 17342 10570 17370 10571
rect 17394 10570 17422 10571
rect 17446 10597 17474 10598
rect 17446 10571 17472 10597
rect 17472 10571 17474 10597
rect 17446 10570 17474 10571
rect 17498 10597 17526 10598
rect 17498 10571 17508 10597
rect 17508 10571 17526 10597
rect 17498 10570 17526 10571
rect 17082 9813 17110 9814
rect 17082 9787 17100 9813
rect 17100 9787 17110 9813
rect 17082 9786 17110 9787
rect 17134 9813 17162 9814
rect 17134 9787 17136 9813
rect 17136 9787 17162 9813
rect 17134 9786 17162 9787
rect 17186 9813 17214 9814
rect 17238 9813 17266 9814
rect 17186 9787 17198 9813
rect 17198 9787 17214 9813
rect 17238 9787 17260 9813
rect 17260 9787 17266 9813
rect 17186 9786 17214 9787
rect 17238 9786 17266 9787
rect 17290 9786 17318 9814
rect 17342 9813 17370 9814
rect 17394 9813 17422 9814
rect 17342 9787 17348 9813
rect 17348 9787 17370 9813
rect 17394 9787 17410 9813
rect 17410 9787 17422 9813
rect 17342 9786 17370 9787
rect 17394 9786 17422 9787
rect 17446 9813 17474 9814
rect 17446 9787 17472 9813
rect 17472 9787 17474 9813
rect 17446 9786 17474 9787
rect 17498 9813 17526 9814
rect 17498 9787 17508 9813
rect 17508 9787 17526 9813
rect 17498 9786 17526 9787
rect 18886 11214 18914 11242
rect 17990 10401 18018 10402
rect 17990 10375 17991 10401
rect 17991 10375 18017 10401
rect 18017 10375 18018 10401
rect 17990 10374 18018 10375
rect 18102 10345 18130 10346
rect 18102 10319 18103 10345
rect 18103 10319 18129 10345
rect 18129 10319 18130 10345
rect 18102 10318 18130 10319
rect 18270 9617 18298 9618
rect 18270 9591 18271 9617
rect 18271 9591 18297 9617
rect 18297 9591 18298 9617
rect 18270 9590 18298 9591
rect 18718 10009 18746 10010
rect 18718 9983 18719 10009
rect 18719 9983 18745 10009
rect 18745 9983 18746 10009
rect 18718 9982 18746 9983
rect 18718 9590 18746 9618
rect 17654 9142 17682 9170
rect 18214 9142 18242 9170
rect 17082 9029 17110 9030
rect 17082 9003 17100 9029
rect 17100 9003 17110 9029
rect 17082 9002 17110 9003
rect 17134 9029 17162 9030
rect 17134 9003 17136 9029
rect 17136 9003 17162 9029
rect 17134 9002 17162 9003
rect 17186 9029 17214 9030
rect 17238 9029 17266 9030
rect 17186 9003 17198 9029
rect 17198 9003 17214 9029
rect 17238 9003 17260 9029
rect 17260 9003 17266 9029
rect 17186 9002 17214 9003
rect 17238 9002 17266 9003
rect 17290 9002 17318 9030
rect 17342 9029 17370 9030
rect 17394 9029 17422 9030
rect 17342 9003 17348 9029
rect 17348 9003 17370 9029
rect 17394 9003 17410 9029
rect 17410 9003 17422 9029
rect 17342 9002 17370 9003
rect 17394 9002 17422 9003
rect 17446 9029 17474 9030
rect 17446 9003 17472 9029
rect 17472 9003 17474 9029
rect 17446 9002 17474 9003
rect 17498 9029 17526 9030
rect 17498 9003 17508 9029
rect 17508 9003 17526 9029
rect 17498 9002 17526 9003
rect 17206 8833 17234 8834
rect 17206 8807 17207 8833
rect 17207 8807 17233 8833
rect 17233 8807 17234 8833
rect 17206 8806 17234 8807
rect 17082 8245 17110 8246
rect 17082 8219 17100 8245
rect 17100 8219 17110 8245
rect 17082 8218 17110 8219
rect 17134 8245 17162 8246
rect 17134 8219 17136 8245
rect 17136 8219 17162 8245
rect 17134 8218 17162 8219
rect 17186 8245 17214 8246
rect 17238 8245 17266 8246
rect 17186 8219 17198 8245
rect 17198 8219 17214 8245
rect 17238 8219 17260 8245
rect 17260 8219 17266 8245
rect 17186 8218 17214 8219
rect 17238 8218 17266 8219
rect 17290 8218 17318 8246
rect 17342 8245 17370 8246
rect 17394 8245 17422 8246
rect 17342 8219 17348 8245
rect 17348 8219 17370 8245
rect 17394 8219 17410 8245
rect 17410 8219 17422 8245
rect 17342 8218 17370 8219
rect 17394 8218 17422 8219
rect 17446 8245 17474 8246
rect 17446 8219 17472 8245
rect 17472 8219 17474 8245
rect 17446 8218 17474 8219
rect 17498 8245 17526 8246
rect 17498 8219 17508 8245
rect 17508 8219 17526 8245
rect 17498 8218 17526 8219
rect 16870 7657 16898 7658
rect 16870 7631 16871 7657
rect 16871 7631 16897 7657
rect 16897 7631 16898 7657
rect 16870 7630 16898 7631
rect 16422 6846 16450 6874
rect 15694 6118 15722 6146
rect 16422 5838 16450 5866
rect 17082 7461 17110 7462
rect 17082 7435 17100 7461
rect 17100 7435 17110 7461
rect 17082 7434 17110 7435
rect 17134 7461 17162 7462
rect 17134 7435 17136 7461
rect 17136 7435 17162 7461
rect 17134 7434 17162 7435
rect 17186 7461 17214 7462
rect 17238 7461 17266 7462
rect 17186 7435 17198 7461
rect 17198 7435 17214 7461
rect 17238 7435 17260 7461
rect 17260 7435 17266 7461
rect 17186 7434 17214 7435
rect 17238 7434 17266 7435
rect 17290 7434 17318 7462
rect 17342 7461 17370 7462
rect 17394 7461 17422 7462
rect 17342 7435 17348 7461
rect 17348 7435 17370 7461
rect 17394 7435 17410 7461
rect 17410 7435 17422 7461
rect 17342 7434 17370 7435
rect 17394 7434 17422 7435
rect 17446 7461 17474 7462
rect 17446 7435 17472 7461
rect 17472 7435 17474 7461
rect 17446 7434 17474 7435
rect 17498 7461 17526 7462
rect 17498 7435 17508 7461
rect 17508 7435 17526 7461
rect 17498 7434 17526 7435
rect 17374 6873 17402 6874
rect 17374 6847 17375 6873
rect 17375 6847 17401 6873
rect 17401 6847 17402 6873
rect 17374 6846 17402 6847
rect 17082 6677 17110 6678
rect 17082 6651 17100 6677
rect 17100 6651 17110 6677
rect 17082 6650 17110 6651
rect 17134 6677 17162 6678
rect 17134 6651 17136 6677
rect 17136 6651 17162 6677
rect 17134 6650 17162 6651
rect 17186 6677 17214 6678
rect 17238 6677 17266 6678
rect 17186 6651 17198 6677
rect 17198 6651 17214 6677
rect 17238 6651 17260 6677
rect 17260 6651 17266 6677
rect 17186 6650 17214 6651
rect 17238 6650 17266 6651
rect 17290 6650 17318 6678
rect 17342 6677 17370 6678
rect 17394 6677 17422 6678
rect 17342 6651 17348 6677
rect 17348 6651 17370 6677
rect 17394 6651 17410 6677
rect 17410 6651 17422 6677
rect 17342 6650 17370 6651
rect 17394 6650 17422 6651
rect 17446 6677 17474 6678
rect 17446 6651 17472 6677
rect 17472 6651 17474 6677
rect 17446 6650 17474 6651
rect 17498 6677 17526 6678
rect 17498 6651 17508 6677
rect 17508 6651 17526 6677
rect 17498 6650 17526 6651
rect 16814 5838 16842 5866
rect 17082 5893 17110 5894
rect 17082 5867 17100 5893
rect 17100 5867 17110 5893
rect 17082 5866 17110 5867
rect 17134 5893 17162 5894
rect 17134 5867 17136 5893
rect 17136 5867 17162 5893
rect 17134 5866 17162 5867
rect 17186 5893 17214 5894
rect 17238 5893 17266 5894
rect 17186 5867 17198 5893
rect 17198 5867 17214 5893
rect 17238 5867 17260 5893
rect 17260 5867 17266 5893
rect 17186 5866 17214 5867
rect 17238 5866 17266 5867
rect 17290 5866 17318 5894
rect 17342 5893 17370 5894
rect 17394 5893 17422 5894
rect 17342 5867 17348 5893
rect 17348 5867 17370 5893
rect 17394 5867 17410 5893
rect 17410 5867 17422 5893
rect 17342 5866 17370 5867
rect 17394 5866 17422 5867
rect 17446 5893 17474 5894
rect 17446 5867 17472 5893
rect 17472 5867 17474 5893
rect 17446 5866 17474 5867
rect 17498 5893 17526 5894
rect 17498 5867 17508 5893
rect 17508 5867 17526 5893
rect 17498 5866 17526 5867
rect 16982 5334 17010 5362
rect 13566 3710 13594 3738
rect 14126 3737 14154 3738
rect 14126 3711 14127 3737
rect 14127 3711 14153 3737
rect 14153 3711 14154 3737
rect 14126 3710 14154 3711
rect 13342 3374 13370 3402
rect 13678 3345 13706 3346
rect 13678 3319 13679 3345
rect 13679 3319 13705 3345
rect 13705 3319 13706 3345
rect 13678 3318 13706 3319
rect 13902 3345 13930 3346
rect 13902 3319 13903 3345
rect 13903 3319 13929 3345
rect 13929 3319 13930 3345
rect 13902 3318 13930 3319
rect 14126 3318 14154 3346
rect 14582 3933 14610 3934
rect 14582 3907 14600 3933
rect 14600 3907 14610 3933
rect 14582 3906 14610 3907
rect 14634 3933 14662 3934
rect 14634 3907 14636 3933
rect 14636 3907 14662 3933
rect 14634 3906 14662 3907
rect 14686 3933 14714 3934
rect 14738 3933 14766 3934
rect 14686 3907 14698 3933
rect 14698 3907 14714 3933
rect 14738 3907 14760 3933
rect 14760 3907 14766 3933
rect 14686 3906 14714 3907
rect 14738 3906 14766 3907
rect 14790 3906 14818 3934
rect 14842 3933 14870 3934
rect 14894 3933 14922 3934
rect 14842 3907 14848 3933
rect 14848 3907 14870 3933
rect 14894 3907 14910 3933
rect 14910 3907 14922 3933
rect 14842 3906 14870 3907
rect 14894 3906 14922 3907
rect 14946 3933 14974 3934
rect 14946 3907 14972 3933
rect 14972 3907 14974 3933
rect 14946 3906 14974 3907
rect 14998 3933 15026 3934
rect 14998 3907 15008 3933
rect 15008 3907 15026 3933
rect 14998 3906 15026 3907
rect 14350 3737 14378 3738
rect 14350 3711 14351 3737
rect 14351 3711 14377 3737
rect 14377 3711 14378 3737
rect 14350 3710 14378 3711
rect 15134 3318 15162 3346
rect 14582 3149 14610 3150
rect 14582 3123 14600 3149
rect 14600 3123 14610 3149
rect 14582 3122 14610 3123
rect 14634 3149 14662 3150
rect 14634 3123 14636 3149
rect 14636 3123 14662 3149
rect 14634 3122 14662 3123
rect 14686 3149 14714 3150
rect 14738 3149 14766 3150
rect 14686 3123 14698 3149
rect 14698 3123 14714 3149
rect 14738 3123 14760 3149
rect 14760 3123 14766 3149
rect 14686 3122 14714 3123
rect 14738 3122 14766 3123
rect 14790 3122 14818 3150
rect 14842 3149 14870 3150
rect 14894 3149 14922 3150
rect 14842 3123 14848 3149
rect 14848 3123 14870 3149
rect 14894 3123 14910 3149
rect 14910 3123 14922 3149
rect 14842 3122 14870 3123
rect 14894 3122 14922 3123
rect 14946 3149 14974 3150
rect 14946 3123 14972 3149
rect 14972 3123 14974 3149
rect 14946 3122 14974 3123
rect 14998 3149 15026 3150
rect 14998 3123 15008 3149
rect 15008 3123 15026 3149
rect 14998 3122 15026 3123
rect 14126 2926 14154 2954
rect 13342 2142 13370 2170
rect 13510 2198 13538 2226
rect 14070 2198 14098 2226
rect 13622 2169 13650 2170
rect 13622 2143 13623 2169
rect 13623 2143 13649 2169
rect 13649 2143 13650 2169
rect 13622 2142 13650 2143
rect 14238 2590 14266 2618
rect 15246 3262 15274 3290
rect 15302 2870 15330 2898
rect 14582 2365 14610 2366
rect 14582 2339 14600 2365
rect 14600 2339 14610 2365
rect 14582 2338 14610 2339
rect 14634 2365 14662 2366
rect 14634 2339 14636 2365
rect 14636 2339 14662 2365
rect 14634 2338 14662 2339
rect 14686 2365 14714 2366
rect 14738 2365 14766 2366
rect 14686 2339 14698 2365
rect 14698 2339 14714 2365
rect 14738 2339 14760 2365
rect 14760 2339 14766 2365
rect 14686 2338 14714 2339
rect 14738 2338 14766 2339
rect 14790 2338 14818 2366
rect 14842 2365 14870 2366
rect 14894 2365 14922 2366
rect 14842 2339 14848 2365
rect 14848 2339 14870 2365
rect 14894 2339 14910 2365
rect 14910 2339 14922 2365
rect 14842 2338 14870 2339
rect 14894 2338 14922 2339
rect 14946 2365 14974 2366
rect 14946 2339 14972 2365
rect 14972 2339 14974 2365
rect 14946 2338 14974 2339
rect 14998 2365 15026 2366
rect 14998 2339 15008 2365
rect 15008 2339 15026 2365
rect 14998 2338 15026 2339
rect 14294 2198 14322 2226
rect 15246 2478 15274 2506
rect 15134 2169 15162 2170
rect 15134 2143 15135 2169
rect 15135 2143 15161 2169
rect 15161 2143 15162 2169
rect 15134 2142 15162 2143
rect 15302 1806 15330 1834
rect 15470 4521 15498 4522
rect 15470 4495 15471 4521
rect 15471 4495 15497 4521
rect 15497 4495 15498 4521
rect 15470 4494 15498 4495
rect 15470 3710 15498 3738
rect 17082 5109 17110 5110
rect 17082 5083 17100 5109
rect 17100 5083 17110 5109
rect 17082 5082 17110 5083
rect 17134 5109 17162 5110
rect 17134 5083 17136 5109
rect 17136 5083 17162 5109
rect 17134 5082 17162 5083
rect 17186 5109 17214 5110
rect 17238 5109 17266 5110
rect 17186 5083 17198 5109
rect 17198 5083 17214 5109
rect 17238 5083 17260 5109
rect 17260 5083 17266 5109
rect 17186 5082 17214 5083
rect 17238 5082 17266 5083
rect 17290 5082 17318 5110
rect 17342 5109 17370 5110
rect 17394 5109 17422 5110
rect 17342 5083 17348 5109
rect 17348 5083 17370 5109
rect 17394 5083 17410 5109
rect 17410 5083 17422 5109
rect 17342 5082 17370 5083
rect 17394 5082 17422 5083
rect 17446 5109 17474 5110
rect 17446 5083 17472 5109
rect 17472 5083 17474 5109
rect 17446 5082 17474 5083
rect 17498 5109 17526 5110
rect 17498 5083 17508 5109
rect 17508 5083 17526 5109
rect 17498 5082 17526 5083
rect 15694 4521 15722 4522
rect 15694 4495 15695 4521
rect 15695 4495 15721 4521
rect 15721 4495 15722 4521
rect 15694 4494 15722 4495
rect 15582 3737 15610 3738
rect 15582 3711 15583 3737
rect 15583 3711 15609 3737
rect 15609 3711 15610 3737
rect 15582 3710 15610 3711
rect 15806 3737 15834 3738
rect 15806 3711 15807 3737
rect 15807 3711 15833 3737
rect 15833 3711 15834 3737
rect 15806 3710 15834 3711
rect 15974 3710 16002 3738
rect 18774 8833 18802 8834
rect 18774 8807 18775 8833
rect 18775 8807 18801 8833
rect 18801 8807 18802 8833
rect 18774 8806 18802 8807
rect 18214 4662 18242 4690
rect 17082 4325 17110 4326
rect 17082 4299 17100 4325
rect 17100 4299 17110 4325
rect 17082 4298 17110 4299
rect 17134 4325 17162 4326
rect 17134 4299 17136 4325
rect 17136 4299 17162 4325
rect 17134 4298 17162 4299
rect 17186 4325 17214 4326
rect 17238 4325 17266 4326
rect 17186 4299 17198 4325
rect 17198 4299 17214 4325
rect 17238 4299 17260 4325
rect 17260 4299 17266 4325
rect 17186 4298 17214 4299
rect 17238 4298 17266 4299
rect 17290 4298 17318 4326
rect 17342 4325 17370 4326
rect 17394 4325 17422 4326
rect 17342 4299 17348 4325
rect 17348 4299 17370 4325
rect 17394 4299 17410 4325
rect 17410 4299 17422 4325
rect 17342 4298 17370 4299
rect 17394 4298 17422 4299
rect 17446 4325 17474 4326
rect 17446 4299 17472 4325
rect 17472 4299 17474 4325
rect 17446 4298 17474 4299
rect 17498 4325 17526 4326
rect 17498 4299 17508 4325
rect 17508 4299 17526 4325
rect 17498 4298 17526 4299
rect 15526 3345 15554 3346
rect 15526 3319 15527 3345
rect 15527 3319 15553 3345
rect 15553 3319 15554 3345
rect 15526 3318 15554 3319
rect 17082 3541 17110 3542
rect 17082 3515 17100 3541
rect 17100 3515 17110 3541
rect 17082 3514 17110 3515
rect 17134 3541 17162 3542
rect 17134 3515 17136 3541
rect 17136 3515 17162 3541
rect 17134 3514 17162 3515
rect 17186 3541 17214 3542
rect 17238 3541 17266 3542
rect 17186 3515 17198 3541
rect 17198 3515 17214 3541
rect 17238 3515 17260 3541
rect 17260 3515 17266 3541
rect 17186 3514 17214 3515
rect 17238 3514 17266 3515
rect 17290 3514 17318 3542
rect 17342 3541 17370 3542
rect 17394 3541 17422 3542
rect 17342 3515 17348 3541
rect 17348 3515 17370 3541
rect 17394 3515 17410 3541
rect 17410 3515 17422 3541
rect 17342 3514 17370 3515
rect 17394 3514 17422 3515
rect 17446 3541 17474 3542
rect 17446 3515 17472 3541
rect 17472 3515 17474 3541
rect 17446 3514 17474 3515
rect 17498 3541 17526 3542
rect 17498 3515 17508 3541
rect 17508 3515 17526 3541
rect 17498 3514 17526 3515
rect 15470 2870 15498 2898
rect 17990 4606 18018 4634
rect 17934 3318 17962 3346
rect 15918 2561 15946 2562
rect 15918 2535 15919 2561
rect 15919 2535 15945 2561
rect 15945 2535 15946 2561
rect 15918 2534 15946 2535
rect 17082 2757 17110 2758
rect 17082 2731 17100 2757
rect 17100 2731 17110 2757
rect 17082 2730 17110 2731
rect 17134 2757 17162 2758
rect 17134 2731 17136 2757
rect 17136 2731 17162 2757
rect 17134 2730 17162 2731
rect 17186 2757 17214 2758
rect 17238 2757 17266 2758
rect 17186 2731 17198 2757
rect 17198 2731 17214 2757
rect 17238 2731 17260 2757
rect 17260 2731 17266 2757
rect 17186 2730 17214 2731
rect 17238 2730 17266 2731
rect 17290 2730 17318 2758
rect 17342 2757 17370 2758
rect 17394 2757 17422 2758
rect 17342 2731 17348 2757
rect 17348 2731 17370 2757
rect 17394 2731 17410 2757
rect 17410 2731 17422 2757
rect 17342 2730 17370 2731
rect 17394 2730 17422 2731
rect 17446 2757 17474 2758
rect 17446 2731 17472 2757
rect 17472 2731 17474 2757
rect 17446 2730 17474 2731
rect 17498 2757 17526 2758
rect 17498 2731 17508 2757
rect 17508 2731 17526 2757
rect 17498 2730 17526 2731
rect 17598 2590 17626 2618
rect 17150 2561 17178 2562
rect 17150 2535 17151 2561
rect 17151 2535 17177 2561
rect 17177 2535 17178 2561
rect 17150 2534 17178 2535
rect 17374 2561 17402 2562
rect 17374 2535 17375 2561
rect 17375 2535 17401 2561
rect 17401 2535 17402 2561
rect 17374 2534 17402 2535
rect 16814 2478 16842 2506
rect 16590 2142 16618 2170
rect 15526 1806 15554 1834
rect 17082 1973 17110 1974
rect 17082 1947 17100 1973
rect 17100 1947 17110 1973
rect 17082 1946 17110 1947
rect 17134 1973 17162 1974
rect 17134 1947 17136 1973
rect 17136 1947 17162 1973
rect 17134 1946 17162 1947
rect 17186 1973 17214 1974
rect 17238 1973 17266 1974
rect 17186 1947 17198 1973
rect 17198 1947 17214 1973
rect 17238 1947 17260 1973
rect 17260 1947 17266 1973
rect 17186 1946 17214 1947
rect 17238 1946 17266 1947
rect 17290 1946 17318 1974
rect 17342 1973 17370 1974
rect 17394 1973 17422 1974
rect 17342 1947 17348 1973
rect 17348 1947 17370 1973
rect 17394 1947 17410 1973
rect 17410 1947 17422 1973
rect 17342 1946 17370 1947
rect 17394 1946 17422 1947
rect 17446 1973 17474 1974
rect 17446 1947 17472 1973
rect 17472 1947 17474 1973
rect 17446 1946 17474 1947
rect 17498 1973 17526 1974
rect 17498 1947 17508 1973
rect 17508 1947 17526 1973
rect 17498 1946 17526 1947
rect 16590 1862 16618 1890
rect 17038 1862 17066 1890
rect 14582 1581 14610 1582
rect 14582 1555 14600 1581
rect 14600 1555 14610 1581
rect 14582 1554 14610 1555
rect 14634 1581 14662 1582
rect 14634 1555 14636 1581
rect 14636 1555 14662 1581
rect 14634 1554 14662 1555
rect 14686 1581 14714 1582
rect 14738 1581 14766 1582
rect 14686 1555 14698 1581
rect 14698 1555 14714 1581
rect 14738 1555 14760 1581
rect 14760 1555 14766 1581
rect 14686 1554 14714 1555
rect 14738 1554 14766 1555
rect 14790 1554 14818 1582
rect 14842 1581 14870 1582
rect 14894 1581 14922 1582
rect 14842 1555 14848 1581
rect 14848 1555 14870 1581
rect 14894 1555 14910 1581
rect 14910 1555 14922 1581
rect 14842 1554 14870 1555
rect 14894 1554 14922 1555
rect 14946 1581 14974 1582
rect 14946 1555 14972 1581
rect 14972 1555 14974 1581
rect 14946 1554 14974 1555
rect 14998 1581 15026 1582
rect 14998 1555 15008 1581
rect 15008 1555 15026 1581
rect 14998 1554 15026 1555
rect 17654 2534 17682 2562
rect 18774 5054 18802 5082
rect 18494 3374 18522 3402
rect 18270 2169 18298 2170
rect 18270 2143 18271 2169
rect 18271 2143 18297 2169
rect 18297 2143 18298 2169
rect 18270 2142 18298 2143
rect 17990 1862 18018 1890
rect 22526 14294 22554 14322
rect 23422 14713 23450 14714
rect 23422 14687 23423 14713
rect 23423 14687 23449 14713
rect 23449 14687 23450 14713
rect 23422 14686 23450 14687
rect 23926 14686 23954 14714
rect 23030 14321 23058 14322
rect 23030 14295 23031 14321
rect 23031 14295 23057 14321
rect 23057 14295 23058 14321
rect 23030 14294 23058 14295
rect 21462 13929 21490 13930
rect 21462 13903 21463 13929
rect 21463 13903 21489 13929
rect 21489 13903 21490 13929
rect 21462 13902 21490 13903
rect 22082 13733 22110 13734
rect 22082 13707 22100 13733
rect 22100 13707 22110 13733
rect 22082 13706 22110 13707
rect 22134 13733 22162 13734
rect 22134 13707 22136 13733
rect 22136 13707 22162 13733
rect 22134 13706 22162 13707
rect 22186 13733 22214 13734
rect 22238 13733 22266 13734
rect 22186 13707 22198 13733
rect 22198 13707 22214 13733
rect 22238 13707 22260 13733
rect 22260 13707 22266 13733
rect 22186 13706 22214 13707
rect 22238 13706 22266 13707
rect 22290 13706 22318 13734
rect 22342 13733 22370 13734
rect 22394 13733 22422 13734
rect 22342 13707 22348 13733
rect 22348 13707 22370 13733
rect 22394 13707 22410 13733
rect 22410 13707 22422 13733
rect 22342 13706 22370 13707
rect 22394 13706 22422 13707
rect 22446 13733 22474 13734
rect 22446 13707 22472 13733
rect 22472 13707 22474 13733
rect 22446 13706 22474 13707
rect 22498 13733 22526 13734
rect 22498 13707 22508 13733
rect 22508 13707 22526 13733
rect 22498 13706 22526 13707
rect 20958 12614 20986 12642
rect 23926 14265 23954 14266
rect 23926 14239 23927 14265
rect 23927 14239 23953 14265
rect 23953 14239 23954 14265
rect 23926 14238 23954 14239
rect 23422 13929 23450 13930
rect 23422 13903 23423 13929
rect 23423 13903 23449 13929
rect 23449 13903 23450 13929
rect 23422 13902 23450 13903
rect 23422 13454 23450 13482
rect 23926 13481 23954 13482
rect 23926 13455 23927 13481
rect 23927 13455 23953 13481
rect 23953 13455 23954 13481
rect 23926 13454 23954 13455
rect 22082 12949 22110 12950
rect 22082 12923 22100 12949
rect 22100 12923 22110 12949
rect 22082 12922 22110 12923
rect 22134 12949 22162 12950
rect 22134 12923 22136 12949
rect 22136 12923 22162 12949
rect 22134 12922 22162 12923
rect 22186 12949 22214 12950
rect 22238 12949 22266 12950
rect 22186 12923 22198 12949
rect 22198 12923 22214 12949
rect 22238 12923 22260 12949
rect 22260 12923 22266 12949
rect 22186 12922 22214 12923
rect 22238 12922 22266 12923
rect 22290 12922 22318 12950
rect 22342 12949 22370 12950
rect 22394 12949 22422 12950
rect 22342 12923 22348 12949
rect 22348 12923 22370 12949
rect 22394 12923 22410 12949
rect 22410 12923 22422 12949
rect 22342 12922 22370 12923
rect 22394 12922 22422 12923
rect 22446 12949 22474 12950
rect 22446 12923 22472 12949
rect 22472 12923 22474 12949
rect 22446 12922 22474 12923
rect 22498 12949 22526 12950
rect 22498 12923 22508 12949
rect 22508 12923 22526 12949
rect 22498 12922 22526 12923
rect 22526 12614 22554 12642
rect 22082 12165 22110 12166
rect 22082 12139 22100 12165
rect 22100 12139 22110 12165
rect 22082 12138 22110 12139
rect 22134 12165 22162 12166
rect 22134 12139 22136 12165
rect 22136 12139 22162 12165
rect 22134 12138 22162 12139
rect 22186 12165 22214 12166
rect 22238 12165 22266 12166
rect 22186 12139 22198 12165
rect 22198 12139 22214 12165
rect 22238 12139 22260 12165
rect 22260 12139 22266 12165
rect 22186 12138 22214 12139
rect 22238 12138 22266 12139
rect 22290 12138 22318 12166
rect 22342 12165 22370 12166
rect 22394 12165 22422 12166
rect 22342 12139 22348 12165
rect 22348 12139 22370 12165
rect 22394 12139 22410 12165
rect 22410 12139 22422 12165
rect 22342 12138 22370 12139
rect 22394 12138 22422 12139
rect 22446 12165 22474 12166
rect 22446 12139 22472 12165
rect 22472 12139 22474 12165
rect 22446 12138 22474 12139
rect 22498 12165 22526 12166
rect 22498 12139 22508 12165
rect 22508 12139 22526 12165
rect 22498 12138 22526 12139
rect 21182 11969 21210 11970
rect 21182 11943 21183 11969
rect 21183 11943 21209 11969
rect 21209 11943 21210 11969
rect 21182 11942 21210 11943
rect 22082 11381 22110 11382
rect 22082 11355 22100 11381
rect 22100 11355 22110 11381
rect 22082 11354 22110 11355
rect 22134 11381 22162 11382
rect 22134 11355 22136 11381
rect 22136 11355 22162 11381
rect 22134 11354 22162 11355
rect 22186 11381 22214 11382
rect 22238 11381 22266 11382
rect 22186 11355 22198 11381
rect 22198 11355 22214 11381
rect 22238 11355 22260 11381
rect 22260 11355 22266 11381
rect 22186 11354 22214 11355
rect 22238 11354 22266 11355
rect 22290 11354 22318 11382
rect 22342 11381 22370 11382
rect 22394 11381 22422 11382
rect 22342 11355 22348 11381
rect 22348 11355 22370 11381
rect 22394 11355 22410 11381
rect 22410 11355 22422 11381
rect 22342 11354 22370 11355
rect 22394 11354 22422 11355
rect 22446 11381 22474 11382
rect 22446 11355 22472 11381
rect 22472 11355 22474 11381
rect 22446 11354 22474 11355
rect 22498 11381 22526 11382
rect 22498 11355 22508 11381
rect 22508 11355 22526 11381
rect 22498 11354 22526 11355
rect 19582 10989 19610 10990
rect 19582 10963 19600 10989
rect 19600 10963 19610 10989
rect 19582 10962 19610 10963
rect 19634 10989 19662 10990
rect 19634 10963 19636 10989
rect 19636 10963 19662 10989
rect 19634 10962 19662 10963
rect 19686 10989 19714 10990
rect 19738 10989 19766 10990
rect 19686 10963 19698 10989
rect 19698 10963 19714 10989
rect 19738 10963 19760 10989
rect 19760 10963 19766 10989
rect 19686 10962 19714 10963
rect 19738 10962 19766 10963
rect 19790 10962 19818 10990
rect 19842 10989 19870 10990
rect 19894 10989 19922 10990
rect 19842 10963 19848 10989
rect 19848 10963 19870 10989
rect 19894 10963 19910 10989
rect 19910 10963 19922 10989
rect 19842 10962 19870 10963
rect 19894 10962 19922 10963
rect 19946 10989 19974 10990
rect 19946 10963 19972 10989
rect 19972 10963 19974 10989
rect 19946 10962 19974 10963
rect 19998 10989 20026 10990
rect 19998 10963 20008 10989
rect 20008 10963 20026 10989
rect 19998 10962 20026 10963
rect 19502 10318 19530 10346
rect 19950 10345 19978 10346
rect 19950 10319 19951 10345
rect 19951 10319 19977 10345
rect 19977 10319 19978 10345
rect 19950 10318 19978 10319
rect 19582 10205 19610 10206
rect 19582 10179 19600 10205
rect 19600 10179 19610 10205
rect 19582 10178 19610 10179
rect 19634 10205 19662 10206
rect 19634 10179 19636 10205
rect 19636 10179 19662 10205
rect 19634 10178 19662 10179
rect 19686 10205 19714 10206
rect 19738 10205 19766 10206
rect 19686 10179 19698 10205
rect 19698 10179 19714 10205
rect 19738 10179 19760 10205
rect 19760 10179 19766 10205
rect 19686 10178 19714 10179
rect 19738 10178 19766 10179
rect 19790 10178 19818 10206
rect 19842 10205 19870 10206
rect 19894 10205 19922 10206
rect 19842 10179 19848 10205
rect 19848 10179 19870 10205
rect 19894 10179 19910 10205
rect 19910 10179 19922 10205
rect 19842 10178 19870 10179
rect 19894 10178 19922 10179
rect 19946 10205 19974 10206
rect 19946 10179 19972 10205
rect 19972 10179 19974 10205
rect 19946 10178 19974 10179
rect 19998 10205 20026 10206
rect 19998 10179 20008 10205
rect 20008 10179 20026 10205
rect 19998 10178 20026 10179
rect 18942 10009 18970 10010
rect 18942 9983 18943 10009
rect 18943 9983 18969 10009
rect 18969 9983 18970 10009
rect 18942 9982 18970 9983
rect 19222 9617 19250 9618
rect 19222 9591 19223 9617
rect 19223 9591 19249 9617
rect 19249 9591 19250 9617
rect 19222 9590 19250 9591
rect 19582 9421 19610 9422
rect 19582 9395 19600 9421
rect 19600 9395 19610 9421
rect 19582 9394 19610 9395
rect 19634 9421 19662 9422
rect 19634 9395 19636 9421
rect 19636 9395 19662 9421
rect 19634 9394 19662 9395
rect 19686 9421 19714 9422
rect 19738 9421 19766 9422
rect 19686 9395 19698 9421
rect 19698 9395 19714 9421
rect 19738 9395 19760 9421
rect 19760 9395 19766 9421
rect 19686 9394 19714 9395
rect 19738 9394 19766 9395
rect 19790 9394 19818 9422
rect 19842 9421 19870 9422
rect 19894 9421 19922 9422
rect 19842 9395 19848 9421
rect 19848 9395 19870 9421
rect 19894 9395 19910 9421
rect 19910 9395 19922 9421
rect 19842 9394 19870 9395
rect 19894 9394 19922 9395
rect 19946 9421 19974 9422
rect 19946 9395 19972 9421
rect 19972 9395 19974 9421
rect 19946 9394 19974 9395
rect 19998 9421 20026 9422
rect 19998 9395 20008 9421
rect 20008 9395 20026 9421
rect 19998 9394 20026 9395
rect 19582 8637 19610 8638
rect 19582 8611 19600 8637
rect 19600 8611 19610 8637
rect 19582 8610 19610 8611
rect 19634 8637 19662 8638
rect 19634 8611 19636 8637
rect 19636 8611 19662 8637
rect 19634 8610 19662 8611
rect 19686 8637 19714 8638
rect 19738 8637 19766 8638
rect 19686 8611 19698 8637
rect 19698 8611 19714 8637
rect 19738 8611 19760 8637
rect 19760 8611 19766 8637
rect 19686 8610 19714 8611
rect 19738 8610 19766 8611
rect 19790 8610 19818 8638
rect 19842 8637 19870 8638
rect 19894 8637 19922 8638
rect 19842 8611 19848 8637
rect 19848 8611 19870 8637
rect 19894 8611 19910 8637
rect 19910 8611 19922 8637
rect 19842 8610 19870 8611
rect 19894 8610 19922 8611
rect 19946 8637 19974 8638
rect 19946 8611 19972 8637
rect 19972 8611 19974 8637
rect 19946 8610 19974 8611
rect 19998 8637 20026 8638
rect 19998 8611 20008 8637
rect 20008 8611 20026 8637
rect 19998 8610 20026 8611
rect 19582 7853 19610 7854
rect 19582 7827 19600 7853
rect 19600 7827 19610 7853
rect 19582 7826 19610 7827
rect 19634 7853 19662 7854
rect 19634 7827 19636 7853
rect 19636 7827 19662 7853
rect 19634 7826 19662 7827
rect 19686 7853 19714 7854
rect 19738 7853 19766 7854
rect 19686 7827 19698 7853
rect 19698 7827 19714 7853
rect 19738 7827 19760 7853
rect 19760 7827 19766 7853
rect 19686 7826 19714 7827
rect 19738 7826 19766 7827
rect 19790 7826 19818 7854
rect 19842 7853 19870 7854
rect 19894 7853 19922 7854
rect 19842 7827 19848 7853
rect 19848 7827 19870 7853
rect 19894 7827 19910 7853
rect 19910 7827 19922 7853
rect 19842 7826 19870 7827
rect 19894 7826 19922 7827
rect 19946 7853 19974 7854
rect 19946 7827 19972 7853
rect 19972 7827 19974 7853
rect 19946 7826 19974 7827
rect 19998 7853 20026 7854
rect 19998 7827 20008 7853
rect 20008 7827 20026 7853
rect 19998 7826 20026 7827
rect 19582 7069 19610 7070
rect 19582 7043 19600 7069
rect 19600 7043 19610 7069
rect 19582 7042 19610 7043
rect 19634 7069 19662 7070
rect 19634 7043 19636 7069
rect 19636 7043 19662 7069
rect 19634 7042 19662 7043
rect 19686 7069 19714 7070
rect 19738 7069 19766 7070
rect 19686 7043 19698 7069
rect 19698 7043 19714 7069
rect 19738 7043 19760 7069
rect 19760 7043 19766 7069
rect 19686 7042 19714 7043
rect 19738 7042 19766 7043
rect 19790 7042 19818 7070
rect 19842 7069 19870 7070
rect 19894 7069 19922 7070
rect 19842 7043 19848 7069
rect 19848 7043 19870 7069
rect 19894 7043 19910 7069
rect 19910 7043 19922 7069
rect 19842 7042 19870 7043
rect 19894 7042 19922 7043
rect 19946 7069 19974 7070
rect 19946 7043 19972 7069
rect 19972 7043 19974 7069
rect 19946 7042 19974 7043
rect 19998 7069 20026 7070
rect 19998 7043 20008 7069
rect 20008 7043 20026 7069
rect 19998 7042 20026 7043
rect 19582 6285 19610 6286
rect 19582 6259 19600 6285
rect 19600 6259 19610 6285
rect 19582 6258 19610 6259
rect 19634 6285 19662 6286
rect 19634 6259 19636 6285
rect 19636 6259 19662 6285
rect 19634 6258 19662 6259
rect 19686 6285 19714 6286
rect 19738 6285 19766 6286
rect 19686 6259 19698 6285
rect 19698 6259 19714 6285
rect 19738 6259 19760 6285
rect 19760 6259 19766 6285
rect 19686 6258 19714 6259
rect 19738 6258 19766 6259
rect 19790 6258 19818 6286
rect 19842 6285 19870 6286
rect 19894 6285 19922 6286
rect 19842 6259 19848 6285
rect 19848 6259 19870 6285
rect 19894 6259 19910 6285
rect 19910 6259 19922 6285
rect 19842 6258 19870 6259
rect 19894 6258 19922 6259
rect 19946 6285 19974 6286
rect 19946 6259 19972 6285
rect 19972 6259 19974 6285
rect 19946 6258 19974 6259
rect 19998 6285 20026 6286
rect 19998 6259 20008 6285
rect 20008 6259 20026 6285
rect 19998 6258 20026 6259
rect 19582 5501 19610 5502
rect 19582 5475 19600 5501
rect 19600 5475 19610 5501
rect 19582 5474 19610 5475
rect 19634 5501 19662 5502
rect 19634 5475 19636 5501
rect 19636 5475 19662 5501
rect 19634 5474 19662 5475
rect 19686 5501 19714 5502
rect 19738 5501 19766 5502
rect 19686 5475 19698 5501
rect 19698 5475 19714 5501
rect 19738 5475 19760 5501
rect 19760 5475 19766 5501
rect 19686 5474 19714 5475
rect 19738 5474 19766 5475
rect 19790 5474 19818 5502
rect 19842 5501 19870 5502
rect 19894 5501 19922 5502
rect 19842 5475 19848 5501
rect 19848 5475 19870 5501
rect 19894 5475 19910 5501
rect 19910 5475 19922 5501
rect 19842 5474 19870 5475
rect 19894 5474 19922 5475
rect 19946 5501 19974 5502
rect 19946 5475 19972 5501
rect 19972 5475 19974 5501
rect 19946 5474 19974 5475
rect 19998 5501 20026 5502
rect 19998 5475 20008 5501
rect 20008 5475 20026 5501
rect 19998 5474 20026 5475
rect 20230 5278 20258 5306
rect 20230 5054 20258 5082
rect 20566 10094 20594 10122
rect 19582 4717 19610 4718
rect 19582 4691 19600 4717
rect 19600 4691 19610 4717
rect 19582 4690 19610 4691
rect 19634 4717 19662 4718
rect 19634 4691 19636 4717
rect 19636 4691 19662 4717
rect 19634 4690 19662 4691
rect 19686 4717 19714 4718
rect 19738 4717 19766 4718
rect 19686 4691 19698 4717
rect 19698 4691 19714 4717
rect 19738 4691 19760 4717
rect 19760 4691 19766 4717
rect 19686 4690 19714 4691
rect 19738 4690 19766 4691
rect 19790 4690 19818 4718
rect 19842 4717 19870 4718
rect 19894 4717 19922 4718
rect 19842 4691 19848 4717
rect 19848 4691 19870 4717
rect 19894 4691 19910 4717
rect 19910 4691 19922 4717
rect 19842 4690 19870 4691
rect 19894 4690 19922 4691
rect 19946 4717 19974 4718
rect 19946 4691 19972 4717
rect 19972 4691 19974 4717
rect 19946 4690 19974 4691
rect 19998 4717 20026 4718
rect 19998 4691 20008 4717
rect 20008 4691 20026 4717
rect 19998 4690 20026 4691
rect 20118 4158 20146 4186
rect 19582 3933 19610 3934
rect 19582 3907 19600 3933
rect 19600 3907 19610 3933
rect 19582 3906 19610 3907
rect 19634 3933 19662 3934
rect 19634 3907 19636 3933
rect 19636 3907 19662 3933
rect 19634 3906 19662 3907
rect 19686 3933 19714 3934
rect 19738 3933 19766 3934
rect 19686 3907 19698 3933
rect 19698 3907 19714 3933
rect 19738 3907 19760 3933
rect 19760 3907 19766 3933
rect 19686 3906 19714 3907
rect 19738 3906 19766 3907
rect 19790 3906 19818 3934
rect 19842 3933 19870 3934
rect 19894 3933 19922 3934
rect 19842 3907 19848 3933
rect 19848 3907 19870 3933
rect 19894 3907 19910 3933
rect 19910 3907 19922 3933
rect 19842 3906 19870 3907
rect 19894 3906 19922 3907
rect 19946 3933 19974 3934
rect 19946 3907 19972 3933
rect 19972 3907 19974 3933
rect 19946 3906 19974 3907
rect 19998 3933 20026 3934
rect 19998 3907 20008 3933
rect 20008 3907 20026 3933
rect 19998 3906 20026 3907
rect 19166 3318 19194 3346
rect 19446 3345 19474 3346
rect 19446 3319 19447 3345
rect 19447 3319 19473 3345
rect 19473 3319 19474 3345
rect 19446 3318 19474 3319
rect 18886 2926 18914 2954
rect 21406 10345 21434 10346
rect 21406 10319 21407 10345
rect 21407 10319 21433 10345
rect 21433 10319 21434 10345
rect 21406 10318 21434 10319
rect 22082 10597 22110 10598
rect 22082 10571 22100 10597
rect 22100 10571 22110 10597
rect 22082 10570 22110 10571
rect 22134 10597 22162 10598
rect 22134 10571 22136 10597
rect 22136 10571 22162 10597
rect 22134 10570 22162 10571
rect 22186 10597 22214 10598
rect 22238 10597 22266 10598
rect 22186 10571 22198 10597
rect 22198 10571 22214 10597
rect 22238 10571 22260 10597
rect 22260 10571 22266 10597
rect 22186 10570 22214 10571
rect 22238 10570 22266 10571
rect 22290 10570 22318 10598
rect 22342 10597 22370 10598
rect 22394 10597 22422 10598
rect 22342 10571 22348 10597
rect 22348 10571 22370 10597
rect 22394 10571 22410 10597
rect 22410 10571 22422 10597
rect 22342 10570 22370 10571
rect 22394 10570 22422 10571
rect 22446 10597 22474 10598
rect 22446 10571 22472 10597
rect 22472 10571 22474 10597
rect 22446 10570 22474 10571
rect 22498 10597 22526 10598
rect 22498 10571 22508 10597
rect 22508 10571 22526 10597
rect 22498 10570 22526 10571
rect 21742 10318 21770 10346
rect 20790 6089 20818 6090
rect 20790 6063 20791 6089
rect 20791 6063 20817 6089
rect 20817 6063 20818 6089
rect 20790 6062 20818 6063
rect 20790 5305 20818 5306
rect 20790 5279 20791 5305
rect 20791 5279 20817 5305
rect 20817 5279 20818 5305
rect 20790 5278 20818 5279
rect 23926 11913 23954 11914
rect 23926 11887 23927 11913
rect 23927 11887 23953 11913
rect 23953 11887 23954 11913
rect 23926 11886 23954 11887
rect 22806 10878 22834 10906
rect 22806 10094 22834 10122
rect 21742 10009 21770 10010
rect 21742 9983 21743 10009
rect 21743 9983 21769 10009
rect 21769 9983 21770 10009
rect 21742 9982 21770 9983
rect 22694 10009 22722 10010
rect 22694 9983 22695 10009
rect 22695 9983 22721 10009
rect 22721 9983 22722 10009
rect 22694 9982 22722 9983
rect 22082 9813 22110 9814
rect 22082 9787 22100 9813
rect 22100 9787 22110 9813
rect 22082 9786 22110 9787
rect 22134 9813 22162 9814
rect 22134 9787 22136 9813
rect 22136 9787 22162 9813
rect 22134 9786 22162 9787
rect 22186 9813 22214 9814
rect 22238 9813 22266 9814
rect 22186 9787 22198 9813
rect 22198 9787 22214 9813
rect 22238 9787 22260 9813
rect 22260 9787 22266 9813
rect 22186 9786 22214 9787
rect 22238 9786 22266 9787
rect 22290 9786 22318 9814
rect 22342 9813 22370 9814
rect 22394 9813 22422 9814
rect 22342 9787 22348 9813
rect 22348 9787 22370 9813
rect 22394 9787 22410 9813
rect 22410 9787 22422 9813
rect 22342 9786 22370 9787
rect 22394 9786 22422 9787
rect 22446 9813 22474 9814
rect 22446 9787 22472 9813
rect 22472 9787 22474 9813
rect 22446 9786 22474 9787
rect 22498 9813 22526 9814
rect 22498 9787 22508 9813
rect 22508 9787 22526 9813
rect 22498 9786 22526 9787
rect 22918 10009 22946 10010
rect 22918 9983 22919 10009
rect 22919 9983 22945 10009
rect 22945 9983 22946 10009
rect 22918 9982 22946 9983
rect 23366 9982 23394 10010
rect 23422 9617 23450 9618
rect 23422 9591 23423 9617
rect 23423 9591 23449 9617
rect 23449 9591 23450 9617
rect 23422 9590 23450 9591
rect 22750 9254 22778 9282
rect 22082 9029 22110 9030
rect 22082 9003 22100 9029
rect 22100 9003 22110 9029
rect 22082 9002 22110 9003
rect 22134 9029 22162 9030
rect 22134 9003 22136 9029
rect 22136 9003 22162 9029
rect 22134 9002 22162 9003
rect 22186 9029 22214 9030
rect 22238 9029 22266 9030
rect 22186 9003 22198 9029
rect 22198 9003 22214 9029
rect 22238 9003 22260 9029
rect 22260 9003 22266 9029
rect 22186 9002 22214 9003
rect 22238 9002 22266 9003
rect 22290 9002 22318 9030
rect 22342 9029 22370 9030
rect 22394 9029 22422 9030
rect 22342 9003 22348 9029
rect 22348 9003 22370 9029
rect 22394 9003 22410 9029
rect 22410 9003 22422 9029
rect 22342 9002 22370 9003
rect 22394 9002 22422 9003
rect 22446 9029 22474 9030
rect 22446 9003 22472 9029
rect 22472 9003 22474 9029
rect 22446 9002 22474 9003
rect 22498 9029 22526 9030
rect 22498 9003 22508 9029
rect 22508 9003 22526 9029
rect 22498 9002 22526 9003
rect 22082 8245 22110 8246
rect 22082 8219 22100 8245
rect 22100 8219 22110 8245
rect 22082 8218 22110 8219
rect 22134 8245 22162 8246
rect 22134 8219 22136 8245
rect 22136 8219 22162 8245
rect 22134 8218 22162 8219
rect 22186 8245 22214 8246
rect 22238 8245 22266 8246
rect 22186 8219 22198 8245
rect 22198 8219 22214 8245
rect 22238 8219 22260 8245
rect 22260 8219 22266 8245
rect 22186 8218 22214 8219
rect 22238 8218 22266 8219
rect 22290 8218 22318 8246
rect 22342 8245 22370 8246
rect 22394 8245 22422 8246
rect 22342 8219 22348 8245
rect 22348 8219 22370 8245
rect 22394 8219 22410 8245
rect 22410 8219 22422 8245
rect 22342 8218 22370 8219
rect 22394 8218 22422 8219
rect 22446 8245 22474 8246
rect 22446 8219 22472 8245
rect 22472 8219 22474 8245
rect 22446 8218 22474 8219
rect 22498 8245 22526 8246
rect 22498 8219 22508 8245
rect 22508 8219 22526 8245
rect 22498 8218 22526 8219
rect 22082 7461 22110 7462
rect 22082 7435 22100 7461
rect 22100 7435 22110 7461
rect 22082 7434 22110 7435
rect 22134 7461 22162 7462
rect 22134 7435 22136 7461
rect 22136 7435 22162 7461
rect 22134 7434 22162 7435
rect 22186 7461 22214 7462
rect 22238 7461 22266 7462
rect 22186 7435 22198 7461
rect 22198 7435 22214 7461
rect 22238 7435 22260 7461
rect 22260 7435 22266 7461
rect 22186 7434 22214 7435
rect 22238 7434 22266 7435
rect 22290 7434 22318 7462
rect 22342 7461 22370 7462
rect 22394 7461 22422 7462
rect 22342 7435 22348 7461
rect 22348 7435 22370 7461
rect 22394 7435 22410 7461
rect 22410 7435 22422 7461
rect 22342 7434 22370 7435
rect 22394 7434 22422 7435
rect 22446 7461 22474 7462
rect 22446 7435 22472 7461
rect 22472 7435 22474 7461
rect 22446 7434 22474 7435
rect 22498 7461 22526 7462
rect 22498 7435 22508 7461
rect 22508 7435 22526 7461
rect 22498 7434 22526 7435
rect 22082 6677 22110 6678
rect 22082 6651 22100 6677
rect 22100 6651 22110 6677
rect 22082 6650 22110 6651
rect 22134 6677 22162 6678
rect 22134 6651 22136 6677
rect 22136 6651 22162 6677
rect 22134 6650 22162 6651
rect 22186 6677 22214 6678
rect 22238 6677 22266 6678
rect 22186 6651 22198 6677
rect 22198 6651 22214 6677
rect 22238 6651 22260 6677
rect 22260 6651 22266 6677
rect 22186 6650 22214 6651
rect 22238 6650 22266 6651
rect 22290 6650 22318 6678
rect 22342 6677 22370 6678
rect 22394 6677 22422 6678
rect 22342 6651 22348 6677
rect 22348 6651 22370 6677
rect 22394 6651 22410 6677
rect 22410 6651 22422 6677
rect 22342 6650 22370 6651
rect 22394 6650 22422 6651
rect 22446 6677 22474 6678
rect 22446 6651 22472 6677
rect 22472 6651 22474 6677
rect 22446 6650 22474 6651
rect 22498 6677 22526 6678
rect 22498 6651 22508 6677
rect 22508 6651 22526 6677
rect 22498 6650 22526 6651
rect 23422 9225 23450 9226
rect 23422 9199 23423 9225
rect 23423 9199 23449 9225
rect 23449 9199 23450 9225
rect 23422 9198 23450 9199
rect 23702 9198 23730 9226
rect 23422 8441 23450 8442
rect 23422 8415 23423 8441
rect 23423 8415 23449 8441
rect 23449 8415 23450 8441
rect 23422 8414 23450 8415
rect 22246 6089 22274 6090
rect 22246 6063 22247 6089
rect 22247 6063 22273 6089
rect 22273 6063 22274 6089
rect 22246 6062 22274 6063
rect 22582 6062 22610 6090
rect 21462 6006 21490 6034
rect 23086 6342 23114 6370
rect 22694 6006 22722 6034
rect 22082 5893 22110 5894
rect 22082 5867 22100 5893
rect 22100 5867 22110 5893
rect 22082 5866 22110 5867
rect 22134 5893 22162 5894
rect 22134 5867 22136 5893
rect 22136 5867 22162 5893
rect 22134 5866 22162 5867
rect 22186 5893 22214 5894
rect 22238 5893 22266 5894
rect 22186 5867 22198 5893
rect 22198 5867 22214 5893
rect 22238 5867 22260 5893
rect 22260 5867 22266 5893
rect 22186 5866 22214 5867
rect 22238 5866 22266 5867
rect 22290 5866 22318 5894
rect 22342 5893 22370 5894
rect 22394 5893 22422 5894
rect 22342 5867 22348 5893
rect 22348 5867 22370 5893
rect 22394 5867 22410 5893
rect 22410 5867 22422 5893
rect 22342 5866 22370 5867
rect 22394 5866 22422 5867
rect 22446 5893 22474 5894
rect 22446 5867 22472 5893
rect 22472 5867 22474 5893
rect 22446 5866 22474 5867
rect 22498 5893 22526 5894
rect 22498 5867 22508 5893
rect 22508 5867 22526 5893
rect 22498 5866 22526 5867
rect 22082 5109 22110 5110
rect 22082 5083 22100 5109
rect 22100 5083 22110 5109
rect 22082 5082 22110 5083
rect 22134 5109 22162 5110
rect 22134 5083 22136 5109
rect 22136 5083 22162 5109
rect 22134 5082 22162 5083
rect 22186 5109 22214 5110
rect 22238 5109 22266 5110
rect 22186 5083 22198 5109
rect 22198 5083 22214 5109
rect 22238 5083 22260 5109
rect 22260 5083 22266 5109
rect 22186 5082 22214 5083
rect 22238 5082 22266 5083
rect 22290 5082 22318 5110
rect 22342 5109 22370 5110
rect 22394 5109 22422 5110
rect 22342 5083 22348 5109
rect 22348 5083 22370 5109
rect 22394 5083 22410 5109
rect 22410 5083 22422 5109
rect 22342 5082 22370 5083
rect 22394 5082 22422 5083
rect 22446 5109 22474 5110
rect 22446 5083 22472 5109
rect 22472 5083 22474 5109
rect 22446 5082 22474 5083
rect 22498 5109 22526 5110
rect 22498 5083 22508 5109
rect 22508 5083 22526 5109
rect 22498 5082 22526 5083
rect 20566 3374 20594 3402
rect 21406 4494 21434 4522
rect 21350 4158 21378 4186
rect 21798 4521 21826 4522
rect 21798 4495 21799 4521
rect 21799 4495 21825 4521
rect 21825 4495 21826 4521
rect 21798 4494 21826 4495
rect 22082 4325 22110 4326
rect 22082 4299 22100 4325
rect 22100 4299 22110 4325
rect 22082 4298 22110 4299
rect 22134 4325 22162 4326
rect 22134 4299 22136 4325
rect 22136 4299 22162 4325
rect 22134 4298 22162 4299
rect 22186 4325 22214 4326
rect 22238 4325 22266 4326
rect 22186 4299 22198 4325
rect 22198 4299 22214 4325
rect 22238 4299 22260 4325
rect 22260 4299 22266 4325
rect 22186 4298 22214 4299
rect 22238 4298 22266 4299
rect 22290 4298 22318 4326
rect 22342 4325 22370 4326
rect 22394 4325 22422 4326
rect 22342 4299 22348 4325
rect 22348 4299 22370 4325
rect 22394 4299 22410 4325
rect 22410 4299 22422 4325
rect 22342 4298 22370 4299
rect 22394 4298 22422 4299
rect 22446 4325 22474 4326
rect 22446 4299 22472 4325
rect 22472 4299 22474 4325
rect 22446 4298 22474 4299
rect 22498 4325 22526 4326
rect 22498 4299 22508 4325
rect 22508 4299 22526 4325
rect 22498 4298 22526 4299
rect 19582 3149 19610 3150
rect 19582 3123 19600 3149
rect 19600 3123 19610 3149
rect 19582 3122 19610 3123
rect 19634 3149 19662 3150
rect 19634 3123 19636 3149
rect 19636 3123 19662 3149
rect 19634 3122 19662 3123
rect 19686 3149 19714 3150
rect 19738 3149 19766 3150
rect 19686 3123 19698 3149
rect 19698 3123 19714 3149
rect 19738 3123 19760 3149
rect 19760 3123 19766 3149
rect 19686 3122 19714 3123
rect 19738 3122 19766 3123
rect 19790 3122 19818 3150
rect 19842 3149 19870 3150
rect 19894 3149 19922 3150
rect 19842 3123 19848 3149
rect 19848 3123 19870 3149
rect 19894 3123 19910 3149
rect 19910 3123 19922 3149
rect 19842 3122 19870 3123
rect 19894 3122 19922 3123
rect 19946 3149 19974 3150
rect 19946 3123 19972 3149
rect 19972 3123 19974 3149
rect 19946 3122 19974 3123
rect 19998 3149 20026 3150
rect 19998 3123 20008 3149
rect 20008 3123 20026 3149
rect 19998 3122 20026 3123
rect 18774 2478 18802 2506
rect 18550 2142 18578 2170
rect 19222 2590 19250 2618
rect 20118 2561 20146 2562
rect 20118 2535 20119 2561
rect 20119 2535 20145 2561
rect 20145 2535 20146 2561
rect 20118 2534 20146 2535
rect 20230 2478 20258 2506
rect 21686 4158 21714 4186
rect 21014 3345 21042 3346
rect 21014 3319 21015 3345
rect 21015 3319 21041 3345
rect 21041 3319 21042 3345
rect 21014 3318 21042 3319
rect 22694 4521 22722 4522
rect 22694 4495 22695 4521
rect 22695 4495 22721 4521
rect 22721 4495 22722 4521
rect 22694 4494 22722 4495
rect 22918 4521 22946 4522
rect 22918 4495 22919 4521
rect 22919 4495 22945 4521
rect 22945 4495 22946 4521
rect 22918 4494 22946 4495
rect 22750 4129 22778 4130
rect 22750 4103 22751 4129
rect 22751 4103 22777 4129
rect 22777 4103 22778 4129
rect 22750 4102 22778 4103
rect 22082 3541 22110 3542
rect 22082 3515 22100 3541
rect 22100 3515 22110 3541
rect 22082 3514 22110 3515
rect 22134 3541 22162 3542
rect 22134 3515 22136 3541
rect 22136 3515 22162 3541
rect 22134 3514 22162 3515
rect 22186 3541 22214 3542
rect 22238 3541 22266 3542
rect 22186 3515 22198 3541
rect 22198 3515 22214 3541
rect 22238 3515 22260 3541
rect 22260 3515 22266 3541
rect 22186 3514 22214 3515
rect 22238 3514 22266 3515
rect 22290 3514 22318 3542
rect 22342 3541 22370 3542
rect 22394 3541 22422 3542
rect 22342 3515 22348 3541
rect 22348 3515 22370 3541
rect 22394 3515 22410 3541
rect 22410 3515 22422 3541
rect 22342 3514 22370 3515
rect 22394 3514 22422 3515
rect 22446 3541 22474 3542
rect 22446 3515 22472 3541
rect 22472 3515 22474 3541
rect 22446 3514 22474 3515
rect 22498 3541 22526 3542
rect 22498 3515 22508 3541
rect 22508 3515 22526 3541
rect 22498 3514 22526 3515
rect 21742 3374 21770 3402
rect 21182 3318 21210 3346
rect 20790 2953 20818 2954
rect 20790 2927 20791 2953
rect 20791 2927 20817 2953
rect 20817 2927 20818 2953
rect 20790 2926 20818 2927
rect 21406 3038 21434 3066
rect 20790 2478 20818 2506
rect 19582 2365 19610 2366
rect 19582 2339 19600 2365
rect 19600 2339 19610 2365
rect 19582 2338 19610 2339
rect 19634 2365 19662 2366
rect 19634 2339 19636 2365
rect 19636 2339 19662 2365
rect 19634 2338 19662 2339
rect 19686 2365 19714 2366
rect 19738 2365 19766 2366
rect 19686 2339 19698 2365
rect 19698 2339 19714 2365
rect 19738 2339 19760 2365
rect 19760 2339 19766 2365
rect 19686 2338 19714 2339
rect 19738 2338 19766 2339
rect 19790 2338 19818 2366
rect 19842 2365 19870 2366
rect 19894 2365 19922 2366
rect 19842 2339 19848 2365
rect 19848 2339 19870 2365
rect 19894 2339 19910 2365
rect 19910 2339 19922 2365
rect 19842 2338 19870 2339
rect 19894 2338 19922 2339
rect 19946 2365 19974 2366
rect 19946 2339 19972 2365
rect 19972 2339 19974 2365
rect 19946 2338 19974 2339
rect 19998 2365 20026 2366
rect 19998 2339 20008 2365
rect 20008 2339 20026 2365
rect 19998 2338 20026 2339
rect 18774 2142 18802 2170
rect 20958 2590 20986 2618
rect 21406 2534 21434 2562
rect 20118 1750 20146 1778
rect 19582 1581 19610 1582
rect 19582 1555 19600 1581
rect 19600 1555 19610 1581
rect 19582 1554 19610 1555
rect 19634 1581 19662 1582
rect 19634 1555 19636 1581
rect 19636 1555 19662 1581
rect 19634 1554 19662 1555
rect 19686 1581 19714 1582
rect 19738 1581 19766 1582
rect 19686 1555 19698 1581
rect 19698 1555 19714 1581
rect 19738 1555 19760 1581
rect 19760 1555 19766 1581
rect 19686 1554 19714 1555
rect 19738 1554 19766 1555
rect 19790 1554 19818 1582
rect 19842 1581 19870 1582
rect 19894 1581 19922 1582
rect 19842 1555 19848 1581
rect 19848 1555 19870 1581
rect 19894 1555 19910 1581
rect 19910 1555 19922 1581
rect 19842 1554 19870 1555
rect 19894 1554 19922 1555
rect 19946 1581 19974 1582
rect 19946 1555 19972 1581
rect 19972 1555 19974 1581
rect 19946 1554 19974 1555
rect 19998 1581 20026 1582
rect 19998 1555 20008 1581
rect 20008 1555 20026 1581
rect 19998 1554 20026 1555
rect 18494 1470 18522 1498
rect 21182 1777 21210 1778
rect 21182 1751 21183 1777
rect 21183 1751 21209 1777
rect 21209 1751 21210 1777
rect 21182 1750 21210 1751
rect 22806 3374 22834 3402
rect 22246 2953 22274 2954
rect 22246 2927 22247 2953
rect 22247 2927 22273 2953
rect 22273 2927 22274 2953
rect 22246 2926 22274 2927
rect 22582 2926 22610 2954
rect 22082 2757 22110 2758
rect 22082 2731 22100 2757
rect 22100 2731 22110 2757
rect 22082 2730 22110 2731
rect 22134 2757 22162 2758
rect 22134 2731 22136 2757
rect 22136 2731 22162 2757
rect 22134 2730 22162 2731
rect 22186 2757 22214 2758
rect 22238 2757 22266 2758
rect 22186 2731 22198 2757
rect 22198 2731 22214 2757
rect 22238 2731 22260 2757
rect 22260 2731 22266 2757
rect 22186 2730 22214 2731
rect 22238 2730 22266 2731
rect 22290 2730 22318 2758
rect 22342 2757 22370 2758
rect 22394 2757 22422 2758
rect 22342 2731 22348 2757
rect 22348 2731 22370 2757
rect 22394 2731 22410 2757
rect 22410 2731 22422 2757
rect 22342 2730 22370 2731
rect 22394 2730 22422 2731
rect 22446 2757 22474 2758
rect 22446 2731 22472 2757
rect 22472 2731 22474 2757
rect 22446 2730 22474 2731
rect 22498 2757 22526 2758
rect 22498 2731 22508 2757
rect 22508 2731 22526 2757
rect 22498 2730 22526 2731
rect 22750 2422 22778 2450
rect 22082 1973 22110 1974
rect 22082 1947 22100 1973
rect 22100 1947 22110 1973
rect 22082 1946 22110 1947
rect 22134 1973 22162 1974
rect 22134 1947 22136 1973
rect 22136 1947 22162 1973
rect 22134 1946 22162 1947
rect 22186 1973 22214 1974
rect 22238 1973 22266 1974
rect 22186 1947 22198 1973
rect 22198 1947 22214 1973
rect 22238 1947 22260 1973
rect 22260 1947 22266 1973
rect 22186 1946 22214 1947
rect 22238 1946 22266 1947
rect 22290 1946 22318 1974
rect 22342 1973 22370 1974
rect 22394 1973 22422 1974
rect 22342 1947 22348 1973
rect 22348 1947 22370 1973
rect 22394 1947 22410 1973
rect 22410 1947 22422 1973
rect 22342 1946 22370 1947
rect 22394 1946 22422 1947
rect 22446 1973 22474 1974
rect 22446 1947 22472 1973
rect 22472 1947 22474 1973
rect 22446 1946 22474 1947
rect 22498 1973 22526 1974
rect 22498 1947 22508 1973
rect 22508 1947 22526 1973
rect 22498 1946 22526 1947
rect 22470 1806 22498 1834
rect 22862 1750 22890 1778
rect 21798 1694 21826 1722
rect 23198 4494 23226 4522
rect 23422 4046 23450 4074
rect 23198 3374 23226 3402
rect 23422 3374 23450 3402
rect 23198 2561 23226 2562
rect 23198 2535 23199 2561
rect 23199 2535 23225 2561
rect 23225 2535 23226 2561
rect 23198 2534 23226 2535
rect 23534 2561 23562 2562
rect 23534 2535 23535 2561
rect 23535 2535 23561 2561
rect 23561 2535 23562 2561
rect 23534 2534 23562 2535
rect 23086 1750 23114 1778
rect 24430 16254 24458 16282
rect 27082 16085 27110 16086
rect 27082 16059 27100 16085
rect 27100 16059 27110 16085
rect 27082 16058 27110 16059
rect 27134 16085 27162 16086
rect 27134 16059 27136 16085
rect 27136 16059 27162 16085
rect 27134 16058 27162 16059
rect 27186 16085 27214 16086
rect 27238 16085 27266 16086
rect 27186 16059 27198 16085
rect 27198 16059 27214 16085
rect 27238 16059 27260 16085
rect 27260 16059 27266 16085
rect 27186 16058 27214 16059
rect 27238 16058 27266 16059
rect 27290 16058 27318 16086
rect 27342 16085 27370 16086
rect 27394 16085 27422 16086
rect 27342 16059 27348 16085
rect 27348 16059 27370 16085
rect 27394 16059 27410 16085
rect 27410 16059 27422 16085
rect 27342 16058 27370 16059
rect 27394 16058 27422 16059
rect 27446 16085 27474 16086
rect 27446 16059 27472 16085
rect 27472 16059 27474 16085
rect 27446 16058 27474 16059
rect 27498 16085 27526 16086
rect 27498 16059 27508 16085
rect 27508 16059 27526 16085
rect 27498 16058 27526 16059
rect 24582 15693 24610 15694
rect 24582 15667 24600 15693
rect 24600 15667 24610 15693
rect 24582 15666 24610 15667
rect 24634 15693 24662 15694
rect 24634 15667 24636 15693
rect 24636 15667 24662 15693
rect 24634 15666 24662 15667
rect 24686 15693 24714 15694
rect 24738 15693 24766 15694
rect 24686 15667 24698 15693
rect 24698 15667 24714 15693
rect 24738 15667 24760 15693
rect 24760 15667 24766 15693
rect 24686 15666 24714 15667
rect 24738 15666 24766 15667
rect 24790 15666 24818 15694
rect 24842 15693 24870 15694
rect 24894 15693 24922 15694
rect 24842 15667 24848 15693
rect 24848 15667 24870 15693
rect 24894 15667 24910 15693
rect 24910 15667 24922 15693
rect 24842 15666 24870 15667
rect 24894 15666 24922 15667
rect 24946 15693 24974 15694
rect 24946 15667 24972 15693
rect 24972 15667 24974 15693
rect 24946 15666 24974 15667
rect 24998 15693 25026 15694
rect 24998 15667 25008 15693
rect 25008 15667 25026 15693
rect 24998 15666 25026 15667
rect 27082 15301 27110 15302
rect 27082 15275 27100 15301
rect 27100 15275 27110 15301
rect 27082 15274 27110 15275
rect 27134 15301 27162 15302
rect 27134 15275 27136 15301
rect 27136 15275 27162 15301
rect 27134 15274 27162 15275
rect 27186 15301 27214 15302
rect 27238 15301 27266 15302
rect 27186 15275 27198 15301
rect 27198 15275 27214 15301
rect 27238 15275 27260 15301
rect 27260 15275 27266 15301
rect 27186 15274 27214 15275
rect 27238 15274 27266 15275
rect 27290 15274 27318 15302
rect 27342 15301 27370 15302
rect 27394 15301 27422 15302
rect 27342 15275 27348 15301
rect 27348 15275 27370 15301
rect 27394 15275 27410 15301
rect 27410 15275 27422 15301
rect 27342 15274 27370 15275
rect 27394 15274 27422 15275
rect 27446 15301 27474 15302
rect 27446 15275 27472 15301
rect 27472 15275 27474 15301
rect 27446 15274 27474 15275
rect 27498 15301 27526 15302
rect 27498 15275 27508 15301
rect 27508 15275 27526 15301
rect 27498 15274 27526 15275
rect 24582 14909 24610 14910
rect 24582 14883 24600 14909
rect 24600 14883 24610 14909
rect 24582 14882 24610 14883
rect 24634 14909 24662 14910
rect 24634 14883 24636 14909
rect 24636 14883 24662 14909
rect 24634 14882 24662 14883
rect 24686 14909 24714 14910
rect 24738 14909 24766 14910
rect 24686 14883 24698 14909
rect 24698 14883 24714 14909
rect 24738 14883 24760 14909
rect 24760 14883 24766 14909
rect 24686 14882 24714 14883
rect 24738 14882 24766 14883
rect 24790 14882 24818 14910
rect 24842 14909 24870 14910
rect 24894 14909 24922 14910
rect 24842 14883 24848 14909
rect 24848 14883 24870 14909
rect 24894 14883 24910 14909
rect 24910 14883 24922 14909
rect 24842 14882 24870 14883
rect 24894 14882 24922 14883
rect 24946 14909 24974 14910
rect 24946 14883 24972 14909
rect 24972 14883 24974 14909
rect 24946 14882 24974 14883
rect 24998 14909 25026 14910
rect 24998 14883 25008 14909
rect 25008 14883 25026 14909
rect 24998 14882 25026 14883
rect 24486 14321 24514 14322
rect 24486 14295 24487 14321
rect 24487 14295 24513 14321
rect 24513 14295 24514 14321
rect 24486 14294 24514 14295
rect 24582 14125 24610 14126
rect 24582 14099 24600 14125
rect 24600 14099 24610 14125
rect 24582 14098 24610 14099
rect 24634 14125 24662 14126
rect 24634 14099 24636 14125
rect 24636 14099 24662 14125
rect 24634 14098 24662 14099
rect 24686 14125 24714 14126
rect 24738 14125 24766 14126
rect 24686 14099 24698 14125
rect 24698 14099 24714 14125
rect 24738 14099 24760 14125
rect 24760 14099 24766 14125
rect 24686 14098 24714 14099
rect 24738 14098 24766 14099
rect 24790 14098 24818 14126
rect 24842 14125 24870 14126
rect 24894 14125 24922 14126
rect 24842 14099 24848 14125
rect 24848 14099 24870 14125
rect 24894 14099 24910 14125
rect 24910 14099 24922 14125
rect 24842 14098 24870 14099
rect 24894 14098 24922 14099
rect 24946 14125 24974 14126
rect 24946 14099 24972 14125
rect 24972 14099 24974 14125
rect 24946 14098 24974 14099
rect 24998 14125 25026 14126
rect 24998 14099 25008 14125
rect 25008 14099 25026 14125
rect 24998 14098 25026 14099
rect 24582 13341 24610 13342
rect 24582 13315 24600 13341
rect 24600 13315 24610 13341
rect 24582 13314 24610 13315
rect 24634 13341 24662 13342
rect 24634 13315 24636 13341
rect 24636 13315 24662 13341
rect 24634 13314 24662 13315
rect 24686 13341 24714 13342
rect 24738 13341 24766 13342
rect 24686 13315 24698 13341
rect 24698 13315 24714 13341
rect 24738 13315 24760 13341
rect 24760 13315 24766 13341
rect 24686 13314 24714 13315
rect 24738 13314 24766 13315
rect 24790 13314 24818 13342
rect 24842 13341 24870 13342
rect 24894 13341 24922 13342
rect 24842 13315 24848 13341
rect 24848 13315 24870 13341
rect 24894 13315 24910 13341
rect 24910 13315 24922 13341
rect 24842 13314 24870 13315
rect 24894 13314 24922 13315
rect 24946 13341 24974 13342
rect 24946 13315 24972 13341
rect 24972 13315 24974 13341
rect 24946 13314 24974 13315
rect 24998 13341 25026 13342
rect 24998 13315 25008 13341
rect 25008 13315 25026 13341
rect 24998 13314 25026 13315
rect 24486 13118 24514 13146
rect 27082 14517 27110 14518
rect 27082 14491 27100 14517
rect 27100 14491 27110 14517
rect 27082 14490 27110 14491
rect 27134 14517 27162 14518
rect 27134 14491 27136 14517
rect 27136 14491 27162 14517
rect 27134 14490 27162 14491
rect 27186 14517 27214 14518
rect 27238 14517 27266 14518
rect 27186 14491 27198 14517
rect 27198 14491 27214 14517
rect 27238 14491 27260 14517
rect 27260 14491 27266 14517
rect 27186 14490 27214 14491
rect 27238 14490 27266 14491
rect 27290 14490 27318 14518
rect 27342 14517 27370 14518
rect 27394 14517 27422 14518
rect 27342 14491 27348 14517
rect 27348 14491 27370 14517
rect 27394 14491 27410 14517
rect 27410 14491 27422 14517
rect 27342 14490 27370 14491
rect 27394 14490 27422 14491
rect 27446 14517 27474 14518
rect 27446 14491 27472 14517
rect 27472 14491 27474 14517
rect 27446 14490 27474 14491
rect 27498 14517 27526 14518
rect 27498 14491 27508 14517
rect 27508 14491 27526 14517
rect 27498 14490 27526 14491
rect 25382 14265 25410 14266
rect 25382 14239 25383 14265
rect 25383 14239 25409 14265
rect 25409 14239 25410 14265
rect 25382 14238 25410 14239
rect 25382 13537 25410 13538
rect 25382 13511 25383 13537
rect 25383 13511 25409 13537
rect 25409 13511 25410 13537
rect 25382 13510 25410 13511
rect 26222 13846 26250 13874
rect 27398 13985 27426 13986
rect 27398 13959 27399 13985
rect 27399 13959 27425 13985
rect 27425 13959 27426 13985
rect 27398 13958 27426 13959
rect 26726 13846 26754 13874
rect 25942 13510 25970 13538
rect 25046 13145 25074 13146
rect 25046 13119 25047 13145
rect 25047 13119 25073 13145
rect 25073 13119 25074 13145
rect 25046 13118 25074 13119
rect 27082 13733 27110 13734
rect 27082 13707 27100 13733
rect 27100 13707 27110 13733
rect 27082 13706 27110 13707
rect 27134 13733 27162 13734
rect 27134 13707 27136 13733
rect 27136 13707 27162 13733
rect 27134 13706 27162 13707
rect 27186 13733 27214 13734
rect 27238 13733 27266 13734
rect 27186 13707 27198 13733
rect 27198 13707 27214 13733
rect 27238 13707 27260 13733
rect 27260 13707 27266 13733
rect 27186 13706 27214 13707
rect 27238 13706 27266 13707
rect 27290 13706 27318 13734
rect 27342 13733 27370 13734
rect 27394 13733 27422 13734
rect 27342 13707 27348 13733
rect 27348 13707 27370 13733
rect 27394 13707 27410 13733
rect 27410 13707 27422 13733
rect 27342 13706 27370 13707
rect 27394 13706 27422 13707
rect 27446 13733 27474 13734
rect 27446 13707 27472 13733
rect 27472 13707 27474 13733
rect 27446 13706 27474 13707
rect 27498 13733 27526 13734
rect 27498 13707 27508 13733
rect 27508 13707 27526 13733
rect 27498 13706 27526 13707
rect 26726 13537 26754 13538
rect 26726 13511 26727 13537
rect 26727 13511 26753 13537
rect 26753 13511 26754 13537
rect 26726 13510 26754 13511
rect 24582 12557 24610 12558
rect 24582 12531 24600 12557
rect 24600 12531 24610 12557
rect 24582 12530 24610 12531
rect 24634 12557 24662 12558
rect 24634 12531 24636 12557
rect 24636 12531 24662 12557
rect 24634 12530 24662 12531
rect 24686 12557 24714 12558
rect 24738 12557 24766 12558
rect 24686 12531 24698 12557
rect 24698 12531 24714 12557
rect 24738 12531 24760 12557
rect 24760 12531 24766 12557
rect 24686 12530 24714 12531
rect 24738 12530 24766 12531
rect 24790 12530 24818 12558
rect 24842 12557 24870 12558
rect 24894 12557 24922 12558
rect 24842 12531 24848 12557
rect 24848 12531 24870 12557
rect 24894 12531 24910 12557
rect 24910 12531 24922 12557
rect 24842 12530 24870 12531
rect 24894 12530 24922 12531
rect 24946 12557 24974 12558
rect 24946 12531 24972 12557
rect 24972 12531 24974 12557
rect 24946 12530 24974 12531
rect 24998 12557 25026 12558
rect 24998 12531 25008 12557
rect 25008 12531 25026 12557
rect 24998 12530 25026 12531
rect 25158 11913 25186 11914
rect 25158 11887 25159 11913
rect 25159 11887 25185 11913
rect 25185 11887 25186 11913
rect 25158 11886 25186 11887
rect 24582 11773 24610 11774
rect 24582 11747 24600 11773
rect 24600 11747 24610 11773
rect 24582 11746 24610 11747
rect 24634 11773 24662 11774
rect 24634 11747 24636 11773
rect 24636 11747 24662 11773
rect 24634 11746 24662 11747
rect 24686 11773 24714 11774
rect 24738 11773 24766 11774
rect 24686 11747 24698 11773
rect 24698 11747 24714 11773
rect 24738 11747 24760 11773
rect 24760 11747 24766 11773
rect 24686 11746 24714 11747
rect 24738 11746 24766 11747
rect 24790 11746 24818 11774
rect 24842 11773 24870 11774
rect 24894 11773 24922 11774
rect 24842 11747 24848 11773
rect 24848 11747 24870 11773
rect 24894 11747 24910 11773
rect 24910 11747 24922 11773
rect 24842 11746 24870 11747
rect 24894 11746 24922 11747
rect 24946 11773 24974 11774
rect 24946 11747 24972 11773
rect 24972 11747 24974 11773
rect 24946 11746 24974 11747
rect 24998 11773 25026 11774
rect 24998 11747 25008 11773
rect 25008 11747 25026 11773
rect 24998 11746 25026 11747
rect 25158 11774 25186 11802
rect 25998 12334 26026 12362
rect 24582 10989 24610 10990
rect 24582 10963 24600 10989
rect 24600 10963 24610 10989
rect 24582 10962 24610 10963
rect 24634 10989 24662 10990
rect 24634 10963 24636 10989
rect 24636 10963 24662 10989
rect 24634 10962 24662 10963
rect 24686 10989 24714 10990
rect 24738 10989 24766 10990
rect 24686 10963 24698 10989
rect 24698 10963 24714 10989
rect 24738 10963 24760 10989
rect 24760 10963 24766 10989
rect 24686 10962 24714 10963
rect 24738 10962 24766 10963
rect 24790 10962 24818 10990
rect 24842 10989 24870 10990
rect 24894 10989 24922 10990
rect 24842 10963 24848 10989
rect 24848 10963 24870 10989
rect 24894 10963 24910 10989
rect 24910 10963 24922 10989
rect 24842 10962 24870 10963
rect 24894 10962 24922 10963
rect 24946 10989 24974 10990
rect 24946 10963 24972 10989
rect 24972 10963 24974 10989
rect 24946 10962 24974 10963
rect 24998 10989 25026 10990
rect 24998 10963 25008 10989
rect 25008 10963 25026 10989
rect 24998 10962 25026 10963
rect 24374 10878 24402 10906
rect 24766 10878 24794 10906
rect 24374 9254 24402 9282
rect 25942 11774 25970 11802
rect 25382 10345 25410 10346
rect 25382 10319 25383 10345
rect 25383 10319 25409 10345
rect 25409 10319 25410 10345
rect 25382 10318 25410 10319
rect 25942 10318 25970 10346
rect 24582 10205 24610 10206
rect 24582 10179 24600 10205
rect 24600 10179 24610 10205
rect 24582 10178 24610 10179
rect 24634 10205 24662 10206
rect 24634 10179 24636 10205
rect 24636 10179 24662 10205
rect 24634 10178 24662 10179
rect 24686 10205 24714 10206
rect 24738 10205 24766 10206
rect 24686 10179 24698 10205
rect 24698 10179 24714 10205
rect 24738 10179 24760 10205
rect 24760 10179 24766 10205
rect 24686 10178 24714 10179
rect 24738 10178 24766 10179
rect 24790 10178 24818 10206
rect 24842 10205 24870 10206
rect 24894 10205 24922 10206
rect 24842 10179 24848 10205
rect 24848 10179 24870 10205
rect 24894 10179 24910 10205
rect 24910 10179 24922 10205
rect 24842 10178 24870 10179
rect 24894 10178 24922 10179
rect 24946 10205 24974 10206
rect 24946 10179 24972 10205
rect 24972 10179 24974 10205
rect 24946 10178 24974 10179
rect 24998 10205 25026 10206
rect 24998 10179 25008 10205
rect 25008 10179 25026 10205
rect 24998 10178 25026 10179
rect 25942 10094 25970 10122
rect 24654 9617 24682 9618
rect 24654 9591 24655 9617
rect 24655 9591 24681 9617
rect 24681 9591 24682 9617
rect 24654 9590 24682 9591
rect 24878 9617 24906 9618
rect 24878 9591 24879 9617
rect 24879 9591 24905 9617
rect 24905 9591 24906 9617
rect 24878 9590 24906 9591
rect 24582 9421 24610 9422
rect 24582 9395 24600 9421
rect 24600 9395 24610 9421
rect 24582 9394 24610 9395
rect 24634 9421 24662 9422
rect 24634 9395 24636 9421
rect 24636 9395 24662 9421
rect 24634 9394 24662 9395
rect 24686 9421 24714 9422
rect 24738 9421 24766 9422
rect 24686 9395 24698 9421
rect 24698 9395 24714 9421
rect 24738 9395 24760 9421
rect 24760 9395 24766 9421
rect 24686 9394 24714 9395
rect 24738 9394 24766 9395
rect 24790 9394 24818 9422
rect 24842 9421 24870 9422
rect 24894 9421 24922 9422
rect 24842 9395 24848 9421
rect 24848 9395 24870 9421
rect 24894 9395 24910 9421
rect 24910 9395 24922 9421
rect 24842 9394 24870 9395
rect 24894 9394 24922 9395
rect 24946 9421 24974 9422
rect 24946 9395 24972 9421
rect 24972 9395 24974 9421
rect 24946 9394 24974 9395
rect 24998 9421 25026 9422
rect 24998 9395 25008 9421
rect 25008 9395 25026 9421
rect 24998 9394 25026 9395
rect 24486 9198 24514 9226
rect 24766 9254 24794 9282
rect 25102 9198 25130 9226
rect 25158 9590 25186 9618
rect 24582 8637 24610 8638
rect 24582 8611 24600 8637
rect 24600 8611 24610 8637
rect 24582 8610 24610 8611
rect 24634 8637 24662 8638
rect 24634 8611 24636 8637
rect 24636 8611 24662 8637
rect 24634 8610 24662 8611
rect 24686 8637 24714 8638
rect 24738 8637 24766 8638
rect 24686 8611 24698 8637
rect 24698 8611 24714 8637
rect 24738 8611 24760 8637
rect 24760 8611 24766 8637
rect 24686 8610 24714 8611
rect 24738 8610 24766 8611
rect 24790 8610 24818 8638
rect 24842 8637 24870 8638
rect 24894 8637 24922 8638
rect 24842 8611 24848 8637
rect 24848 8611 24870 8637
rect 24894 8611 24910 8637
rect 24910 8611 24922 8637
rect 24842 8610 24870 8611
rect 24894 8610 24922 8611
rect 24946 8637 24974 8638
rect 24946 8611 24972 8637
rect 24972 8611 24974 8637
rect 24946 8610 24974 8611
rect 24998 8637 25026 8638
rect 24998 8611 25008 8637
rect 25008 8611 25026 8637
rect 24998 8610 25026 8611
rect 24878 8414 24906 8442
rect 24582 7853 24610 7854
rect 24582 7827 24600 7853
rect 24600 7827 24610 7853
rect 24582 7826 24610 7827
rect 24634 7853 24662 7854
rect 24634 7827 24636 7853
rect 24636 7827 24662 7853
rect 24634 7826 24662 7827
rect 24686 7853 24714 7854
rect 24738 7853 24766 7854
rect 24686 7827 24698 7853
rect 24698 7827 24714 7853
rect 24738 7827 24760 7853
rect 24760 7827 24766 7853
rect 24686 7826 24714 7827
rect 24738 7826 24766 7827
rect 24790 7826 24818 7854
rect 24842 7853 24870 7854
rect 24894 7853 24922 7854
rect 24842 7827 24848 7853
rect 24848 7827 24870 7853
rect 24894 7827 24910 7853
rect 24910 7827 24922 7853
rect 24842 7826 24870 7827
rect 24894 7826 24922 7827
rect 24946 7853 24974 7854
rect 24946 7827 24972 7853
rect 24972 7827 24974 7853
rect 24946 7826 24974 7827
rect 24998 7853 25026 7854
rect 24998 7827 25008 7853
rect 25008 7827 25026 7853
rect 24998 7826 25026 7827
rect 25438 9086 25466 9114
rect 26502 13145 26530 13146
rect 26502 13119 26503 13145
rect 26503 13119 26529 13145
rect 26529 13119 26530 13145
rect 26502 13118 26530 13119
rect 27082 12949 27110 12950
rect 27082 12923 27100 12949
rect 27100 12923 27110 12949
rect 27082 12922 27110 12923
rect 27134 12949 27162 12950
rect 27134 12923 27136 12949
rect 27136 12923 27162 12949
rect 27134 12922 27162 12923
rect 27186 12949 27214 12950
rect 27238 12949 27266 12950
rect 27186 12923 27198 12949
rect 27198 12923 27214 12949
rect 27238 12923 27260 12949
rect 27260 12923 27266 12949
rect 27186 12922 27214 12923
rect 27238 12922 27266 12923
rect 27290 12922 27318 12950
rect 27342 12949 27370 12950
rect 27394 12949 27422 12950
rect 27342 12923 27348 12949
rect 27348 12923 27370 12949
rect 27394 12923 27410 12949
rect 27410 12923 27422 12949
rect 27342 12922 27370 12923
rect 27394 12922 27422 12923
rect 27446 12949 27474 12950
rect 27446 12923 27472 12949
rect 27472 12923 27474 12949
rect 27446 12922 27474 12923
rect 27498 12949 27526 12950
rect 27498 12923 27508 12949
rect 27508 12923 27526 12949
rect 27498 12922 27526 12923
rect 26894 12361 26922 12362
rect 26894 12335 26895 12361
rect 26895 12335 26921 12361
rect 26921 12335 26922 12361
rect 26894 12334 26922 12335
rect 27174 12334 27202 12362
rect 27082 12165 27110 12166
rect 27082 12139 27100 12165
rect 27100 12139 27110 12165
rect 27082 12138 27110 12139
rect 27134 12165 27162 12166
rect 27134 12139 27136 12165
rect 27136 12139 27162 12165
rect 27134 12138 27162 12139
rect 27186 12165 27214 12166
rect 27238 12165 27266 12166
rect 27186 12139 27198 12165
rect 27198 12139 27214 12165
rect 27238 12139 27260 12165
rect 27260 12139 27266 12165
rect 27186 12138 27214 12139
rect 27238 12138 27266 12139
rect 27290 12138 27318 12166
rect 27342 12165 27370 12166
rect 27394 12165 27422 12166
rect 27342 12139 27348 12165
rect 27348 12139 27370 12165
rect 27394 12139 27410 12165
rect 27410 12139 27422 12165
rect 27342 12138 27370 12139
rect 27394 12138 27422 12139
rect 27446 12165 27474 12166
rect 27446 12139 27472 12165
rect 27472 12139 27474 12165
rect 27446 12138 27474 12139
rect 27498 12165 27526 12166
rect 27498 12139 27508 12165
rect 27508 12139 27526 12165
rect 27498 12138 27526 12139
rect 27006 11969 27034 11970
rect 27006 11943 27007 11969
rect 27007 11943 27033 11969
rect 27033 11943 27034 11969
rect 27006 11942 27034 11943
rect 29582 18045 29610 18046
rect 29582 18019 29600 18045
rect 29600 18019 29610 18045
rect 29582 18018 29610 18019
rect 29634 18045 29662 18046
rect 29634 18019 29636 18045
rect 29636 18019 29662 18045
rect 29634 18018 29662 18019
rect 29686 18045 29714 18046
rect 29738 18045 29766 18046
rect 29686 18019 29698 18045
rect 29698 18019 29714 18045
rect 29738 18019 29760 18045
rect 29760 18019 29766 18045
rect 29686 18018 29714 18019
rect 29738 18018 29766 18019
rect 29790 18018 29818 18046
rect 29842 18045 29870 18046
rect 29894 18045 29922 18046
rect 29842 18019 29848 18045
rect 29848 18019 29870 18045
rect 29894 18019 29910 18045
rect 29910 18019 29922 18045
rect 29842 18018 29870 18019
rect 29894 18018 29922 18019
rect 29946 18045 29974 18046
rect 29946 18019 29972 18045
rect 29972 18019 29974 18045
rect 29946 18018 29974 18019
rect 29998 18045 30026 18046
rect 29998 18019 30008 18045
rect 30008 18019 30026 18045
rect 29998 18018 30026 18019
rect 29582 17261 29610 17262
rect 29582 17235 29600 17261
rect 29600 17235 29610 17261
rect 29582 17234 29610 17235
rect 29634 17261 29662 17262
rect 29634 17235 29636 17261
rect 29636 17235 29662 17261
rect 29634 17234 29662 17235
rect 29686 17261 29714 17262
rect 29738 17261 29766 17262
rect 29686 17235 29698 17261
rect 29698 17235 29714 17261
rect 29738 17235 29760 17261
rect 29760 17235 29766 17261
rect 29686 17234 29714 17235
rect 29738 17234 29766 17235
rect 29790 17234 29818 17262
rect 29842 17261 29870 17262
rect 29894 17261 29922 17262
rect 29842 17235 29848 17261
rect 29848 17235 29870 17261
rect 29894 17235 29910 17261
rect 29910 17235 29922 17261
rect 29842 17234 29870 17235
rect 29894 17234 29922 17235
rect 29946 17261 29974 17262
rect 29946 17235 29972 17261
rect 29972 17235 29974 17261
rect 29946 17234 29974 17235
rect 29998 17261 30026 17262
rect 29998 17235 30008 17261
rect 30008 17235 30026 17261
rect 29998 17234 30026 17235
rect 29582 16477 29610 16478
rect 29582 16451 29600 16477
rect 29600 16451 29610 16477
rect 29582 16450 29610 16451
rect 29634 16477 29662 16478
rect 29634 16451 29636 16477
rect 29636 16451 29662 16477
rect 29634 16450 29662 16451
rect 29686 16477 29714 16478
rect 29738 16477 29766 16478
rect 29686 16451 29698 16477
rect 29698 16451 29714 16477
rect 29738 16451 29760 16477
rect 29760 16451 29766 16477
rect 29686 16450 29714 16451
rect 29738 16450 29766 16451
rect 29790 16450 29818 16478
rect 29842 16477 29870 16478
rect 29894 16477 29922 16478
rect 29842 16451 29848 16477
rect 29848 16451 29870 16477
rect 29894 16451 29910 16477
rect 29910 16451 29922 16477
rect 29842 16450 29870 16451
rect 29894 16450 29922 16451
rect 29946 16477 29974 16478
rect 29946 16451 29972 16477
rect 29972 16451 29974 16477
rect 29946 16450 29974 16451
rect 29998 16477 30026 16478
rect 29998 16451 30008 16477
rect 30008 16451 30026 16477
rect 29998 16450 30026 16451
rect 29582 15693 29610 15694
rect 29582 15667 29600 15693
rect 29600 15667 29610 15693
rect 29582 15666 29610 15667
rect 29634 15693 29662 15694
rect 29634 15667 29636 15693
rect 29636 15667 29662 15693
rect 29634 15666 29662 15667
rect 29686 15693 29714 15694
rect 29738 15693 29766 15694
rect 29686 15667 29698 15693
rect 29698 15667 29714 15693
rect 29738 15667 29760 15693
rect 29760 15667 29766 15693
rect 29686 15666 29714 15667
rect 29738 15666 29766 15667
rect 29790 15666 29818 15694
rect 29842 15693 29870 15694
rect 29894 15693 29922 15694
rect 29842 15667 29848 15693
rect 29848 15667 29870 15693
rect 29894 15667 29910 15693
rect 29910 15667 29922 15693
rect 29842 15666 29870 15667
rect 29894 15666 29922 15667
rect 29946 15693 29974 15694
rect 29946 15667 29972 15693
rect 29972 15667 29974 15693
rect 29946 15666 29974 15667
rect 29998 15693 30026 15694
rect 29998 15667 30008 15693
rect 30008 15667 30026 15693
rect 29998 15666 30026 15667
rect 29582 14909 29610 14910
rect 29582 14883 29600 14909
rect 29600 14883 29610 14909
rect 29582 14882 29610 14883
rect 29634 14909 29662 14910
rect 29634 14883 29636 14909
rect 29636 14883 29662 14909
rect 29634 14882 29662 14883
rect 29686 14909 29714 14910
rect 29738 14909 29766 14910
rect 29686 14883 29698 14909
rect 29698 14883 29714 14909
rect 29738 14883 29760 14909
rect 29760 14883 29766 14909
rect 29686 14882 29714 14883
rect 29738 14882 29766 14883
rect 29790 14882 29818 14910
rect 29842 14909 29870 14910
rect 29894 14909 29922 14910
rect 29842 14883 29848 14909
rect 29848 14883 29870 14909
rect 29894 14883 29910 14909
rect 29910 14883 29922 14909
rect 29842 14882 29870 14883
rect 29894 14882 29922 14883
rect 29946 14909 29974 14910
rect 29946 14883 29972 14909
rect 29972 14883 29974 14909
rect 29946 14882 29974 14883
rect 29998 14909 30026 14910
rect 29998 14883 30008 14909
rect 30008 14883 30026 14909
rect 29998 14882 30026 14883
rect 27678 13958 27706 13986
rect 27678 13481 27706 13482
rect 27678 13455 27679 13481
rect 27679 13455 27705 13481
rect 27705 13455 27706 13481
rect 27678 13454 27706 13455
rect 28462 13537 28490 13538
rect 28462 13511 28463 13537
rect 28463 13511 28489 13537
rect 28489 13511 28490 13537
rect 28462 13510 28490 13511
rect 28462 12614 28490 12642
rect 29022 12614 29050 12642
rect 27622 12334 27650 12362
rect 29582 14125 29610 14126
rect 29582 14099 29600 14125
rect 29600 14099 29610 14125
rect 29582 14098 29610 14099
rect 29634 14125 29662 14126
rect 29634 14099 29636 14125
rect 29636 14099 29662 14125
rect 29634 14098 29662 14099
rect 29686 14125 29714 14126
rect 29738 14125 29766 14126
rect 29686 14099 29698 14125
rect 29698 14099 29714 14125
rect 29738 14099 29760 14125
rect 29760 14099 29766 14125
rect 29686 14098 29714 14099
rect 29738 14098 29766 14099
rect 29790 14098 29818 14126
rect 29842 14125 29870 14126
rect 29894 14125 29922 14126
rect 29842 14099 29848 14125
rect 29848 14099 29870 14125
rect 29894 14099 29910 14125
rect 29910 14099 29922 14125
rect 29842 14098 29870 14099
rect 29894 14098 29922 14099
rect 29946 14125 29974 14126
rect 29946 14099 29972 14125
rect 29972 14099 29974 14125
rect 29946 14098 29974 14099
rect 29998 14125 30026 14126
rect 29998 14099 30008 14125
rect 30008 14099 30026 14125
rect 29998 14098 30026 14099
rect 29358 13481 29386 13482
rect 29358 13455 29359 13481
rect 29359 13455 29385 13481
rect 29385 13455 29386 13481
rect 29358 13454 29386 13455
rect 29582 13341 29610 13342
rect 29582 13315 29600 13341
rect 29600 13315 29610 13341
rect 29582 13314 29610 13315
rect 29634 13341 29662 13342
rect 29634 13315 29636 13341
rect 29636 13315 29662 13341
rect 29634 13314 29662 13315
rect 29686 13341 29714 13342
rect 29738 13341 29766 13342
rect 29686 13315 29698 13341
rect 29698 13315 29714 13341
rect 29738 13315 29760 13341
rect 29760 13315 29766 13341
rect 29686 13314 29714 13315
rect 29738 13314 29766 13315
rect 29790 13314 29818 13342
rect 29842 13341 29870 13342
rect 29894 13341 29922 13342
rect 29842 13315 29848 13341
rect 29848 13315 29870 13341
rect 29894 13315 29910 13341
rect 29910 13315 29922 13341
rect 29842 13314 29870 13315
rect 29894 13314 29922 13315
rect 29946 13341 29974 13342
rect 29946 13315 29972 13341
rect 29972 13315 29974 13341
rect 29946 13314 29974 13315
rect 29998 13341 30026 13342
rect 29998 13315 30008 13341
rect 30008 13315 30026 13341
rect 29998 13314 30026 13315
rect 29246 12334 29274 12362
rect 30478 12614 30506 12642
rect 29582 12557 29610 12558
rect 29582 12531 29600 12557
rect 29600 12531 29610 12557
rect 29582 12530 29610 12531
rect 29634 12557 29662 12558
rect 29634 12531 29636 12557
rect 29636 12531 29662 12557
rect 29634 12530 29662 12531
rect 29686 12557 29714 12558
rect 29738 12557 29766 12558
rect 29686 12531 29698 12557
rect 29698 12531 29714 12557
rect 29738 12531 29760 12557
rect 29760 12531 29766 12557
rect 29686 12530 29714 12531
rect 29738 12530 29766 12531
rect 29790 12530 29818 12558
rect 29842 12557 29870 12558
rect 29894 12557 29922 12558
rect 29842 12531 29848 12557
rect 29848 12531 29870 12557
rect 29894 12531 29910 12557
rect 29910 12531 29922 12557
rect 29842 12530 29870 12531
rect 29894 12530 29922 12531
rect 29946 12557 29974 12558
rect 29946 12531 29972 12557
rect 29972 12531 29974 12557
rect 29946 12530 29974 12531
rect 29998 12557 30026 12558
rect 29998 12531 30008 12557
rect 30008 12531 30026 12557
rect 29998 12530 30026 12531
rect 27622 12054 27650 12082
rect 29246 12054 29274 12082
rect 27678 11774 27706 11802
rect 27398 11577 27426 11578
rect 27398 11551 27399 11577
rect 27399 11551 27425 11577
rect 27425 11551 27426 11577
rect 27398 11550 27426 11551
rect 27082 11381 27110 11382
rect 27082 11355 27100 11381
rect 27100 11355 27110 11381
rect 27082 11354 27110 11355
rect 27134 11381 27162 11382
rect 27134 11355 27136 11381
rect 27136 11355 27162 11381
rect 27134 11354 27162 11355
rect 27186 11381 27214 11382
rect 27238 11381 27266 11382
rect 27186 11355 27198 11381
rect 27198 11355 27214 11381
rect 27238 11355 27260 11381
rect 27260 11355 27266 11381
rect 27186 11354 27214 11355
rect 27238 11354 27266 11355
rect 27290 11354 27318 11382
rect 27342 11381 27370 11382
rect 27394 11381 27422 11382
rect 27342 11355 27348 11381
rect 27348 11355 27370 11381
rect 27394 11355 27410 11381
rect 27410 11355 27422 11381
rect 27342 11354 27370 11355
rect 27394 11354 27422 11355
rect 27446 11381 27474 11382
rect 27446 11355 27472 11381
rect 27472 11355 27474 11381
rect 27446 11354 27474 11355
rect 27498 11381 27526 11382
rect 27498 11355 27508 11381
rect 27508 11355 27526 11381
rect 27498 11354 27526 11355
rect 26950 11046 26978 11074
rect 27230 11046 27258 11074
rect 28462 11969 28490 11970
rect 28462 11943 28463 11969
rect 28463 11943 28489 11969
rect 28489 11943 28490 11969
rect 28462 11942 28490 11943
rect 27678 11102 27706 11130
rect 27846 11550 27874 11578
rect 27454 11046 27482 11074
rect 26222 10878 26250 10906
rect 26726 10878 26754 10906
rect 27286 10793 27314 10794
rect 27286 10767 27287 10793
rect 27287 10767 27313 10793
rect 27313 10767 27314 10793
rect 27286 10766 27314 10767
rect 27566 10766 27594 10794
rect 27082 10597 27110 10598
rect 27082 10571 27100 10597
rect 27100 10571 27110 10597
rect 27082 10570 27110 10571
rect 27134 10597 27162 10598
rect 27134 10571 27136 10597
rect 27136 10571 27162 10597
rect 27134 10570 27162 10571
rect 27186 10597 27214 10598
rect 27238 10597 27266 10598
rect 27186 10571 27198 10597
rect 27198 10571 27214 10597
rect 27238 10571 27260 10597
rect 27260 10571 27266 10597
rect 27186 10570 27214 10571
rect 27238 10570 27266 10571
rect 27290 10570 27318 10598
rect 27342 10597 27370 10598
rect 27394 10597 27422 10598
rect 27342 10571 27348 10597
rect 27348 10571 27370 10597
rect 27394 10571 27410 10597
rect 27410 10571 27422 10597
rect 27342 10570 27370 10571
rect 27394 10570 27422 10571
rect 27446 10597 27474 10598
rect 27446 10571 27472 10597
rect 27472 10571 27474 10597
rect 27446 10570 27474 10571
rect 27498 10597 27526 10598
rect 27498 10571 27508 10597
rect 27508 10571 27526 10597
rect 27498 10570 27526 10571
rect 26726 10401 26754 10402
rect 26726 10375 26727 10401
rect 26727 10375 26753 10401
rect 26753 10375 26754 10401
rect 26726 10374 26754 10375
rect 28462 11185 28490 11186
rect 28462 11159 28463 11185
rect 28463 11159 28489 11185
rect 28489 11159 28490 11185
rect 28462 11158 28490 11159
rect 28630 11102 28658 11130
rect 28854 11102 28882 11130
rect 28406 10374 28434 10402
rect 28630 10318 28658 10346
rect 27566 10038 27594 10066
rect 27398 10009 27426 10010
rect 27398 9983 27399 10009
rect 27399 9983 27425 10009
rect 27425 9983 27426 10009
rect 27398 9982 27426 9983
rect 27082 9813 27110 9814
rect 27082 9787 27100 9813
rect 27100 9787 27110 9813
rect 27082 9786 27110 9787
rect 27134 9813 27162 9814
rect 27134 9787 27136 9813
rect 27136 9787 27162 9813
rect 27134 9786 27162 9787
rect 27186 9813 27214 9814
rect 27238 9813 27266 9814
rect 27186 9787 27198 9813
rect 27198 9787 27214 9813
rect 27238 9787 27260 9813
rect 27260 9787 27266 9813
rect 27186 9786 27214 9787
rect 27238 9786 27266 9787
rect 27290 9786 27318 9814
rect 27342 9813 27370 9814
rect 27394 9813 27422 9814
rect 27342 9787 27348 9813
rect 27348 9787 27370 9813
rect 27394 9787 27410 9813
rect 27410 9787 27422 9813
rect 27342 9786 27370 9787
rect 27394 9786 27422 9787
rect 27446 9813 27474 9814
rect 27446 9787 27472 9813
rect 27472 9787 27474 9813
rect 27446 9786 27474 9787
rect 27498 9813 27526 9814
rect 27498 9787 27508 9813
rect 27508 9787 27526 9813
rect 27498 9786 27526 9787
rect 26950 9590 26978 9618
rect 27230 9617 27258 9618
rect 27230 9591 27231 9617
rect 27231 9591 27257 9617
rect 27257 9591 27258 9617
rect 27230 9590 27258 9591
rect 27454 9617 27482 9618
rect 27454 9591 27455 9617
rect 27455 9591 27481 9617
rect 27481 9591 27482 9617
rect 27454 9590 27482 9591
rect 26502 9225 26530 9226
rect 26502 9199 26503 9225
rect 26503 9199 26529 9225
rect 26529 9199 26530 9225
rect 26502 9198 26530 9199
rect 25998 9086 26026 9114
rect 27082 9029 27110 9030
rect 27082 9003 27100 9029
rect 27100 9003 27110 9029
rect 27082 9002 27110 9003
rect 27134 9029 27162 9030
rect 27134 9003 27136 9029
rect 27136 9003 27162 9029
rect 27134 9002 27162 9003
rect 27186 9029 27214 9030
rect 27238 9029 27266 9030
rect 27186 9003 27198 9029
rect 27198 9003 27214 9029
rect 27238 9003 27260 9029
rect 27260 9003 27266 9029
rect 27186 9002 27214 9003
rect 27238 9002 27266 9003
rect 27290 9002 27318 9030
rect 27342 9029 27370 9030
rect 27394 9029 27422 9030
rect 27342 9003 27348 9029
rect 27348 9003 27370 9029
rect 27394 9003 27410 9029
rect 27410 9003 27422 9029
rect 27342 9002 27370 9003
rect 27394 9002 27422 9003
rect 27446 9029 27474 9030
rect 27446 9003 27472 9029
rect 27472 9003 27474 9029
rect 27446 9002 27474 9003
rect 27498 9029 27526 9030
rect 27498 9003 27508 9029
rect 27508 9003 27526 9029
rect 27498 9002 27526 9003
rect 25158 8414 25186 8442
rect 25438 8441 25466 8442
rect 25438 8415 25439 8441
rect 25439 8415 25465 8441
rect 25465 8415 25466 8441
rect 25438 8414 25466 8415
rect 25158 7238 25186 7266
rect 24582 7069 24610 7070
rect 24582 7043 24600 7069
rect 24600 7043 24610 7069
rect 24582 7042 24610 7043
rect 24634 7069 24662 7070
rect 24634 7043 24636 7069
rect 24636 7043 24662 7069
rect 24634 7042 24662 7043
rect 24686 7069 24714 7070
rect 24738 7069 24766 7070
rect 24686 7043 24698 7069
rect 24698 7043 24714 7069
rect 24738 7043 24760 7069
rect 24760 7043 24766 7069
rect 24686 7042 24714 7043
rect 24738 7042 24766 7043
rect 24790 7042 24818 7070
rect 24842 7069 24870 7070
rect 24894 7069 24922 7070
rect 24842 7043 24848 7069
rect 24848 7043 24870 7069
rect 24894 7043 24910 7069
rect 24910 7043 24922 7069
rect 24842 7042 24870 7043
rect 24894 7042 24922 7043
rect 24946 7069 24974 7070
rect 24946 7043 24972 7069
rect 24972 7043 24974 7069
rect 24946 7042 24974 7043
rect 24998 7069 25026 7070
rect 24998 7043 25008 7069
rect 25008 7043 25026 7069
rect 24998 7042 25026 7043
rect 24374 6481 24402 6482
rect 24374 6455 24375 6481
rect 24375 6455 24401 6481
rect 24401 6455 24402 6481
rect 24374 6454 24402 6455
rect 24766 6454 24794 6482
rect 25214 6873 25242 6874
rect 25214 6847 25215 6873
rect 25215 6847 25241 6873
rect 25241 6847 25242 6873
rect 25214 6846 25242 6847
rect 24582 6285 24610 6286
rect 24582 6259 24600 6285
rect 24600 6259 24610 6285
rect 24582 6258 24610 6259
rect 24634 6285 24662 6286
rect 24634 6259 24636 6285
rect 24636 6259 24662 6285
rect 24634 6258 24662 6259
rect 24686 6285 24714 6286
rect 24738 6285 24766 6286
rect 24686 6259 24698 6285
rect 24698 6259 24714 6285
rect 24738 6259 24760 6285
rect 24760 6259 24766 6285
rect 24686 6258 24714 6259
rect 24738 6258 24766 6259
rect 24790 6258 24818 6286
rect 24842 6285 24870 6286
rect 24894 6285 24922 6286
rect 24842 6259 24848 6285
rect 24848 6259 24870 6285
rect 24894 6259 24910 6285
rect 24910 6259 24922 6285
rect 24842 6258 24870 6259
rect 24894 6258 24922 6259
rect 24946 6285 24974 6286
rect 24946 6259 24972 6285
rect 24972 6259 24974 6285
rect 24946 6258 24974 6259
rect 24998 6285 25026 6286
rect 24998 6259 25008 6285
rect 25008 6259 25026 6285
rect 24998 6258 25026 6259
rect 24374 6062 24402 6090
rect 24766 6089 24794 6090
rect 24766 6063 24767 6089
rect 24767 6063 24793 6089
rect 24793 6063 24794 6089
rect 24766 6062 24794 6063
rect 25382 7126 25410 7154
rect 24582 5501 24610 5502
rect 24582 5475 24600 5501
rect 24600 5475 24610 5501
rect 24582 5474 24610 5475
rect 24634 5501 24662 5502
rect 24634 5475 24636 5501
rect 24636 5475 24662 5501
rect 24634 5474 24662 5475
rect 24686 5501 24714 5502
rect 24738 5501 24766 5502
rect 24686 5475 24698 5501
rect 24698 5475 24714 5501
rect 24738 5475 24760 5501
rect 24760 5475 24766 5501
rect 24686 5474 24714 5475
rect 24738 5474 24766 5475
rect 24790 5474 24818 5502
rect 24842 5501 24870 5502
rect 24894 5501 24922 5502
rect 24842 5475 24848 5501
rect 24848 5475 24870 5501
rect 24894 5475 24910 5501
rect 24910 5475 24922 5501
rect 24842 5474 24870 5475
rect 24894 5474 24922 5475
rect 24946 5501 24974 5502
rect 24946 5475 24972 5501
rect 24972 5475 24974 5501
rect 24946 5474 24974 5475
rect 24998 5501 25026 5502
rect 24998 5475 25008 5501
rect 25008 5475 25026 5501
rect 24998 5474 25026 5475
rect 24374 4129 24402 4130
rect 24374 4103 24375 4129
rect 24375 4103 24401 4129
rect 24401 4103 24402 4129
rect 24374 4102 24402 4103
rect 24430 5334 24458 5362
rect 24094 2478 24122 2506
rect 24374 3710 24402 3738
rect 24374 2422 24402 2450
rect 24582 4717 24610 4718
rect 24582 4691 24600 4717
rect 24600 4691 24610 4717
rect 24582 4690 24610 4691
rect 24634 4717 24662 4718
rect 24634 4691 24636 4717
rect 24636 4691 24662 4717
rect 24634 4690 24662 4691
rect 24686 4717 24714 4718
rect 24738 4717 24766 4718
rect 24686 4691 24698 4717
rect 24698 4691 24714 4717
rect 24738 4691 24760 4717
rect 24760 4691 24766 4717
rect 24686 4690 24714 4691
rect 24738 4690 24766 4691
rect 24790 4690 24818 4718
rect 24842 4717 24870 4718
rect 24894 4717 24922 4718
rect 24842 4691 24848 4717
rect 24848 4691 24870 4717
rect 24894 4691 24910 4717
rect 24910 4691 24922 4717
rect 24842 4690 24870 4691
rect 24894 4690 24922 4691
rect 24946 4717 24974 4718
rect 24946 4691 24972 4717
rect 24972 4691 24974 4717
rect 24946 4690 24974 4691
rect 24998 4717 25026 4718
rect 24998 4691 25008 4717
rect 25008 4691 25026 4717
rect 24998 4690 25026 4691
rect 24766 4102 24794 4130
rect 24654 4046 24682 4074
rect 24878 4046 24906 4074
rect 25438 6873 25466 6874
rect 25438 6847 25439 6873
rect 25439 6847 25465 6873
rect 25465 6847 25466 6873
rect 25438 6846 25466 6847
rect 26222 6089 26250 6090
rect 26222 6063 26223 6089
rect 26223 6063 26249 6089
rect 26249 6063 26250 6089
rect 26222 6062 26250 6063
rect 25942 5222 25970 5250
rect 26054 5278 26082 5306
rect 26894 8441 26922 8442
rect 26894 8415 26895 8441
rect 26895 8415 26921 8441
rect 26921 8415 26922 8441
rect 26894 8414 26922 8415
rect 26670 5950 26698 5978
rect 27174 8414 27202 8442
rect 27082 8245 27110 8246
rect 27082 8219 27100 8245
rect 27100 8219 27110 8245
rect 27082 8218 27110 8219
rect 27134 8245 27162 8246
rect 27134 8219 27136 8245
rect 27136 8219 27162 8245
rect 27134 8218 27162 8219
rect 27186 8245 27214 8246
rect 27238 8245 27266 8246
rect 27186 8219 27198 8245
rect 27198 8219 27214 8245
rect 27238 8219 27260 8245
rect 27260 8219 27266 8245
rect 27186 8218 27214 8219
rect 27238 8218 27266 8219
rect 27290 8218 27318 8246
rect 27342 8245 27370 8246
rect 27394 8245 27422 8246
rect 27342 8219 27348 8245
rect 27348 8219 27370 8245
rect 27394 8219 27410 8245
rect 27410 8219 27422 8245
rect 27342 8218 27370 8219
rect 27394 8218 27422 8219
rect 27446 8245 27474 8246
rect 27446 8219 27472 8245
rect 27472 8219 27474 8245
rect 27446 8218 27474 8219
rect 27498 8245 27526 8246
rect 27498 8219 27508 8245
rect 27508 8219 27526 8245
rect 27498 8218 27526 8219
rect 26726 6846 26754 6874
rect 27082 7461 27110 7462
rect 27082 7435 27100 7461
rect 27100 7435 27110 7461
rect 27082 7434 27110 7435
rect 27134 7461 27162 7462
rect 27134 7435 27136 7461
rect 27136 7435 27162 7461
rect 27134 7434 27162 7435
rect 27186 7461 27214 7462
rect 27238 7461 27266 7462
rect 27186 7435 27198 7461
rect 27198 7435 27214 7461
rect 27238 7435 27260 7461
rect 27260 7435 27266 7461
rect 27186 7434 27214 7435
rect 27238 7434 27266 7435
rect 27290 7434 27318 7462
rect 27342 7461 27370 7462
rect 27394 7461 27422 7462
rect 27342 7435 27348 7461
rect 27348 7435 27370 7461
rect 27394 7435 27410 7461
rect 27410 7435 27422 7461
rect 27342 7434 27370 7435
rect 27394 7434 27422 7435
rect 27446 7461 27474 7462
rect 27446 7435 27472 7461
rect 27472 7435 27474 7461
rect 27446 7434 27474 7435
rect 27498 7461 27526 7462
rect 27498 7435 27508 7461
rect 27508 7435 27526 7461
rect 27498 7434 27526 7435
rect 27174 7265 27202 7266
rect 27174 7239 27175 7265
rect 27175 7239 27201 7265
rect 27201 7239 27202 7265
rect 27174 7238 27202 7239
rect 27398 7265 27426 7266
rect 27398 7239 27399 7265
rect 27399 7239 27425 7265
rect 27425 7239 27426 7265
rect 27398 7238 27426 7239
rect 26726 6062 26754 6090
rect 26894 6734 26922 6762
rect 27006 7182 27034 7210
rect 27902 9982 27930 10010
rect 27902 9534 27930 9562
rect 28406 9534 28434 9562
rect 29582 11773 29610 11774
rect 29582 11747 29600 11773
rect 29600 11747 29610 11773
rect 29582 11746 29610 11747
rect 29634 11773 29662 11774
rect 29634 11747 29636 11773
rect 29636 11747 29662 11773
rect 29634 11746 29662 11747
rect 29686 11773 29714 11774
rect 29738 11773 29766 11774
rect 29686 11747 29698 11773
rect 29698 11747 29714 11773
rect 29738 11747 29760 11773
rect 29760 11747 29766 11773
rect 29686 11746 29714 11747
rect 29738 11746 29766 11747
rect 29790 11746 29818 11774
rect 29842 11773 29870 11774
rect 29894 11773 29922 11774
rect 29842 11747 29848 11773
rect 29848 11747 29870 11773
rect 29894 11747 29910 11773
rect 29910 11747 29922 11773
rect 29842 11746 29870 11747
rect 29894 11746 29922 11747
rect 29946 11773 29974 11774
rect 29946 11747 29972 11773
rect 29972 11747 29974 11773
rect 29946 11746 29974 11747
rect 29998 11773 30026 11774
rect 29998 11747 30008 11773
rect 30008 11747 30026 11773
rect 29998 11746 30026 11747
rect 31094 12361 31122 12362
rect 31094 12335 31095 12361
rect 31095 12335 31121 12361
rect 31121 12335 31122 12361
rect 31094 12334 31122 12335
rect 29470 11494 29498 11522
rect 29022 11158 29050 11186
rect 29414 11382 29442 11410
rect 29414 11046 29442 11074
rect 28966 10038 28994 10066
rect 28574 9982 28602 10010
rect 28574 9590 28602 9618
rect 28462 9198 28490 9226
rect 28462 8049 28490 8050
rect 28462 8023 28463 8049
rect 28463 8023 28489 8049
rect 28489 8023 28490 8049
rect 28462 8022 28490 8023
rect 27678 7182 27706 7210
rect 28462 6846 28490 6874
rect 27082 6677 27110 6678
rect 27082 6651 27100 6677
rect 27100 6651 27110 6677
rect 27082 6650 27110 6651
rect 27134 6677 27162 6678
rect 27134 6651 27136 6677
rect 27136 6651 27162 6677
rect 27134 6650 27162 6651
rect 27186 6677 27214 6678
rect 27238 6677 27266 6678
rect 27186 6651 27198 6677
rect 27198 6651 27214 6677
rect 27238 6651 27260 6677
rect 27260 6651 27266 6677
rect 27186 6650 27214 6651
rect 27238 6650 27266 6651
rect 27290 6650 27318 6678
rect 27342 6677 27370 6678
rect 27394 6677 27422 6678
rect 27342 6651 27348 6677
rect 27348 6651 27370 6677
rect 27394 6651 27410 6677
rect 27410 6651 27422 6677
rect 27342 6650 27370 6651
rect 27394 6650 27422 6651
rect 27446 6677 27474 6678
rect 27446 6651 27472 6677
rect 27472 6651 27474 6677
rect 27446 6650 27474 6651
rect 27498 6677 27526 6678
rect 27498 6651 27508 6677
rect 27508 6651 27526 6677
rect 27498 6650 27526 6651
rect 26894 6118 26922 6146
rect 27174 6145 27202 6146
rect 27174 6119 27175 6145
rect 27175 6119 27201 6145
rect 27201 6119 27202 6145
rect 27174 6118 27202 6119
rect 26782 5222 26810 5250
rect 26054 5166 26082 5194
rect 25214 4046 25242 4074
rect 24582 3933 24610 3934
rect 24582 3907 24600 3933
rect 24600 3907 24610 3933
rect 24582 3906 24610 3907
rect 24634 3933 24662 3934
rect 24634 3907 24636 3933
rect 24636 3907 24662 3933
rect 24634 3906 24662 3907
rect 24686 3933 24714 3934
rect 24738 3933 24766 3934
rect 24686 3907 24698 3933
rect 24698 3907 24714 3933
rect 24738 3907 24760 3933
rect 24760 3907 24766 3933
rect 24686 3906 24714 3907
rect 24738 3906 24766 3907
rect 24790 3906 24818 3934
rect 24842 3933 24870 3934
rect 24894 3933 24922 3934
rect 24842 3907 24848 3933
rect 24848 3907 24870 3933
rect 24894 3907 24910 3933
rect 24910 3907 24922 3933
rect 24842 3906 24870 3907
rect 24894 3906 24922 3907
rect 24946 3933 24974 3934
rect 24946 3907 24972 3933
rect 24972 3907 24974 3933
rect 24946 3906 24974 3907
rect 24998 3933 25026 3934
rect 24998 3907 25008 3933
rect 25008 3907 25026 3933
rect 24998 3906 25026 3907
rect 24766 3737 24794 3738
rect 24766 3711 24767 3737
rect 24767 3711 24793 3737
rect 24793 3711 24794 3737
rect 24766 3710 24794 3711
rect 25214 3737 25242 3738
rect 25214 3711 25215 3737
rect 25215 3711 25241 3737
rect 25241 3711 25242 3737
rect 25214 3710 25242 3711
rect 24582 3149 24610 3150
rect 24582 3123 24600 3149
rect 24600 3123 24610 3149
rect 24582 3122 24610 3123
rect 24634 3149 24662 3150
rect 24634 3123 24636 3149
rect 24636 3123 24662 3149
rect 24634 3122 24662 3123
rect 24686 3149 24714 3150
rect 24738 3149 24766 3150
rect 24686 3123 24698 3149
rect 24698 3123 24714 3149
rect 24738 3123 24760 3149
rect 24760 3123 24766 3149
rect 24686 3122 24714 3123
rect 24738 3122 24766 3123
rect 24790 3122 24818 3150
rect 24842 3149 24870 3150
rect 24894 3149 24922 3150
rect 24842 3123 24848 3149
rect 24848 3123 24870 3149
rect 24894 3123 24910 3149
rect 24910 3123 24922 3149
rect 24842 3122 24870 3123
rect 24894 3122 24922 3123
rect 24946 3149 24974 3150
rect 24946 3123 24972 3149
rect 24972 3123 24974 3149
rect 24946 3122 24974 3123
rect 24998 3149 25026 3150
rect 24998 3123 25008 3149
rect 25008 3123 25026 3149
rect 24998 3122 25026 3123
rect 24654 2561 24682 2562
rect 24654 2535 24655 2561
rect 24655 2535 24681 2561
rect 24681 2535 24682 2561
rect 24654 2534 24682 2535
rect 24486 2422 24514 2450
rect 24878 2561 24906 2562
rect 24878 2535 24879 2561
rect 24879 2535 24905 2561
rect 24905 2535 24906 2561
rect 24878 2534 24906 2535
rect 25214 2534 25242 2562
rect 24766 2422 24794 2450
rect 24582 2365 24610 2366
rect 24582 2339 24600 2365
rect 24600 2339 24610 2365
rect 24582 2338 24610 2339
rect 24634 2365 24662 2366
rect 24634 2339 24636 2365
rect 24636 2339 24662 2365
rect 24634 2338 24662 2339
rect 24686 2365 24714 2366
rect 24738 2365 24766 2366
rect 24686 2339 24698 2365
rect 24698 2339 24714 2365
rect 24738 2339 24760 2365
rect 24760 2339 24766 2365
rect 24686 2338 24714 2339
rect 24738 2338 24766 2339
rect 24790 2338 24818 2366
rect 24842 2365 24870 2366
rect 24894 2365 24922 2366
rect 24842 2339 24848 2365
rect 24848 2339 24870 2365
rect 24894 2339 24910 2365
rect 24910 2339 24922 2365
rect 24842 2338 24870 2339
rect 24894 2338 24922 2339
rect 24946 2365 24974 2366
rect 24946 2339 24972 2365
rect 24972 2339 24974 2365
rect 24946 2338 24974 2339
rect 24998 2365 25026 2366
rect 24998 2339 25008 2365
rect 25008 2339 25026 2365
rect 24998 2338 25026 2339
rect 24486 2142 24514 2170
rect 24318 1862 24346 1890
rect 22918 1414 22946 1442
rect 24766 2169 24794 2170
rect 24766 2143 24767 2169
rect 24767 2143 24793 2169
rect 24793 2143 24794 2169
rect 24766 2142 24794 2143
rect 25438 3737 25466 3738
rect 25438 3711 25439 3737
rect 25439 3711 25465 3737
rect 25465 3711 25466 3737
rect 25438 3710 25466 3711
rect 25438 2534 25466 2562
rect 26334 4494 26362 4522
rect 26278 2534 26306 2562
rect 26054 2505 26082 2506
rect 26054 2479 26055 2505
rect 26055 2479 26081 2505
rect 26081 2479 26082 2505
rect 26054 2478 26082 2479
rect 26222 2505 26250 2506
rect 26222 2479 26223 2505
rect 26223 2479 26249 2505
rect 26249 2479 26250 2505
rect 26222 2478 26250 2479
rect 26894 3737 26922 3738
rect 26894 3711 26895 3737
rect 26895 3711 26921 3737
rect 26921 3711 26922 3737
rect 26894 3710 26922 3711
rect 26894 3374 26922 3402
rect 26726 2561 26754 2562
rect 26726 2535 26727 2561
rect 26727 2535 26753 2561
rect 26753 2535 26754 2561
rect 26726 2534 26754 2535
rect 26894 2646 26922 2674
rect 26334 2422 26362 2450
rect 26222 2169 26250 2170
rect 26222 2143 26223 2169
rect 26223 2143 26249 2169
rect 26249 2143 26250 2169
rect 26222 2142 26250 2143
rect 24582 1581 24610 1582
rect 24582 1555 24600 1581
rect 24600 1555 24610 1581
rect 24582 1554 24610 1555
rect 24634 1581 24662 1582
rect 24634 1555 24636 1581
rect 24636 1555 24662 1581
rect 24634 1554 24662 1555
rect 24686 1581 24714 1582
rect 24738 1581 24766 1582
rect 24686 1555 24698 1581
rect 24698 1555 24714 1581
rect 24738 1555 24760 1581
rect 24760 1555 24766 1581
rect 24686 1554 24714 1555
rect 24738 1554 24766 1555
rect 24790 1554 24818 1582
rect 24842 1581 24870 1582
rect 24894 1581 24922 1582
rect 24842 1555 24848 1581
rect 24848 1555 24870 1581
rect 24894 1555 24910 1581
rect 24910 1555 24922 1581
rect 24842 1554 24870 1555
rect 24894 1554 24922 1555
rect 24946 1581 24974 1582
rect 24946 1555 24972 1581
rect 24972 1555 24974 1581
rect 24946 1554 24974 1555
rect 24998 1581 25026 1582
rect 24998 1555 25008 1581
rect 25008 1555 25026 1581
rect 24998 1554 25026 1555
rect 27082 5893 27110 5894
rect 27082 5867 27100 5893
rect 27100 5867 27110 5893
rect 27082 5866 27110 5867
rect 27134 5893 27162 5894
rect 27134 5867 27136 5893
rect 27136 5867 27162 5893
rect 27134 5866 27162 5867
rect 27186 5893 27214 5894
rect 27238 5893 27266 5894
rect 27186 5867 27198 5893
rect 27198 5867 27214 5893
rect 27238 5867 27260 5893
rect 27260 5867 27266 5893
rect 27186 5866 27214 5867
rect 27238 5866 27266 5867
rect 27290 5866 27318 5894
rect 27342 5893 27370 5894
rect 27394 5893 27422 5894
rect 27342 5867 27348 5893
rect 27348 5867 27370 5893
rect 27394 5867 27410 5893
rect 27410 5867 27422 5893
rect 27342 5866 27370 5867
rect 27394 5866 27422 5867
rect 27446 5893 27474 5894
rect 27446 5867 27472 5893
rect 27472 5867 27474 5893
rect 27446 5866 27474 5867
rect 27498 5893 27526 5894
rect 27498 5867 27508 5893
rect 27508 5867 27526 5893
rect 27498 5866 27526 5867
rect 28070 5782 28098 5810
rect 28070 5361 28098 5362
rect 28070 5335 28071 5361
rect 28071 5335 28097 5361
rect 28097 5335 28098 5361
rect 28070 5334 28098 5335
rect 28014 5278 28042 5306
rect 28182 5305 28210 5306
rect 28182 5279 28183 5305
rect 28183 5279 28209 5305
rect 28209 5279 28210 5305
rect 28182 5278 28210 5279
rect 28014 5166 28042 5194
rect 27082 5109 27110 5110
rect 27082 5083 27100 5109
rect 27100 5083 27110 5109
rect 27082 5082 27110 5083
rect 27134 5109 27162 5110
rect 27134 5083 27136 5109
rect 27136 5083 27162 5109
rect 27134 5082 27162 5083
rect 27186 5109 27214 5110
rect 27238 5109 27266 5110
rect 27186 5083 27198 5109
rect 27198 5083 27214 5109
rect 27238 5083 27260 5109
rect 27260 5083 27266 5109
rect 27186 5082 27214 5083
rect 27238 5082 27266 5083
rect 27290 5082 27318 5110
rect 27342 5109 27370 5110
rect 27394 5109 27422 5110
rect 27342 5083 27348 5109
rect 27348 5083 27370 5109
rect 27394 5083 27410 5109
rect 27410 5083 27422 5109
rect 27342 5082 27370 5083
rect 27394 5082 27422 5083
rect 27446 5109 27474 5110
rect 27446 5083 27472 5109
rect 27472 5083 27474 5109
rect 27446 5082 27474 5083
rect 27498 5109 27526 5110
rect 27498 5083 27508 5109
rect 27508 5083 27526 5109
rect 27498 5082 27526 5083
rect 27082 4325 27110 4326
rect 27082 4299 27100 4325
rect 27100 4299 27110 4325
rect 27082 4298 27110 4299
rect 27134 4325 27162 4326
rect 27134 4299 27136 4325
rect 27136 4299 27162 4325
rect 27134 4298 27162 4299
rect 27186 4325 27214 4326
rect 27238 4325 27266 4326
rect 27186 4299 27198 4325
rect 27198 4299 27214 4325
rect 27238 4299 27260 4325
rect 27260 4299 27266 4325
rect 27186 4298 27214 4299
rect 27238 4298 27266 4299
rect 27290 4298 27318 4326
rect 27342 4325 27370 4326
rect 27394 4325 27422 4326
rect 27342 4299 27348 4325
rect 27348 4299 27370 4325
rect 27394 4299 27410 4325
rect 27410 4299 27422 4325
rect 27342 4298 27370 4299
rect 27394 4298 27422 4299
rect 27446 4325 27474 4326
rect 27446 4299 27472 4325
rect 27472 4299 27474 4325
rect 27446 4298 27474 4299
rect 27498 4325 27526 4326
rect 27498 4299 27508 4325
rect 27508 4299 27526 4325
rect 27498 4298 27526 4299
rect 27398 4129 27426 4130
rect 27398 4103 27399 4129
rect 27399 4103 27425 4129
rect 27425 4103 27426 4129
rect 27398 4102 27426 4103
rect 27678 4102 27706 4130
rect 27174 3710 27202 3738
rect 27082 3541 27110 3542
rect 27082 3515 27100 3541
rect 27100 3515 27110 3541
rect 27082 3514 27110 3515
rect 27134 3541 27162 3542
rect 27134 3515 27136 3541
rect 27136 3515 27162 3541
rect 27134 3514 27162 3515
rect 27186 3541 27214 3542
rect 27238 3541 27266 3542
rect 27186 3515 27198 3541
rect 27198 3515 27214 3541
rect 27238 3515 27260 3541
rect 27260 3515 27266 3541
rect 27186 3514 27214 3515
rect 27238 3514 27266 3515
rect 27290 3514 27318 3542
rect 27342 3541 27370 3542
rect 27394 3541 27422 3542
rect 27342 3515 27348 3541
rect 27348 3515 27370 3541
rect 27394 3515 27410 3541
rect 27410 3515 27422 3541
rect 27342 3514 27370 3515
rect 27394 3514 27422 3515
rect 27446 3541 27474 3542
rect 27446 3515 27472 3541
rect 27472 3515 27474 3541
rect 27446 3514 27474 3515
rect 27498 3541 27526 3542
rect 27498 3515 27508 3541
rect 27508 3515 27526 3541
rect 27498 3514 27526 3515
rect 27174 3374 27202 3402
rect 27398 3374 27426 3402
rect 28406 5305 28434 5306
rect 28406 5279 28407 5305
rect 28407 5279 28433 5305
rect 28433 5279 28434 5305
rect 28406 5278 28434 5279
rect 28126 4521 28154 4522
rect 28126 4495 28127 4521
rect 28127 4495 28153 4521
rect 28153 4495 28154 4521
rect 28126 4494 28154 4495
rect 28350 3793 28378 3794
rect 28350 3767 28351 3793
rect 28351 3767 28377 3793
rect 28377 3767 28378 3793
rect 28350 3766 28378 3767
rect 27082 2757 27110 2758
rect 27082 2731 27100 2757
rect 27100 2731 27110 2757
rect 27082 2730 27110 2731
rect 27134 2757 27162 2758
rect 27134 2731 27136 2757
rect 27136 2731 27162 2757
rect 27134 2730 27162 2731
rect 27186 2757 27214 2758
rect 27238 2757 27266 2758
rect 27186 2731 27198 2757
rect 27198 2731 27214 2757
rect 27238 2731 27260 2757
rect 27260 2731 27266 2757
rect 27186 2730 27214 2731
rect 27238 2730 27266 2731
rect 27290 2730 27318 2758
rect 27342 2757 27370 2758
rect 27394 2757 27422 2758
rect 27342 2731 27348 2757
rect 27348 2731 27370 2757
rect 27394 2731 27410 2757
rect 27410 2731 27422 2757
rect 27342 2730 27370 2731
rect 27394 2730 27422 2731
rect 27446 2757 27474 2758
rect 27446 2731 27472 2757
rect 27472 2731 27474 2757
rect 27446 2730 27474 2731
rect 27498 2757 27526 2758
rect 27498 2731 27508 2757
rect 27508 2731 27526 2757
rect 27498 2730 27526 2731
rect 27174 2646 27202 2674
rect 28238 2478 28266 2506
rect 28350 3262 28378 3290
rect 28966 9617 28994 9618
rect 28966 9591 28967 9617
rect 28967 9591 28993 9617
rect 28993 9591 28994 9617
rect 28966 9590 28994 9591
rect 29022 9225 29050 9226
rect 29022 9199 29023 9225
rect 29023 9199 29049 9225
rect 29049 9199 29050 9225
rect 29022 9198 29050 9199
rect 29134 10345 29162 10346
rect 29134 10319 29135 10345
rect 29135 10319 29161 10345
rect 29161 10319 29162 10345
rect 29134 10318 29162 10319
rect 29582 10989 29610 10990
rect 29582 10963 29600 10989
rect 29600 10963 29610 10989
rect 29582 10962 29610 10963
rect 29634 10989 29662 10990
rect 29634 10963 29636 10989
rect 29636 10963 29662 10989
rect 29634 10962 29662 10963
rect 29686 10989 29714 10990
rect 29738 10989 29766 10990
rect 29686 10963 29698 10989
rect 29698 10963 29714 10989
rect 29738 10963 29760 10989
rect 29760 10963 29766 10989
rect 29686 10962 29714 10963
rect 29738 10962 29766 10963
rect 29790 10962 29818 10990
rect 29842 10989 29870 10990
rect 29894 10989 29922 10990
rect 29842 10963 29848 10989
rect 29848 10963 29870 10989
rect 29894 10963 29910 10989
rect 29910 10963 29922 10989
rect 29842 10962 29870 10963
rect 29894 10962 29922 10963
rect 29946 10989 29974 10990
rect 29946 10963 29972 10989
rect 29972 10963 29974 10989
rect 29946 10962 29974 10963
rect 29998 10989 30026 10990
rect 29998 10963 30008 10989
rect 30008 10963 30026 10989
rect 29998 10962 30026 10963
rect 29918 10793 29946 10794
rect 29918 10767 29919 10793
rect 29919 10767 29945 10793
rect 29945 10767 29946 10793
rect 29918 10766 29946 10767
rect 30478 11577 30506 11578
rect 30478 11551 30479 11577
rect 30479 11551 30505 11577
rect 30505 11551 30506 11577
rect 30478 11550 30506 11551
rect 31374 11969 31402 11970
rect 31374 11943 31375 11969
rect 31375 11943 31401 11969
rect 31401 11943 31402 11969
rect 31374 11942 31402 11943
rect 30982 11550 31010 11578
rect 30702 11214 30730 11242
rect 31374 11494 31402 11522
rect 32082 18437 32110 18438
rect 32082 18411 32100 18437
rect 32100 18411 32110 18437
rect 32082 18410 32110 18411
rect 32134 18437 32162 18438
rect 32134 18411 32136 18437
rect 32136 18411 32162 18437
rect 32134 18410 32162 18411
rect 32186 18437 32214 18438
rect 32238 18437 32266 18438
rect 32186 18411 32198 18437
rect 32198 18411 32214 18437
rect 32238 18411 32260 18437
rect 32260 18411 32266 18437
rect 32186 18410 32214 18411
rect 32238 18410 32266 18411
rect 32290 18410 32318 18438
rect 32342 18437 32370 18438
rect 32394 18437 32422 18438
rect 32342 18411 32348 18437
rect 32348 18411 32370 18437
rect 32394 18411 32410 18437
rect 32410 18411 32422 18437
rect 32342 18410 32370 18411
rect 32394 18410 32422 18411
rect 32446 18437 32474 18438
rect 32446 18411 32472 18437
rect 32472 18411 32474 18437
rect 32446 18410 32474 18411
rect 32498 18437 32526 18438
rect 32498 18411 32508 18437
rect 32508 18411 32526 18437
rect 32498 18410 32526 18411
rect 34582 18045 34610 18046
rect 34582 18019 34600 18045
rect 34600 18019 34610 18045
rect 34582 18018 34610 18019
rect 34634 18045 34662 18046
rect 34634 18019 34636 18045
rect 34636 18019 34662 18045
rect 34634 18018 34662 18019
rect 34686 18045 34714 18046
rect 34738 18045 34766 18046
rect 34686 18019 34698 18045
rect 34698 18019 34714 18045
rect 34738 18019 34760 18045
rect 34760 18019 34766 18045
rect 34686 18018 34714 18019
rect 34738 18018 34766 18019
rect 34790 18018 34818 18046
rect 34842 18045 34870 18046
rect 34894 18045 34922 18046
rect 34842 18019 34848 18045
rect 34848 18019 34870 18045
rect 34894 18019 34910 18045
rect 34910 18019 34922 18045
rect 34842 18018 34870 18019
rect 34894 18018 34922 18019
rect 34946 18045 34974 18046
rect 34946 18019 34972 18045
rect 34972 18019 34974 18045
rect 34946 18018 34974 18019
rect 34998 18045 35026 18046
rect 34998 18019 35008 18045
rect 35008 18019 35026 18045
rect 34998 18018 35026 18019
rect 32082 17653 32110 17654
rect 32082 17627 32100 17653
rect 32100 17627 32110 17653
rect 32082 17626 32110 17627
rect 32134 17653 32162 17654
rect 32134 17627 32136 17653
rect 32136 17627 32162 17653
rect 32134 17626 32162 17627
rect 32186 17653 32214 17654
rect 32238 17653 32266 17654
rect 32186 17627 32198 17653
rect 32198 17627 32214 17653
rect 32238 17627 32260 17653
rect 32260 17627 32266 17653
rect 32186 17626 32214 17627
rect 32238 17626 32266 17627
rect 32290 17626 32318 17654
rect 32342 17653 32370 17654
rect 32394 17653 32422 17654
rect 32342 17627 32348 17653
rect 32348 17627 32370 17653
rect 32394 17627 32410 17653
rect 32410 17627 32422 17653
rect 32342 17626 32370 17627
rect 32394 17626 32422 17627
rect 32446 17653 32474 17654
rect 32446 17627 32472 17653
rect 32472 17627 32474 17653
rect 32446 17626 32474 17627
rect 32498 17653 32526 17654
rect 32498 17627 32508 17653
rect 32508 17627 32526 17653
rect 32498 17626 32526 17627
rect 34582 17261 34610 17262
rect 34582 17235 34600 17261
rect 34600 17235 34610 17261
rect 34582 17234 34610 17235
rect 34634 17261 34662 17262
rect 34634 17235 34636 17261
rect 34636 17235 34662 17261
rect 34634 17234 34662 17235
rect 34686 17261 34714 17262
rect 34738 17261 34766 17262
rect 34686 17235 34698 17261
rect 34698 17235 34714 17261
rect 34738 17235 34760 17261
rect 34760 17235 34766 17261
rect 34686 17234 34714 17235
rect 34738 17234 34766 17235
rect 34790 17234 34818 17262
rect 34842 17261 34870 17262
rect 34894 17261 34922 17262
rect 34842 17235 34848 17261
rect 34848 17235 34870 17261
rect 34894 17235 34910 17261
rect 34910 17235 34922 17261
rect 34842 17234 34870 17235
rect 34894 17234 34922 17235
rect 34946 17261 34974 17262
rect 34946 17235 34972 17261
rect 34972 17235 34974 17261
rect 34946 17234 34974 17235
rect 34998 17261 35026 17262
rect 34998 17235 35008 17261
rect 35008 17235 35026 17261
rect 34998 17234 35026 17235
rect 32082 16869 32110 16870
rect 32082 16843 32100 16869
rect 32100 16843 32110 16869
rect 32082 16842 32110 16843
rect 32134 16869 32162 16870
rect 32134 16843 32136 16869
rect 32136 16843 32162 16869
rect 32134 16842 32162 16843
rect 32186 16869 32214 16870
rect 32238 16869 32266 16870
rect 32186 16843 32198 16869
rect 32198 16843 32214 16869
rect 32238 16843 32260 16869
rect 32260 16843 32266 16869
rect 32186 16842 32214 16843
rect 32238 16842 32266 16843
rect 32290 16842 32318 16870
rect 32342 16869 32370 16870
rect 32394 16869 32422 16870
rect 32342 16843 32348 16869
rect 32348 16843 32370 16869
rect 32394 16843 32410 16869
rect 32410 16843 32422 16869
rect 32342 16842 32370 16843
rect 32394 16842 32422 16843
rect 32446 16869 32474 16870
rect 32446 16843 32472 16869
rect 32472 16843 32474 16869
rect 32446 16842 32474 16843
rect 32498 16869 32526 16870
rect 32498 16843 32508 16869
rect 32508 16843 32526 16869
rect 32498 16842 32526 16843
rect 34582 16477 34610 16478
rect 34582 16451 34600 16477
rect 34600 16451 34610 16477
rect 34582 16450 34610 16451
rect 34634 16477 34662 16478
rect 34634 16451 34636 16477
rect 34636 16451 34662 16477
rect 34634 16450 34662 16451
rect 34686 16477 34714 16478
rect 34738 16477 34766 16478
rect 34686 16451 34698 16477
rect 34698 16451 34714 16477
rect 34738 16451 34760 16477
rect 34760 16451 34766 16477
rect 34686 16450 34714 16451
rect 34738 16450 34766 16451
rect 34790 16450 34818 16478
rect 34842 16477 34870 16478
rect 34894 16477 34922 16478
rect 34842 16451 34848 16477
rect 34848 16451 34870 16477
rect 34894 16451 34910 16477
rect 34910 16451 34922 16477
rect 34842 16450 34870 16451
rect 34894 16450 34922 16451
rect 34946 16477 34974 16478
rect 34946 16451 34972 16477
rect 34972 16451 34974 16477
rect 34946 16450 34974 16451
rect 34998 16477 35026 16478
rect 34998 16451 35008 16477
rect 35008 16451 35026 16477
rect 34998 16450 35026 16451
rect 32082 16085 32110 16086
rect 32082 16059 32100 16085
rect 32100 16059 32110 16085
rect 32082 16058 32110 16059
rect 32134 16085 32162 16086
rect 32134 16059 32136 16085
rect 32136 16059 32162 16085
rect 32134 16058 32162 16059
rect 32186 16085 32214 16086
rect 32238 16085 32266 16086
rect 32186 16059 32198 16085
rect 32198 16059 32214 16085
rect 32238 16059 32260 16085
rect 32260 16059 32266 16085
rect 32186 16058 32214 16059
rect 32238 16058 32266 16059
rect 32290 16058 32318 16086
rect 32342 16085 32370 16086
rect 32394 16085 32422 16086
rect 32342 16059 32348 16085
rect 32348 16059 32370 16085
rect 32394 16059 32410 16085
rect 32410 16059 32422 16085
rect 32342 16058 32370 16059
rect 32394 16058 32422 16059
rect 32446 16085 32474 16086
rect 32446 16059 32472 16085
rect 32472 16059 32474 16085
rect 32446 16058 32474 16059
rect 32498 16085 32526 16086
rect 32498 16059 32508 16085
rect 32508 16059 32526 16085
rect 32498 16058 32526 16059
rect 34582 15693 34610 15694
rect 34582 15667 34600 15693
rect 34600 15667 34610 15693
rect 34582 15666 34610 15667
rect 34634 15693 34662 15694
rect 34634 15667 34636 15693
rect 34636 15667 34662 15693
rect 34634 15666 34662 15667
rect 34686 15693 34714 15694
rect 34738 15693 34766 15694
rect 34686 15667 34698 15693
rect 34698 15667 34714 15693
rect 34738 15667 34760 15693
rect 34760 15667 34766 15693
rect 34686 15666 34714 15667
rect 34738 15666 34766 15667
rect 34790 15666 34818 15694
rect 34842 15693 34870 15694
rect 34894 15693 34922 15694
rect 34842 15667 34848 15693
rect 34848 15667 34870 15693
rect 34894 15667 34910 15693
rect 34910 15667 34922 15693
rect 34842 15666 34870 15667
rect 34894 15666 34922 15667
rect 34946 15693 34974 15694
rect 34946 15667 34972 15693
rect 34972 15667 34974 15693
rect 34946 15666 34974 15667
rect 34998 15693 35026 15694
rect 34998 15667 35008 15693
rect 35008 15667 35026 15693
rect 34998 15666 35026 15667
rect 32082 15301 32110 15302
rect 32082 15275 32100 15301
rect 32100 15275 32110 15301
rect 32082 15274 32110 15275
rect 32134 15301 32162 15302
rect 32134 15275 32136 15301
rect 32136 15275 32162 15301
rect 32134 15274 32162 15275
rect 32186 15301 32214 15302
rect 32238 15301 32266 15302
rect 32186 15275 32198 15301
rect 32198 15275 32214 15301
rect 32238 15275 32260 15301
rect 32260 15275 32266 15301
rect 32186 15274 32214 15275
rect 32238 15274 32266 15275
rect 32290 15274 32318 15302
rect 32342 15301 32370 15302
rect 32394 15301 32422 15302
rect 32342 15275 32348 15301
rect 32348 15275 32370 15301
rect 32394 15275 32410 15301
rect 32410 15275 32422 15301
rect 32342 15274 32370 15275
rect 32394 15274 32422 15275
rect 32446 15301 32474 15302
rect 32446 15275 32472 15301
rect 32472 15275 32474 15301
rect 32446 15274 32474 15275
rect 32498 15301 32526 15302
rect 32498 15275 32508 15301
rect 32508 15275 32526 15301
rect 32498 15274 32526 15275
rect 34582 14909 34610 14910
rect 34582 14883 34600 14909
rect 34600 14883 34610 14909
rect 34582 14882 34610 14883
rect 34634 14909 34662 14910
rect 34634 14883 34636 14909
rect 34636 14883 34662 14909
rect 34634 14882 34662 14883
rect 34686 14909 34714 14910
rect 34738 14909 34766 14910
rect 34686 14883 34698 14909
rect 34698 14883 34714 14909
rect 34738 14883 34760 14909
rect 34760 14883 34766 14909
rect 34686 14882 34714 14883
rect 34738 14882 34766 14883
rect 34790 14882 34818 14910
rect 34842 14909 34870 14910
rect 34894 14909 34922 14910
rect 34842 14883 34848 14909
rect 34848 14883 34870 14909
rect 34894 14883 34910 14909
rect 34910 14883 34922 14909
rect 34842 14882 34870 14883
rect 34894 14882 34922 14883
rect 34946 14909 34974 14910
rect 34946 14883 34972 14909
rect 34972 14883 34974 14909
rect 34946 14882 34974 14883
rect 34998 14909 35026 14910
rect 34998 14883 35008 14909
rect 35008 14883 35026 14909
rect 34998 14882 35026 14883
rect 32082 14517 32110 14518
rect 32082 14491 32100 14517
rect 32100 14491 32110 14517
rect 32082 14490 32110 14491
rect 32134 14517 32162 14518
rect 32134 14491 32136 14517
rect 32136 14491 32162 14517
rect 32134 14490 32162 14491
rect 32186 14517 32214 14518
rect 32238 14517 32266 14518
rect 32186 14491 32198 14517
rect 32198 14491 32214 14517
rect 32238 14491 32260 14517
rect 32260 14491 32266 14517
rect 32186 14490 32214 14491
rect 32238 14490 32266 14491
rect 32290 14490 32318 14518
rect 32342 14517 32370 14518
rect 32394 14517 32422 14518
rect 32342 14491 32348 14517
rect 32348 14491 32370 14517
rect 32394 14491 32410 14517
rect 32410 14491 32422 14517
rect 32342 14490 32370 14491
rect 32394 14490 32422 14491
rect 32446 14517 32474 14518
rect 32446 14491 32472 14517
rect 32472 14491 32474 14517
rect 32446 14490 32474 14491
rect 32498 14517 32526 14518
rect 32498 14491 32508 14517
rect 32508 14491 32526 14517
rect 32498 14490 32526 14491
rect 34582 14125 34610 14126
rect 34582 14099 34600 14125
rect 34600 14099 34610 14125
rect 34582 14098 34610 14099
rect 34634 14125 34662 14126
rect 34634 14099 34636 14125
rect 34636 14099 34662 14125
rect 34634 14098 34662 14099
rect 34686 14125 34714 14126
rect 34738 14125 34766 14126
rect 34686 14099 34698 14125
rect 34698 14099 34714 14125
rect 34738 14099 34760 14125
rect 34760 14099 34766 14125
rect 34686 14098 34714 14099
rect 34738 14098 34766 14099
rect 34790 14098 34818 14126
rect 34842 14125 34870 14126
rect 34894 14125 34922 14126
rect 34842 14099 34848 14125
rect 34848 14099 34870 14125
rect 34894 14099 34910 14125
rect 34910 14099 34922 14125
rect 34842 14098 34870 14099
rect 34894 14098 34922 14099
rect 34946 14125 34974 14126
rect 34946 14099 34972 14125
rect 34972 14099 34974 14125
rect 34946 14098 34974 14099
rect 34998 14125 35026 14126
rect 34998 14099 35008 14125
rect 35008 14099 35026 14125
rect 34998 14098 35026 14099
rect 32082 13733 32110 13734
rect 32082 13707 32100 13733
rect 32100 13707 32110 13733
rect 32082 13706 32110 13707
rect 32134 13733 32162 13734
rect 32134 13707 32136 13733
rect 32136 13707 32162 13733
rect 32134 13706 32162 13707
rect 32186 13733 32214 13734
rect 32238 13733 32266 13734
rect 32186 13707 32198 13733
rect 32198 13707 32214 13733
rect 32238 13707 32260 13733
rect 32260 13707 32266 13733
rect 32186 13706 32214 13707
rect 32238 13706 32266 13707
rect 32290 13706 32318 13734
rect 32342 13733 32370 13734
rect 32394 13733 32422 13734
rect 32342 13707 32348 13733
rect 32348 13707 32370 13733
rect 32394 13707 32410 13733
rect 32410 13707 32422 13733
rect 32342 13706 32370 13707
rect 32394 13706 32422 13707
rect 32446 13733 32474 13734
rect 32446 13707 32472 13733
rect 32472 13707 32474 13733
rect 32446 13706 32474 13707
rect 32498 13733 32526 13734
rect 32498 13707 32508 13733
rect 32508 13707 32526 13733
rect 32498 13706 32526 13707
rect 34582 13341 34610 13342
rect 34582 13315 34600 13341
rect 34600 13315 34610 13341
rect 34582 13314 34610 13315
rect 34634 13341 34662 13342
rect 34634 13315 34636 13341
rect 34636 13315 34662 13341
rect 34634 13314 34662 13315
rect 34686 13341 34714 13342
rect 34738 13341 34766 13342
rect 34686 13315 34698 13341
rect 34698 13315 34714 13341
rect 34738 13315 34760 13341
rect 34760 13315 34766 13341
rect 34686 13314 34714 13315
rect 34738 13314 34766 13315
rect 34790 13314 34818 13342
rect 34842 13341 34870 13342
rect 34894 13341 34922 13342
rect 34842 13315 34848 13341
rect 34848 13315 34870 13341
rect 34894 13315 34910 13341
rect 34910 13315 34922 13341
rect 34842 13314 34870 13315
rect 34894 13314 34922 13315
rect 34946 13341 34974 13342
rect 34946 13315 34972 13341
rect 34972 13315 34974 13341
rect 34946 13314 34974 13315
rect 34998 13341 35026 13342
rect 34998 13315 35008 13341
rect 35008 13315 35026 13341
rect 34998 13314 35026 13315
rect 32082 12949 32110 12950
rect 32082 12923 32100 12949
rect 32100 12923 32110 12949
rect 32082 12922 32110 12923
rect 32134 12949 32162 12950
rect 32134 12923 32136 12949
rect 32136 12923 32162 12949
rect 32134 12922 32162 12923
rect 32186 12949 32214 12950
rect 32238 12949 32266 12950
rect 32186 12923 32198 12949
rect 32198 12923 32214 12949
rect 32238 12923 32260 12949
rect 32260 12923 32266 12949
rect 32186 12922 32214 12923
rect 32238 12922 32266 12923
rect 32290 12922 32318 12950
rect 32342 12949 32370 12950
rect 32394 12949 32422 12950
rect 32342 12923 32348 12949
rect 32348 12923 32370 12949
rect 32394 12923 32410 12949
rect 32410 12923 32422 12949
rect 32342 12922 32370 12923
rect 32394 12922 32422 12923
rect 32446 12949 32474 12950
rect 32446 12923 32472 12949
rect 32472 12923 32474 12949
rect 32446 12922 32474 12923
rect 32498 12949 32526 12950
rect 32498 12923 32508 12949
rect 32508 12923 32526 12949
rect 32498 12922 32526 12923
rect 34582 12557 34610 12558
rect 34582 12531 34600 12557
rect 34600 12531 34610 12557
rect 34582 12530 34610 12531
rect 34634 12557 34662 12558
rect 34634 12531 34636 12557
rect 34636 12531 34662 12557
rect 34634 12530 34662 12531
rect 34686 12557 34714 12558
rect 34738 12557 34766 12558
rect 34686 12531 34698 12557
rect 34698 12531 34714 12557
rect 34738 12531 34760 12557
rect 34760 12531 34766 12557
rect 34686 12530 34714 12531
rect 34738 12530 34766 12531
rect 34790 12530 34818 12558
rect 34842 12557 34870 12558
rect 34894 12557 34922 12558
rect 34842 12531 34848 12557
rect 34848 12531 34870 12557
rect 34894 12531 34910 12557
rect 34910 12531 34922 12557
rect 34842 12530 34870 12531
rect 34894 12530 34922 12531
rect 34946 12557 34974 12558
rect 34946 12531 34972 12557
rect 34972 12531 34974 12557
rect 34946 12530 34974 12531
rect 34998 12557 35026 12558
rect 34998 12531 35008 12557
rect 35008 12531 35026 12557
rect 34998 12530 35026 12531
rect 32082 12165 32110 12166
rect 32082 12139 32100 12165
rect 32100 12139 32110 12165
rect 32082 12138 32110 12139
rect 32134 12165 32162 12166
rect 32134 12139 32136 12165
rect 32136 12139 32162 12165
rect 32134 12138 32162 12139
rect 32186 12165 32214 12166
rect 32238 12165 32266 12166
rect 32186 12139 32198 12165
rect 32198 12139 32214 12165
rect 32238 12139 32260 12165
rect 32260 12139 32266 12165
rect 32186 12138 32214 12139
rect 32238 12138 32266 12139
rect 32290 12138 32318 12166
rect 32342 12165 32370 12166
rect 32394 12165 32422 12166
rect 32342 12139 32348 12165
rect 32348 12139 32370 12165
rect 32394 12139 32410 12165
rect 32410 12139 32422 12165
rect 32342 12138 32370 12139
rect 32394 12138 32422 12139
rect 32446 12165 32474 12166
rect 32446 12139 32472 12165
rect 32472 12139 32474 12165
rect 32446 12138 32474 12139
rect 32498 12165 32526 12166
rect 32498 12139 32508 12165
rect 32508 12139 32526 12165
rect 32498 12138 32526 12139
rect 31934 11382 31962 11410
rect 32830 11969 32858 11970
rect 32830 11943 32831 11969
rect 32831 11943 32857 11969
rect 32857 11943 32858 11969
rect 32830 11942 32858 11943
rect 33110 11942 33138 11970
rect 31990 11550 32018 11578
rect 31934 11214 31962 11242
rect 30982 11158 31010 11186
rect 31094 11102 31122 11130
rect 30086 10766 30114 10794
rect 30254 10710 30282 10738
rect 30702 10710 30730 10738
rect 30702 10401 30730 10402
rect 30702 10375 30703 10401
rect 30703 10375 30729 10401
rect 30729 10375 30730 10401
rect 30702 10374 30730 10375
rect 29582 10205 29610 10206
rect 29582 10179 29600 10205
rect 29600 10179 29610 10205
rect 29582 10178 29610 10179
rect 29634 10205 29662 10206
rect 29634 10179 29636 10205
rect 29636 10179 29662 10205
rect 29634 10178 29662 10179
rect 29686 10205 29714 10206
rect 29738 10205 29766 10206
rect 29686 10179 29698 10205
rect 29698 10179 29714 10205
rect 29738 10179 29760 10205
rect 29760 10179 29766 10205
rect 29686 10178 29714 10179
rect 29738 10178 29766 10179
rect 29790 10178 29818 10206
rect 29842 10205 29870 10206
rect 29894 10205 29922 10206
rect 29842 10179 29848 10205
rect 29848 10179 29870 10205
rect 29894 10179 29910 10205
rect 29910 10179 29922 10205
rect 29842 10178 29870 10179
rect 29894 10178 29922 10179
rect 29946 10205 29974 10206
rect 29946 10179 29972 10205
rect 29972 10179 29974 10205
rect 29946 10178 29974 10179
rect 29998 10205 30026 10206
rect 29998 10179 30008 10205
rect 30008 10179 30026 10205
rect 29998 10178 30026 10179
rect 31374 10766 31402 10794
rect 31934 10430 31962 10458
rect 29302 10009 29330 10010
rect 29302 9983 29303 10009
rect 29303 9983 29329 10009
rect 29329 9983 29330 10009
rect 29302 9982 29330 9983
rect 29078 9086 29106 9114
rect 29414 9590 29442 9618
rect 29414 9254 29442 9282
rect 29358 8470 29386 8498
rect 29022 8022 29050 8050
rect 31094 10038 31122 10066
rect 29582 9421 29610 9422
rect 29582 9395 29600 9421
rect 29600 9395 29610 9421
rect 29582 9394 29610 9395
rect 29634 9421 29662 9422
rect 29634 9395 29636 9421
rect 29636 9395 29662 9421
rect 29634 9394 29662 9395
rect 29686 9421 29714 9422
rect 29738 9421 29766 9422
rect 29686 9395 29698 9421
rect 29698 9395 29714 9421
rect 29738 9395 29760 9421
rect 29760 9395 29766 9421
rect 29686 9394 29714 9395
rect 29738 9394 29766 9395
rect 29790 9394 29818 9422
rect 29842 9421 29870 9422
rect 29894 9421 29922 9422
rect 29842 9395 29848 9421
rect 29848 9395 29870 9421
rect 29894 9395 29910 9421
rect 29910 9395 29922 9421
rect 29842 9394 29870 9395
rect 29894 9394 29922 9395
rect 29946 9421 29974 9422
rect 29946 9395 29972 9421
rect 29972 9395 29974 9421
rect 29946 9394 29974 9395
rect 29998 9421 30026 9422
rect 29998 9395 30008 9421
rect 30008 9395 30026 9421
rect 29998 9394 30026 9395
rect 29694 9281 29722 9282
rect 29694 9255 29695 9281
rect 29695 9255 29721 9281
rect 29721 9255 29722 9281
rect 29694 9254 29722 9255
rect 31038 9702 31066 9730
rect 30422 9086 30450 9114
rect 30478 9198 30506 9226
rect 29582 8637 29610 8638
rect 29582 8611 29600 8637
rect 29600 8611 29610 8637
rect 29582 8610 29610 8611
rect 29634 8637 29662 8638
rect 29634 8611 29636 8637
rect 29636 8611 29662 8637
rect 29634 8610 29662 8611
rect 29686 8637 29714 8638
rect 29738 8637 29766 8638
rect 29686 8611 29698 8637
rect 29698 8611 29714 8637
rect 29738 8611 29760 8637
rect 29760 8611 29766 8637
rect 29686 8610 29714 8611
rect 29738 8610 29766 8611
rect 29790 8610 29818 8638
rect 29842 8637 29870 8638
rect 29894 8637 29922 8638
rect 29842 8611 29848 8637
rect 29848 8611 29870 8637
rect 29894 8611 29910 8637
rect 29910 8611 29922 8637
rect 29842 8610 29870 8611
rect 29894 8610 29922 8611
rect 29946 8637 29974 8638
rect 29946 8611 29972 8637
rect 29972 8611 29974 8637
rect 29946 8610 29974 8611
rect 29998 8637 30026 8638
rect 29998 8611 30008 8637
rect 30008 8611 30026 8637
rect 29998 8610 30026 8611
rect 29918 8497 29946 8498
rect 29918 8471 29919 8497
rect 29919 8471 29945 8497
rect 29945 8471 29946 8497
rect 29918 8470 29946 8471
rect 28742 6873 28770 6874
rect 28742 6847 28743 6873
rect 28743 6847 28769 6873
rect 28769 6847 28770 6873
rect 28742 6846 28770 6847
rect 29582 7853 29610 7854
rect 29582 7827 29600 7853
rect 29600 7827 29610 7853
rect 29582 7826 29610 7827
rect 29634 7853 29662 7854
rect 29634 7827 29636 7853
rect 29636 7827 29662 7853
rect 29634 7826 29662 7827
rect 29686 7853 29714 7854
rect 29738 7853 29766 7854
rect 29686 7827 29698 7853
rect 29698 7827 29714 7853
rect 29738 7827 29760 7853
rect 29760 7827 29766 7853
rect 29686 7826 29714 7827
rect 29738 7826 29766 7827
rect 29790 7826 29818 7854
rect 29842 7853 29870 7854
rect 29894 7853 29922 7854
rect 29842 7827 29848 7853
rect 29848 7827 29870 7853
rect 29894 7827 29910 7853
rect 29910 7827 29922 7853
rect 29842 7826 29870 7827
rect 29894 7826 29922 7827
rect 29946 7853 29974 7854
rect 29946 7827 29972 7853
rect 29972 7827 29974 7853
rect 29946 7826 29974 7827
rect 29998 7853 30026 7854
rect 29998 7827 30008 7853
rect 30008 7827 30026 7853
rect 29998 7826 30026 7827
rect 29022 6790 29050 6818
rect 28686 6734 28714 6762
rect 29190 6734 29218 6762
rect 30982 9086 31010 9114
rect 31094 9590 31122 9618
rect 31038 8862 31066 8890
rect 30982 8414 31010 8442
rect 31262 10065 31290 10066
rect 31262 10039 31263 10065
rect 31263 10039 31289 10065
rect 31289 10039 31290 10065
rect 31262 10038 31290 10039
rect 31374 9617 31402 9618
rect 31374 9591 31375 9617
rect 31375 9591 31401 9617
rect 31401 9591 31402 9617
rect 31374 9590 31402 9591
rect 32774 11577 32802 11578
rect 32774 11551 32775 11577
rect 32775 11551 32801 11577
rect 32801 11551 32802 11577
rect 32774 11550 32802 11551
rect 32082 11381 32110 11382
rect 32082 11355 32100 11381
rect 32100 11355 32110 11381
rect 32082 11354 32110 11355
rect 32134 11381 32162 11382
rect 32134 11355 32136 11381
rect 32136 11355 32162 11381
rect 32134 11354 32162 11355
rect 32186 11381 32214 11382
rect 32238 11381 32266 11382
rect 32186 11355 32198 11381
rect 32198 11355 32214 11381
rect 32238 11355 32260 11381
rect 32260 11355 32266 11381
rect 32186 11354 32214 11355
rect 32238 11354 32266 11355
rect 32290 11354 32318 11382
rect 32342 11381 32370 11382
rect 32394 11381 32422 11382
rect 32342 11355 32348 11381
rect 32348 11355 32370 11381
rect 32394 11355 32410 11381
rect 32410 11355 32422 11381
rect 32342 11354 32370 11355
rect 32394 11354 32422 11355
rect 32446 11381 32474 11382
rect 32446 11355 32472 11381
rect 32472 11355 32474 11381
rect 32446 11354 32474 11355
rect 32498 11381 32526 11382
rect 32498 11355 32508 11381
rect 32508 11355 32526 11381
rect 32498 11354 32526 11355
rect 32438 11185 32466 11186
rect 32438 11159 32439 11185
rect 32439 11159 32465 11185
rect 32465 11159 32466 11185
rect 32438 11158 32466 11159
rect 32998 11158 33026 11186
rect 34582 11773 34610 11774
rect 34582 11747 34600 11773
rect 34600 11747 34610 11773
rect 34582 11746 34610 11747
rect 34634 11773 34662 11774
rect 34634 11747 34636 11773
rect 34636 11747 34662 11773
rect 34634 11746 34662 11747
rect 34686 11773 34714 11774
rect 34738 11773 34766 11774
rect 34686 11747 34698 11773
rect 34698 11747 34714 11773
rect 34738 11747 34760 11773
rect 34760 11747 34766 11773
rect 34686 11746 34714 11747
rect 34738 11746 34766 11747
rect 34790 11746 34818 11774
rect 34842 11773 34870 11774
rect 34894 11773 34922 11774
rect 34842 11747 34848 11773
rect 34848 11747 34870 11773
rect 34894 11747 34910 11773
rect 34910 11747 34922 11773
rect 34842 11746 34870 11747
rect 34894 11746 34922 11747
rect 34946 11773 34974 11774
rect 34946 11747 34972 11773
rect 34972 11747 34974 11773
rect 34946 11746 34974 11747
rect 34998 11773 35026 11774
rect 34998 11747 35008 11773
rect 35008 11747 35026 11773
rect 34998 11746 35026 11747
rect 33110 11129 33138 11130
rect 33110 11103 33111 11129
rect 33111 11103 33137 11129
rect 33137 11103 33138 11129
rect 33110 11102 33138 11103
rect 35294 11494 35322 11522
rect 34958 11185 34986 11186
rect 34958 11159 34959 11185
rect 34959 11159 34985 11185
rect 34985 11159 34986 11185
rect 34958 11158 34986 11159
rect 37082 18437 37110 18438
rect 37082 18411 37100 18437
rect 37100 18411 37110 18437
rect 37082 18410 37110 18411
rect 37134 18437 37162 18438
rect 37134 18411 37136 18437
rect 37136 18411 37162 18437
rect 37134 18410 37162 18411
rect 37186 18437 37214 18438
rect 37238 18437 37266 18438
rect 37186 18411 37198 18437
rect 37198 18411 37214 18437
rect 37238 18411 37260 18437
rect 37260 18411 37266 18437
rect 37186 18410 37214 18411
rect 37238 18410 37266 18411
rect 37290 18410 37318 18438
rect 37342 18437 37370 18438
rect 37394 18437 37422 18438
rect 37342 18411 37348 18437
rect 37348 18411 37370 18437
rect 37394 18411 37410 18437
rect 37410 18411 37422 18437
rect 37342 18410 37370 18411
rect 37394 18410 37422 18411
rect 37446 18437 37474 18438
rect 37446 18411 37472 18437
rect 37472 18411 37474 18437
rect 37446 18410 37474 18411
rect 37498 18437 37526 18438
rect 37498 18411 37508 18437
rect 37508 18411 37526 18437
rect 37498 18410 37526 18411
rect 37082 17653 37110 17654
rect 37082 17627 37100 17653
rect 37100 17627 37110 17653
rect 37082 17626 37110 17627
rect 37134 17653 37162 17654
rect 37134 17627 37136 17653
rect 37136 17627 37162 17653
rect 37134 17626 37162 17627
rect 37186 17653 37214 17654
rect 37238 17653 37266 17654
rect 37186 17627 37198 17653
rect 37198 17627 37214 17653
rect 37238 17627 37260 17653
rect 37260 17627 37266 17653
rect 37186 17626 37214 17627
rect 37238 17626 37266 17627
rect 37290 17626 37318 17654
rect 37342 17653 37370 17654
rect 37394 17653 37422 17654
rect 37342 17627 37348 17653
rect 37348 17627 37370 17653
rect 37394 17627 37410 17653
rect 37410 17627 37422 17653
rect 37342 17626 37370 17627
rect 37394 17626 37422 17627
rect 37446 17653 37474 17654
rect 37446 17627 37472 17653
rect 37472 17627 37474 17653
rect 37446 17626 37474 17627
rect 37498 17653 37526 17654
rect 37498 17627 37508 17653
rect 37508 17627 37526 17653
rect 37498 17626 37526 17627
rect 37082 16869 37110 16870
rect 37082 16843 37100 16869
rect 37100 16843 37110 16869
rect 37082 16842 37110 16843
rect 37134 16869 37162 16870
rect 37134 16843 37136 16869
rect 37136 16843 37162 16869
rect 37134 16842 37162 16843
rect 37186 16869 37214 16870
rect 37238 16869 37266 16870
rect 37186 16843 37198 16869
rect 37198 16843 37214 16869
rect 37238 16843 37260 16869
rect 37260 16843 37266 16869
rect 37186 16842 37214 16843
rect 37238 16842 37266 16843
rect 37290 16842 37318 16870
rect 37342 16869 37370 16870
rect 37394 16869 37422 16870
rect 37342 16843 37348 16869
rect 37348 16843 37370 16869
rect 37394 16843 37410 16869
rect 37410 16843 37422 16869
rect 37342 16842 37370 16843
rect 37394 16842 37422 16843
rect 37446 16869 37474 16870
rect 37446 16843 37472 16869
rect 37472 16843 37474 16869
rect 37446 16842 37474 16843
rect 37498 16869 37526 16870
rect 37498 16843 37508 16869
rect 37508 16843 37526 16869
rect 37498 16842 37526 16843
rect 37082 16085 37110 16086
rect 37082 16059 37100 16085
rect 37100 16059 37110 16085
rect 37082 16058 37110 16059
rect 37134 16085 37162 16086
rect 37134 16059 37136 16085
rect 37136 16059 37162 16085
rect 37134 16058 37162 16059
rect 37186 16085 37214 16086
rect 37238 16085 37266 16086
rect 37186 16059 37198 16085
rect 37198 16059 37214 16085
rect 37238 16059 37260 16085
rect 37260 16059 37266 16085
rect 37186 16058 37214 16059
rect 37238 16058 37266 16059
rect 37290 16058 37318 16086
rect 37342 16085 37370 16086
rect 37394 16085 37422 16086
rect 37342 16059 37348 16085
rect 37348 16059 37370 16085
rect 37394 16059 37410 16085
rect 37410 16059 37422 16085
rect 37342 16058 37370 16059
rect 37394 16058 37422 16059
rect 37446 16085 37474 16086
rect 37446 16059 37472 16085
rect 37472 16059 37474 16085
rect 37446 16058 37474 16059
rect 37498 16085 37526 16086
rect 37498 16059 37508 16085
rect 37508 16059 37526 16085
rect 37498 16058 37526 16059
rect 37082 15301 37110 15302
rect 37082 15275 37100 15301
rect 37100 15275 37110 15301
rect 37082 15274 37110 15275
rect 37134 15301 37162 15302
rect 37134 15275 37136 15301
rect 37136 15275 37162 15301
rect 37134 15274 37162 15275
rect 37186 15301 37214 15302
rect 37238 15301 37266 15302
rect 37186 15275 37198 15301
rect 37198 15275 37214 15301
rect 37238 15275 37260 15301
rect 37260 15275 37266 15301
rect 37186 15274 37214 15275
rect 37238 15274 37266 15275
rect 37290 15274 37318 15302
rect 37342 15301 37370 15302
rect 37394 15301 37422 15302
rect 37342 15275 37348 15301
rect 37348 15275 37370 15301
rect 37394 15275 37410 15301
rect 37410 15275 37422 15301
rect 37342 15274 37370 15275
rect 37394 15274 37422 15275
rect 37446 15301 37474 15302
rect 37446 15275 37472 15301
rect 37472 15275 37474 15301
rect 37446 15274 37474 15275
rect 37498 15301 37526 15302
rect 37498 15275 37508 15301
rect 37508 15275 37526 15301
rect 37498 15274 37526 15275
rect 37082 14517 37110 14518
rect 37082 14491 37100 14517
rect 37100 14491 37110 14517
rect 37082 14490 37110 14491
rect 37134 14517 37162 14518
rect 37134 14491 37136 14517
rect 37136 14491 37162 14517
rect 37134 14490 37162 14491
rect 37186 14517 37214 14518
rect 37238 14517 37266 14518
rect 37186 14491 37198 14517
rect 37198 14491 37214 14517
rect 37238 14491 37260 14517
rect 37260 14491 37266 14517
rect 37186 14490 37214 14491
rect 37238 14490 37266 14491
rect 37290 14490 37318 14518
rect 37342 14517 37370 14518
rect 37394 14517 37422 14518
rect 37342 14491 37348 14517
rect 37348 14491 37370 14517
rect 37394 14491 37410 14517
rect 37410 14491 37422 14517
rect 37342 14490 37370 14491
rect 37394 14490 37422 14491
rect 37446 14517 37474 14518
rect 37446 14491 37472 14517
rect 37472 14491 37474 14517
rect 37446 14490 37474 14491
rect 37498 14517 37526 14518
rect 37498 14491 37508 14517
rect 37508 14491 37526 14517
rect 37498 14490 37526 14491
rect 37082 13733 37110 13734
rect 37082 13707 37100 13733
rect 37100 13707 37110 13733
rect 37082 13706 37110 13707
rect 37134 13733 37162 13734
rect 37134 13707 37136 13733
rect 37136 13707 37162 13733
rect 37134 13706 37162 13707
rect 37186 13733 37214 13734
rect 37238 13733 37266 13734
rect 37186 13707 37198 13733
rect 37198 13707 37214 13733
rect 37238 13707 37260 13733
rect 37260 13707 37266 13733
rect 37186 13706 37214 13707
rect 37238 13706 37266 13707
rect 37290 13706 37318 13734
rect 37342 13733 37370 13734
rect 37394 13733 37422 13734
rect 37342 13707 37348 13733
rect 37348 13707 37370 13733
rect 37394 13707 37410 13733
rect 37410 13707 37422 13733
rect 37342 13706 37370 13707
rect 37394 13706 37422 13707
rect 37446 13733 37474 13734
rect 37446 13707 37472 13733
rect 37472 13707 37474 13733
rect 37446 13706 37474 13707
rect 37498 13733 37526 13734
rect 37498 13707 37508 13733
rect 37508 13707 37526 13733
rect 37498 13706 37526 13707
rect 37082 12949 37110 12950
rect 37082 12923 37100 12949
rect 37100 12923 37110 12949
rect 37082 12922 37110 12923
rect 37134 12949 37162 12950
rect 37134 12923 37136 12949
rect 37136 12923 37162 12949
rect 37134 12922 37162 12923
rect 37186 12949 37214 12950
rect 37238 12949 37266 12950
rect 37186 12923 37198 12949
rect 37198 12923 37214 12949
rect 37238 12923 37260 12949
rect 37260 12923 37266 12949
rect 37186 12922 37214 12923
rect 37238 12922 37266 12923
rect 37290 12922 37318 12950
rect 37342 12949 37370 12950
rect 37394 12949 37422 12950
rect 37342 12923 37348 12949
rect 37348 12923 37370 12949
rect 37394 12923 37410 12949
rect 37410 12923 37422 12949
rect 37342 12922 37370 12923
rect 37394 12922 37422 12923
rect 37446 12949 37474 12950
rect 37446 12923 37472 12949
rect 37472 12923 37474 12949
rect 37446 12922 37474 12923
rect 37498 12949 37526 12950
rect 37498 12923 37508 12949
rect 37508 12923 37526 12949
rect 37498 12922 37526 12923
rect 37082 12165 37110 12166
rect 37082 12139 37100 12165
rect 37100 12139 37110 12165
rect 37082 12138 37110 12139
rect 37134 12165 37162 12166
rect 37134 12139 37136 12165
rect 37136 12139 37162 12165
rect 37134 12138 37162 12139
rect 37186 12165 37214 12166
rect 37238 12165 37266 12166
rect 37186 12139 37198 12165
rect 37198 12139 37214 12165
rect 37238 12139 37260 12165
rect 37260 12139 37266 12165
rect 37186 12138 37214 12139
rect 37238 12138 37266 12139
rect 37290 12138 37318 12166
rect 37342 12165 37370 12166
rect 37394 12165 37422 12166
rect 37342 12139 37348 12165
rect 37348 12139 37370 12165
rect 37394 12139 37410 12165
rect 37410 12139 37422 12165
rect 37342 12138 37370 12139
rect 37394 12138 37422 12139
rect 37446 12165 37474 12166
rect 37446 12139 37472 12165
rect 37472 12139 37474 12165
rect 37446 12138 37474 12139
rect 37498 12165 37526 12166
rect 37498 12139 37508 12165
rect 37508 12139 37526 12165
rect 37498 12138 37526 12139
rect 37082 11381 37110 11382
rect 37082 11355 37100 11381
rect 37100 11355 37110 11381
rect 37082 11354 37110 11355
rect 37134 11381 37162 11382
rect 37134 11355 37136 11381
rect 37136 11355 37162 11381
rect 37134 11354 37162 11355
rect 37186 11381 37214 11382
rect 37238 11381 37266 11382
rect 37186 11355 37198 11381
rect 37198 11355 37214 11381
rect 37238 11355 37260 11381
rect 37260 11355 37266 11381
rect 37186 11354 37214 11355
rect 37238 11354 37266 11355
rect 37290 11354 37318 11382
rect 37342 11381 37370 11382
rect 37394 11381 37422 11382
rect 37342 11355 37348 11381
rect 37348 11355 37370 11381
rect 37394 11355 37410 11381
rect 37410 11355 37422 11381
rect 37342 11354 37370 11355
rect 37394 11354 37422 11355
rect 37446 11381 37474 11382
rect 37446 11355 37472 11381
rect 37472 11355 37474 11381
rect 37446 11354 37474 11355
rect 37498 11381 37526 11382
rect 37498 11355 37508 11381
rect 37508 11355 37526 11381
rect 37498 11354 37526 11355
rect 33894 11102 33922 11130
rect 32082 10597 32110 10598
rect 32082 10571 32100 10597
rect 32100 10571 32110 10597
rect 32082 10570 32110 10571
rect 32134 10597 32162 10598
rect 32134 10571 32136 10597
rect 32136 10571 32162 10597
rect 32134 10570 32162 10571
rect 32186 10597 32214 10598
rect 32238 10597 32266 10598
rect 32186 10571 32198 10597
rect 32198 10571 32214 10597
rect 32238 10571 32260 10597
rect 32260 10571 32266 10597
rect 32186 10570 32214 10571
rect 32238 10570 32266 10571
rect 32290 10570 32318 10598
rect 32342 10597 32370 10598
rect 32394 10597 32422 10598
rect 32342 10571 32348 10597
rect 32348 10571 32370 10597
rect 32394 10571 32410 10597
rect 32410 10571 32422 10597
rect 32342 10570 32370 10571
rect 32394 10570 32422 10571
rect 32446 10597 32474 10598
rect 32446 10571 32472 10597
rect 32472 10571 32474 10597
rect 32446 10570 32474 10571
rect 32498 10597 32526 10598
rect 32498 10571 32508 10597
rect 32508 10571 32526 10597
rect 32498 10570 32526 10571
rect 32158 10430 32186 10458
rect 32606 10374 32634 10402
rect 31990 10038 32018 10066
rect 32082 9813 32110 9814
rect 32082 9787 32100 9813
rect 32100 9787 32110 9813
rect 32082 9786 32110 9787
rect 32134 9813 32162 9814
rect 32134 9787 32136 9813
rect 32136 9787 32162 9813
rect 32134 9786 32162 9787
rect 32186 9813 32214 9814
rect 32238 9813 32266 9814
rect 32186 9787 32198 9813
rect 32198 9787 32214 9813
rect 32238 9787 32260 9813
rect 32260 9787 32266 9813
rect 32186 9786 32214 9787
rect 32238 9786 32266 9787
rect 32290 9786 32318 9814
rect 32342 9813 32370 9814
rect 32394 9813 32422 9814
rect 32342 9787 32348 9813
rect 32348 9787 32370 9813
rect 32394 9787 32410 9813
rect 32410 9787 32422 9813
rect 32342 9786 32370 9787
rect 32394 9786 32422 9787
rect 32446 9813 32474 9814
rect 32446 9787 32472 9813
rect 32472 9787 32474 9813
rect 32446 9786 32474 9787
rect 32498 9813 32526 9814
rect 32498 9787 32508 9813
rect 32508 9787 32526 9813
rect 32498 9786 32526 9787
rect 31990 9702 32018 9730
rect 32438 9198 32466 9226
rect 32774 9142 32802 9170
rect 32830 9617 32858 9618
rect 32830 9591 32831 9617
rect 32831 9591 32857 9617
rect 32857 9591 32858 9617
rect 32830 9590 32858 9591
rect 32082 9029 32110 9030
rect 32082 9003 32100 9029
rect 32100 9003 32110 9029
rect 32082 9002 32110 9003
rect 32134 9029 32162 9030
rect 32134 9003 32136 9029
rect 32136 9003 32162 9029
rect 32134 9002 32162 9003
rect 32186 9029 32214 9030
rect 32238 9029 32266 9030
rect 32186 9003 32198 9029
rect 32198 9003 32214 9029
rect 32238 9003 32260 9029
rect 32260 9003 32266 9029
rect 32186 9002 32214 9003
rect 32238 9002 32266 9003
rect 32290 9002 32318 9030
rect 32342 9029 32370 9030
rect 32394 9029 32422 9030
rect 32342 9003 32348 9029
rect 32348 9003 32370 9029
rect 32394 9003 32410 9029
rect 32410 9003 32422 9029
rect 32342 9002 32370 9003
rect 32394 9002 32422 9003
rect 32446 9029 32474 9030
rect 32446 9003 32472 9029
rect 32472 9003 32474 9029
rect 32446 9002 32474 9003
rect 32498 9029 32526 9030
rect 32498 9003 32508 9029
rect 32508 9003 32526 9029
rect 32498 9002 32526 9003
rect 31374 8358 31402 8386
rect 31878 8358 31906 8386
rect 32942 9225 32970 9226
rect 32942 9199 32943 9225
rect 32943 9199 32969 9225
rect 32969 9199 32970 9225
rect 32942 9198 32970 9199
rect 32158 8414 32186 8442
rect 32214 8526 32242 8554
rect 31878 8022 31906 8050
rect 29582 7069 29610 7070
rect 29582 7043 29600 7069
rect 29600 7043 29610 7069
rect 29582 7042 29610 7043
rect 29634 7069 29662 7070
rect 29634 7043 29636 7069
rect 29636 7043 29662 7069
rect 29634 7042 29662 7043
rect 29686 7069 29714 7070
rect 29738 7069 29766 7070
rect 29686 7043 29698 7069
rect 29698 7043 29714 7069
rect 29738 7043 29760 7069
rect 29760 7043 29766 7069
rect 29686 7042 29714 7043
rect 29738 7042 29766 7043
rect 29790 7042 29818 7070
rect 29842 7069 29870 7070
rect 29894 7069 29922 7070
rect 29842 7043 29848 7069
rect 29848 7043 29870 7069
rect 29894 7043 29910 7069
rect 29910 7043 29922 7069
rect 29842 7042 29870 7043
rect 29894 7042 29922 7043
rect 29946 7069 29974 7070
rect 29946 7043 29972 7069
rect 29972 7043 29974 7069
rect 29946 7042 29974 7043
rect 29998 7069 30026 7070
rect 29998 7043 30008 7069
rect 30008 7043 30026 7069
rect 29998 7042 30026 7043
rect 29470 6846 29498 6874
rect 30646 6873 30674 6874
rect 30646 6847 30647 6873
rect 30647 6847 30673 6873
rect 30673 6847 30674 6873
rect 30646 6846 30674 6847
rect 30478 6790 30506 6818
rect 30926 6790 30954 6818
rect 29414 6734 29442 6762
rect 30310 6734 30338 6762
rect 29582 6285 29610 6286
rect 29582 6259 29600 6285
rect 29600 6259 29610 6285
rect 29582 6258 29610 6259
rect 29634 6285 29662 6286
rect 29634 6259 29636 6285
rect 29636 6259 29662 6285
rect 29634 6258 29662 6259
rect 29686 6285 29714 6286
rect 29738 6285 29766 6286
rect 29686 6259 29698 6285
rect 29698 6259 29714 6285
rect 29738 6259 29760 6285
rect 29760 6259 29766 6285
rect 29686 6258 29714 6259
rect 29738 6258 29766 6259
rect 29790 6258 29818 6286
rect 29842 6285 29870 6286
rect 29894 6285 29922 6286
rect 29842 6259 29848 6285
rect 29848 6259 29870 6285
rect 29894 6259 29910 6285
rect 29910 6259 29922 6285
rect 29842 6258 29870 6259
rect 29894 6258 29922 6259
rect 29946 6285 29974 6286
rect 29946 6259 29972 6285
rect 29972 6259 29974 6285
rect 29946 6258 29974 6259
rect 29998 6285 30026 6286
rect 29998 6259 30008 6285
rect 30008 6259 30026 6285
rect 29998 6258 30026 6259
rect 30086 6174 30114 6202
rect 29470 6118 29498 6146
rect 28742 5838 28770 5866
rect 29918 6145 29946 6146
rect 29918 6119 29919 6145
rect 29919 6119 29945 6145
rect 29945 6119 29946 6145
rect 29918 6118 29946 6119
rect 30142 5782 30170 5810
rect 29582 5501 29610 5502
rect 29582 5475 29600 5501
rect 29600 5475 29610 5501
rect 29582 5474 29610 5475
rect 29634 5501 29662 5502
rect 29634 5475 29636 5501
rect 29636 5475 29662 5501
rect 29634 5474 29662 5475
rect 29686 5501 29714 5502
rect 29738 5501 29766 5502
rect 29686 5475 29698 5501
rect 29698 5475 29714 5501
rect 29738 5475 29760 5501
rect 29760 5475 29766 5501
rect 29686 5474 29714 5475
rect 29738 5474 29766 5475
rect 29790 5474 29818 5502
rect 29842 5501 29870 5502
rect 29894 5501 29922 5502
rect 29842 5475 29848 5501
rect 29848 5475 29870 5501
rect 29894 5475 29910 5501
rect 29910 5475 29922 5501
rect 29842 5474 29870 5475
rect 29894 5474 29922 5475
rect 29946 5501 29974 5502
rect 29946 5475 29972 5501
rect 29972 5475 29974 5501
rect 29946 5474 29974 5475
rect 29998 5501 30026 5502
rect 29998 5475 30008 5501
rect 30008 5475 30026 5501
rect 29998 5474 30026 5475
rect 30142 5278 30170 5306
rect 29582 4717 29610 4718
rect 29582 4691 29600 4717
rect 29600 4691 29610 4717
rect 29582 4690 29610 4691
rect 29634 4717 29662 4718
rect 29634 4691 29636 4717
rect 29636 4691 29662 4717
rect 29634 4690 29662 4691
rect 29686 4717 29714 4718
rect 29738 4717 29766 4718
rect 29686 4691 29698 4717
rect 29698 4691 29714 4717
rect 29738 4691 29760 4717
rect 29760 4691 29766 4717
rect 29686 4690 29714 4691
rect 29738 4690 29766 4691
rect 29790 4690 29818 4718
rect 29842 4717 29870 4718
rect 29894 4717 29922 4718
rect 29842 4691 29848 4717
rect 29848 4691 29870 4717
rect 29894 4691 29910 4717
rect 29910 4691 29922 4717
rect 29842 4690 29870 4691
rect 29894 4690 29922 4691
rect 29946 4717 29974 4718
rect 29946 4691 29972 4717
rect 29972 4691 29974 4717
rect 29946 4690 29974 4691
rect 29998 4717 30026 4718
rect 29998 4691 30008 4717
rect 30008 4691 30026 4717
rect 29998 4690 30026 4691
rect 28630 3038 28658 3066
rect 30030 3990 30058 4018
rect 29582 3933 29610 3934
rect 29582 3907 29600 3933
rect 29600 3907 29610 3933
rect 29582 3906 29610 3907
rect 29634 3933 29662 3934
rect 29634 3907 29636 3933
rect 29636 3907 29662 3933
rect 29634 3906 29662 3907
rect 29686 3933 29714 3934
rect 29738 3933 29766 3934
rect 29686 3907 29698 3933
rect 29698 3907 29714 3933
rect 29738 3907 29760 3933
rect 29760 3907 29766 3933
rect 29686 3906 29714 3907
rect 29738 3906 29766 3907
rect 29790 3906 29818 3934
rect 29842 3933 29870 3934
rect 29894 3933 29922 3934
rect 29842 3907 29848 3933
rect 29848 3907 29870 3933
rect 29894 3907 29910 3933
rect 29910 3907 29922 3933
rect 29842 3906 29870 3907
rect 29894 3906 29922 3907
rect 29946 3933 29974 3934
rect 29946 3907 29972 3933
rect 29972 3907 29974 3933
rect 29946 3906 29974 3907
rect 29998 3933 30026 3934
rect 29998 3907 30008 3933
rect 30008 3907 30026 3933
rect 29998 3906 30026 3907
rect 30030 3822 30058 3850
rect 29470 3710 29498 3738
rect 29358 3374 29386 3402
rect 29918 3737 29946 3738
rect 29918 3711 29919 3737
rect 29919 3711 29945 3737
rect 29945 3711 29946 3737
rect 29918 3710 29946 3711
rect 28686 2646 28714 2674
rect 28462 2561 28490 2562
rect 28462 2535 28463 2561
rect 28463 2535 28489 2561
rect 28489 2535 28490 2561
rect 28462 2534 28490 2535
rect 28630 2534 28658 2562
rect 27082 1973 27110 1974
rect 27082 1947 27100 1973
rect 27100 1947 27110 1973
rect 27082 1946 27110 1947
rect 27134 1973 27162 1974
rect 27134 1947 27136 1973
rect 27136 1947 27162 1973
rect 27134 1946 27162 1947
rect 27186 1973 27214 1974
rect 27238 1973 27266 1974
rect 27186 1947 27198 1973
rect 27198 1947 27214 1973
rect 27238 1947 27260 1973
rect 27260 1947 27266 1973
rect 27186 1946 27214 1947
rect 27238 1946 27266 1947
rect 27290 1946 27318 1974
rect 27342 1973 27370 1974
rect 27394 1973 27422 1974
rect 27342 1947 27348 1973
rect 27348 1947 27370 1973
rect 27394 1947 27410 1973
rect 27410 1947 27422 1973
rect 27342 1946 27370 1947
rect 27394 1946 27422 1947
rect 27446 1973 27474 1974
rect 27446 1947 27472 1973
rect 27472 1947 27474 1973
rect 27446 1946 27474 1947
rect 27498 1973 27526 1974
rect 27498 1947 27508 1973
rect 27508 1947 27526 1973
rect 27498 1946 27526 1947
rect 30198 4913 30226 4914
rect 30198 4887 30199 4913
rect 30199 4887 30225 4913
rect 30225 4887 30226 4913
rect 30198 4886 30226 4887
rect 30086 3766 30114 3794
rect 30254 5278 30282 5306
rect 30310 4913 30338 4914
rect 30310 4887 30311 4913
rect 30311 4887 30337 4913
rect 30337 4887 30338 4913
rect 30310 4886 30338 4887
rect 30030 3289 30058 3290
rect 30030 3263 30031 3289
rect 30031 3263 30057 3289
rect 30057 3263 30058 3289
rect 30030 3262 30058 3263
rect 29582 3149 29610 3150
rect 29582 3123 29600 3149
rect 29600 3123 29610 3149
rect 29582 3122 29610 3123
rect 29634 3149 29662 3150
rect 29634 3123 29636 3149
rect 29636 3123 29662 3149
rect 29634 3122 29662 3123
rect 29686 3149 29714 3150
rect 29738 3149 29766 3150
rect 29686 3123 29698 3149
rect 29698 3123 29714 3149
rect 29738 3123 29760 3149
rect 29760 3123 29766 3149
rect 29686 3122 29714 3123
rect 29738 3122 29766 3123
rect 29790 3122 29818 3150
rect 29842 3149 29870 3150
rect 29894 3149 29922 3150
rect 29842 3123 29848 3149
rect 29848 3123 29870 3149
rect 29894 3123 29910 3149
rect 29910 3123 29922 3149
rect 29842 3122 29870 3123
rect 29894 3122 29922 3123
rect 29946 3149 29974 3150
rect 29946 3123 29972 3149
rect 29972 3123 29974 3149
rect 29946 3122 29974 3123
rect 29998 3149 30026 3150
rect 29998 3123 30008 3149
rect 30008 3123 30026 3149
rect 29998 3122 30026 3123
rect 29022 2534 29050 2562
rect 30310 2982 30338 3010
rect 30366 2534 30394 2562
rect 30030 2478 30058 2506
rect 29582 2365 29610 2366
rect 29582 2339 29600 2365
rect 29600 2339 29610 2365
rect 29582 2338 29610 2339
rect 29634 2365 29662 2366
rect 29634 2339 29636 2365
rect 29636 2339 29662 2365
rect 29634 2338 29662 2339
rect 29686 2365 29714 2366
rect 29738 2365 29766 2366
rect 29686 2339 29698 2365
rect 29698 2339 29714 2365
rect 29738 2339 29760 2365
rect 29760 2339 29766 2365
rect 29686 2338 29714 2339
rect 29738 2338 29766 2339
rect 29790 2338 29818 2366
rect 29842 2365 29870 2366
rect 29894 2365 29922 2366
rect 29842 2339 29848 2365
rect 29848 2339 29870 2365
rect 29894 2339 29910 2365
rect 29910 2339 29922 2365
rect 29842 2338 29870 2339
rect 29894 2338 29922 2339
rect 29946 2365 29974 2366
rect 29946 2339 29972 2365
rect 29972 2339 29974 2365
rect 29946 2338 29974 2339
rect 29998 2365 30026 2366
rect 29998 2339 30008 2365
rect 30008 2339 30026 2365
rect 29998 2338 30026 2339
rect 29414 2198 29442 2226
rect 28798 1638 28826 1666
rect 30254 2142 30282 2170
rect 31374 6790 31402 6818
rect 30982 6454 31010 6482
rect 30926 5670 30954 5698
rect 31374 6145 31402 6146
rect 31374 6119 31375 6145
rect 31375 6119 31401 6145
rect 31401 6119 31402 6145
rect 31374 6118 31402 6119
rect 31878 6790 31906 6818
rect 32082 8245 32110 8246
rect 32082 8219 32100 8245
rect 32100 8219 32110 8245
rect 32082 8218 32110 8219
rect 32134 8245 32162 8246
rect 32134 8219 32136 8245
rect 32136 8219 32162 8245
rect 32134 8218 32162 8219
rect 32186 8245 32214 8246
rect 32238 8245 32266 8246
rect 32186 8219 32198 8245
rect 32198 8219 32214 8245
rect 32238 8219 32260 8245
rect 32260 8219 32266 8245
rect 32186 8218 32214 8219
rect 32238 8218 32266 8219
rect 32290 8218 32318 8246
rect 32342 8245 32370 8246
rect 32394 8245 32422 8246
rect 32342 8219 32348 8245
rect 32348 8219 32370 8245
rect 32394 8219 32410 8245
rect 32410 8219 32422 8245
rect 32342 8218 32370 8219
rect 32394 8218 32422 8219
rect 32446 8245 32474 8246
rect 32446 8219 32472 8245
rect 32472 8219 32474 8245
rect 32446 8218 32474 8219
rect 32498 8245 32526 8246
rect 32498 8219 32508 8245
rect 32508 8219 32526 8245
rect 32498 8218 32526 8219
rect 32438 8134 32466 8162
rect 32158 7657 32186 7658
rect 32158 7631 32159 7657
rect 32159 7631 32185 7657
rect 32185 7631 32186 7657
rect 32158 7630 32186 7631
rect 32326 7657 32354 7658
rect 32326 7631 32327 7657
rect 32327 7631 32353 7657
rect 32353 7631 32354 7657
rect 32326 7630 32354 7631
rect 32438 7630 32466 7658
rect 35294 11102 35322 11130
rect 35854 11102 35882 11130
rect 36134 11158 36162 11186
rect 34582 10989 34610 10990
rect 34582 10963 34600 10989
rect 34600 10963 34610 10989
rect 34582 10962 34610 10963
rect 34634 10989 34662 10990
rect 34634 10963 34636 10989
rect 34636 10963 34662 10989
rect 34634 10962 34662 10963
rect 34686 10989 34714 10990
rect 34738 10989 34766 10990
rect 34686 10963 34698 10989
rect 34698 10963 34714 10989
rect 34738 10963 34760 10989
rect 34760 10963 34766 10989
rect 34686 10962 34714 10963
rect 34738 10962 34766 10963
rect 34790 10962 34818 10990
rect 34842 10989 34870 10990
rect 34894 10989 34922 10990
rect 34842 10963 34848 10989
rect 34848 10963 34870 10989
rect 34894 10963 34910 10989
rect 34910 10963 34922 10989
rect 34842 10962 34870 10963
rect 34894 10962 34922 10963
rect 34946 10989 34974 10990
rect 34946 10963 34972 10989
rect 34972 10963 34974 10989
rect 34946 10962 34974 10963
rect 34998 10989 35026 10990
rect 34998 10963 35008 10989
rect 35008 10963 35026 10989
rect 34998 10962 35026 10963
rect 33894 10793 33922 10794
rect 33894 10767 33895 10793
rect 33895 10767 33921 10793
rect 33921 10767 33922 10793
rect 33894 10766 33922 10767
rect 35350 10793 35378 10794
rect 35350 10767 35351 10793
rect 35351 10767 35377 10793
rect 35377 10767 35378 10793
rect 35350 10766 35378 10767
rect 34582 10205 34610 10206
rect 34582 10179 34600 10205
rect 34600 10179 34610 10205
rect 34582 10178 34610 10179
rect 34634 10205 34662 10206
rect 34634 10179 34636 10205
rect 34636 10179 34662 10205
rect 34634 10178 34662 10179
rect 34686 10205 34714 10206
rect 34738 10205 34766 10206
rect 34686 10179 34698 10205
rect 34698 10179 34714 10205
rect 34738 10179 34760 10205
rect 34760 10179 34766 10205
rect 34686 10178 34714 10179
rect 34738 10178 34766 10179
rect 34790 10178 34818 10206
rect 34842 10205 34870 10206
rect 34894 10205 34922 10206
rect 34842 10179 34848 10205
rect 34848 10179 34870 10205
rect 34894 10179 34910 10205
rect 34910 10179 34922 10205
rect 34842 10178 34870 10179
rect 34894 10178 34922 10179
rect 34946 10205 34974 10206
rect 34946 10179 34972 10205
rect 34972 10179 34974 10205
rect 34946 10178 34974 10179
rect 34998 10205 35026 10206
rect 34998 10179 35008 10205
rect 35008 10179 35026 10205
rect 34998 10178 35026 10179
rect 33110 9590 33138 9618
rect 34230 10038 34258 10066
rect 33390 9254 33418 9282
rect 32998 8750 33026 8778
rect 32942 8414 32970 8442
rect 33334 8049 33362 8050
rect 33334 8023 33335 8049
rect 33335 8023 33361 8049
rect 33361 8023 33362 8049
rect 33334 8022 33362 8023
rect 33334 7686 33362 7714
rect 32102 7518 32130 7546
rect 32082 7461 32110 7462
rect 32082 7435 32100 7461
rect 32100 7435 32110 7461
rect 32082 7434 32110 7435
rect 32134 7461 32162 7462
rect 32134 7435 32136 7461
rect 32136 7435 32162 7461
rect 32134 7434 32162 7435
rect 32186 7461 32214 7462
rect 32238 7461 32266 7462
rect 32186 7435 32198 7461
rect 32198 7435 32214 7461
rect 32238 7435 32260 7461
rect 32260 7435 32266 7461
rect 32186 7434 32214 7435
rect 32238 7434 32266 7435
rect 32290 7434 32318 7462
rect 32342 7461 32370 7462
rect 32394 7461 32422 7462
rect 32342 7435 32348 7461
rect 32348 7435 32370 7461
rect 32394 7435 32410 7461
rect 32410 7435 32422 7461
rect 32342 7434 32370 7435
rect 32394 7434 32422 7435
rect 32446 7461 32474 7462
rect 32446 7435 32472 7461
rect 32472 7435 32474 7461
rect 32446 7434 32474 7435
rect 32498 7461 32526 7462
rect 32498 7435 32508 7461
rect 32508 7435 32526 7461
rect 32498 7434 32526 7435
rect 32606 7462 32634 7490
rect 32438 7265 32466 7266
rect 32438 7239 32439 7265
rect 32439 7239 32465 7265
rect 32465 7239 32466 7265
rect 32438 7238 32466 7239
rect 32158 6734 32186 6762
rect 32438 6734 32466 6762
rect 32082 6677 32110 6678
rect 32082 6651 32100 6677
rect 32100 6651 32110 6677
rect 32082 6650 32110 6651
rect 32134 6677 32162 6678
rect 32134 6651 32136 6677
rect 32136 6651 32162 6677
rect 32134 6650 32162 6651
rect 32186 6677 32214 6678
rect 32238 6677 32266 6678
rect 32186 6651 32198 6677
rect 32198 6651 32214 6677
rect 32238 6651 32260 6677
rect 32260 6651 32266 6677
rect 32186 6650 32214 6651
rect 32238 6650 32266 6651
rect 32290 6650 32318 6678
rect 32342 6677 32370 6678
rect 32394 6677 32422 6678
rect 32342 6651 32348 6677
rect 32348 6651 32370 6677
rect 32394 6651 32410 6677
rect 32410 6651 32422 6677
rect 32342 6650 32370 6651
rect 32394 6650 32422 6651
rect 32446 6677 32474 6678
rect 32446 6651 32472 6677
rect 32472 6651 32474 6677
rect 32446 6650 32474 6651
rect 32498 6677 32526 6678
rect 32498 6651 32508 6677
rect 32508 6651 32526 6677
rect 32498 6650 32526 6651
rect 32158 6481 32186 6482
rect 32158 6455 32159 6481
rect 32159 6455 32185 6481
rect 32185 6455 32186 6481
rect 32158 6454 32186 6455
rect 31990 6174 32018 6202
rect 31934 5782 31962 5810
rect 31318 4102 31346 4130
rect 31318 3737 31346 3738
rect 31318 3711 31319 3737
rect 31319 3711 31345 3737
rect 31345 3711 31346 3737
rect 31318 3710 31346 3711
rect 30702 3345 30730 3346
rect 30702 3319 30703 3345
rect 30703 3319 30729 3345
rect 30729 3319 30730 3345
rect 30702 3318 30730 3319
rect 31878 3374 31906 3402
rect 31934 5278 31962 5306
rect 30702 2561 30730 2562
rect 30702 2535 30703 2561
rect 30703 2535 30729 2561
rect 30729 2535 30730 2561
rect 30702 2534 30730 2535
rect 31262 2225 31290 2226
rect 31262 2199 31263 2225
rect 31263 2199 31289 2225
rect 31289 2199 31290 2225
rect 31262 2198 31290 2199
rect 29022 1638 29050 1666
rect 29582 1581 29610 1582
rect 29582 1555 29600 1581
rect 29600 1555 29610 1581
rect 29582 1554 29610 1555
rect 29634 1581 29662 1582
rect 29634 1555 29636 1581
rect 29636 1555 29662 1581
rect 29634 1554 29662 1555
rect 29686 1581 29714 1582
rect 29738 1581 29766 1582
rect 29686 1555 29698 1581
rect 29698 1555 29714 1581
rect 29738 1555 29760 1581
rect 29760 1555 29766 1581
rect 29686 1554 29714 1555
rect 29738 1554 29766 1555
rect 29790 1554 29818 1582
rect 29842 1581 29870 1582
rect 29894 1581 29922 1582
rect 29842 1555 29848 1581
rect 29848 1555 29870 1581
rect 29894 1555 29910 1581
rect 29910 1555 29922 1581
rect 29842 1554 29870 1555
rect 29894 1554 29922 1555
rect 29946 1581 29974 1582
rect 29946 1555 29972 1581
rect 29972 1555 29974 1581
rect 29946 1554 29974 1555
rect 29998 1581 30026 1582
rect 29998 1555 30008 1581
rect 30008 1555 30026 1581
rect 29998 1554 30026 1555
rect 31598 2422 31626 2450
rect 32158 6089 32186 6090
rect 32158 6063 32159 6089
rect 32159 6063 32185 6089
rect 32185 6063 32186 6089
rect 32158 6062 32186 6063
rect 32326 6089 32354 6090
rect 32326 6063 32327 6089
rect 32327 6063 32353 6089
rect 32353 6063 32354 6089
rect 32326 6062 32354 6063
rect 32082 5893 32110 5894
rect 32082 5867 32100 5893
rect 32100 5867 32110 5893
rect 32082 5866 32110 5867
rect 32134 5893 32162 5894
rect 32134 5867 32136 5893
rect 32136 5867 32162 5893
rect 32134 5866 32162 5867
rect 32186 5893 32214 5894
rect 32238 5893 32266 5894
rect 32186 5867 32198 5893
rect 32198 5867 32214 5893
rect 32238 5867 32260 5893
rect 32260 5867 32266 5893
rect 32186 5866 32214 5867
rect 32238 5866 32266 5867
rect 32290 5866 32318 5894
rect 32342 5893 32370 5894
rect 32394 5893 32422 5894
rect 32342 5867 32348 5893
rect 32348 5867 32370 5893
rect 32394 5867 32410 5893
rect 32410 5867 32422 5893
rect 32342 5866 32370 5867
rect 32394 5866 32422 5867
rect 32446 5893 32474 5894
rect 32446 5867 32472 5893
rect 32472 5867 32474 5893
rect 32446 5866 32474 5867
rect 32498 5893 32526 5894
rect 32498 5867 32508 5893
rect 32508 5867 32526 5893
rect 32498 5866 32526 5867
rect 32158 5697 32186 5698
rect 32158 5671 32159 5697
rect 32159 5671 32185 5697
rect 32185 5671 32186 5697
rect 32158 5670 32186 5671
rect 32158 5305 32186 5306
rect 32158 5279 32159 5305
rect 32159 5279 32185 5305
rect 32185 5279 32186 5305
rect 32158 5278 32186 5279
rect 32326 5305 32354 5306
rect 32326 5279 32327 5305
rect 32327 5279 32353 5305
rect 32353 5279 32354 5305
rect 32326 5278 32354 5279
rect 32082 5109 32110 5110
rect 32082 5083 32100 5109
rect 32100 5083 32110 5109
rect 32082 5082 32110 5083
rect 32134 5109 32162 5110
rect 32134 5083 32136 5109
rect 32136 5083 32162 5109
rect 32134 5082 32162 5083
rect 32186 5109 32214 5110
rect 32238 5109 32266 5110
rect 32186 5083 32198 5109
rect 32198 5083 32214 5109
rect 32238 5083 32260 5109
rect 32260 5083 32266 5109
rect 32186 5082 32214 5083
rect 32238 5082 32266 5083
rect 32290 5082 32318 5110
rect 32342 5109 32370 5110
rect 32394 5109 32422 5110
rect 32342 5083 32348 5109
rect 32348 5083 32370 5109
rect 32394 5083 32410 5109
rect 32410 5083 32422 5109
rect 32342 5082 32370 5083
rect 32394 5082 32422 5083
rect 32446 5109 32474 5110
rect 32446 5083 32472 5109
rect 32472 5083 32474 5109
rect 32446 5082 32474 5083
rect 32498 5109 32526 5110
rect 32498 5083 32508 5109
rect 32508 5083 32526 5109
rect 32498 5082 32526 5083
rect 32158 4913 32186 4914
rect 32158 4887 32159 4913
rect 32159 4887 32185 4913
rect 32185 4887 32186 4913
rect 32158 4886 32186 4887
rect 32886 7518 32914 7546
rect 32942 7657 32970 7658
rect 32942 7631 32943 7657
rect 32943 7631 32969 7657
rect 32969 7631 32970 7657
rect 32942 7630 32970 7631
rect 32774 7126 32802 7154
rect 32886 7238 32914 7266
rect 32718 6454 32746 6482
rect 32886 6342 32914 6370
rect 32606 4662 32634 4690
rect 32662 5670 32690 5698
rect 32774 5305 32802 5306
rect 32774 5279 32775 5305
rect 32775 5279 32801 5305
rect 32801 5279 32802 5305
rect 32774 5278 32802 5279
rect 33726 7574 33754 7602
rect 33670 7462 33698 7490
rect 33726 7182 33754 7210
rect 34454 9590 34482 9618
rect 34958 9617 34986 9618
rect 34958 9591 34959 9617
rect 34959 9591 34985 9617
rect 34985 9591 34986 9617
rect 34958 9590 34986 9591
rect 35350 9534 35378 9562
rect 34582 9421 34610 9422
rect 34582 9395 34600 9421
rect 34600 9395 34610 9421
rect 34582 9394 34610 9395
rect 34634 9421 34662 9422
rect 34634 9395 34636 9421
rect 34636 9395 34662 9421
rect 34634 9394 34662 9395
rect 34686 9421 34714 9422
rect 34738 9421 34766 9422
rect 34686 9395 34698 9421
rect 34698 9395 34714 9421
rect 34738 9395 34760 9421
rect 34760 9395 34766 9421
rect 34686 9394 34714 9395
rect 34738 9394 34766 9395
rect 34790 9394 34818 9422
rect 34842 9421 34870 9422
rect 34894 9421 34922 9422
rect 34842 9395 34848 9421
rect 34848 9395 34870 9421
rect 34894 9395 34910 9421
rect 34910 9395 34922 9421
rect 34842 9394 34870 9395
rect 34894 9394 34922 9395
rect 34946 9421 34974 9422
rect 34946 9395 34972 9421
rect 34972 9395 34974 9421
rect 34946 9394 34974 9395
rect 34998 9421 35026 9422
rect 34998 9395 35008 9421
rect 35008 9395 35026 9421
rect 34998 9394 35026 9395
rect 34622 9254 34650 9282
rect 34174 9225 34202 9226
rect 34174 9199 34175 9225
rect 34175 9199 34201 9225
rect 34201 9199 34202 9225
rect 34174 9198 34202 9199
rect 34846 9254 34874 9282
rect 35070 9254 35098 9282
rect 34958 8833 34986 8834
rect 34958 8807 34959 8833
rect 34959 8807 34985 8833
rect 34985 8807 34986 8833
rect 34958 8806 34986 8807
rect 34582 8637 34610 8638
rect 34582 8611 34600 8637
rect 34600 8611 34610 8637
rect 34582 8610 34610 8611
rect 34634 8637 34662 8638
rect 34634 8611 34636 8637
rect 34636 8611 34662 8637
rect 34634 8610 34662 8611
rect 34686 8637 34714 8638
rect 34738 8637 34766 8638
rect 34686 8611 34698 8637
rect 34698 8611 34714 8637
rect 34738 8611 34760 8637
rect 34760 8611 34766 8637
rect 34686 8610 34714 8611
rect 34738 8610 34766 8611
rect 34790 8610 34818 8638
rect 34842 8637 34870 8638
rect 34894 8637 34922 8638
rect 34842 8611 34848 8637
rect 34848 8611 34870 8637
rect 34894 8611 34910 8637
rect 34910 8611 34922 8637
rect 34842 8610 34870 8611
rect 34894 8610 34922 8611
rect 34946 8637 34974 8638
rect 34946 8611 34972 8637
rect 34972 8611 34974 8637
rect 34946 8610 34974 8611
rect 34998 8637 35026 8638
rect 34998 8611 35008 8637
rect 35008 8611 35026 8637
rect 34998 8610 35026 8611
rect 33894 8497 33922 8498
rect 33894 8471 33895 8497
rect 33895 8471 33921 8497
rect 33921 8471 33922 8497
rect 33894 8470 33922 8471
rect 36078 10374 36106 10402
rect 35854 9561 35882 9562
rect 35854 9535 35855 9561
rect 35855 9535 35881 9561
rect 35881 9535 35882 9561
rect 35854 9534 35882 9535
rect 35630 9198 35658 9226
rect 35854 9198 35882 9226
rect 35238 9086 35266 9114
rect 33838 7713 33866 7714
rect 33838 7687 33839 7713
rect 33839 7687 33865 7713
rect 33865 7687 33866 7713
rect 33838 7686 33866 7687
rect 33670 7126 33698 7154
rect 33334 6790 33362 6818
rect 32998 6734 33026 6762
rect 33670 6678 33698 6706
rect 33614 6174 33642 6202
rect 33278 5838 33306 5866
rect 33334 5894 33362 5922
rect 32942 4942 32970 4970
rect 33054 5782 33082 5810
rect 32082 4325 32110 4326
rect 32082 4299 32100 4325
rect 32100 4299 32110 4325
rect 32082 4298 32110 4299
rect 32134 4325 32162 4326
rect 32134 4299 32136 4325
rect 32136 4299 32162 4325
rect 32134 4298 32162 4299
rect 32186 4325 32214 4326
rect 32238 4325 32266 4326
rect 32186 4299 32198 4325
rect 32198 4299 32214 4325
rect 32238 4299 32260 4325
rect 32260 4299 32266 4325
rect 32186 4298 32214 4299
rect 32238 4298 32266 4299
rect 32290 4298 32318 4326
rect 32342 4325 32370 4326
rect 32394 4325 32422 4326
rect 32342 4299 32348 4325
rect 32348 4299 32370 4325
rect 32394 4299 32410 4325
rect 32410 4299 32422 4325
rect 32342 4298 32370 4299
rect 32394 4298 32422 4299
rect 32446 4325 32474 4326
rect 32446 4299 32472 4325
rect 32472 4299 32474 4325
rect 32446 4298 32474 4299
rect 32498 4325 32526 4326
rect 32498 4299 32508 4325
rect 32508 4299 32526 4325
rect 32498 4298 32526 4299
rect 32158 4046 32186 4074
rect 32082 3541 32110 3542
rect 32082 3515 32100 3541
rect 32100 3515 32110 3541
rect 32082 3514 32110 3515
rect 32134 3541 32162 3542
rect 32134 3515 32136 3541
rect 32136 3515 32162 3541
rect 32134 3514 32162 3515
rect 32186 3541 32214 3542
rect 32238 3541 32266 3542
rect 32186 3515 32198 3541
rect 32198 3515 32214 3541
rect 32238 3515 32260 3541
rect 32260 3515 32266 3541
rect 32186 3514 32214 3515
rect 32238 3514 32266 3515
rect 32290 3514 32318 3542
rect 32342 3541 32370 3542
rect 32394 3541 32422 3542
rect 32342 3515 32348 3541
rect 32348 3515 32370 3541
rect 32394 3515 32410 3541
rect 32410 3515 32422 3541
rect 32342 3514 32370 3515
rect 32394 3514 32422 3515
rect 32446 3541 32474 3542
rect 32446 3515 32472 3541
rect 32472 3515 32474 3541
rect 32446 3514 32474 3515
rect 32498 3541 32526 3542
rect 32498 3515 32508 3541
rect 32508 3515 32526 3541
rect 32498 3514 32526 3515
rect 32158 3345 32186 3346
rect 32158 3319 32159 3345
rect 32159 3319 32185 3345
rect 32185 3319 32186 3345
rect 32158 3318 32186 3319
rect 31990 3262 32018 3290
rect 32046 3009 32074 3010
rect 32046 2983 32047 3009
rect 32047 2983 32073 3009
rect 32073 2983 32074 3009
rect 32046 2982 32074 2983
rect 32214 2953 32242 2954
rect 32214 2927 32215 2953
rect 32215 2927 32241 2953
rect 32241 2927 32242 2953
rect 32214 2926 32242 2927
rect 32382 2953 32410 2954
rect 32382 2927 32383 2953
rect 32383 2927 32409 2953
rect 32409 2927 32410 2953
rect 32382 2926 32410 2927
rect 32606 2926 32634 2954
rect 32774 3737 32802 3738
rect 32774 3711 32775 3737
rect 32775 3711 32801 3737
rect 32801 3711 32802 3737
rect 32774 3710 32802 3711
rect 32082 2757 32110 2758
rect 32082 2731 32100 2757
rect 32100 2731 32110 2757
rect 32082 2730 32110 2731
rect 32134 2757 32162 2758
rect 32134 2731 32136 2757
rect 32136 2731 32162 2757
rect 32134 2730 32162 2731
rect 32186 2757 32214 2758
rect 32238 2757 32266 2758
rect 32186 2731 32198 2757
rect 32198 2731 32214 2757
rect 32238 2731 32260 2757
rect 32260 2731 32266 2757
rect 32186 2730 32214 2731
rect 32238 2730 32266 2731
rect 32290 2730 32318 2758
rect 32342 2757 32370 2758
rect 32394 2757 32422 2758
rect 32342 2731 32348 2757
rect 32348 2731 32370 2757
rect 32394 2731 32410 2757
rect 32410 2731 32422 2757
rect 32342 2730 32370 2731
rect 32394 2730 32422 2731
rect 32446 2757 32474 2758
rect 32446 2731 32472 2757
rect 32472 2731 32474 2757
rect 32446 2730 32474 2731
rect 32498 2757 32526 2758
rect 32498 2731 32508 2757
rect 32508 2731 32526 2757
rect 32498 2730 32526 2731
rect 32438 2646 32466 2674
rect 31654 2169 31682 2170
rect 31654 2143 31655 2169
rect 31655 2143 31681 2169
rect 31681 2143 31682 2169
rect 31654 2142 31682 2143
rect 32082 1973 32110 1974
rect 32082 1947 32100 1973
rect 32100 1947 32110 1973
rect 32082 1946 32110 1947
rect 32134 1973 32162 1974
rect 32134 1947 32136 1973
rect 32136 1947 32162 1973
rect 32134 1946 32162 1947
rect 32186 1973 32214 1974
rect 32238 1973 32266 1974
rect 32186 1947 32198 1973
rect 32198 1947 32214 1973
rect 32238 1947 32260 1973
rect 32260 1947 32266 1973
rect 32186 1946 32214 1947
rect 32238 1946 32266 1947
rect 32290 1946 32318 1974
rect 32342 1973 32370 1974
rect 32394 1973 32422 1974
rect 32342 1947 32348 1973
rect 32348 1947 32370 1973
rect 32394 1947 32410 1973
rect 32410 1947 32422 1973
rect 32342 1946 32370 1947
rect 32394 1946 32422 1947
rect 32446 1973 32474 1974
rect 32446 1947 32472 1973
rect 32472 1947 32474 1973
rect 32446 1946 32474 1947
rect 32498 1973 32526 1974
rect 32498 1947 32508 1973
rect 32508 1947 32526 1973
rect 32498 1946 32526 1947
rect 31598 1806 31626 1834
rect 33670 5894 33698 5922
rect 33726 6425 33754 6426
rect 33726 6399 33727 6425
rect 33727 6399 33753 6425
rect 33753 6399 33754 6425
rect 33726 6398 33754 6399
rect 33614 5838 33642 5866
rect 33334 5334 33362 5362
rect 33614 5334 33642 5362
rect 33334 3374 33362 3402
rect 33782 5838 33810 5866
rect 33726 5641 33754 5642
rect 33726 5615 33727 5641
rect 33727 5615 33753 5641
rect 33753 5615 33754 5641
rect 33726 5614 33754 5615
rect 34398 8441 34426 8442
rect 34398 8415 34399 8441
rect 34399 8415 34425 8441
rect 34425 8415 34426 8441
rect 34398 8414 34426 8415
rect 34958 8414 34986 8442
rect 35238 8470 35266 8498
rect 34582 7853 34610 7854
rect 34582 7827 34600 7853
rect 34600 7827 34610 7853
rect 34582 7826 34610 7827
rect 34634 7853 34662 7854
rect 34634 7827 34636 7853
rect 34636 7827 34662 7853
rect 34634 7826 34662 7827
rect 34686 7853 34714 7854
rect 34738 7853 34766 7854
rect 34686 7827 34698 7853
rect 34698 7827 34714 7853
rect 34738 7827 34760 7853
rect 34760 7827 34766 7853
rect 34686 7826 34714 7827
rect 34738 7826 34766 7827
rect 34790 7826 34818 7854
rect 34842 7853 34870 7854
rect 34894 7853 34922 7854
rect 34842 7827 34848 7853
rect 34848 7827 34870 7853
rect 34894 7827 34910 7853
rect 34910 7827 34922 7853
rect 34842 7826 34870 7827
rect 34894 7826 34922 7827
rect 34946 7853 34974 7854
rect 34946 7827 34972 7853
rect 34972 7827 34974 7853
rect 34946 7826 34974 7827
rect 34998 7853 35026 7854
rect 34998 7827 35008 7853
rect 35008 7827 35026 7853
rect 34998 7826 35026 7827
rect 33894 7294 33922 7322
rect 33894 7209 33922 7210
rect 33894 7183 33895 7209
rect 33895 7183 33921 7209
rect 33921 7183 33922 7209
rect 33894 7182 33922 7183
rect 33950 6790 33978 6818
rect 33894 6425 33922 6426
rect 33894 6399 33895 6425
rect 33895 6399 33921 6425
rect 33921 6399 33922 6425
rect 33894 6398 33922 6399
rect 33838 5054 33866 5082
rect 33894 5641 33922 5642
rect 33894 5615 33895 5641
rect 33895 5615 33921 5641
rect 33921 5615 33922 5641
rect 33894 5614 33922 5615
rect 33894 5222 33922 5250
rect 34398 7518 34426 7546
rect 34678 7265 34706 7266
rect 34678 7239 34679 7265
rect 34679 7239 34705 7265
rect 34705 7239 34706 7265
rect 34678 7238 34706 7239
rect 34582 7069 34610 7070
rect 34582 7043 34600 7069
rect 34600 7043 34610 7069
rect 34582 7042 34610 7043
rect 34634 7069 34662 7070
rect 34634 7043 34636 7069
rect 34636 7043 34662 7069
rect 34634 7042 34662 7043
rect 34686 7069 34714 7070
rect 34738 7069 34766 7070
rect 34686 7043 34698 7069
rect 34698 7043 34714 7069
rect 34738 7043 34760 7069
rect 34760 7043 34766 7069
rect 34686 7042 34714 7043
rect 34738 7042 34766 7043
rect 34790 7042 34818 7070
rect 34842 7069 34870 7070
rect 34894 7069 34922 7070
rect 34842 7043 34848 7069
rect 34848 7043 34870 7069
rect 34894 7043 34910 7069
rect 34910 7043 34922 7069
rect 34842 7042 34870 7043
rect 34894 7042 34922 7043
rect 34946 7069 34974 7070
rect 34946 7043 34972 7069
rect 34972 7043 34974 7069
rect 34946 7042 34974 7043
rect 34998 7069 35026 7070
rect 34998 7043 35008 7069
rect 35008 7043 35026 7069
rect 34998 7042 35026 7043
rect 34398 6873 34426 6874
rect 34398 6847 34399 6873
rect 34399 6847 34425 6873
rect 34425 6847 34426 6873
rect 34398 6846 34426 6847
rect 34678 6846 34706 6874
rect 34006 6678 34034 6706
rect 34398 6734 34426 6762
rect 35630 7294 35658 7322
rect 35126 6790 35154 6818
rect 35350 6790 35378 6818
rect 35070 6734 35098 6762
rect 35518 7126 35546 7154
rect 34582 6285 34610 6286
rect 34582 6259 34600 6285
rect 34600 6259 34610 6285
rect 34582 6258 34610 6259
rect 34634 6285 34662 6286
rect 34634 6259 34636 6285
rect 34636 6259 34662 6285
rect 34634 6258 34662 6259
rect 34686 6285 34714 6286
rect 34738 6285 34766 6286
rect 34686 6259 34698 6285
rect 34698 6259 34714 6285
rect 34738 6259 34760 6285
rect 34760 6259 34766 6285
rect 34686 6258 34714 6259
rect 34738 6258 34766 6259
rect 34790 6258 34818 6286
rect 34842 6285 34870 6286
rect 34894 6285 34922 6286
rect 34842 6259 34848 6285
rect 34848 6259 34870 6285
rect 34894 6259 34910 6285
rect 34910 6259 34922 6285
rect 34842 6258 34870 6259
rect 34894 6258 34922 6259
rect 34946 6285 34974 6286
rect 34946 6259 34972 6285
rect 34972 6259 34974 6285
rect 34946 6258 34974 6259
rect 34998 6285 35026 6286
rect 34998 6259 35008 6285
rect 35008 6259 35026 6285
rect 34998 6258 35026 6259
rect 35126 5894 35154 5922
rect 35742 7182 35770 7210
rect 34582 5501 34610 5502
rect 34582 5475 34600 5501
rect 34600 5475 34610 5501
rect 34582 5474 34610 5475
rect 34634 5501 34662 5502
rect 34634 5475 34636 5501
rect 34636 5475 34662 5501
rect 34634 5474 34662 5475
rect 34686 5501 34714 5502
rect 34738 5501 34766 5502
rect 34686 5475 34698 5501
rect 34698 5475 34714 5501
rect 34738 5475 34760 5501
rect 34760 5475 34766 5501
rect 34686 5474 34714 5475
rect 34738 5474 34766 5475
rect 34790 5474 34818 5502
rect 34842 5501 34870 5502
rect 34894 5501 34922 5502
rect 34842 5475 34848 5501
rect 34848 5475 34870 5501
rect 34894 5475 34910 5501
rect 34910 5475 34922 5501
rect 34842 5474 34870 5475
rect 34894 5474 34922 5475
rect 34946 5501 34974 5502
rect 34946 5475 34972 5501
rect 34972 5475 34974 5501
rect 34946 5474 34974 5475
rect 34998 5501 35026 5502
rect 34998 5475 35008 5501
rect 35008 5475 35026 5501
rect 34998 5474 35026 5475
rect 34174 5305 34202 5306
rect 34174 5279 34175 5305
rect 34175 5279 34201 5305
rect 34201 5279 34202 5305
rect 34174 5278 34202 5279
rect 34174 4886 34202 4914
rect 33670 2982 33698 3010
rect 33334 2870 33362 2898
rect 33334 2590 33362 2618
rect 33670 2561 33698 2562
rect 33670 2535 33671 2561
rect 33671 2535 33697 2561
rect 33697 2535 33698 2561
rect 33670 2534 33698 2535
rect 34174 4521 34202 4522
rect 34174 4495 34175 4521
rect 34175 4495 34201 4521
rect 34201 4495 34202 4521
rect 34174 4494 34202 4495
rect 34510 5054 34538 5082
rect 34678 4913 34706 4914
rect 34678 4887 34679 4913
rect 34679 4887 34705 4913
rect 34705 4887 34706 4913
rect 34678 4886 34706 4887
rect 34582 4717 34610 4718
rect 34582 4691 34600 4717
rect 34600 4691 34610 4717
rect 34582 4690 34610 4691
rect 34634 4717 34662 4718
rect 34634 4691 34636 4717
rect 34636 4691 34662 4717
rect 34634 4690 34662 4691
rect 34686 4717 34714 4718
rect 34738 4717 34766 4718
rect 34686 4691 34698 4717
rect 34698 4691 34714 4717
rect 34738 4691 34760 4717
rect 34760 4691 34766 4717
rect 34686 4690 34714 4691
rect 34738 4690 34766 4691
rect 34790 4690 34818 4718
rect 34842 4717 34870 4718
rect 34894 4717 34922 4718
rect 34842 4691 34848 4717
rect 34848 4691 34870 4717
rect 34894 4691 34910 4717
rect 34910 4691 34922 4717
rect 34842 4690 34870 4691
rect 34894 4690 34922 4691
rect 34946 4717 34974 4718
rect 34946 4691 34972 4717
rect 34972 4691 34974 4717
rect 34946 4690 34974 4691
rect 34998 4717 35026 4718
rect 34998 4691 35008 4717
rect 35008 4691 35026 4717
rect 34998 4690 35026 4691
rect 34678 4494 34706 4522
rect 33782 3345 33810 3346
rect 33782 3319 33783 3345
rect 33783 3319 33809 3345
rect 33809 3319 33810 3345
rect 33782 3318 33810 3319
rect 33782 2926 33810 2954
rect 34174 3737 34202 3738
rect 34174 3711 34175 3737
rect 34175 3711 34201 3737
rect 34201 3711 34202 3737
rect 34174 3710 34202 3711
rect 35070 4382 35098 4410
rect 34846 4102 34874 4130
rect 34582 3933 34610 3934
rect 34582 3907 34600 3933
rect 34600 3907 34610 3933
rect 34582 3906 34610 3907
rect 34634 3933 34662 3934
rect 34634 3907 34636 3933
rect 34636 3907 34662 3933
rect 34634 3906 34662 3907
rect 34686 3933 34714 3934
rect 34738 3933 34766 3934
rect 34686 3907 34698 3933
rect 34698 3907 34714 3933
rect 34738 3907 34760 3933
rect 34760 3907 34766 3933
rect 34686 3906 34714 3907
rect 34738 3906 34766 3907
rect 34790 3906 34818 3934
rect 34842 3933 34870 3934
rect 34894 3933 34922 3934
rect 34842 3907 34848 3933
rect 34848 3907 34870 3933
rect 34894 3907 34910 3933
rect 34910 3907 34922 3933
rect 34842 3906 34870 3907
rect 34894 3906 34922 3907
rect 34946 3933 34974 3934
rect 34946 3907 34972 3933
rect 34972 3907 34974 3933
rect 34946 3906 34974 3907
rect 34998 3933 35026 3934
rect 34998 3907 35008 3933
rect 35008 3907 35026 3933
rect 34998 3906 35026 3907
rect 35238 5305 35266 5306
rect 35238 5279 35239 5305
rect 35239 5279 35265 5305
rect 35265 5279 35266 5305
rect 35238 5278 35266 5279
rect 35182 4129 35210 4130
rect 35182 4103 35183 4129
rect 35183 4103 35209 4129
rect 35209 4103 35210 4129
rect 35182 4102 35210 4103
rect 33950 3345 33978 3346
rect 33950 3319 33951 3345
rect 33951 3319 33977 3345
rect 33977 3319 33978 3345
rect 33950 3318 33978 3319
rect 33894 3262 33922 3290
rect 33894 2870 33922 2898
rect 34582 3149 34610 3150
rect 34582 3123 34600 3149
rect 34600 3123 34610 3149
rect 34582 3122 34610 3123
rect 34634 3149 34662 3150
rect 34634 3123 34636 3149
rect 34636 3123 34662 3149
rect 34634 3122 34662 3123
rect 34686 3149 34714 3150
rect 34738 3149 34766 3150
rect 34686 3123 34698 3149
rect 34698 3123 34714 3149
rect 34738 3123 34760 3149
rect 34760 3123 34766 3149
rect 34686 3122 34714 3123
rect 34738 3122 34766 3123
rect 34790 3122 34818 3150
rect 34842 3149 34870 3150
rect 34894 3149 34922 3150
rect 34842 3123 34848 3149
rect 34848 3123 34870 3149
rect 34894 3123 34910 3149
rect 34910 3123 34922 3149
rect 34842 3122 34870 3123
rect 34894 3122 34922 3123
rect 34946 3149 34974 3150
rect 34946 3123 34972 3149
rect 34972 3123 34974 3149
rect 34946 3122 34974 3123
rect 34998 3149 35026 3150
rect 34998 3123 35008 3149
rect 35008 3123 35026 3149
rect 34998 3122 35026 3123
rect 34678 2590 34706 2618
rect 34510 2422 34538 2450
rect 33446 1721 33474 1722
rect 33446 1695 33447 1721
rect 33447 1695 33473 1721
rect 33473 1695 33474 1721
rect 33446 1694 33474 1695
rect 34582 2365 34610 2366
rect 34582 2339 34600 2365
rect 34600 2339 34610 2365
rect 34582 2338 34610 2339
rect 34634 2365 34662 2366
rect 34634 2339 34636 2365
rect 34636 2339 34662 2365
rect 34634 2338 34662 2339
rect 34686 2365 34714 2366
rect 34738 2365 34766 2366
rect 34686 2339 34698 2365
rect 34698 2339 34714 2365
rect 34738 2339 34760 2365
rect 34760 2339 34766 2365
rect 34686 2338 34714 2339
rect 34738 2338 34766 2339
rect 34790 2338 34818 2366
rect 34842 2365 34870 2366
rect 34894 2365 34922 2366
rect 34842 2339 34848 2365
rect 34848 2339 34870 2365
rect 34894 2339 34910 2365
rect 34910 2339 34922 2365
rect 34842 2338 34870 2339
rect 34894 2338 34922 2339
rect 34946 2365 34974 2366
rect 34946 2339 34972 2365
rect 34972 2339 34974 2365
rect 34946 2338 34974 2339
rect 34998 2365 35026 2366
rect 34998 2339 35008 2365
rect 35008 2339 35026 2365
rect 34998 2338 35026 2339
rect 35070 1694 35098 1722
rect 35350 4129 35378 4130
rect 35350 4103 35351 4129
rect 35351 4103 35377 4129
rect 35377 4103 35378 4129
rect 35350 4102 35378 4103
rect 35294 3374 35322 3402
rect 35630 5950 35658 5978
rect 35686 4886 35714 4914
rect 36694 11102 36722 11130
rect 37082 10597 37110 10598
rect 37082 10571 37100 10597
rect 37100 10571 37110 10597
rect 37082 10570 37110 10571
rect 37134 10597 37162 10598
rect 37134 10571 37136 10597
rect 37136 10571 37162 10597
rect 37134 10570 37162 10571
rect 37186 10597 37214 10598
rect 37238 10597 37266 10598
rect 37186 10571 37198 10597
rect 37198 10571 37214 10597
rect 37238 10571 37260 10597
rect 37260 10571 37266 10597
rect 37186 10570 37214 10571
rect 37238 10570 37266 10571
rect 37290 10570 37318 10598
rect 37342 10597 37370 10598
rect 37394 10597 37422 10598
rect 37342 10571 37348 10597
rect 37348 10571 37370 10597
rect 37394 10571 37410 10597
rect 37410 10571 37422 10597
rect 37342 10570 37370 10571
rect 37394 10570 37422 10571
rect 37446 10597 37474 10598
rect 37446 10571 37472 10597
rect 37472 10571 37474 10597
rect 37446 10570 37474 10571
rect 37498 10597 37526 10598
rect 37498 10571 37508 10597
rect 37508 10571 37526 10597
rect 37498 10570 37526 10571
rect 36190 9926 36218 9954
rect 36694 9926 36722 9954
rect 36134 9142 36162 9170
rect 36358 9590 36386 9618
rect 36862 9534 36890 9562
rect 36694 9142 36722 9170
rect 36414 8806 36442 8834
rect 36134 8078 36162 8106
rect 37082 9813 37110 9814
rect 37082 9787 37100 9813
rect 37100 9787 37110 9813
rect 37082 9786 37110 9787
rect 37134 9813 37162 9814
rect 37134 9787 37136 9813
rect 37136 9787 37162 9813
rect 37134 9786 37162 9787
rect 37186 9813 37214 9814
rect 37238 9813 37266 9814
rect 37186 9787 37198 9813
rect 37198 9787 37214 9813
rect 37238 9787 37260 9813
rect 37260 9787 37266 9813
rect 37186 9786 37214 9787
rect 37238 9786 37266 9787
rect 37290 9786 37318 9814
rect 37342 9813 37370 9814
rect 37394 9813 37422 9814
rect 37342 9787 37348 9813
rect 37348 9787 37370 9813
rect 37394 9787 37410 9813
rect 37410 9787 37422 9813
rect 37342 9786 37370 9787
rect 37394 9786 37422 9787
rect 37446 9813 37474 9814
rect 37446 9787 37472 9813
rect 37472 9787 37474 9813
rect 37446 9786 37474 9787
rect 37498 9813 37526 9814
rect 37498 9787 37508 9813
rect 37508 9787 37526 9813
rect 37498 9786 37526 9787
rect 37310 9198 37338 9226
rect 37590 9225 37618 9226
rect 37590 9199 37591 9225
rect 37591 9199 37617 9225
rect 37617 9199 37618 9225
rect 37590 9198 37618 9199
rect 36918 9086 36946 9114
rect 37082 9029 37110 9030
rect 37082 9003 37100 9029
rect 37100 9003 37110 9029
rect 37082 9002 37110 9003
rect 37134 9029 37162 9030
rect 37134 9003 37136 9029
rect 37136 9003 37162 9029
rect 37134 9002 37162 9003
rect 37186 9029 37214 9030
rect 37238 9029 37266 9030
rect 37186 9003 37198 9029
rect 37198 9003 37214 9029
rect 37238 9003 37260 9029
rect 37260 9003 37266 9029
rect 37186 9002 37214 9003
rect 37238 9002 37266 9003
rect 37290 9002 37318 9030
rect 37342 9029 37370 9030
rect 37394 9029 37422 9030
rect 37342 9003 37348 9029
rect 37348 9003 37370 9029
rect 37394 9003 37410 9029
rect 37410 9003 37422 9029
rect 37342 9002 37370 9003
rect 37394 9002 37422 9003
rect 37446 9029 37474 9030
rect 37446 9003 37472 9029
rect 37472 9003 37474 9029
rect 37446 9002 37474 9003
rect 37498 9029 37526 9030
rect 37498 9003 37508 9029
rect 37508 9003 37526 9029
rect 37498 9002 37526 9003
rect 36862 8750 36890 8778
rect 37310 8777 37338 8778
rect 37310 8751 37311 8777
rect 37311 8751 37337 8777
rect 37337 8751 37338 8777
rect 37310 8750 37338 8751
rect 37082 8245 37110 8246
rect 37082 8219 37100 8245
rect 37100 8219 37110 8245
rect 37082 8218 37110 8219
rect 37134 8245 37162 8246
rect 37134 8219 37136 8245
rect 37136 8219 37162 8245
rect 37134 8218 37162 8219
rect 37186 8245 37214 8246
rect 37238 8245 37266 8246
rect 37186 8219 37198 8245
rect 37198 8219 37214 8245
rect 37238 8219 37260 8245
rect 37260 8219 37266 8245
rect 37186 8218 37214 8219
rect 37238 8218 37266 8219
rect 37290 8218 37318 8246
rect 37342 8245 37370 8246
rect 37394 8245 37422 8246
rect 37342 8219 37348 8245
rect 37348 8219 37370 8245
rect 37394 8219 37410 8245
rect 37410 8219 37422 8245
rect 37342 8218 37370 8219
rect 37394 8218 37422 8219
rect 37446 8245 37474 8246
rect 37446 8219 37472 8245
rect 37472 8219 37474 8245
rect 37446 8218 37474 8219
rect 37498 8245 37526 8246
rect 37498 8219 37508 8245
rect 37508 8219 37526 8245
rect 37498 8218 37526 8219
rect 37646 8750 37674 8778
rect 37082 7461 37110 7462
rect 37082 7435 37100 7461
rect 37100 7435 37110 7461
rect 37082 7434 37110 7435
rect 37134 7461 37162 7462
rect 37134 7435 37136 7461
rect 37136 7435 37162 7461
rect 37134 7434 37162 7435
rect 37186 7461 37214 7462
rect 37238 7461 37266 7462
rect 37186 7435 37198 7461
rect 37198 7435 37214 7461
rect 37238 7435 37260 7461
rect 37260 7435 37266 7461
rect 37186 7434 37214 7435
rect 37238 7434 37266 7435
rect 37290 7434 37318 7462
rect 37342 7461 37370 7462
rect 37394 7461 37422 7462
rect 37342 7435 37348 7461
rect 37348 7435 37370 7461
rect 37394 7435 37410 7461
rect 37410 7435 37422 7461
rect 37342 7434 37370 7435
rect 37394 7434 37422 7435
rect 37446 7461 37474 7462
rect 37446 7435 37472 7461
rect 37472 7435 37474 7461
rect 37446 7434 37474 7435
rect 37498 7461 37526 7462
rect 37498 7435 37508 7461
rect 37508 7435 37526 7461
rect 37498 7434 37526 7435
rect 36078 7238 36106 7266
rect 36414 7265 36442 7266
rect 36414 7239 36415 7265
rect 36415 7239 36441 7265
rect 36441 7239 36442 7265
rect 36414 7238 36442 7239
rect 36694 7238 36722 7266
rect 36134 6734 36162 6762
rect 36694 6734 36722 6762
rect 37082 6677 37110 6678
rect 37082 6651 37100 6677
rect 37100 6651 37110 6677
rect 37082 6650 37110 6651
rect 37134 6677 37162 6678
rect 37134 6651 37136 6677
rect 37136 6651 37162 6677
rect 37134 6650 37162 6651
rect 37186 6677 37214 6678
rect 37238 6677 37266 6678
rect 37186 6651 37198 6677
rect 37198 6651 37214 6677
rect 37238 6651 37260 6677
rect 37260 6651 37266 6677
rect 37186 6650 37214 6651
rect 37238 6650 37266 6651
rect 37290 6650 37318 6678
rect 37342 6677 37370 6678
rect 37394 6677 37422 6678
rect 37342 6651 37348 6677
rect 37348 6651 37370 6677
rect 37394 6651 37410 6677
rect 37410 6651 37422 6677
rect 37342 6650 37370 6651
rect 37394 6650 37422 6651
rect 37446 6677 37474 6678
rect 37446 6651 37472 6677
rect 37472 6651 37474 6677
rect 37446 6650 37474 6651
rect 37498 6677 37526 6678
rect 37498 6651 37508 6677
rect 37508 6651 37526 6677
rect 37498 6650 37526 6651
rect 37082 5893 37110 5894
rect 37082 5867 37100 5893
rect 37100 5867 37110 5893
rect 37082 5866 37110 5867
rect 37134 5893 37162 5894
rect 37134 5867 37136 5893
rect 37136 5867 37162 5893
rect 37134 5866 37162 5867
rect 37186 5893 37214 5894
rect 37238 5893 37266 5894
rect 37186 5867 37198 5893
rect 37198 5867 37214 5893
rect 37238 5867 37260 5893
rect 37260 5867 37266 5893
rect 37186 5866 37214 5867
rect 37238 5866 37266 5867
rect 37290 5866 37318 5894
rect 37342 5893 37370 5894
rect 37394 5893 37422 5894
rect 37342 5867 37348 5893
rect 37348 5867 37370 5893
rect 37394 5867 37410 5893
rect 37410 5867 37422 5893
rect 37342 5866 37370 5867
rect 37394 5866 37422 5867
rect 37446 5893 37474 5894
rect 37446 5867 37472 5893
rect 37472 5867 37474 5893
rect 37446 5866 37474 5867
rect 37498 5893 37526 5894
rect 37498 5867 37508 5893
rect 37508 5867 37526 5893
rect 37498 5866 37526 5867
rect 35966 5670 35994 5698
rect 35742 5222 35770 5250
rect 35686 4438 35714 4466
rect 35910 5222 35938 5250
rect 35966 5278 35994 5306
rect 37142 5697 37170 5698
rect 37142 5671 37143 5697
rect 37143 5671 37169 5697
rect 37169 5671 37170 5697
rect 37142 5670 37170 5671
rect 36134 4942 36162 4970
rect 36078 4886 36106 4914
rect 35742 3793 35770 3794
rect 35742 3767 35743 3793
rect 35743 3767 35769 3793
rect 35769 3767 35770 3793
rect 35742 3766 35770 3767
rect 35518 2478 35546 2506
rect 35742 3374 35770 3402
rect 35742 3009 35770 3010
rect 35742 2983 35743 3009
rect 35743 2983 35769 3009
rect 35769 2983 35770 3009
rect 35742 2982 35770 2983
rect 35686 2534 35714 2562
rect 35910 3793 35938 3794
rect 35910 3767 35911 3793
rect 35911 3767 35937 3793
rect 35937 3767 35938 3793
rect 35910 3766 35938 3767
rect 35854 3318 35882 3346
rect 35910 3009 35938 3010
rect 35910 2983 35911 3009
rect 35911 2983 35937 3009
rect 35937 2983 35938 3009
rect 35910 2982 35938 2983
rect 35686 1750 35714 1778
rect 37082 5109 37110 5110
rect 37082 5083 37100 5109
rect 37100 5083 37110 5109
rect 37082 5082 37110 5083
rect 37134 5109 37162 5110
rect 37134 5083 37136 5109
rect 37136 5083 37162 5109
rect 37134 5082 37162 5083
rect 37186 5109 37214 5110
rect 37238 5109 37266 5110
rect 37186 5083 37198 5109
rect 37198 5083 37214 5109
rect 37238 5083 37260 5109
rect 37260 5083 37266 5109
rect 37186 5082 37214 5083
rect 37238 5082 37266 5083
rect 37290 5082 37318 5110
rect 37342 5109 37370 5110
rect 37394 5109 37422 5110
rect 37342 5083 37348 5109
rect 37348 5083 37370 5109
rect 37394 5083 37410 5109
rect 37410 5083 37422 5109
rect 37342 5082 37370 5083
rect 37394 5082 37422 5083
rect 37446 5109 37474 5110
rect 37446 5083 37472 5109
rect 37472 5083 37474 5109
rect 37446 5082 37474 5083
rect 37498 5109 37526 5110
rect 37498 5083 37508 5109
rect 37508 5083 37526 5109
rect 37498 5082 37526 5083
rect 36694 4942 36722 4970
rect 36862 4942 36890 4970
rect 36694 3374 36722 3402
rect 37310 4942 37338 4970
rect 37590 4913 37618 4914
rect 37590 4887 37591 4913
rect 37591 4887 37617 4913
rect 37617 4887 37618 4913
rect 37590 4886 37618 4887
rect 37702 5222 37730 5250
rect 37646 4942 37674 4970
rect 38262 5222 38290 5250
rect 38430 5222 38458 5250
rect 38598 5222 38626 5250
rect 38150 4886 38178 4914
rect 37870 4550 37898 4578
rect 37590 4438 37618 4466
rect 37082 4325 37110 4326
rect 37082 4299 37100 4325
rect 37100 4299 37110 4325
rect 37082 4298 37110 4299
rect 37134 4325 37162 4326
rect 37134 4299 37136 4325
rect 37136 4299 37162 4325
rect 37134 4298 37162 4299
rect 37186 4325 37214 4326
rect 37238 4325 37266 4326
rect 37186 4299 37198 4325
rect 37198 4299 37214 4325
rect 37238 4299 37260 4325
rect 37260 4299 37266 4325
rect 37186 4298 37214 4299
rect 37238 4298 37266 4299
rect 37290 4298 37318 4326
rect 37342 4325 37370 4326
rect 37394 4325 37422 4326
rect 37342 4299 37348 4325
rect 37348 4299 37370 4325
rect 37394 4299 37410 4325
rect 37410 4299 37422 4325
rect 37342 4298 37370 4299
rect 37394 4298 37422 4299
rect 37446 4325 37474 4326
rect 37446 4299 37472 4325
rect 37472 4299 37474 4325
rect 37446 4298 37474 4299
rect 37498 4325 37526 4326
rect 37498 4299 37508 4325
rect 37508 4299 37526 4325
rect 37498 4298 37526 4299
rect 37082 3541 37110 3542
rect 37082 3515 37100 3541
rect 37100 3515 37110 3541
rect 37082 3514 37110 3515
rect 37134 3541 37162 3542
rect 37134 3515 37136 3541
rect 37136 3515 37162 3541
rect 37134 3514 37162 3515
rect 37186 3541 37214 3542
rect 37238 3541 37266 3542
rect 37186 3515 37198 3541
rect 37198 3515 37214 3541
rect 37238 3515 37260 3541
rect 37260 3515 37266 3541
rect 37186 3514 37214 3515
rect 37238 3514 37266 3515
rect 37290 3514 37318 3542
rect 37342 3541 37370 3542
rect 37394 3541 37422 3542
rect 37342 3515 37348 3541
rect 37348 3515 37370 3541
rect 37394 3515 37410 3541
rect 37410 3515 37422 3541
rect 37342 3514 37370 3515
rect 37394 3514 37422 3515
rect 37446 3541 37474 3542
rect 37446 3515 37472 3541
rect 37472 3515 37474 3541
rect 37446 3514 37474 3515
rect 37498 3541 37526 3542
rect 37498 3515 37508 3541
rect 37508 3515 37526 3541
rect 37498 3514 37526 3515
rect 36134 2926 36162 2954
rect 36694 2953 36722 2954
rect 36694 2927 36695 2953
rect 36695 2927 36721 2953
rect 36721 2927 36722 2953
rect 36694 2926 36722 2927
rect 37030 3262 37058 3290
rect 36862 2926 36890 2954
rect 36134 2590 36162 2618
rect 37646 4382 37674 4410
rect 37702 4129 37730 4130
rect 37702 4103 37703 4129
rect 37703 4103 37729 4129
rect 37729 4103 37730 4129
rect 37702 4102 37730 4103
rect 37870 4129 37898 4130
rect 37870 4103 37871 4129
rect 37871 4103 37897 4129
rect 37897 4103 37898 4129
rect 37870 4102 37898 4103
rect 37590 3345 37618 3346
rect 37590 3319 37591 3345
rect 37591 3319 37617 3345
rect 37617 3319 37618 3345
rect 37590 3318 37618 3319
rect 37142 2953 37170 2954
rect 37142 2927 37143 2953
rect 37143 2927 37169 2953
rect 37169 2927 37170 2953
rect 37142 2926 37170 2927
rect 37366 2953 37394 2954
rect 37366 2927 37367 2953
rect 37367 2927 37393 2953
rect 37393 2927 37394 2953
rect 37366 2926 37394 2927
rect 37082 2757 37110 2758
rect 37082 2731 37100 2757
rect 37100 2731 37110 2757
rect 37082 2730 37110 2731
rect 37134 2757 37162 2758
rect 37134 2731 37136 2757
rect 37136 2731 37162 2757
rect 37134 2730 37162 2731
rect 37186 2757 37214 2758
rect 37238 2757 37266 2758
rect 37186 2731 37198 2757
rect 37198 2731 37214 2757
rect 37238 2731 37260 2757
rect 37260 2731 37266 2757
rect 37186 2730 37214 2731
rect 37238 2730 37266 2731
rect 37290 2730 37318 2758
rect 37342 2757 37370 2758
rect 37394 2757 37422 2758
rect 37342 2731 37348 2757
rect 37348 2731 37370 2757
rect 37394 2731 37410 2757
rect 37410 2731 37422 2757
rect 37342 2730 37370 2731
rect 37394 2730 37422 2731
rect 37446 2757 37474 2758
rect 37446 2731 37472 2757
rect 37472 2731 37474 2757
rect 37446 2730 37474 2731
rect 37498 2757 37526 2758
rect 37498 2731 37508 2757
rect 37508 2731 37526 2757
rect 37498 2730 37526 2731
rect 38262 4577 38290 4578
rect 38262 4551 38263 4577
rect 38263 4551 38289 4577
rect 38289 4551 38290 4577
rect 38262 4550 38290 4551
rect 38430 4577 38458 4578
rect 38430 4551 38431 4577
rect 38431 4551 38457 4577
rect 38457 4551 38458 4577
rect 38430 4550 38458 4551
rect 38878 4913 38906 4914
rect 38878 4887 38879 4913
rect 38879 4887 38905 4913
rect 38905 4887 38906 4913
rect 38878 4886 38906 4887
rect 38262 4102 38290 4130
rect 38654 4129 38682 4130
rect 38654 4103 38655 4129
rect 38655 4103 38681 4129
rect 38681 4103 38682 4129
rect 38654 4102 38682 4103
rect 37702 3289 37730 3290
rect 37702 3263 37703 3289
rect 37703 3263 37729 3289
rect 37729 3263 37730 3289
rect 37702 3262 37730 3263
rect 37926 3262 37954 3290
rect 38150 3318 38178 3346
rect 37702 2982 37730 3010
rect 38150 2534 38178 2562
rect 38262 3262 38290 3290
rect 37082 1973 37110 1974
rect 37082 1947 37100 1973
rect 37100 1947 37110 1973
rect 37082 1946 37110 1947
rect 37134 1973 37162 1974
rect 37134 1947 37136 1973
rect 37136 1947 37162 1973
rect 37134 1946 37162 1947
rect 37186 1973 37214 1974
rect 37238 1973 37266 1974
rect 37186 1947 37198 1973
rect 37198 1947 37214 1973
rect 37238 1947 37260 1973
rect 37260 1947 37266 1973
rect 37186 1946 37214 1947
rect 37238 1946 37266 1947
rect 37290 1946 37318 1974
rect 37342 1973 37370 1974
rect 37394 1973 37422 1974
rect 37342 1947 37348 1973
rect 37348 1947 37370 1973
rect 37394 1947 37410 1973
rect 37410 1947 37422 1973
rect 37342 1946 37370 1947
rect 37394 1946 37422 1947
rect 37446 1973 37474 1974
rect 37446 1947 37472 1973
rect 37472 1947 37474 1973
rect 37446 1946 37474 1947
rect 37498 1973 37526 1974
rect 37498 1947 37508 1973
rect 37508 1947 37526 1973
rect 37498 1946 37526 1947
rect 36190 1862 36218 1890
rect 37590 1862 37618 1890
rect 38150 1806 38178 1834
rect 37142 1721 37170 1722
rect 37142 1695 37143 1721
rect 37143 1695 37169 1721
rect 37169 1695 37170 1721
rect 37142 1694 37170 1695
rect 37422 1750 37450 1778
rect 34582 1581 34610 1582
rect 34582 1555 34600 1581
rect 34600 1555 34610 1581
rect 34582 1554 34610 1555
rect 34634 1581 34662 1582
rect 34634 1555 34636 1581
rect 34636 1555 34662 1581
rect 34634 1554 34662 1555
rect 34686 1581 34714 1582
rect 34738 1581 34766 1582
rect 34686 1555 34698 1581
rect 34698 1555 34714 1581
rect 34738 1555 34760 1581
rect 34760 1555 34766 1581
rect 34686 1554 34714 1555
rect 34738 1554 34766 1555
rect 34790 1554 34818 1582
rect 34842 1581 34870 1582
rect 34894 1581 34922 1582
rect 34842 1555 34848 1581
rect 34848 1555 34870 1581
rect 34894 1555 34910 1581
rect 34910 1555 34922 1581
rect 34842 1554 34870 1555
rect 34894 1554 34922 1555
rect 34946 1581 34974 1582
rect 34946 1555 34972 1581
rect 34972 1555 34974 1581
rect 34946 1554 34974 1555
rect 34998 1581 35026 1582
rect 34998 1555 35008 1581
rect 35008 1555 35026 1581
rect 34998 1554 35026 1555
rect 38430 2590 38458 2618
rect 38822 2590 38850 2618
rect 38878 2561 38906 2562
rect 38878 2535 38879 2561
rect 38879 2535 38905 2561
rect 38905 2535 38906 2561
rect 38878 2534 38906 2535
rect 38990 2478 39018 2506
rect 38934 1806 38962 1834
rect 38654 1777 38682 1778
rect 38654 1751 38655 1777
rect 38655 1751 38681 1777
rect 38681 1751 38682 1777
rect 38654 1750 38682 1751
rect 38822 1777 38850 1778
rect 38822 1751 38823 1777
rect 38823 1751 38849 1777
rect 38849 1751 38850 1777
rect 38822 1750 38850 1751
<< metal3 >>
rect 2077 18410 2082 18438
rect 2110 18410 2134 18438
rect 2162 18410 2186 18438
rect 2214 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2394 18438
rect 2422 18410 2446 18438
rect 2474 18410 2498 18438
rect 2526 18410 2531 18438
rect 7077 18410 7082 18438
rect 7110 18410 7134 18438
rect 7162 18410 7186 18438
rect 7214 18410 7238 18438
rect 7266 18410 7290 18438
rect 7318 18410 7342 18438
rect 7370 18410 7394 18438
rect 7422 18410 7446 18438
rect 7474 18410 7498 18438
rect 7526 18410 7531 18438
rect 12077 18410 12082 18438
rect 12110 18410 12134 18438
rect 12162 18410 12186 18438
rect 12214 18410 12238 18438
rect 12266 18410 12290 18438
rect 12318 18410 12342 18438
rect 12370 18410 12394 18438
rect 12422 18410 12446 18438
rect 12474 18410 12498 18438
rect 12526 18410 12531 18438
rect 17077 18410 17082 18438
rect 17110 18410 17134 18438
rect 17162 18410 17186 18438
rect 17214 18410 17238 18438
rect 17266 18410 17290 18438
rect 17318 18410 17342 18438
rect 17370 18410 17394 18438
rect 17422 18410 17446 18438
rect 17474 18410 17498 18438
rect 17526 18410 17531 18438
rect 22077 18410 22082 18438
rect 22110 18410 22134 18438
rect 22162 18410 22186 18438
rect 22214 18410 22238 18438
rect 22266 18410 22290 18438
rect 22318 18410 22342 18438
rect 22370 18410 22394 18438
rect 22422 18410 22446 18438
rect 22474 18410 22498 18438
rect 22526 18410 22531 18438
rect 27077 18410 27082 18438
rect 27110 18410 27134 18438
rect 27162 18410 27186 18438
rect 27214 18410 27238 18438
rect 27266 18410 27290 18438
rect 27318 18410 27342 18438
rect 27370 18410 27394 18438
rect 27422 18410 27446 18438
rect 27474 18410 27498 18438
rect 27526 18410 27531 18438
rect 32077 18410 32082 18438
rect 32110 18410 32134 18438
rect 32162 18410 32186 18438
rect 32214 18410 32238 18438
rect 32266 18410 32290 18438
rect 32318 18410 32342 18438
rect 32370 18410 32394 18438
rect 32422 18410 32446 18438
rect 32474 18410 32498 18438
rect 32526 18410 32531 18438
rect 37077 18410 37082 18438
rect 37110 18410 37134 18438
rect 37162 18410 37186 18438
rect 37214 18410 37238 18438
rect 37266 18410 37290 18438
rect 37318 18410 37342 18438
rect 37370 18410 37394 18438
rect 37422 18410 37446 18438
rect 37474 18410 37498 18438
rect 37526 18410 37531 18438
rect 13393 18214 13398 18242
rect 13426 18214 14630 18242
rect 14658 18214 15078 18242
rect 15106 18214 15111 18242
rect 4577 18018 4582 18046
rect 4610 18018 4634 18046
rect 4662 18018 4686 18046
rect 4714 18018 4738 18046
rect 4766 18018 4790 18046
rect 4818 18018 4842 18046
rect 4870 18018 4894 18046
rect 4922 18018 4946 18046
rect 4974 18018 4998 18046
rect 5026 18018 5031 18046
rect 9577 18018 9582 18046
rect 9610 18018 9634 18046
rect 9662 18018 9686 18046
rect 9714 18018 9738 18046
rect 9766 18018 9790 18046
rect 9818 18018 9842 18046
rect 9870 18018 9894 18046
rect 9922 18018 9946 18046
rect 9974 18018 9998 18046
rect 10026 18018 10031 18046
rect 14577 18018 14582 18046
rect 14610 18018 14634 18046
rect 14662 18018 14686 18046
rect 14714 18018 14738 18046
rect 14766 18018 14790 18046
rect 14818 18018 14842 18046
rect 14870 18018 14894 18046
rect 14922 18018 14946 18046
rect 14974 18018 14998 18046
rect 15026 18018 15031 18046
rect 19577 18018 19582 18046
rect 19610 18018 19634 18046
rect 19662 18018 19686 18046
rect 19714 18018 19738 18046
rect 19766 18018 19790 18046
rect 19818 18018 19842 18046
rect 19870 18018 19894 18046
rect 19922 18018 19946 18046
rect 19974 18018 19998 18046
rect 20026 18018 20031 18046
rect 24577 18018 24582 18046
rect 24610 18018 24634 18046
rect 24662 18018 24686 18046
rect 24714 18018 24738 18046
rect 24766 18018 24790 18046
rect 24818 18018 24842 18046
rect 24870 18018 24894 18046
rect 24922 18018 24946 18046
rect 24974 18018 24998 18046
rect 25026 18018 25031 18046
rect 29577 18018 29582 18046
rect 29610 18018 29634 18046
rect 29662 18018 29686 18046
rect 29714 18018 29738 18046
rect 29766 18018 29790 18046
rect 29818 18018 29842 18046
rect 29870 18018 29894 18046
rect 29922 18018 29946 18046
rect 29974 18018 29998 18046
rect 30026 18018 30031 18046
rect 34577 18018 34582 18046
rect 34610 18018 34634 18046
rect 34662 18018 34686 18046
rect 34714 18018 34738 18046
rect 34766 18018 34790 18046
rect 34818 18018 34842 18046
rect 34870 18018 34894 18046
rect 34922 18018 34946 18046
rect 34974 18018 34998 18046
rect 35026 18018 35031 18046
rect 9249 17822 9254 17850
rect 9282 17822 9814 17850
rect 9842 17822 11102 17850
rect 11130 17822 11135 17850
rect 14233 17822 14238 17850
rect 14266 17822 14574 17850
rect 14602 17822 15806 17850
rect 15834 17822 15839 17850
rect 2077 17626 2082 17654
rect 2110 17626 2134 17654
rect 2162 17626 2186 17654
rect 2214 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2394 17654
rect 2422 17626 2446 17654
rect 2474 17626 2498 17654
rect 2526 17626 2531 17654
rect 7077 17626 7082 17654
rect 7110 17626 7134 17654
rect 7162 17626 7186 17654
rect 7214 17626 7238 17654
rect 7266 17626 7290 17654
rect 7318 17626 7342 17654
rect 7370 17626 7394 17654
rect 7422 17626 7446 17654
rect 7474 17626 7498 17654
rect 7526 17626 7531 17654
rect 12077 17626 12082 17654
rect 12110 17626 12134 17654
rect 12162 17626 12186 17654
rect 12214 17626 12238 17654
rect 12266 17626 12290 17654
rect 12318 17626 12342 17654
rect 12370 17626 12394 17654
rect 12422 17626 12446 17654
rect 12474 17626 12498 17654
rect 12526 17626 12531 17654
rect 17077 17626 17082 17654
rect 17110 17626 17134 17654
rect 17162 17626 17186 17654
rect 17214 17626 17238 17654
rect 17266 17626 17290 17654
rect 17318 17626 17342 17654
rect 17370 17626 17394 17654
rect 17422 17626 17446 17654
rect 17474 17626 17498 17654
rect 17526 17626 17531 17654
rect 22077 17626 22082 17654
rect 22110 17626 22134 17654
rect 22162 17626 22186 17654
rect 22214 17626 22238 17654
rect 22266 17626 22290 17654
rect 22318 17626 22342 17654
rect 22370 17626 22394 17654
rect 22422 17626 22446 17654
rect 22474 17626 22498 17654
rect 22526 17626 22531 17654
rect 27077 17626 27082 17654
rect 27110 17626 27134 17654
rect 27162 17626 27186 17654
rect 27214 17626 27238 17654
rect 27266 17626 27290 17654
rect 27318 17626 27342 17654
rect 27370 17626 27394 17654
rect 27422 17626 27446 17654
rect 27474 17626 27498 17654
rect 27526 17626 27531 17654
rect 32077 17626 32082 17654
rect 32110 17626 32134 17654
rect 32162 17626 32186 17654
rect 32214 17626 32238 17654
rect 32266 17626 32290 17654
rect 32318 17626 32342 17654
rect 32370 17626 32394 17654
rect 32422 17626 32446 17654
rect 32474 17626 32498 17654
rect 32526 17626 32531 17654
rect 37077 17626 37082 17654
rect 37110 17626 37134 17654
rect 37162 17626 37186 17654
rect 37214 17626 37238 17654
rect 37266 17626 37290 17654
rect 37318 17626 37342 17654
rect 37370 17626 37394 17654
rect 37422 17626 37446 17654
rect 37474 17626 37498 17654
rect 37526 17626 37531 17654
rect 12609 17318 12614 17346
rect 12642 17318 18494 17346
rect 18522 17318 18527 17346
rect 4577 17234 4582 17262
rect 4610 17234 4634 17262
rect 4662 17234 4686 17262
rect 4714 17234 4738 17262
rect 4766 17234 4790 17262
rect 4818 17234 4842 17262
rect 4870 17234 4894 17262
rect 4922 17234 4946 17262
rect 4974 17234 4998 17262
rect 5026 17234 5031 17262
rect 9577 17234 9582 17262
rect 9610 17234 9634 17262
rect 9662 17234 9686 17262
rect 9714 17234 9738 17262
rect 9766 17234 9790 17262
rect 9818 17234 9842 17262
rect 9870 17234 9894 17262
rect 9922 17234 9946 17262
rect 9974 17234 9998 17262
rect 10026 17234 10031 17262
rect 14577 17234 14582 17262
rect 14610 17234 14634 17262
rect 14662 17234 14686 17262
rect 14714 17234 14738 17262
rect 14766 17234 14790 17262
rect 14818 17234 14842 17262
rect 14870 17234 14894 17262
rect 14922 17234 14946 17262
rect 14974 17234 14998 17262
rect 15026 17234 15031 17262
rect 19577 17234 19582 17262
rect 19610 17234 19634 17262
rect 19662 17234 19686 17262
rect 19714 17234 19738 17262
rect 19766 17234 19790 17262
rect 19818 17234 19842 17262
rect 19870 17234 19894 17262
rect 19922 17234 19946 17262
rect 19974 17234 19998 17262
rect 20026 17234 20031 17262
rect 24577 17234 24582 17262
rect 24610 17234 24634 17262
rect 24662 17234 24686 17262
rect 24714 17234 24738 17262
rect 24766 17234 24790 17262
rect 24818 17234 24842 17262
rect 24870 17234 24894 17262
rect 24922 17234 24946 17262
rect 24974 17234 24998 17262
rect 25026 17234 25031 17262
rect 29577 17234 29582 17262
rect 29610 17234 29634 17262
rect 29662 17234 29686 17262
rect 29714 17234 29738 17262
rect 29766 17234 29790 17262
rect 29818 17234 29842 17262
rect 29870 17234 29894 17262
rect 29922 17234 29946 17262
rect 29974 17234 29998 17262
rect 30026 17234 30031 17262
rect 34577 17234 34582 17262
rect 34610 17234 34634 17262
rect 34662 17234 34686 17262
rect 34714 17234 34738 17262
rect 34766 17234 34790 17262
rect 34818 17234 34842 17262
rect 34870 17234 34894 17262
rect 34922 17234 34946 17262
rect 34974 17234 34998 17262
rect 35026 17234 35031 17262
rect 2077 16842 2082 16870
rect 2110 16842 2134 16870
rect 2162 16842 2186 16870
rect 2214 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2394 16870
rect 2422 16842 2446 16870
rect 2474 16842 2498 16870
rect 2526 16842 2531 16870
rect 7077 16842 7082 16870
rect 7110 16842 7134 16870
rect 7162 16842 7186 16870
rect 7214 16842 7238 16870
rect 7266 16842 7290 16870
rect 7318 16842 7342 16870
rect 7370 16842 7394 16870
rect 7422 16842 7446 16870
rect 7474 16842 7498 16870
rect 7526 16842 7531 16870
rect 12077 16842 12082 16870
rect 12110 16842 12134 16870
rect 12162 16842 12186 16870
rect 12214 16842 12238 16870
rect 12266 16842 12290 16870
rect 12318 16842 12342 16870
rect 12370 16842 12394 16870
rect 12422 16842 12446 16870
rect 12474 16842 12498 16870
rect 12526 16842 12531 16870
rect 17077 16842 17082 16870
rect 17110 16842 17134 16870
rect 17162 16842 17186 16870
rect 17214 16842 17238 16870
rect 17266 16842 17290 16870
rect 17318 16842 17342 16870
rect 17370 16842 17394 16870
rect 17422 16842 17446 16870
rect 17474 16842 17498 16870
rect 17526 16842 17531 16870
rect 22077 16842 22082 16870
rect 22110 16842 22134 16870
rect 22162 16842 22186 16870
rect 22214 16842 22238 16870
rect 22266 16842 22290 16870
rect 22318 16842 22342 16870
rect 22370 16842 22394 16870
rect 22422 16842 22446 16870
rect 22474 16842 22498 16870
rect 22526 16842 22531 16870
rect 27077 16842 27082 16870
rect 27110 16842 27134 16870
rect 27162 16842 27186 16870
rect 27214 16842 27238 16870
rect 27266 16842 27290 16870
rect 27318 16842 27342 16870
rect 27370 16842 27394 16870
rect 27422 16842 27446 16870
rect 27474 16842 27498 16870
rect 27526 16842 27531 16870
rect 32077 16842 32082 16870
rect 32110 16842 32134 16870
rect 32162 16842 32186 16870
rect 32214 16842 32238 16870
rect 32266 16842 32290 16870
rect 32318 16842 32342 16870
rect 32370 16842 32394 16870
rect 32422 16842 32446 16870
rect 32474 16842 32498 16870
rect 32526 16842 32531 16870
rect 37077 16842 37082 16870
rect 37110 16842 37134 16870
rect 37162 16842 37186 16870
rect 37214 16842 37238 16870
rect 37266 16842 37290 16870
rect 37318 16842 37342 16870
rect 37370 16842 37394 16870
rect 37422 16842 37446 16870
rect 37474 16842 37498 16870
rect 37526 16842 37531 16870
rect 7793 16646 7798 16674
rect 7826 16646 9254 16674
rect 9282 16646 9287 16674
rect 11825 16646 11830 16674
rect 11858 16646 12222 16674
rect 12250 16646 12446 16674
rect 12474 16646 14238 16674
rect 14266 16646 14271 16674
rect 16753 16646 16758 16674
rect 16786 16646 16926 16674
rect 16954 16646 16959 16674
rect 4577 16450 4582 16478
rect 4610 16450 4634 16478
rect 4662 16450 4686 16478
rect 4714 16450 4738 16478
rect 4766 16450 4790 16478
rect 4818 16450 4842 16478
rect 4870 16450 4894 16478
rect 4922 16450 4946 16478
rect 4974 16450 4998 16478
rect 5026 16450 5031 16478
rect 9577 16450 9582 16478
rect 9610 16450 9634 16478
rect 9662 16450 9686 16478
rect 9714 16450 9738 16478
rect 9766 16450 9790 16478
rect 9818 16450 9842 16478
rect 9870 16450 9894 16478
rect 9922 16450 9946 16478
rect 9974 16450 9998 16478
rect 10026 16450 10031 16478
rect 14577 16450 14582 16478
rect 14610 16450 14634 16478
rect 14662 16450 14686 16478
rect 14714 16450 14738 16478
rect 14766 16450 14790 16478
rect 14818 16450 14842 16478
rect 14870 16450 14894 16478
rect 14922 16450 14946 16478
rect 14974 16450 14998 16478
rect 15026 16450 15031 16478
rect 19577 16450 19582 16478
rect 19610 16450 19634 16478
rect 19662 16450 19686 16478
rect 19714 16450 19738 16478
rect 19766 16450 19790 16478
rect 19818 16450 19842 16478
rect 19870 16450 19894 16478
rect 19922 16450 19946 16478
rect 19974 16450 19998 16478
rect 20026 16450 20031 16478
rect 24577 16450 24582 16478
rect 24610 16450 24634 16478
rect 24662 16450 24686 16478
rect 24714 16450 24738 16478
rect 24766 16450 24790 16478
rect 24818 16450 24842 16478
rect 24870 16450 24894 16478
rect 24922 16450 24946 16478
rect 24974 16450 24998 16478
rect 25026 16450 25031 16478
rect 29577 16450 29582 16478
rect 29610 16450 29634 16478
rect 29662 16450 29686 16478
rect 29714 16450 29738 16478
rect 29766 16450 29790 16478
rect 29818 16450 29842 16478
rect 29870 16450 29894 16478
rect 29922 16450 29946 16478
rect 29974 16450 29998 16478
rect 30026 16450 30031 16478
rect 34577 16450 34582 16478
rect 34610 16450 34634 16478
rect 34662 16450 34686 16478
rect 34714 16450 34738 16478
rect 34766 16450 34790 16478
rect 34818 16450 34842 16478
rect 34870 16450 34894 16478
rect 34922 16450 34946 16478
rect 34974 16450 34998 16478
rect 35026 16450 35031 16478
rect 18489 16366 18494 16394
rect 18522 16366 24094 16394
rect 24122 16366 24127 16394
rect 10075 16254 10094 16282
rect 10122 16254 10127 16282
rect 10985 16254 10990 16282
rect 11018 16254 11830 16282
rect 11858 16254 11942 16282
rect 11970 16254 11975 16282
rect 16249 16254 16254 16282
rect 16282 16254 16814 16282
rect 16842 16254 16847 16282
rect 22577 16254 22582 16282
rect 22610 16254 24430 16282
rect 24458 16254 24463 16282
rect 15969 16142 15974 16170
rect 16002 16142 16310 16170
rect 16338 16142 16814 16170
rect 16842 16142 16847 16170
rect 2077 16058 2082 16086
rect 2110 16058 2134 16086
rect 2162 16058 2186 16086
rect 2214 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2394 16086
rect 2422 16058 2446 16086
rect 2474 16058 2498 16086
rect 2526 16058 2531 16086
rect 7077 16058 7082 16086
rect 7110 16058 7134 16086
rect 7162 16058 7186 16086
rect 7214 16058 7238 16086
rect 7266 16058 7290 16086
rect 7318 16058 7342 16086
rect 7370 16058 7394 16086
rect 7422 16058 7446 16086
rect 7474 16058 7498 16086
rect 7526 16058 7531 16086
rect 12077 16058 12082 16086
rect 12110 16058 12134 16086
rect 12162 16058 12186 16086
rect 12214 16058 12238 16086
rect 12266 16058 12290 16086
rect 12318 16058 12342 16086
rect 12370 16058 12394 16086
rect 12422 16058 12446 16086
rect 12474 16058 12498 16086
rect 12526 16058 12531 16086
rect 17077 16058 17082 16086
rect 17110 16058 17134 16086
rect 17162 16058 17186 16086
rect 17214 16058 17238 16086
rect 17266 16058 17290 16086
rect 17318 16058 17342 16086
rect 17370 16058 17394 16086
rect 17422 16058 17446 16086
rect 17474 16058 17498 16086
rect 17526 16058 17531 16086
rect 22077 16058 22082 16086
rect 22110 16058 22134 16086
rect 22162 16058 22186 16086
rect 22214 16058 22238 16086
rect 22266 16058 22290 16086
rect 22318 16058 22342 16086
rect 22370 16058 22394 16086
rect 22422 16058 22446 16086
rect 22474 16058 22498 16086
rect 22526 16058 22531 16086
rect 27077 16058 27082 16086
rect 27110 16058 27134 16086
rect 27162 16058 27186 16086
rect 27214 16058 27238 16086
rect 27266 16058 27290 16086
rect 27318 16058 27342 16086
rect 27370 16058 27394 16086
rect 27422 16058 27446 16086
rect 27474 16058 27498 16086
rect 27526 16058 27531 16086
rect 32077 16058 32082 16086
rect 32110 16058 32134 16086
rect 32162 16058 32186 16086
rect 32214 16058 32238 16086
rect 32266 16058 32290 16086
rect 32318 16058 32342 16086
rect 32370 16058 32394 16086
rect 32422 16058 32446 16086
rect 32474 16058 32498 16086
rect 32526 16058 32531 16086
rect 37077 16058 37082 16086
rect 37110 16058 37134 16086
rect 37162 16058 37186 16086
rect 37214 16058 37238 16086
rect 37266 16058 37290 16086
rect 37318 16058 37342 16086
rect 37370 16058 37394 16086
rect 37422 16058 37446 16086
rect 37474 16058 37498 16086
rect 37526 16058 37531 16086
rect 11825 15974 11830 16002
rect 11858 15974 12222 16002
rect 12250 15974 12446 16002
rect 12474 15974 12479 16002
rect 17873 15974 17878 16002
rect 17906 15974 18718 16002
rect 18746 15974 19222 16002
rect 19250 15974 19255 16002
rect 13281 15918 13286 15946
rect 13314 15918 13734 15946
rect 13762 15918 13767 15946
rect 18265 15862 18270 15890
rect 18298 15862 18774 15890
rect 18802 15862 18807 15890
rect 10425 15806 10430 15834
rect 10458 15806 10990 15834
rect 11018 15806 11023 15834
rect 4577 15666 4582 15694
rect 4610 15666 4634 15694
rect 4662 15666 4686 15694
rect 4714 15666 4738 15694
rect 4766 15666 4790 15694
rect 4818 15666 4842 15694
rect 4870 15666 4894 15694
rect 4922 15666 4946 15694
rect 4974 15666 4998 15694
rect 5026 15666 5031 15694
rect 9577 15666 9582 15694
rect 9610 15666 9634 15694
rect 9662 15666 9686 15694
rect 9714 15666 9738 15694
rect 9766 15666 9790 15694
rect 9818 15666 9842 15694
rect 9870 15666 9894 15694
rect 9922 15666 9946 15694
rect 9974 15666 9998 15694
rect 10026 15666 10031 15694
rect 14577 15666 14582 15694
rect 14610 15666 14634 15694
rect 14662 15666 14686 15694
rect 14714 15666 14738 15694
rect 14766 15666 14790 15694
rect 14818 15666 14842 15694
rect 14870 15666 14894 15694
rect 14922 15666 14946 15694
rect 14974 15666 14998 15694
rect 15026 15666 15031 15694
rect 19577 15666 19582 15694
rect 19610 15666 19634 15694
rect 19662 15666 19686 15694
rect 19714 15666 19738 15694
rect 19766 15666 19790 15694
rect 19818 15666 19842 15694
rect 19870 15666 19894 15694
rect 19922 15666 19946 15694
rect 19974 15666 19998 15694
rect 20026 15666 20031 15694
rect 24577 15666 24582 15694
rect 24610 15666 24634 15694
rect 24662 15666 24686 15694
rect 24714 15666 24738 15694
rect 24766 15666 24790 15694
rect 24818 15666 24842 15694
rect 24870 15666 24894 15694
rect 24922 15666 24946 15694
rect 24974 15666 24998 15694
rect 25026 15666 25031 15694
rect 29577 15666 29582 15694
rect 29610 15666 29634 15694
rect 29662 15666 29686 15694
rect 29714 15666 29738 15694
rect 29766 15666 29790 15694
rect 29818 15666 29842 15694
rect 29870 15666 29894 15694
rect 29922 15666 29946 15694
rect 29974 15666 29998 15694
rect 30026 15666 30031 15694
rect 34577 15666 34582 15694
rect 34610 15666 34634 15694
rect 34662 15666 34686 15694
rect 34714 15666 34738 15694
rect 34766 15666 34790 15694
rect 34818 15666 34842 15694
rect 34870 15666 34894 15694
rect 34922 15666 34946 15694
rect 34974 15666 34998 15694
rect 35026 15666 35031 15694
rect 10033 15470 10038 15498
rect 10066 15470 10094 15498
rect 10122 15470 11270 15498
rect 11298 15470 11303 15498
rect 2077 15274 2082 15302
rect 2110 15274 2134 15302
rect 2162 15274 2186 15302
rect 2214 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2394 15302
rect 2422 15274 2446 15302
rect 2474 15274 2498 15302
rect 2526 15274 2531 15302
rect 7077 15274 7082 15302
rect 7110 15274 7134 15302
rect 7162 15274 7186 15302
rect 7214 15274 7238 15302
rect 7266 15274 7290 15302
rect 7318 15274 7342 15302
rect 7370 15274 7394 15302
rect 7422 15274 7446 15302
rect 7474 15274 7498 15302
rect 7526 15274 7531 15302
rect 12077 15274 12082 15302
rect 12110 15274 12134 15302
rect 12162 15274 12186 15302
rect 12214 15274 12238 15302
rect 12266 15274 12290 15302
rect 12318 15274 12342 15302
rect 12370 15274 12394 15302
rect 12422 15274 12446 15302
rect 12474 15274 12498 15302
rect 12526 15274 12531 15302
rect 17077 15274 17082 15302
rect 17110 15274 17134 15302
rect 17162 15274 17186 15302
rect 17214 15274 17238 15302
rect 17266 15274 17290 15302
rect 17318 15274 17342 15302
rect 17370 15274 17394 15302
rect 17422 15274 17446 15302
rect 17474 15274 17498 15302
rect 17526 15274 17531 15302
rect 22077 15274 22082 15302
rect 22110 15274 22134 15302
rect 22162 15274 22186 15302
rect 22214 15274 22238 15302
rect 22266 15274 22290 15302
rect 22318 15274 22342 15302
rect 22370 15274 22394 15302
rect 22422 15274 22446 15302
rect 22474 15274 22498 15302
rect 22526 15274 22531 15302
rect 27077 15274 27082 15302
rect 27110 15274 27134 15302
rect 27162 15274 27186 15302
rect 27214 15274 27238 15302
rect 27266 15274 27290 15302
rect 27318 15274 27342 15302
rect 27370 15274 27394 15302
rect 27422 15274 27446 15302
rect 27474 15274 27498 15302
rect 27526 15274 27531 15302
rect 32077 15274 32082 15302
rect 32110 15274 32134 15302
rect 32162 15274 32186 15302
rect 32214 15274 32238 15302
rect 32266 15274 32290 15302
rect 32318 15274 32342 15302
rect 32370 15274 32394 15302
rect 32422 15274 32446 15302
rect 32474 15274 32498 15302
rect 32526 15274 32531 15302
rect 37077 15274 37082 15302
rect 37110 15274 37134 15302
rect 37162 15274 37186 15302
rect 37214 15274 37238 15302
rect 37266 15274 37290 15302
rect 37318 15274 37342 15302
rect 37370 15274 37394 15302
rect 37422 15274 37446 15302
rect 37474 15274 37498 15302
rect 37526 15274 37531 15302
rect 16305 15134 16310 15162
rect 16338 15134 16926 15162
rect 16954 15134 16959 15162
rect 3817 15078 3822 15106
rect 3850 15078 5558 15106
rect 5586 15078 6118 15106
rect 6146 15078 6151 15106
rect 4577 14882 4582 14910
rect 4610 14882 4634 14910
rect 4662 14882 4686 14910
rect 4714 14882 4738 14910
rect 4766 14882 4790 14910
rect 4818 14882 4842 14910
rect 4870 14882 4894 14910
rect 4922 14882 4946 14910
rect 4974 14882 4998 14910
rect 5026 14882 5031 14910
rect 9577 14882 9582 14910
rect 9610 14882 9634 14910
rect 9662 14882 9686 14910
rect 9714 14882 9738 14910
rect 9766 14882 9790 14910
rect 9818 14882 9842 14910
rect 9870 14882 9894 14910
rect 9922 14882 9946 14910
rect 9974 14882 9998 14910
rect 10026 14882 10031 14910
rect 14577 14882 14582 14910
rect 14610 14882 14634 14910
rect 14662 14882 14686 14910
rect 14714 14882 14738 14910
rect 14766 14882 14790 14910
rect 14818 14882 14842 14910
rect 14870 14882 14894 14910
rect 14922 14882 14946 14910
rect 14974 14882 14998 14910
rect 15026 14882 15031 14910
rect 19577 14882 19582 14910
rect 19610 14882 19634 14910
rect 19662 14882 19686 14910
rect 19714 14882 19738 14910
rect 19766 14882 19790 14910
rect 19818 14882 19842 14910
rect 19870 14882 19894 14910
rect 19922 14882 19946 14910
rect 19974 14882 19998 14910
rect 20026 14882 20031 14910
rect 24577 14882 24582 14910
rect 24610 14882 24634 14910
rect 24662 14882 24686 14910
rect 24714 14882 24738 14910
rect 24766 14882 24790 14910
rect 24818 14882 24842 14910
rect 24870 14882 24894 14910
rect 24922 14882 24946 14910
rect 24974 14882 24998 14910
rect 25026 14882 25031 14910
rect 29577 14882 29582 14910
rect 29610 14882 29634 14910
rect 29662 14882 29686 14910
rect 29714 14882 29738 14910
rect 29766 14882 29790 14910
rect 29818 14882 29842 14910
rect 29870 14882 29894 14910
rect 29922 14882 29946 14910
rect 29974 14882 29998 14910
rect 30026 14882 30031 14910
rect 34577 14882 34582 14910
rect 34610 14882 34634 14910
rect 34662 14882 34686 14910
rect 34714 14882 34738 14910
rect 34766 14882 34790 14910
rect 34818 14882 34842 14910
rect 34870 14882 34894 14910
rect 34922 14882 34946 14910
rect 34974 14882 34998 14910
rect 35026 14882 35031 14910
rect 6113 14798 6118 14826
rect 6146 14798 6902 14826
rect 6930 14798 6935 14826
rect 1969 14686 1974 14714
rect 2002 14686 2478 14714
rect 2506 14686 2646 14714
rect 2674 14686 2679 14714
rect 5553 14686 5558 14714
rect 5586 14686 6118 14714
rect 6146 14686 7798 14714
rect 7826 14686 7831 14714
rect 8465 14686 8470 14714
rect 8498 14686 8974 14714
rect 9002 14686 9007 14714
rect 23417 14686 23422 14714
rect 23450 14686 23926 14714
rect 23954 14686 23959 14714
rect 6897 14630 6902 14658
rect 6930 14630 20790 14658
rect 20818 14630 22582 14658
rect 22610 14630 22615 14658
rect 2077 14490 2082 14518
rect 2110 14490 2134 14518
rect 2162 14490 2186 14518
rect 2214 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2394 14518
rect 2422 14490 2446 14518
rect 2474 14490 2498 14518
rect 2526 14490 2531 14518
rect 7077 14490 7082 14518
rect 7110 14490 7134 14518
rect 7162 14490 7186 14518
rect 7214 14490 7238 14518
rect 7266 14490 7290 14518
rect 7318 14490 7342 14518
rect 7370 14490 7394 14518
rect 7422 14490 7446 14518
rect 7474 14490 7498 14518
rect 7526 14490 7531 14518
rect 12077 14490 12082 14518
rect 12110 14490 12134 14518
rect 12162 14490 12186 14518
rect 12214 14490 12238 14518
rect 12266 14490 12290 14518
rect 12318 14490 12342 14518
rect 12370 14490 12394 14518
rect 12422 14490 12446 14518
rect 12474 14490 12498 14518
rect 12526 14490 12531 14518
rect 17077 14490 17082 14518
rect 17110 14490 17134 14518
rect 17162 14490 17186 14518
rect 17214 14490 17238 14518
rect 17266 14490 17290 14518
rect 17318 14490 17342 14518
rect 17370 14490 17394 14518
rect 17422 14490 17446 14518
rect 17474 14490 17498 14518
rect 17526 14490 17531 14518
rect 22077 14490 22082 14518
rect 22110 14490 22134 14518
rect 22162 14490 22186 14518
rect 22214 14490 22238 14518
rect 22266 14490 22290 14518
rect 22318 14490 22342 14518
rect 22370 14490 22394 14518
rect 22422 14490 22446 14518
rect 22474 14490 22498 14518
rect 22526 14490 22531 14518
rect 27077 14490 27082 14518
rect 27110 14490 27134 14518
rect 27162 14490 27186 14518
rect 27214 14490 27238 14518
rect 27266 14490 27290 14518
rect 27318 14490 27342 14518
rect 27370 14490 27394 14518
rect 27422 14490 27446 14518
rect 27474 14490 27498 14518
rect 27526 14490 27531 14518
rect 32077 14490 32082 14518
rect 32110 14490 32134 14518
rect 32162 14490 32186 14518
rect 32214 14490 32238 14518
rect 32266 14490 32290 14518
rect 32318 14490 32342 14518
rect 32370 14490 32394 14518
rect 32422 14490 32446 14518
rect 32474 14490 32498 14518
rect 32526 14490 32531 14518
rect 37077 14490 37082 14518
rect 37110 14490 37134 14518
rect 37162 14490 37186 14518
rect 37214 14490 37238 14518
rect 37266 14490 37290 14518
rect 37318 14490 37342 14518
rect 37370 14490 37394 14518
rect 37422 14490 37446 14518
rect 37474 14490 37498 14518
rect 37526 14490 37531 14518
rect 2753 14294 2758 14322
rect 2786 14294 3318 14322
rect 3346 14294 3822 14322
rect 3850 14294 3855 14322
rect 8969 14294 8974 14322
rect 9002 14294 10374 14322
rect 10402 14294 10407 14322
rect 15185 14294 15190 14322
rect 15218 14294 16254 14322
rect 16282 14294 16814 14322
rect 16842 14294 18270 14322
rect 18298 14294 18303 14322
rect 19441 14294 19446 14322
rect 19474 14294 20678 14322
rect 20706 14294 21014 14322
rect 21042 14294 21047 14322
rect 22521 14294 22526 14322
rect 22554 14294 23030 14322
rect 23058 14294 24486 14322
rect 24514 14294 24519 14322
rect 15969 14238 15974 14266
rect 16002 14238 16366 14266
rect 16394 14238 16982 14266
rect 17010 14238 17430 14266
rect 17458 14238 17934 14266
rect 17962 14238 17967 14266
rect 23921 14238 23926 14266
rect 23954 14238 25382 14266
rect 25410 14238 25415 14266
rect 4577 14098 4582 14126
rect 4610 14098 4634 14126
rect 4662 14098 4686 14126
rect 4714 14098 4738 14126
rect 4766 14098 4790 14126
rect 4818 14098 4842 14126
rect 4870 14098 4894 14126
rect 4922 14098 4946 14126
rect 4974 14098 4998 14126
rect 5026 14098 5031 14126
rect 9577 14098 9582 14126
rect 9610 14098 9634 14126
rect 9662 14098 9686 14126
rect 9714 14098 9738 14126
rect 9766 14098 9790 14126
rect 9818 14098 9842 14126
rect 9870 14098 9894 14126
rect 9922 14098 9946 14126
rect 9974 14098 9998 14126
rect 10026 14098 10031 14126
rect 14577 14098 14582 14126
rect 14610 14098 14634 14126
rect 14662 14098 14686 14126
rect 14714 14098 14738 14126
rect 14766 14098 14790 14126
rect 14818 14098 14842 14126
rect 14870 14098 14894 14126
rect 14922 14098 14946 14126
rect 14974 14098 14998 14126
rect 15026 14098 15031 14126
rect 19577 14098 19582 14126
rect 19610 14098 19634 14126
rect 19662 14098 19686 14126
rect 19714 14098 19738 14126
rect 19766 14098 19790 14126
rect 19818 14098 19842 14126
rect 19870 14098 19894 14126
rect 19922 14098 19946 14126
rect 19974 14098 19998 14126
rect 20026 14098 20031 14126
rect 24577 14098 24582 14126
rect 24610 14098 24634 14126
rect 24662 14098 24686 14126
rect 24714 14098 24738 14126
rect 24766 14098 24790 14126
rect 24818 14098 24842 14126
rect 24870 14098 24894 14126
rect 24922 14098 24946 14126
rect 24974 14098 24998 14126
rect 25026 14098 25031 14126
rect 29577 14098 29582 14126
rect 29610 14098 29634 14126
rect 29662 14098 29686 14126
rect 29714 14098 29738 14126
rect 29766 14098 29790 14126
rect 29818 14098 29842 14126
rect 29870 14098 29894 14126
rect 29922 14098 29946 14126
rect 29974 14098 29998 14126
rect 30026 14098 30031 14126
rect 34577 14098 34582 14126
rect 34610 14098 34634 14126
rect 34662 14098 34686 14126
rect 34714 14098 34738 14126
rect 34766 14098 34790 14126
rect 34818 14098 34842 14126
rect 34870 14098 34894 14126
rect 34922 14098 34946 14126
rect 34974 14098 34998 14126
rect 35026 14098 35031 14126
rect 27393 13958 27398 13986
rect 27426 13958 27678 13986
rect 27706 13958 27711 13986
rect 11993 13902 11998 13930
rect 12026 13902 12446 13930
rect 12474 13902 12479 13930
rect 14457 13902 14462 13930
rect 14490 13902 14910 13930
rect 14938 13902 15974 13930
rect 16002 13902 16007 13930
rect 21457 13902 21462 13930
rect 21490 13902 23422 13930
rect 23450 13902 23455 13930
rect 8857 13846 8862 13874
rect 8890 13846 26222 13874
rect 26250 13846 26726 13874
rect 26754 13846 26759 13874
rect 2077 13706 2082 13734
rect 2110 13706 2134 13734
rect 2162 13706 2186 13734
rect 2214 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2394 13734
rect 2422 13706 2446 13734
rect 2474 13706 2498 13734
rect 2526 13706 2531 13734
rect 7077 13706 7082 13734
rect 7110 13706 7134 13734
rect 7162 13706 7186 13734
rect 7214 13706 7238 13734
rect 7266 13706 7290 13734
rect 7318 13706 7342 13734
rect 7370 13706 7394 13734
rect 7422 13706 7446 13734
rect 7474 13706 7498 13734
rect 7526 13706 7531 13734
rect 12077 13706 12082 13734
rect 12110 13706 12134 13734
rect 12162 13706 12186 13734
rect 12214 13706 12238 13734
rect 12266 13706 12290 13734
rect 12318 13706 12342 13734
rect 12370 13706 12394 13734
rect 12422 13706 12446 13734
rect 12474 13706 12498 13734
rect 12526 13706 12531 13734
rect 17077 13706 17082 13734
rect 17110 13706 17134 13734
rect 17162 13706 17186 13734
rect 17214 13706 17238 13734
rect 17266 13706 17290 13734
rect 17318 13706 17342 13734
rect 17370 13706 17394 13734
rect 17422 13706 17446 13734
rect 17474 13706 17498 13734
rect 17526 13706 17531 13734
rect 22077 13706 22082 13734
rect 22110 13706 22134 13734
rect 22162 13706 22186 13734
rect 22214 13706 22238 13734
rect 22266 13706 22290 13734
rect 22318 13706 22342 13734
rect 22370 13706 22394 13734
rect 22422 13706 22446 13734
rect 22474 13706 22498 13734
rect 22526 13706 22531 13734
rect 27077 13706 27082 13734
rect 27110 13706 27134 13734
rect 27162 13706 27186 13734
rect 27214 13706 27238 13734
rect 27266 13706 27290 13734
rect 27318 13706 27342 13734
rect 27370 13706 27394 13734
rect 27422 13706 27446 13734
rect 27474 13706 27498 13734
rect 27526 13706 27531 13734
rect 32077 13706 32082 13734
rect 32110 13706 32134 13734
rect 32162 13706 32186 13734
rect 32214 13706 32238 13734
rect 32266 13706 32290 13734
rect 32318 13706 32342 13734
rect 32370 13706 32394 13734
rect 32422 13706 32446 13734
rect 32474 13706 32498 13734
rect 32526 13706 32531 13734
rect 37077 13706 37082 13734
rect 37110 13706 37134 13734
rect 37162 13706 37186 13734
rect 37214 13706 37238 13734
rect 37266 13706 37290 13734
rect 37318 13706 37342 13734
rect 37370 13706 37394 13734
rect 37422 13706 37446 13734
rect 37474 13706 37498 13734
rect 37526 13706 37531 13734
rect 5889 13510 5894 13538
rect 5922 13510 6454 13538
rect 6482 13510 6487 13538
rect 10425 13510 10430 13538
rect 10458 13510 10766 13538
rect 10794 13510 10799 13538
rect 12217 13510 12222 13538
rect 12250 13510 12950 13538
rect 12978 13510 13678 13538
rect 13706 13510 14406 13538
rect 14434 13510 14439 13538
rect 25377 13510 25382 13538
rect 25410 13510 25942 13538
rect 25970 13510 25975 13538
rect 26721 13510 26726 13538
rect 26754 13510 28462 13538
rect 28490 13510 28495 13538
rect 13785 13454 13790 13482
rect 13818 13454 14126 13482
rect 14154 13454 14159 13482
rect 16814 13454 17598 13482
rect 17626 13454 17631 13482
rect 23417 13454 23422 13482
rect 23450 13454 23926 13482
rect 23954 13454 27678 13482
rect 27706 13454 29358 13482
rect 29386 13454 29391 13482
rect 16809 13426 16814 13454
rect 16842 13426 16847 13454
rect 13225 13398 13230 13426
rect 13258 13398 13734 13426
rect 13762 13398 13767 13426
rect 18545 13398 18550 13426
rect 18578 13398 19054 13426
rect 19082 13398 19087 13426
rect 4577 13314 4582 13342
rect 4610 13314 4634 13342
rect 4662 13314 4686 13342
rect 4714 13314 4738 13342
rect 4766 13314 4790 13342
rect 4818 13314 4842 13342
rect 4870 13314 4894 13342
rect 4922 13314 4946 13342
rect 4974 13314 4998 13342
rect 5026 13314 5031 13342
rect 9577 13314 9582 13342
rect 9610 13314 9634 13342
rect 9662 13314 9686 13342
rect 9714 13314 9738 13342
rect 9766 13314 9790 13342
rect 9818 13314 9842 13342
rect 9870 13314 9894 13342
rect 9922 13314 9946 13342
rect 9974 13314 9998 13342
rect 10026 13314 10031 13342
rect 14577 13314 14582 13342
rect 14610 13314 14634 13342
rect 14662 13314 14686 13342
rect 14714 13314 14738 13342
rect 14766 13314 14790 13342
rect 14818 13314 14842 13342
rect 14870 13314 14894 13342
rect 14922 13314 14946 13342
rect 14974 13314 14998 13342
rect 15026 13314 15031 13342
rect 19577 13314 19582 13342
rect 19610 13314 19634 13342
rect 19662 13314 19686 13342
rect 19714 13314 19738 13342
rect 19766 13314 19790 13342
rect 19818 13314 19842 13342
rect 19870 13314 19894 13342
rect 19922 13314 19946 13342
rect 19974 13314 19998 13342
rect 20026 13314 20031 13342
rect 24577 13314 24582 13342
rect 24610 13314 24634 13342
rect 24662 13314 24686 13342
rect 24714 13314 24738 13342
rect 24766 13314 24790 13342
rect 24818 13314 24842 13342
rect 24870 13314 24894 13342
rect 24922 13314 24946 13342
rect 24974 13314 24998 13342
rect 25026 13314 25031 13342
rect 29577 13314 29582 13342
rect 29610 13314 29634 13342
rect 29662 13314 29686 13342
rect 29714 13314 29738 13342
rect 29766 13314 29790 13342
rect 29818 13314 29842 13342
rect 29870 13314 29894 13342
rect 29922 13314 29946 13342
rect 29974 13314 29998 13342
rect 30026 13314 30031 13342
rect 34577 13314 34582 13342
rect 34610 13314 34634 13342
rect 34662 13314 34686 13342
rect 34714 13314 34738 13342
rect 34766 13314 34790 13342
rect 34818 13314 34842 13342
rect 34870 13314 34894 13342
rect 34922 13314 34946 13342
rect 34974 13314 34998 13342
rect 35026 13314 35031 13342
rect 1969 13118 1974 13146
rect 2002 13118 2366 13146
rect 2394 13118 2399 13146
rect 15129 13118 15134 13146
rect 15162 13118 15470 13146
rect 15498 13118 15750 13146
rect 15778 13118 15783 13146
rect 17985 13118 17990 13146
rect 18018 13118 19446 13146
rect 19474 13118 19479 13146
rect 24481 13118 24486 13146
rect 24514 13118 25046 13146
rect 25074 13118 26502 13146
rect 26530 13118 26535 13146
rect 2077 12922 2082 12950
rect 2110 12922 2134 12950
rect 2162 12922 2186 12950
rect 2214 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2394 12950
rect 2422 12922 2446 12950
rect 2474 12922 2498 12950
rect 2526 12922 2531 12950
rect 7077 12922 7082 12950
rect 7110 12922 7134 12950
rect 7162 12922 7186 12950
rect 7214 12922 7238 12950
rect 7266 12922 7290 12950
rect 7318 12922 7342 12950
rect 7370 12922 7394 12950
rect 7422 12922 7446 12950
rect 7474 12922 7498 12950
rect 7526 12922 7531 12950
rect 12077 12922 12082 12950
rect 12110 12922 12134 12950
rect 12162 12922 12186 12950
rect 12214 12922 12238 12950
rect 12266 12922 12290 12950
rect 12318 12922 12342 12950
rect 12370 12922 12394 12950
rect 12422 12922 12446 12950
rect 12474 12922 12498 12950
rect 12526 12922 12531 12950
rect 17077 12922 17082 12950
rect 17110 12922 17134 12950
rect 17162 12922 17186 12950
rect 17214 12922 17238 12950
rect 17266 12922 17290 12950
rect 17318 12922 17342 12950
rect 17370 12922 17394 12950
rect 17422 12922 17446 12950
rect 17474 12922 17498 12950
rect 17526 12922 17531 12950
rect 22077 12922 22082 12950
rect 22110 12922 22134 12950
rect 22162 12922 22186 12950
rect 22214 12922 22238 12950
rect 22266 12922 22290 12950
rect 22318 12922 22342 12950
rect 22370 12922 22394 12950
rect 22422 12922 22446 12950
rect 22474 12922 22498 12950
rect 22526 12922 22531 12950
rect 27077 12922 27082 12950
rect 27110 12922 27134 12950
rect 27162 12922 27186 12950
rect 27214 12922 27238 12950
rect 27266 12922 27290 12950
rect 27318 12922 27342 12950
rect 27370 12922 27394 12950
rect 27422 12922 27446 12950
rect 27474 12922 27498 12950
rect 27526 12922 27531 12950
rect 32077 12922 32082 12950
rect 32110 12922 32134 12950
rect 32162 12922 32186 12950
rect 32214 12922 32238 12950
rect 32266 12922 32290 12950
rect 32318 12922 32342 12950
rect 32370 12922 32394 12950
rect 32422 12922 32446 12950
rect 32474 12922 32498 12950
rect 32526 12922 32531 12950
rect 37077 12922 37082 12950
rect 37110 12922 37134 12950
rect 37162 12922 37186 12950
rect 37214 12922 37238 12950
rect 37266 12922 37290 12950
rect 37318 12922 37342 12950
rect 37370 12922 37394 12950
rect 37422 12922 37446 12950
rect 37474 12922 37498 12950
rect 37526 12922 37531 12950
rect 2473 12726 2478 12754
rect 2506 12726 2758 12754
rect 2786 12726 2791 12754
rect 5553 12726 5558 12754
rect 5586 12726 6118 12754
rect 6146 12726 6151 12754
rect 11769 12726 11774 12754
rect 11802 12726 13230 12754
rect 13258 12726 13263 12754
rect 6449 12670 6454 12698
rect 6482 12670 7014 12698
rect 7042 12670 7047 12698
rect 19441 12670 19446 12698
rect 19474 12670 19950 12698
rect 19978 12670 19983 12698
rect 18769 12614 18774 12642
rect 18802 12614 20510 12642
rect 20538 12614 20958 12642
rect 20986 12614 22526 12642
rect 22554 12614 22559 12642
rect 28457 12614 28462 12642
rect 28490 12614 29022 12642
rect 29050 12614 30478 12642
rect 30506 12614 30511 12642
rect 4577 12530 4582 12558
rect 4610 12530 4634 12558
rect 4662 12530 4686 12558
rect 4714 12530 4738 12558
rect 4766 12530 4790 12558
rect 4818 12530 4842 12558
rect 4870 12530 4894 12558
rect 4922 12530 4946 12558
rect 4974 12530 4998 12558
rect 5026 12530 5031 12558
rect 9577 12530 9582 12558
rect 9610 12530 9634 12558
rect 9662 12530 9686 12558
rect 9714 12530 9738 12558
rect 9766 12530 9790 12558
rect 9818 12530 9842 12558
rect 9870 12530 9894 12558
rect 9922 12530 9946 12558
rect 9974 12530 9998 12558
rect 10026 12530 10031 12558
rect 14577 12530 14582 12558
rect 14610 12530 14634 12558
rect 14662 12530 14686 12558
rect 14714 12530 14738 12558
rect 14766 12530 14790 12558
rect 14818 12530 14842 12558
rect 14870 12530 14894 12558
rect 14922 12530 14946 12558
rect 14974 12530 14998 12558
rect 15026 12530 15031 12558
rect 19577 12530 19582 12558
rect 19610 12530 19634 12558
rect 19662 12530 19686 12558
rect 19714 12530 19738 12558
rect 19766 12530 19790 12558
rect 19818 12530 19842 12558
rect 19870 12530 19894 12558
rect 19922 12530 19946 12558
rect 19974 12530 19998 12558
rect 20026 12530 20031 12558
rect 24577 12530 24582 12558
rect 24610 12530 24634 12558
rect 24662 12530 24686 12558
rect 24714 12530 24738 12558
rect 24766 12530 24790 12558
rect 24818 12530 24842 12558
rect 24870 12530 24894 12558
rect 24922 12530 24946 12558
rect 24974 12530 24998 12558
rect 25026 12530 25031 12558
rect 29577 12530 29582 12558
rect 29610 12530 29634 12558
rect 29662 12530 29686 12558
rect 29714 12530 29738 12558
rect 29766 12530 29790 12558
rect 29818 12530 29842 12558
rect 29870 12530 29894 12558
rect 29922 12530 29946 12558
rect 29974 12530 29998 12558
rect 30026 12530 30031 12558
rect 34577 12530 34582 12558
rect 34610 12530 34634 12558
rect 34662 12530 34686 12558
rect 34714 12530 34738 12558
rect 34766 12530 34790 12558
rect 34818 12530 34842 12558
rect 34870 12530 34894 12558
rect 34922 12530 34946 12558
rect 34974 12530 34998 12558
rect 35026 12530 35031 12558
rect 7009 12390 7014 12418
rect 7042 12390 8358 12418
rect 8386 12390 8391 12418
rect 16025 12390 16030 12418
rect 16058 12390 16422 12418
rect 16450 12390 16455 12418
rect 6113 12334 6118 12362
rect 6146 12334 7574 12362
rect 7602 12334 7607 12362
rect 9529 12334 9534 12362
rect 9562 12334 10094 12362
rect 10122 12334 11270 12362
rect 11298 12334 11303 12362
rect 25993 12334 25998 12362
rect 26026 12334 26894 12362
rect 26922 12334 27174 12362
rect 27202 12334 27622 12362
rect 27650 12334 27655 12362
rect 29241 12334 29246 12362
rect 29274 12334 31094 12362
rect 31122 12334 31127 12362
rect 2077 12138 2082 12166
rect 2110 12138 2134 12166
rect 2162 12138 2186 12166
rect 2214 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2394 12166
rect 2422 12138 2446 12166
rect 2474 12138 2498 12166
rect 2526 12138 2531 12166
rect 7077 12138 7082 12166
rect 7110 12138 7134 12166
rect 7162 12138 7186 12166
rect 7214 12138 7238 12166
rect 7266 12138 7290 12166
rect 7318 12138 7342 12166
rect 7370 12138 7394 12166
rect 7422 12138 7446 12166
rect 7474 12138 7498 12166
rect 7526 12138 7531 12166
rect 12077 12138 12082 12166
rect 12110 12138 12134 12166
rect 12162 12138 12186 12166
rect 12214 12138 12238 12166
rect 12266 12138 12290 12166
rect 12318 12138 12342 12166
rect 12370 12138 12394 12166
rect 12422 12138 12446 12166
rect 12474 12138 12498 12166
rect 12526 12138 12531 12166
rect 17077 12138 17082 12166
rect 17110 12138 17134 12166
rect 17162 12138 17186 12166
rect 17214 12138 17238 12166
rect 17266 12138 17290 12166
rect 17318 12138 17342 12166
rect 17370 12138 17394 12166
rect 17422 12138 17446 12166
rect 17474 12138 17498 12166
rect 17526 12138 17531 12166
rect 22077 12138 22082 12166
rect 22110 12138 22134 12166
rect 22162 12138 22186 12166
rect 22214 12138 22238 12166
rect 22266 12138 22290 12166
rect 22318 12138 22342 12166
rect 22370 12138 22394 12166
rect 22422 12138 22446 12166
rect 22474 12138 22498 12166
rect 22526 12138 22531 12166
rect 27077 12138 27082 12166
rect 27110 12138 27134 12166
rect 27162 12138 27186 12166
rect 27214 12138 27238 12166
rect 27266 12138 27290 12166
rect 27318 12138 27342 12166
rect 27370 12138 27394 12166
rect 27422 12138 27446 12166
rect 27474 12138 27498 12166
rect 27526 12138 27531 12166
rect 32077 12138 32082 12166
rect 32110 12138 32134 12166
rect 32162 12138 32186 12166
rect 32214 12138 32238 12166
rect 32266 12138 32290 12166
rect 32318 12138 32342 12166
rect 32370 12138 32394 12166
rect 32422 12138 32446 12166
rect 32474 12138 32498 12166
rect 32526 12138 32531 12166
rect 37077 12138 37082 12166
rect 37110 12138 37134 12166
rect 37162 12138 37186 12166
rect 37214 12138 37238 12166
rect 37266 12138 37290 12166
rect 37318 12138 37342 12166
rect 37370 12138 37394 12166
rect 37422 12138 37446 12166
rect 37474 12138 37498 12166
rect 37526 12138 37531 12166
rect 27617 12054 27622 12082
rect 27650 12054 29246 12082
rect 29274 12054 29279 12082
rect 8969 11942 8974 11970
rect 9002 11942 9702 11970
rect 9730 11942 10374 11970
rect 10402 11942 10407 11970
rect 11265 11942 11270 11970
rect 11298 11942 11718 11970
rect 11746 11942 11751 11970
rect 15857 11942 15862 11970
rect 15890 11942 16926 11970
rect 16954 11942 16959 11970
rect 19945 11942 19950 11970
rect 19978 11942 20118 11970
rect 20146 11942 21182 11970
rect 21210 11942 21215 11970
rect 27001 11942 27006 11970
rect 27034 11942 28462 11970
rect 28490 11942 28495 11970
rect 31369 11942 31374 11970
rect 31402 11942 32830 11970
rect 32858 11942 33110 11970
rect 33138 11942 33143 11970
rect 23921 11886 23926 11914
rect 23954 11886 25158 11914
rect 25186 11886 25191 11914
rect 7569 11774 7574 11802
rect 7602 11774 8078 11802
rect 8106 11774 9478 11802
rect 9506 11774 9511 11802
rect 25153 11774 25158 11802
rect 25186 11774 25942 11802
rect 25970 11774 27678 11802
rect 27706 11774 27711 11802
rect 4577 11746 4582 11774
rect 4610 11746 4634 11774
rect 4662 11746 4686 11774
rect 4714 11746 4738 11774
rect 4766 11746 4790 11774
rect 4818 11746 4842 11774
rect 4870 11746 4894 11774
rect 4922 11746 4946 11774
rect 4974 11746 4998 11774
rect 5026 11746 5031 11774
rect 9577 11746 9582 11774
rect 9610 11746 9634 11774
rect 9662 11746 9686 11774
rect 9714 11746 9738 11774
rect 9766 11746 9790 11774
rect 9818 11746 9842 11774
rect 9870 11746 9894 11774
rect 9922 11746 9946 11774
rect 9974 11746 9998 11774
rect 10026 11746 10031 11774
rect 14577 11746 14582 11774
rect 14610 11746 14634 11774
rect 14662 11746 14686 11774
rect 14714 11746 14738 11774
rect 14766 11746 14790 11774
rect 14818 11746 14842 11774
rect 14870 11746 14894 11774
rect 14922 11746 14946 11774
rect 14974 11746 14998 11774
rect 15026 11746 15031 11774
rect 19577 11746 19582 11774
rect 19610 11746 19634 11774
rect 19662 11746 19686 11774
rect 19714 11746 19738 11774
rect 19766 11746 19790 11774
rect 19818 11746 19842 11774
rect 19870 11746 19894 11774
rect 19922 11746 19946 11774
rect 19974 11746 19998 11774
rect 20026 11746 20031 11774
rect 24577 11746 24582 11774
rect 24610 11746 24634 11774
rect 24662 11746 24686 11774
rect 24714 11746 24738 11774
rect 24766 11746 24790 11774
rect 24818 11746 24842 11774
rect 24870 11746 24894 11774
rect 24922 11746 24946 11774
rect 24974 11746 24998 11774
rect 25026 11746 25031 11774
rect 29577 11746 29582 11774
rect 29610 11746 29634 11774
rect 29662 11746 29686 11774
rect 29714 11746 29738 11774
rect 29766 11746 29790 11774
rect 29818 11746 29842 11774
rect 29870 11746 29894 11774
rect 29922 11746 29946 11774
rect 29974 11746 29998 11774
rect 30026 11746 30031 11774
rect 34577 11746 34582 11774
rect 34610 11746 34634 11774
rect 34662 11746 34686 11774
rect 34714 11746 34738 11774
rect 34766 11746 34790 11774
rect 34818 11746 34842 11774
rect 34870 11746 34894 11774
rect 34922 11746 34946 11774
rect 34974 11746 34998 11774
rect 35026 11746 35031 11774
rect 15073 11606 15078 11634
rect 15106 11606 16198 11634
rect 16226 11606 16758 11634
rect 16786 11606 16791 11634
rect 27393 11550 27398 11578
rect 27426 11550 27846 11578
rect 27874 11550 27879 11578
rect 30473 11550 30478 11578
rect 30506 11550 30982 11578
rect 31010 11550 31015 11578
rect 31985 11550 31990 11578
rect 32018 11550 32774 11578
rect 32802 11550 32807 11578
rect 29465 11494 29470 11522
rect 29498 11494 31374 11522
rect 31402 11494 35294 11522
rect 35322 11494 35327 11522
rect 29409 11382 29414 11410
rect 29442 11382 31934 11410
rect 31962 11382 31967 11410
rect 2077 11354 2082 11382
rect 2110 11354 2134 11382
rect 2162 11354 2186 11382
rect 2214 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2394 11382
rect 2422 11354 2446 11382
rect 2474 11354 2498 11382
rect 2526 11354 2531 11382
rect 7077 11354 7082 11382
rect 7110 11354 7134 11382
rect 7162 11354 7186 11382
rect 7214 11354 7238 11382
rect 7266 11354 7290 11382
rect 7318 11354 7342 11382
rect 7370 11354 7394 11382
rect 7422 11354 7446 11382
rect 7474 11354 7498 11382
rect 7526 11354 7531 11382
rect 12077 11354 12082 11382
rect 12110 11354 12134 11382
rect 12162 11354 12186 11382
rect 12214 11354 12238 11382
rect 12266 11354 12290 11382
rect 12318 11354 12342 11382
rect 12370 11354 12394 11382
rect 12422 11354 12446 11382
rect 12474 11354 12498 11382
rect 12526 11354 12531 11382
rect 17077 11354 17082 11382
rect 17110 11354 17134 11382
rect 17162 11354 17186 11382
rect 17214 11354 17238 11382
rect 17266 11354 17290 11382
rect 17318 11354 17342 11382
rect 17370 11354 17394 11382
rect 17422 11354 17446 11382
rect 17474 11354 17498 11382
rect 17526 11354 17531 11382
rect 22077 11354 22082 11382
rect 22110 11354 22134 11382
rect 22162 11354 22186 11382
rect 22214 11354 22238 11382
rect 22266 11354 22290 11382
rect 22318 11354 22342 11382
rect 22370 11354 22394 11382
rect 22422 11354 22446 11382
rect 22474 11354 22498 11382
rect 22526 11354 22531 11382
rect 27077 11354 27082 11382
rect 27110 11354 27134 11382
rect 27162 11354 27186 11382
rect 27214 11354 27238 11382
rect 27266 11354 27290 11382
rect 27318 11354 27342 11382
rect 27370 11354 27394 11382
rect 27422 11354 27446 11382
rect 27474 11354 27498 11382
rect 27526 11354 27531 11382
rect 32077 11354 32082 11382
rect 32110 11354 32134 11382
rect 32162 11354 32186 11382
rect 32214 11354 32238 11382
rect 32266 11354 32290 11382
rect 32318 11354 32342 11382
rect 32370 11354 32394 11382
rect 32422 11354 32446 11382
rect 32474 11354 32498 11382
rect 32526 11354 32531 11382
rect 37077 11354 37082 11382
rect 37110 11354 37134 11382
rect 37162 11354 37186 11382
rect 37214 11354 37238 11382
rect 37266 11354 37290 11382
rect 37318 11354 37342 11382
rect 37370 11354 37394 11382
rect 37422 11354 37446 11382
rect 37474 11354 37498 11382
rect 37526 11354 37531 11382
rect 18881 11214 18886 11242
rect 18914 11214 30702 11242
rect 30730 11214 31934 11242
rect 31962 11214 31967 11242
rect 13225 11158 13230 11186
rect 13258 11158 13510 11186
rect 13538 11158 13543 11186
rect 28457 11158 28462 11186
rect 28490 11158 29022 11186
rect 29050 11158 29055 11186
rect 30977 11158 30982 11186
rect 31010 11158 32438 11186
rect 32466 11158 32998 11186
rect 33026 11158 33031 11186
rect 34953 11158 34958 11186
rect 34986 11158 36134 11186
rect 36162 11158 36167 11186
rect 8465 11102 8470 11130
rect 8498 11102 8974 11130
rect 9002 11102 10374 11130
rect 10402 11102 10407 11130
rect 27673 11102 27678 11130
rect 27706 11102 28630 11130
rect 28658 11102 28854 11130
rect 28882 11102 31094 11130
rect 31122 11102 31127 11130
rect 33105 11102 33110 11130
rect 33138 11102 33894 11130
rect 33922 11102 33927 11130
rect 35289 11102 35294 11130
rect 35322 11102 35854 11130
rect 35882 11102 36694 11130
rect 36722 11102 36727 11130
rect 26945 11046 26950 11074
rect 26978 11046 27230 11074
rect 27258 11046 27454 11074
rect 27482 11046 29414 11074
rect 29442 11046 29447 11074
rect 4577 10962 4582 10990
rect 4610 10962 4634 10990
rect 4662 10962 4686 10990
rect 4714 10962 4738 10990
rect 4766 10962 4790 10990
rect 4818 10962 4842 10990
rect 4870 10962 4894 10990
rect 4922 10962 4946 10990
rect 4974 10962 4998 10990
rect 5026 10962 5031 10990
rect 9577 10962 9582 10990
rect 9610 10962 9634 10990
rect 9662 10962 9686 10990
rect 9714 10962 9738 10990
rect 9766 10962 9790 10990
rect 9818 10962 9842 10990
rect 9870 10962 9894 10990
rect 9922 10962 9946 10990
rect 9974 10962 9998 10990
rect 10026 10962 10031 10990
rect 14577 10962 14582 10990
rect 14610 10962 14634 10990
rect 14662 10962 14686 10990
rect 14714 10962 14738 10990
rect 14766 10962 14790 10990
rect 14818 10962 14842 10990
rect 14870 10962 14894 10990
rect 14922 10962 14946 10990
rect 14974 10962 14998 10990
rect 15026 10962 15031 10990
rect 19577 10962 19582 10990
rect 19610 10962 19634 10990
rect 19662 10962 19686 10990
rect 19714 10962 19738 10990
rect 19766 10962 19790 10990
rect 19818 10962 19842 10990
rect 19870 10962 19894 10990
rect 19922 10962 19946 10990
rect 19974 10962 19998 10990
rect 20026 10962 20031 10990
rect 24577 10962 24582 10990
rect 24610 10962 24634 10990
rect 24662 10962 24686 10990
rect 24714 10962 24738 10990
rect 24766 10962 24790 10990
rect 24818 10962 24842 10990
rect 24870 10962 24894 10990
rect 24922 10962 24946 10990
rect 24974 10962 24998 10990
rect 25026 10962 25031 10990
rect 29577 10962 29582 10990
rect 29610 10962 29634 10990
rect 29662 10962 29686 10990
rect 29714 10962 29738 10990
rect 29766 10962 29790 10990
rect 29818 10962 29842 10990
rect 29870 10962 29894 10990
rect 29922 10962 29946 10990
rect 29974 10962 29998 10990
rect 30026 10962 30031 10990
rect 34577 10962 34582 10990
rect 34610 10962 34634 10990
rect 34662 10962 34686 10990
rect 34714 10962 34738 10990
rect 34766 10962 34790 10990
rect 34818 10962 34842 10990
rect 34870 10962 34894 10990
rect 34922 10962 34946 10990
rect 34974 10962 34998 10990
rect 35026 10962 35031 10990
rect 22801 10878 22806 10906
rect 22834 10878 24374 10906
rect 24402 10878 24766 10906
rect 24794 10878 26222 10906
rect 26250 10878 26726 10906
rect 26754 10878 26759 10906
rect 27281 10766 27286 10794
rect 27314 10766 27566 10794
rect 27594 10766 27599 10794
rect 29913 10766 29918 10794
rect 29946 10766 30086 10794
rect 30114 10766 31374 10794
rect 31402 10766 31407 10794
rect 33889 10766 33894 10794
rect 33922 10766 35350 10794
rect 35378 10766 35383 10794
rect 17649 10710 17654 10738
rect 17682 10710 30254 10738
rect 30282 10710 30702 10738
rect 30730 10710 30735 10738
rect 2077 10570 2082 10598
rect 2110 10570 2134 10598
rect 2162 10570 2186 10598
rect 2214 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2394 10598
rect 2422 10570 2446 10598
rect 2474 10570 2498 10598
rect 2526 10570 2531 10598
rect 7077 10570 7082 10598
rect 7110 10570 7134 10598
rect 7162 10570 7186 10598
rect 7214 10570 7238 10598
rect 7266 10570 7290 10598
rect 7318 10570 7342 10598
rect 7370 10570 7394 10598
rect 7422 10570 7446 10598
rect 7474 10570 7498 10598
rect 7526 10570 7531 10598
rect 12077 10570 12082 10598
rect 12110 10570 12134 10598
rect 12162 10570 12186 10598
rect 12214 10570 12238 10598
rect 12266 10570 12290 10598
rect 12318 10570 12342 10598
rect 12370 10570 12394 10598
rect 12422 10570 12446 10598
rect 12474 10570 12498 10598
rect 12526 10570 12531 10598
rect 17077 10570 17082 10598
rect 17110 10570 17134 10598
rect 17162 10570 17186 10598
rect 17214 10570 17238 10598
rect 17266 10570 17290 10598
rect 17318 10570 17342 10598
rect 17370 10570 17394 10598
rect 17422 10570 17446 10598
rect 17474 10570 17498 10598
rect 17526 10570 17531 10598
rect 22077 10570 22082 10598
rect 22110 10570 22134 10598
rect 22162 10570 22186 10598
rect 22214 10570 22238 10598
rect 22266 10570 22290 10598
rect 22318 10570 22342 10598
rect 22370 10570 22394 10598
rect 22422 10570 22446 10598
rect 22474 10570 22498 10598
rect 22526 10570 22531 10598
rect 27077 10570 27082 10598
rect 27110 10570 27134 10598
rect 27162 10570 27186 10598
rect 27214 10570 27238 10598
rect 27266 10570 27290 10598
rect 27318 10570 27342 10598
rect 27370 10570 27394 10598
rect 27422 10570 27446 10598
rect 27474 10570 27498 10598
rect 27526 10570 27531 10598
rect 32077 10570 32082 10598
rect 32110 10570 32134 10598
rect 32162 10570 32186 10598
rect 32214 10570 32238 10598
rect 32266 10570 32290 10598
rect 32318 10570 32342 10598
rect 32370 10570 32394 10598
rect 32422 10570 32446 10598
rect 32474 10570 32498 10598
rect 32526 10570 32531 10598
rect 37077 10570 37082 10598
rect 37110 10570 37134 10598
rect 37162 10570 37186 10598
rect 37214 10570 37238 10598
rect 37266 10570 37290 10598
rect 37318 10570 37342 10598
rect 37370 10570 37394 10598
rect 37422 10570 37446 10598
rect 37474 10570 37498 10598
rect 37526 10570 37531 10598
rect 31929 10430 31934 10458
rect 31962 10430 32158 10458
rect 32186 10430 33614 10458
rect 33586 10402 33614 10430
rect 16361 10374 16366 10402
rect 16394 10374 17990 10402
rect 18018 10374 18023 10402
rect 26721 10374 26726 10402
rect 26754 10374 28406 10402
rect 28434 10374 28439 10402
rect 30697 10374 30702 10402
rect 30730 10374 32606 10402
rect 32634 10374 32639 10402
rect 33586 10374 36078 10402
rect 36106 10374 36111 10402
rect 18097 10318 18102 10346
rect 18130 10318 19502 10346
rect 19530 10318 19950 10346
rect 19978 10318 21406 10346
rect 21434 10318 21742 10346
rect 21770 10318 21775 10346
rect 25377 10318 25382 10346
rect 25410 10318 25942 10346
rect 25970 10318 25975 10346
rect 28625 10318 28630 10346
rect 28658 10318 29134 10346
rect 29162 10318 29167 10346
rect 4577 10178 4582 10206
rect 4610 10178 4634 10206
rect 4662 10178 4686 10206
rect 4714 10178 4738 10206
rect 4766 10178 4790 10206
rect 4818 10178 4842 10206
rect 4870 10178 4894 10206
rect 4922 10178 4946 10206
rect 4974 10178 4998 10206
rect 5026 10178 5031 10206
rect 9577 10178 9582 10206
rect 9610 10178 9634 10206
rect 9662 10178 9686 10206
rect 9714 10178 9738 10206
rect 9766 10178 9790 10206
rect 9818 10178 9842 10206
rect 9870 10178 9894 10206
rect 9922 10178 9946 10206
rect 9974 10178 9998 10206
rect 10026 10178 10031 10206
rect 14577 10178 14582 10206
rect 14610 10178 14634 10206
rect 14662 10178 14686 10206
rect 14714 10178 14738 10206
rect 14766 10178 14790 10206
rect 14818 10178 14842 10206
rect 14870 10178 14894 10206
rect 14922 10178 14946 10206
rect 14974 10178 14998 10206
rect 15026 10178 15031 10206
rect 19577 10178 19582 10206
rect 19610 10178 19634 10206
rect 19662 10178 19686 10206
rect 19714 10178 19738 10206
rect 19766 10178 19790 10206
rect 19818 10178 19842 10206
rect 19870 10178 19894 10206
rect 19922 10178 19946 10206
rect 19974 10178 19998 10206
rect 20026 10178 20031 10206
rect 24577 10178 24582 10206
rect 24610 10178 24634 10206
rect 24662 10178 24686 10206
rect 24714 10178 24738 10206
rect 24766 10178 24790 10206
rect 24818 10178 24842 10206
rect 24870 10178 24894 10206
rect 24922 10178 24946 10206
rect 24974 10178 24998 10206
rect 25026 10178 25031 10206
rect 29577 10178 29582 10206
rect 29610 10178 29634 10206
rect 29662 10178 29686 10206
rect 29714 10178 29738 10206
rect 29766 10178 29790 10206
rect 29818 10178 29842 10206
rect 29870 10178 29894 10206
rect 29922 10178 29946 10206
rect 29974 10178 29998 10206
rect 30026 10178 30031 10206
rect 34577 10178 34582 10206
rect 34610 10178 34634 10206
rect 34662 10178 34686 10206
rect 34714 10178 34738 10206
rect 34766 10178 34790 10206
rect 34818 10178 34842 10206
rect 34870 10178 34894 10206
rect 34922 10178 34946 10206
rect 34974 10178 34998 10206
rect 35026 10178 35031 10206
rect 20561 10094 20566 10122
rect 20594 10094 22806 10122
rect 22834 10094 22839 10122
rect 25937 10094 25942 10122
rect 25970 10094 27594 10122
rect 27566 10066 27594 10094
rect 27528 10038 27566 10066
rect 27594 10038 28966 10066
rect 28994 10038 28999 10066
rect 31089 10038 31094 10066
rect 31122 10038 31262 10066
rect 31290 10038 31295 10066
rect 31985 10038 31990 10066
rect 32018 10038 34230 10066
rect 34258 10038 34263 10066
rect 12441 9982 12446 10010
rect 12474 9982 12950 10010
rect 12978 9982 12983 10010
rect 18713 9982 18718 10010
rect 18746 9982 18942 10010
rect 18970 9982 18975 10010
rect 21737 9982 21742 10010
rect 21770 9982 22694 10010
rect 22722 9982 22918 10010
rect 22946 9982 23366 10010
rect 23394 9982 23399 10010
rect 27393 9982 27398 10010
rect 27426 9982 27902 10010
rect 27930 9982 27935 10010
rect 28569 9982 28574 10010
rect 28602 9982 29302 10010
rect 29330 9982 29335 10010
rect 5889 9926 5894 9954
rect 5922 9926 36190 9954
rect 36218 9926 36694 9954
rect 36722 9926 36727 9954
rect 2077 9786 2082 9814
rect 2110 9786 2134 9814
rect 2162 9786 2186 9814
rect 2214 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2394 9814
rect 2422 9786 2446 9814
rect 2474 9786 2498 9814
rect 2526 9786 2531 9814
rect 7077 9786 7082 9814
rect 7110 9786 7134 9814
rect 7162 9786 7186 9814
rect 7214 9786 7238 9814
rect 7266 9786 7290 9814
rect 7318 9786 7342 9814
rect 7370 9786 7394 9814
rect 7422 9786 7446 9814
rect 7474 9786 7498 9814
rect 7526 9786 7531 9814
rect 12077 9786 12082 9814
rect 12110 9786 12134 9814
rect 12162 9786 12186 9814
rect 12214 9786 12238 9814
rect 12266 9786 12290 9814
rect 12318 9786 12342 9814
rect 12370 9786 12394 9814
rect 12422 9786 12446 9814
rect 12474 9786 12498 9814
rect 12526 9786 12531 9814
rect 17077 9786 17082 9814
rect 17110 9786 17134 9814
rect 17162 9786 17186 9814
rect 17214 9786 17238 9814
rect 17266 9786 17290 9814
rect 17318 9786 17342 9814
rect 17370 9786 17394 9814
rect 17422 9786 17446 9814
rect 17474 9786 17498 9814
rect 17526 9786 17531 9814
rect 22077 9786 22082 9814
rect 22110 9786 22134 9814
rect 22162 9786 22186 9814
rect 22214 9786 22238 9814
rect 22266 9786 22290 9814
rect 22318 9786 22342 9814
rect 22370 9786 22394 9814
rect 22422 9786 22446 9814
rect 22474 9786 22498 9814
rect 22526 9786 22531 9814
rect 27077 9786 27082 9814
rect 27110 9786 27134 9814
rect 27162 9786 27186 9814
rect 27214 9786 27238 9814
rect 27266 9786 27290 9814
rect 27318 9786 27342 9814
rect 27370 9786 27394 9814
rect 27422 9786 27446 9814
rect 27474 9786 27498 9814
rect 27526 9786 27531 9814
rect 32077 9786 32082 9814
rect 32110 9786 32134 9814
rect 32162 9786 32186 9814
rect 32214 9786 32238 9814
rect 32266 9786 32290 9814
rect 32318 9786 32342 9814
rect 32370 9786 32394 9814
rect 32422 9786 32446 9814
rect 32474 9786 32498 9814
rect 32526 9786 32531 9814
rect 37077 9786 37082 9814
rect 37110 9786 37134 9814
rect 37162 9786 37186 9814
rect 37214 9786 37238 9814
rect 37266 9786 37290 9814
rect 37318 9786 37342 9814
rect 37370 9786 37394 9814
rect 37422 9786 37446 9814
rect 37474 9786 37498 9814
rect 37526 9786 37531 9814
rect 31033 9702 31038 9730
rect 31066 9702 31990 9730
rect 32018 9702 32023 9730
rect 11881 9646 11886 9674
rect 11914 9646 12054 9674
rect 12082 9646 13510 9674
rect 13538 9646 13543 9674
rect 18265 9590 18270 9618
rect 18298 9590 18718 9618
rect 18746 9590 19222 9618
rect 19250 9590 19255 9618
rect 23417 9590 23422 9618
rect 23450 9590 24654 9618
rect 24682 9590 24878 9618
rect 24906 9590 25158 9618
rect 25186 9590 25191 9618
rect 26945 9590 26950 9618
rect 26978 9590 27230 9618
rect 27258 9590 27454 9618
rect 27482 9590 28574 9618
rect 28602 9590 28607 9618
rect 28961 9590 28966 9618
rect 28994 9590 29414 9618
rect 29442 9590 31094 9618
rect 31122 9590 31374 9618
rect 31402 9590 32830 9618
rect 32858 9590 33110 9618
rect 33138 9590 33143 9618
rect 34449 9590 34454 9618
rect 34482 9590 34958 9618
rect 34986 9590 36358 9618
rect 36386 9590 36391 9618
rect 4993 9534 4998 9562
rect 5026 9534 6454 9562
rect 6482 9534 7014 9562
rect 7042 9534 7047 9562
rect 12945 9534 12950 9562
rect 12978 9534 14406 9562
rect 14434 9534 14439 9562
rect 27897 9534 27902 9562
rect 27930 9534 28406 9562
rect 28434 9534 28439 9562
rect 35345 9534 35350 9562
rect 35378 9534 35854 9562
rect 35882 9534 36862 9562
rect 36890 9534 36895 9562
rect 4577 9394 4582 9422
rect 4610 9394 4634 9422
rect 4662 9394 4686 9422
rect 4714 9394 4738 9422
rect 4766 9394 4790 9422
rect 4818 9394 4842 9422
rect 4870 9394 4894 9422
rect 4922 9394 4946 9422
rect 4974 9394 4998 9422
rect 5026 9394 5031 9422
rect 9577 9394 9582 9422
rect 9610 9394 9634 9422
rect 9662 9394 9686 9422
rect 9714 9394 9738 9422
rect 9766 9394 9790 9422
rect 9818 9394 9842 9422
rect 9870 9394 9894 9422
rect 9922 9394 9946 9422
rect 9974 9394 9998 9422
rect 10026 9394 10031 9422
rect 14577 9394 14582 9422
rect 14610 9394 14634 9422
rect 14662 9394 14686 9422
rect 14714 9394 14738 9422
rect 14766 9394 14790 9422
rect 14818 9394 14842 9422
rect 14870 9394 14894 9422
rect 14922 9394 14946 9422
rect 14974 9394 14998 9422
rect 15026 9394 15031 9422
rect 19577 9394 19582 9422
rect 19610 9394 19634 9422
rect 19662 9394 19686 9422
rect 19714 9394 19738 9422
rect 19766 9394 19790 9422
rect 19818 9394 19842 9422
rect 19870 9394 19894 9422
rect 19922 9394 19946 9422
rect 19974 9394 19998 9422
rect 20026 9394 20031 9422
rect 24577 9394 24582 9422
rect 24610 9394 24634 9422
rect 24662 9394 24686 9422
rect 24714 9394 24738 9422
rect 24766 9394 24790 9422
rect 24818 9394 24842 9422
rect 24870 9394 24894 9422
rect 24922 9394 24946 9422
rect 24974 9394 24998 9422
rect 25026 9394 25031 9422
rect 29577 9394 29582 9422
rect 29610 9394 29634 9422
rect 29662 9394 29686 9422
rect 29714 9394 29738 9422
rect 29766 9394 29790 9422
rect 29818 9394 29842 9422
rect 29870 9394 29894 9422
rect 29922 9394 29946 9422
rect 29974 9394 29998 9422
rect 30026 9394 30031 9422
rect 34577 9394 34582 9422
rect 34610 9394 34634 9422
rect 34662 9394 34686 9422
rect 34714 9394 34738 9422
rect 34766 9394 34790 9422
rect 34818 9394 34842 9422
rect 34870 9394 34894 9422
rect 34922 9394 34946 9422
rect 34974 9394 34998 9422
rect 35026 9394 35031 9422
rect 22745 9254 22750 9282
rect 22778 9254 24374 9282
rect 24402 9254 24766 9282
rect 24794 9254 24799 9282
rect 29409 9254 29414 9282
rect 29442 9254 29694 9282
rect 29722 9254 29727 9282
rect 33385 9254 33390 9282
rect 33418 9254 34622 9282
rect 34650 9254 34846 9282
rect 34874 9254 35070 9282
rect 35098 9254 35103 9282
rect 1577 9198 1582 9226
rect 1610 9198 1918 9226
rect 1946 9198 1951 9226
rect 2473 9198 2478 9226
rect 2506 9198 3038 9226
rect 3066 9198 4494 9226
rect 4522 9198 4527 9226
rect 9473 9198 9478 9226
rect 9506 9198 9814 9226
rect 9842 9198 9847 9226
rect 23417 9198 23422 9226
rect 23450 9198 23702 9226
rect 23730 9198 23735 9226
rect 24481 9198 24486 9226
rect 24514 9198 25102 9226
rect 25130 9198 26502 9226
rect 26530 9198 26535 9226
rect 28457 9198 28462 9226
rect 28490 9198 29022 9226
rect 29050 9198 30478 9226
rect 30506 9198 30511 9226
rect 32433 9198 32438 9226
rect 32466 9198 32942 9226
rect 32970 9198 32975 9226
rect 33586 9198 34174 9226
rect 34202 9198 34207 9226
rect 35625 9198 35630 9226
rect 35658 9198 35854 9226
rect 35882 9198 37310 9226
rect 37338 9198 37590 9226
rect 37618 9198 37623 9226
rect 33586 9170 33614 9198
rect 15521 9142 15526 9170
rect 15554 9142 17654 9170
rect 17682 9142 17687 9170
rect 18209 9142 18214 9170
rect 18242 9142 32774 9170
rect 32802 9142 33614 9170
rect 36129 9142 36134 9170
rect 36162 9142 36694 9170
rect 36722 9142 36727 9170
rect 25433 9086 25438 9114
rect 25466 9086 25998 9114
rect 26026 9086 26031 9114
rect 29073 9086 29078 9114
rect 29106 9086 30422 9114
rect 30450 9086 30982 9114
rect 31010 9086 31015 9114
rect 35233 9086 35238 9114
rect 35266 9086 36918 9114
rect 36946 9086 36951 9114
rect 2077 9002 2082 9030
rect 2110 9002 2134 9030
rect 2162 9002 2186 9030
rect 2214 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2394 9030
rect 2422 9002 2446 9030
rect 2474 9002 2498 9030
rect 2526 9002 2531 9030
rect 7077 9002 7082 9030
rect 7110 9002 7134 9030
rect 7162 9002 7186 9030
rect 7214 9002 7238 9030
rect 7266 9002 7290 9030
rect 7318 9002 7342 9030
rect 7370 9002 7394 9030
rect 7422 9002 7446 9030
rect 7474 9002 7498 9030
rect 7526 9002 7531 9030
rect 12077 9002 12082 9030
rect 12110 9002 12134 9030
rect 12162 9002 12186 9030
rect 12214 9002 12238 9030
rect 12266 9002 12290 9030
rect 12318 9002 12342 9030
rect 12370 9002 12394 9030
rect 12422 9002 12446 9030
rect 12474 9002 12498 9030
rect 12526 9002 12531 9030
rect 17077 9002 17082 9030
rect 17110 9002 17134 9030
rect 17162 9002 17186 9030
rect 17214 9002 17238 9030
rect 17266 9002 17290 9030
rect 17318 9002 17342 9030
rect 17370 9002 17394 9030
rect 17422 9002 17446 9030
rect 17474 9002 17498 9030
rect 17526 9002 17531 9030
rect 22077 9002 22082 9030
rect 22110 9002 22134 9030
rect 22162 9002 22186 9030
rect 22214 9002 22238 9030
rect 22266 9002 22290 9030
rect 22318 9002 22342 9030
rect 22370 9002 22394 9030
rect 22422 9002 22446 9030
rect 22474 9002 22498 9030
rect 22526 9002 22531 9030
rect 27077 9002 27082 9030
rect 27110 9002 27134 9030
rect 27162 9002 27186 9030
rect 27214 9002 27238 9030
rect 27266 9002 27290 9030
rect 27318 9002 27342 9030
rect 27370 9002 27394 9030
rect 27422 9002 27446 9030
rect 27474 9002 27498 9030
rect 27526 9002 27531 9030
rect 32077 9002 32082 9030
rect 32110 9002 32134 9030
rect 32162 9002 32186 9030
rect 32214 9002 32238 9030
rect 32266 9002 32290 9030
rect 32318 9002 32342 9030
rect 32370 9002 32394 9030
rect 32422 9002 32446 9030
rect 32474 9002 32498 9030
rect 32526 9002 32531 9030
rect 37077 9002 37082 9030
rect 37110 9002 37134 9030
rect 37162 9002 37186 9030
rect 37214 9002 37238 9030
rect 37266 9002 37290 9030
rect 37318 9002 37342 9030
rect 37370 9002 37394 9030
rect 37422 9002 37446 9030
rect 37474 9002 37498 9030
rect 37526 9002 37531 9030
rect 3705 8862 3710 8890
rect 3738 8862 31038 8890
rect 31066 8862 31071 8890
rect 1745 8806 1750 8834
rect 1778 8806 1974 8834
rect 2002 8806 2310 8834
rect 2338 8806 2343 8834
rect 4489 8806 4494 8834
rect 4522 8806 5950 8834
rect 5978 8806 6230 8834
rect 6258 8806 6790 8834
rect 6818 8806 6823 8834
rect 13505 8806 13510 8834
rect 13538 8806 14070 8834
rect 14098 8806 14103 8834
rect 17201 8806 17206 8834
rect 17234 8806 18774 8834
rect 18802 8806 18807 8834
rect 34953 8806 34958 8834
rect 34986 8806 36414 8834
rect 36442 8806 36447 8834
rect 34958 8778 34986 8806
rect 32993 8750 32998 8778
rect 33026 8750 34986 8778
rect 36857 8750 36862 8778
rect 36890 8750 37310 8778
rect 37338 8750 37646 8778
rect 37674 8750 37679 8778
rect 4577 8610 4582 8638
rect 4610 8610 4634 8638
rect 4662 8610 4686 8638
rect 4714 8610 4738 8638
rect 4766 8610 4790 8638
rect 4818 8610 4842 8638
rect 4870 8610 4894 8638
rect 4922 8610 4946 8638
rect 4974 8610 4998 8638
rect 5026 8610 5031 8638
rect 9577 8610 9582 8638
rect 9610 8610 9634 8638
rect 9662 8610 9686 8638
rect 9714 8610 9738 8638
rect 9766 8610 9790 8638
rect 9818 8610 9842 8638
rect 9870 8610 9894 8638
rect 9922 8610 9946 8638
rect 9974 8610 9998 8638
rect 10026 8610 10031 8638
rect 14577 8610 14582 8638
rect 14610 8610 14634 8638
rect 14662 8610 14686 8638
rect 14714 8610 14738 8638
rect 14766 8610 14790 8638
rect 14818 8610 14842 8638
rect 14870 8610 14894 8638
rect 14922 8610 14946 8638
rect 14974 8610 14998 8638
rect 15026 8610 15031 8638
rect 19577 8610 19582 8638
rect 19610 8610 19634 8638
rect 19662 8610 19686 8638
rect 19714 8610 19738 8638
rect 19766 8610 19790 8638
rect 19818 8610 19842 8638
rect 19870 8610 19894 8638
rect 19922 8610 19946 8638
rect 19974 8610 19998 8638
rect 20026 8610 20031 8638
rect 24577 8610 24582 8638
rect 24610 8610 24634 8638
rect 24662 8610 24686 8638
rect 24714 8610 24738 8638
rect 24766 8610 24790 8638
rect 24818 8610 24842 8638
rect 24870 8610 24894 8638
rect 24922 8610 24946 8638
rect 24974 8610 24998 8638
rect 25026 8610 25031 8638
rect 29577 8610 29582 8638
rect 29610 8610 29634 8638
rect 29662 8610 29686 8638
rect 29714 8610 29738 8638
rect 29766 8610 29790 8638
rect 29818 8610 29842 8638
rect 29870 8610 29894 8638
rect 29922 8610 29946 8638
rect 29974 8610 29998 8638
rect 30026 8610 30031 8638
rect 34577 8610 34582 8638
rect 34610 8610 34634 8638
rect 34662 8610 34686 8638
rect 34714 8610 34738 8638
rect 34766 8610 34790 8638
rect 34818 8610 34842 8638
rect 34870 8610 34894 8638
rect 34922 8610 34946 8638
rect 34974 8610 34998 8638
rect 35026 8610 35031 8638
rect 31929 8526 31934 8554
rect 31962 8526 32214 8554
rect 32242 8526 32247 8554
rect 2529 8470 2534 8498
rect 2562 8470 4214 8498
rect 4242 8470 4247 8498
rect 8353 8470 8358 8498
rect 8386 8470 10262 8498
rect 10290 8470 10295 8498
rect 29353 8470 29358 8498
rect 29386 8470 29918 8498
rect 29946 8470 33894 8498
rect 33922 8470 35238 8498
rect 35266 8470 35271 8498
rect 1913 8414 1918 8442
rect 1946 8414 2142 8442
rect 2170 8414 3598 8442
rect 3626 8414 3631 8442
rect 9249 8414 9254 8442
rect 9282 8414 9814 8442
rect 9842 8414 9847 8442
rect 11545 8414 11550 8442
rect 11578 8414 11998 8442
rect 12026 8414 12031 8442
rect 14401 8414 14406 8442
rect 14434 8414 14966 8442
rect 14994 8414 15694 8442
rect 15722 8414 15918 8442
rect 15946 8414 15951 8442
rect 23417 8414 23422 8442
rect 23450 8414 24878 8442
rect 24906 8414 25158 8442
rect 25186 8414 25438 8442
rect 25466 8414 26894 8442
rect 26922 8414 27174 8442
rect 27202 8414 27207 8442
rect 30977 8414 30982 8442
rect 31010 8414 32158 8442
rect 32186 8414 32191 8442
rect 32937 8414 32942 8442
rect 32970 8414 34398 8442
rect 34426 8414 34958 8442
rect 34986 8414 34991 8442
rect 11937 8358 11942 8386
rect 11970 8358 12222 8386
rect 12250 8358 12255 8386
rect 31369 8358 31374 8386
rect 31402 8358 31878 8386
rect 31906 8358 31911 8386
rect 2077 8218 2082 8246
rect 2110 8218 2134 8246
rect 2162 8218 2186 8246
rect 2214 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2394 8246
rect 2422 8218 2446 8246
rect 2474 8218 2498 8246
rect 2526 8218 2531 8246
rect 7077 8218 7082 8246
rect 7110 8218 7134 8246
rect 7162 8218 7186 8246
rect 7214 8218 7238 8246
rect 7266 8218 7290 8246
rect 7318 8218 7342 8246
rect 7370 8218 7394 8246
rect 7422 8218 7446 8246
rect 7474 8218 7498 8246
rect 7526 8218 7531 8246
rect 12077 8218 12082 8246
rect 12110 8218 12134 8246
rect 12162 8218 12186 8246
rect 12214 8218 12238 8246
rect 12266 8218 12290 8246
rect 12318 8218 12342 8246
rect 12370 8218 12394 8246
rect 12422 8218 12446 8246
rect 12474 8218 12498 8246
rect 12526 8218 12531 8246
rect 17077 8218 17082 8246
rect 17110 8218 17134 8246
rect 17162 8218 17186 8246
rect 17214 8218 17238 8246
rect 17266 8218 17290 8246
rect 17318 8218 17342 8246
rect 17370 8218 17394 8246
rect 17422 8218 17446 8246
rect 17474 8218 17498 8246
rect 17526 8218 17531 8246
rect 22077 8218 22082 8246
rect 22110 8218 22134 8246
rect 22162 8218 22186 8246
rect 22214 8218 22238 8246
rect 22266 8218 22290 8246
rect 22318 8218 22342 8246
rect 22370 8218 22394 8246
rect 22422 8218 22446 8246
rect 22474 8218 22498 8246
rect 22526 8218 22531 8246
rect 27077 8218 27082 8246
rect 27110 8218 27134 8246
rect 27162 8218 27186 8246
rect 27214 8218 27238 8246
rect 27266 8218 27290 8246
rect 27318 8218 27342 8246
rect 27370 8218 27394 8246
rect 27422 8218 27446 8246
rect 27474 8218 27498 8246
rect 27526 8218 27531 8246
rect 31990 8162 32018 8414
rect 32077 8218 32082 8246
rect 32110 8218 32134 8246
rect 32162 8218 32186 8246
rect 32214 8218 32238 8246
rect 32266 8218 32290 8246
rect 32318 8218 32342 8246
rect 32370 8218 32394 8246
rect 32422 8218 32446 8246
rect 32474 8218 32498 8246
rect 32526 8218 32531 8246
rect 37077 8218 37082 8246
rect 37110 8218 37134 8246
rect 37162 8218 37186 8246
rect 37214 8218 37238 8246
rect 37266 8218 37290 8246
rect 37318 8218 37342 8246
rect 37370 8218 37394 8246
rect 37422 8218 37446 8246
rect 37474 8218 37498 8246
rect 37526 8218 37531 8246
rect 31990 8134 32438 8162
rect 32466 8134 32471 8162
rect 2921 8078 2926 8106
rect 2954 8078 36134 8106
rect 36162 8078 36167 8106
rect 12049 8022 12054 8050
rect 12082 8022 13398 8050
rect 13426 8022 13431 8050
rect 28457 8022 28462 8050
rect 28490 8022 29022 8050
rect 29050 8022 29055 8050
rect 31873 8022 31878 8050
rect 31906 8022 33334 8050
rect 33362 8022 33367 8050
rect 1017 7966 1022 7994
rect 1050 7966 5894 7994
rect 5922 7966 5927 7994
rect 12441 7966 12446 7994
rect 12474 7966 14182 7994
rect 14210 7966 14215 7994
rect 4577 7826 4582 7854
rect 4610 7826 4634 7854
rect 4662 7826 4686 7854
rect 4714 7826 4738 7854
rect 4766 7826 4790 7854
rect 4818 7826 4842 7854
rect 4870 7826 4894 7854
rect 4922 7826 4946 7854
rect 4974 7826 4998 7854
rect 5026 7826 5031 7854
rect 9577 7826 9582 7854
rect 9610 7826 9634 7854
rect 9662 7826 9686 7854
rect 9714 7826 9738 7854
rect 9766 7826 9790 7854
rect 9818 7826 9842 7854
rect 9870 7826 9894 7854
rect 9922 7826 9946 7854
rect 9974 7826 9998 7854
rect 10026 7826 10031 7854
rect 14577 7826 14582 7854
rect 14610 7826 14634 7854
rect 14662 7826 14686 7854
rect 14714 7826 14738 7854
rect 14766 7826 14790 7854
rect 14818 7826 14842 7854
rect 14870 7826 14894 7854
rect 14922 7826 14946 7854
rect 14974 7826 14998 7854
rect 15026 7826 15031 7854
rect 19577 7826 19582 7854
rect 19610 7826 19634 7854
rect 19662 7826 19686 7854
rect 19714 7826 19738 7854
rect 19766 7826 19790 7854
rect 19818 7826 19842 7854
rect 19870 7826 19894 7854
rect 19922 7826 19946 7854
rect 19974 7826 19998 7854
rect 20026 7826 20031 7854
rect 24577 7826 24582 7854
rect 24610 7826 24634 7854
rect 24662 7826 24686 7854
rect 24714 7826 24738 7854
rect 24766 7826 24790 7854
rect 24818 7826 24842 7854
rect 24870 7826 24894 7854
rect 24922 7826 24946 7854
rect 24974 7826 24998 7854
rect 25026 7826 25031 7854
rect 29577 7826 29582 7854
rect 29610 7826 29634 7854
rect 29662 7826 29686 7854
rect 29714 7826 29738 7854
rect 29766 7826 29790 7854
rect 29818 7826 29842 7854
rect 29870 7826 29894 7854
rect 29922 7826 29946 7854
rect 29974 7826 29998 7854
rect 30026 7826 30031 7854
rect 34577 7826 34582 7854
rect 34610 7826 34634 7854
rect 34662 7826 34686 7854
rect 34714 7826 34738 7854
rect 34766 7826 34790 7854
rect 34818 7826 34842 7854
rect 34870 7826 34894 7854
rect 34922 7826 34946 7854
rect 34974 7826 34998 7854
rect 35026 7826 35031 7854
rect 33329 7686 33334 7714
rect 33362 7686 33838 7714
rect 33866 7686 33871 7714
rect 2585 7630 2590 7658
rect 2618 7630 3038 7658
rect 3066 7630 3071 7658
rect 6225 7630 6230 7658
rect 6258 7630 7014 7658
rect 7042 7630 7742 7658
rect 7770 7630 7966 7658
rect 7994 7630 8470 7658
rect 8498 7630 8503 7658
rect 9249 7630 9254 7658
rect 9282 7630 9814 7658
rect 9842 7630 9847 7658
rect 14065 7630 14070 7658
rect 14098 7630 15190 7658
rect 15218 7630 15223 7658
rect 16753 7630 16758 7658
rect 16786 7630 16870 7658
rect 16898 7630 16903 7658
rect 31985 7630 31990 7658
rect 32018 7630 32158 7658
rect 32186 7630 32326 7658
rect 32354 7630 32359 7658
rect 32433 7630 32438 7658
rect 32466 7630 32942 7658
rect 32970 7630 32975 7658
rect 32326 7602 32354 7630
rect 10318 7574 10878 7602
rect 10906 7574 11774 7602
rect 11802 7574 11942 7602
rect 11970 7574 12222 7602
rect 12250 7574 12255 7602
rect 32326 7574 33726 7602
rect 33754 7574 33759 7602
rect 10318 7546 10346 7574
rect 10201 7518 10206 7546
rect 10234 7518 10346 7546
rect 32097 7518 32102 7546
rect 32130 7518 32634 7546
rect 32881 7518 32886 7546
rect 32914 7518 34398 7546
rect 34426 7518 34431 7546
rect 32606 7490 32634 7518
rect 32601 7462 32606 7490
rect 32634 7462 33670 7490
rect 33698 7462 33703 7490
rect 2077 7434 2082 7462
rect 2110 7434 2134 7462
rect 2162 7434 2186 7462
rect 2214 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2394 7462
rect 2422 7434 2446 7462
rect 2474 7434 2498 7462
rect 2526 7434 2531 7462
rect 7077 7434 7082 7462
rect 7110 7434 7134 7462
rect 7162 7434 7186 7462
rect 7214 7434 7238 7462
rect 7266 7434 7290 7462
rect 7318 7434 7342 7462
rect 7370 7434 7394 7462
rect 7422 7434 7446 7462
rect 7474 7434 7498 7462
rect 7526 7434 7531 7462
rect 12077 7434 12082 7462
rect 12110 7434 12134 7462
rect 12162 7434 12186 7462
rect 12214 7434 12238 7462
rect 12266 7434 12290 7462
rect 12318 7434 12342 7462
rect 12370 7434 12394 7462
rect 12422 7434 12446 7462
rect 12474 7434 12498 7462
rect 12526 7434 12531 7462
rect 17077 7434 17082 7462
rect 17110 7434 17134 7462
rect 17162 7434 17186 7462
rect 17214 7434 17238 7462
rect 17266 7434 17290 7462
rect 17318 7434 17342 7462
rect 17370 7434 17394 7462
rect 17422 7434 17446 7462
rect 17474 7434 17498 7462
rect 17526 7434 17531 7462
rect 22077 7434 22082 7462
rect 22110 7434 22134 7462
rect 22162 7434 22186 7462
rect 22214 7434 22238 7462
rect 22266 7434 22290 7462
rect 22318 7434 22342 7462
rect 22370 7434 22394 7462
rect 22422 7434 22446 7462
rect 22474 7434 22498 7462
rect 22526 7434 22531 7462
rect 27077 7434 27082 7462
rect 27110 7434 27134 7462
rect 27162 7434 27186 7462
rect 27214 7434 27238 7462
rect 27266 7434 27290 7462
rect 27318 7434 27342 7462
rect 27370 7434 27394 7462
rect 27422 7434 27446 7462
rect 27474 7434 27498 7462
rect 27526 7434 27531 7462
rect 32077 7434 32082 7462
rect 32110 7434 32134 7462
rect 32162 7434 32186 7462
rect 32214 7434 32238 7462
rect 32266 7434 32290 7462
rect 32318 7434 32342 7462
rect 32370 7434 32394 7462
rect 32422 7434 32446 7462
rect 32474 7434 32498 7462
rect 32526 7434 32531 7462
rect 37077 7434 37082 7462
rect 37110 7434 37134 7462
rect 37162 7434 37186 7462
rect 37214 7434 37238 7462
rect 37266 7434 37290 7462
rect 37318 7434 37342 7462
rect 37370 7434 37394 7462
rect 37422 7434 37446 7462
rect 37474 7434 37498 7462
rect 37526 7434 37531 7462
rect 33889 7294 33894 7322
rect 33922 7294 35630 7322
rect 35658 7294 35663 7322
rect 1801 7238 1806 7266
rect 1834 7238 2030 7266
rect 2058 7238 2366 7266
rect 2394 7238 2399 7266
rect 25153 7238 25158 7266
rect 25186 7238 27174 7266
rect 27202 7238 27398 7266
rect 27426 7238 27431 7266
rect 31066 7238 32438 7266
rect 32466 7238 32471 7266
rect 32881 7238 32886 7266
rect 32914 7238 34678 7266
rect 34706 7238 34711 7266
rect 36073 7238 36078 7266
rect 36106 7238 36414 7266
rect 36442 7238 36694 7266
rect 36722 7238 36727 7266
rect 31066 7210 31094 7238
rect 27001 7182 27006 7210
rect 27034 7182 27678 7210
rect 27706 7182 31094 7210
rect 33721 7182 33726 7210
rect 33754 7182 33894 7210
rect 33922 7182 35742 7210
rect 35770 7182 35775 7210
rect 25377 7126 25382 7154
rect 25410 7126 32774 7154
rect 32802 7126 32807 7154
rect 33665 7126 33670 7154
rect 33698 7126 35518 7154
rect 35546 7126 35551 7154
rect 4577 7042 4582 7070
rect 4610 7042 4634 7070
rect 4662 7042 4686 7070
rect 4714 7042 4738 7070
rect 4766 7042 4790 7070
rect 4818 7042 4842 7070
rect 4870 7042 4894 7070
rect 4922 7042 4946 7070
rect 4974 7042 4998 7070
rect 5026 7042 5031 7070
rect 9577 7042 9582 7070
rect 9610 7042 9634 7070
rect 9662 7042 9686 7070
rect 9714 7042 9738 7070
rect 9766 7042 9790 7070
rect 9818 7042 9842 7070
rect 9870 7042 9894 7070
rect 9922 7042 9946 7070
rect 9974 7042 9998 7070
rect 10026 7042 10031 7070
rect 14577 7042 14582 7070
rect 14610 7042 14634 7070
rect 14662 7042 14686 7070
rect 14714 7042 14738 7070
rect 14766 7042 14790 7070
rect 14818 7042 14842 7070
rect 14870 7042 14894 7070
rect 14922 7042 14946 7070
rect 14974 7042 14998 7070
rect 15026 7042 15031 7070
rect 19577 7042 19582 7070
rect 19610 7042 19634 7070
rect 19662 7042 19686 7070
rect 19714 7042 19738 7070
rect 19766 7042 19790 7070
rect 19818 7042 19842 7070
rect 19870 7042 19894 7070
rect 19922 7042 19946 7070
rect 19974 7042 19998 7070
rect 20026 7042 20031 7070
rect 24577 7042 24582 7070
rect 24610 7042 24634 7070
rect 24662 7042 24686 7070
rect 24714 7042 24738 7070
rect 24766 7042 24790 7070
rect 24818 7042 24842 7070
rect 24870 7042 24894 7070
rect 24922 7042 24946 7070
rect 24974 7042 24998 7070
rect 25026 7042 25031 7070
rect 29577 7042 29582 7070
rect 29610 7042 29634 7070
rect 29662 7042 29686 7070
rect 29714 7042 29738 7070
rect 29766 7042 29790 7070
rect 29818 7042 29842 7070
rect 29870 7042 29894 7070
rect 29922 7042 29946 7070
rect 29974 7042 29998 7070
rect 30026 7042 30031 7070
rect 34577 7042 34582 7070
rect 34610 7042 34634 7070
rect 34662 7042 34686 7070
rect 34714 7042 34738 7070
rect 34766 7042 34790 7070
rect 34818 7042 34842 7070
rect 34870 7042 34894 7070
rect 34922 7042 34946 7070
rect 34974 7042 34998 7070
rect 35026 7042 35031 7070
rect 11769 6846 11774 6874
rect 11802 6846 11998 6874
rect 12026 6846 12222 6874
rect 12250 6846 12255 6874
rect 14289 6846 14294 6874
rect 14322 6846 14406 6874
rect 14434 6846 15078 6874
rect 15106 6846 16198 6874
rect 16226 6846 16422 6874
rect 16450 6846 17374 6874
rect 17402 6846 17407 6874
rect 25209 6846 25214 6874
rect 25242 6846 25438 6874
rect 25466 6846 25471 6874
rect 26721 6846 26726 6874
rect 26754 6846 28462 6874
rect 28490 6846 28742 6874
rect 28770 6846 28775 6874
rect 29465 6846 29470 6874
rect 29498 6846 30646 6874
rect 30674 6846 31094 6874
rect 34393 6846 34398 6874
rect 34426 6846 34678 6874
rect 34706 6846 34711 6874
rect 31066 6818 31094 6846
rect 3593 6790 3598 6818
rect 3626 6790 4102 6818
rect 4130 6790 5278 6818
rect 5306 6790 5311 6818
rect 29017 6790 29022 6818
rect 29050 6790 30478 6818
rect 30506 6790 30926 6818
rect 30954 6790 30959 6818
rect 31066 6790 31374 6818
rect 31402 6790 31878 6818
rect 31906 6790 33334 6818
rect 33362 6790 33950 6818
rect 33978 6790 35126 6818
rect 35154 6790 35350 6818
rect 35378 6790 35383 6818
rect 26889 6734 26894 6762
rect 26922 6734 28686 6762
rect 28714 6734 29190 6762
rect 29218 6734 29414 6762
rect 29442 6734 29447 6762
rect 30305 6734 30310 6762
rect 30338 6734 31990 6762
rect 32018 6734 32158 6762
rect 32186 6734 32191 6762
rect 32433 6734 32438 6762
rect 32466 6734 32998 6762
rect 33026 6734 34398 6762
rect 34426 6734 34431 6762
rect 35065 6734 35070 6762
rect 35098 6734 36134 6762
rect 36162 6734 36694 6762
rect 36722 6734 36727 6762
rect 33665 6678 33670 6706
rect 33698 6678 34006 6706
rect 34034 6678 34039 6706
rect 2077 6650 2082 6678
rect 2110 6650 2134 6678
rect 2162 6650 2186 6678
rect 2214 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2394 6678
rect 2422 6650 2446 6678
rect 2474 6650 2498 6678
rect 2526 6650 2531 6678
rect 7077 6650 7082 6678
rect 7110 6650 7134 6678
rect 7162 6650 7186 6678
rect 7214 6650 7238 6678
rect 7266 6650 7290 6678
rect 7318 6650 7342 6678
rect 7370 6650 7394 6678
rect 7422 6650 7446 6678
rect 7474 6650 7498 6678
rect 7526 6650 7531 6678
rect 12077 6650 12082 6678
rect 12110 6650 12134 6678
rect 12162 6650 12186 6678
rect 12214 6650 12238 6678
rect 12266 6650 12290 6678
rect 12318 6650 12342 6678
rect 12370 6650 12394 6678
rect 12422 6650 12446 6678
rect 12474 6650 12498 6678
rect 12526 6650 12531 6678
rect 17077 6650 17082 6678
rect 17110 6650 17134 6678
rect 17162 6650 17186 6678
rect 17214 6650 17238 6678
rect 17266 6650 17290 6678
rect 17318 6650 17342 6678
rect 17370 6650 17394 6678
rect 17422 6650 17446 6678
rect 17474 6650 17498 6678
rect 17526 6650 17531 6678
rect 22077 6650 22082 6678
rect 22110 6650 22134 6678
rect 22162 6650 22186 6678
rect 22214 6650 22238 6678
rect 22266 6650 22290 6678
rect 22318 6650 22342 6678
rect 22370 6650 22394 6678
rect 22422 6650 22446 6678
rect 22474 6650 22498 6678
rect 22526 6650 22531 6678
rect 27077 6650 27082 6678
rect 27110 6650 27134 6678
rect 27162 6650 27186 6678
rect 27214 6650 27238 6678
rect 27266 6650 27290 6678
rect 27318 6650 27342 6678
rect 27370 6650 27394 6678
rect 27422 6650 27446 6678
rect 27474 6650 27498 6678
rect 27526 6650 27531 6678
rect 32077 6650 32082 6678
rect 32110 6650 32134 6678
rect 32162 6650 32186 6678
rect 32214 6650 32238 6678
rect 32266 6650 32290 6678
rect 32318 6650 32342 6678
rect 32370 6650 32394 6678
rect 32422 6650 32446 6678
rect 32474 6650 32498 6678
rect 32526 6650 32531 6678
rect 37077 6650 37082 6678
rect 37110 6650 37134 6678
rect 37162 6650 37186 6678
rect 37214 6650 37238 6678
rect 37266 6650 37290 6678
rect 37318 6650 37342 6678
rect 37370 6650 37394 6678
rect 37422 6650 37446 6678
rect 37474 6650 37498 6678
rect 37526 6650 37531 6678
rect 10201 6454 10206 6482
rect 10234 6454 10318 6482
rect 10346 6454 10351 6482
rect 11993 6454 11998 6482
rect 12026 6454 12334 6482
rect 12362 6454 12367 6482
rect 24369 6454 24374 6482
rect 24402 6454 24766 6482
rect 24794 6454 24799 6482
rect 30977 6454 30982 6482
rect 31010 6454 32158 6482
rect 32186 6454 32718 6482
rect 32746 6454 32751 6482
rect 33721 6398 33726 6426
rect 33754 6398 33894 6426
rect 33922 6398 33927 6426
rect 23081 6342 23086 6370
rect 23114 6342 32886 6370
rect 32914 6342 32919 6370
rect 4577 6258 4582 6286
rect 4610 6258 4634 6286
rect 4662 6258 4686 6286
rect 4714 6258 4738 6286
rect 4766 6258 4790 6286
rect 4818 6258 4842 6286
rect 4870 6258 4894 6286
rect 4922 6258 4946 6286
rect 4974 6258 4998 6286
rect 5026 6258 5031 6286
rect 9577 6258 9582 6286
rect 9610 6258 9634 6286
rect 9662 6258 9686 6286
rect 9714 6258 9738 6286
rect 9766 6258 9790 6286
rect 9818 6258 9842 6286
rect 9870 6258 9894 6286
rect 9922 6258 9946 6286
rect 9974 6258 9998 6286
rect 10026 6258 10031 6286
rect 14577 6258 14582 6286
rect 14610 6258 14634 6286
rect 14662 6258 14686 6286
rect 14714 6258 14738 6286
rect 14766 6258 14790 6286
rect 14818 6258 14842 6286
rect 14870 6258 14894 6286
rect 14922 6258 14946 6286
rect 14974 6258 14998 6286
rect 15026 6258 15031 6286
rect 19577 6258 19582 6286
rect 19610 6258 19634 6286
rect 19662 6258 19686 6286
rect 19714 6258 19738 6286
rect 19766 6258 19790 6286
rect 19818 6258 19842 6286
rect 19870 6258 19894 6286
rect 19922 6258 19946 6286
rect 19974 6258 19998 6286
rect 20026 6258 20031 6286
rect 24577 6258 24582 6286
rect 24610 6258 24634 6286
rect 24662 6258 24686 6286
rect 24714 6258 24738 6286
rect 24766 6258 24790 6286
rect 24818 6258 24842 6286
rect 24870 6258 24894 6286
rect 24922 6258 24946 6286
rect 24974 6258 24998 6286
rect 25026 6258 25031 6286
rect 29577 6258 29582 6286
rect 29610 6258 29634 6286
rect 29662 6258 29686 6286
rect 29714 6258 29738 6286
rect 29766 6258 29790 6286
rect 29818 6258 29842 6286
rect 29870 6258 29894 6286
rect 29922 6258 29946 6286
rect 29974 6258 29998 6286
rect 30026 6258 30031 6286
rect 34577 6258 34582 6286
rect 34610 6258 34634 6286
rect 34662 6258 34686 6286
rect 34714 6258 34738 6286
rect 34766 6258 34790 6286
rect 34818 6258 34842 6286
rect 34870 6258 34894 6286
rect 34922 6258 34946 6286
rect 34974 6258 34998 6286
rect 35026 6258 35031 6286
rect 30081 6174 30086 6202
rect 30114 6174 31990 6202
rect 32018 6174 33614 6202
rect 33642 6174 33647 6202
rect 14457 6118 14462 6146
rect 14490 6118 14854 6146
rect 14882 6118 15694 6146
rect 15722 6118 15727 6146
rect 26889 6118 26894 6146
rect 26922 6118 27174 6146
rect 27202 6118 27207 6146
rect 29465 6118 29470 6146
rect 29498 6118 29918 6146
rect 29946 6118 31374 6146
rect 31402 6118 31407 6146
rect 2585 6062 2590 6090
rect 2618 6062 3038 6090
rect 3066 6062 3598 6090
rect 3626 6062 4102 6090
rect 4130 6062 4135 6090
rect 6449 6062 6454 6090
rect 6482 6062 7014 6090
rect 7042 6062 8358 6090
rect 8386 6062 8391 6090
rect 12441 6062 12446 6090
rect 12474 6062 12950 6090
rect 12978 6062 12983 6090
rect 13337 6062 13342 6090
rect 13370 6062 13510 6090
rect 13538 6062 13958 6090
rect 13986 6062 15190 6090
rect 15218 6062 15223 6090
rect 20785 6062 20790 6090
rect 20818 6062 22246 6090
rect 22274 6062 22582 6090
rect 22610 6062 22615 6090
rect 24369 6062 24374 6090
rect 24402 6062 24766 6090
rect 24794 6062 26222 6090
rect 26250 6062 26726 6090
rect 26754 6062 26759 6090
rect 31985 6062 31990 6090
rect 32018 6062 32158 6090
rect 32186 6062 32326 6090
rect 32354 6062 32359 6090
rect 21457 6006 21462 6034
rect 21490 6006 22694 6034
rect 22722 6006 22727 6034
rect 33614 5978 33642 6174
rect 26665 5950 26670 5978
rect 26698 5950 27734 5978
rect 33614 5950 35630 5978
rect 35658 5950 35663 5978
rect 2077 5866 2082 5894
rect 2110 5866 2134 5894
rect 2162 5866 2186 5894
rect 2214 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2394 5894
rect 2422 5866 2446 5894
rect 2474 5866 2498 5894
rect 2526 5866 2531 5894
rect 7077 5866 7082 5894
rect 7110 5866 7134 5894
rect 7162 5866 7186 5894
rect 7214 5866 7238 5894
rect 7266 5866 7290 5894
rect 7318 5866 7342 5894
rect 7370 5866 7394 5894
rect 7422 5866 7446 5894
rect 7474 5866 7498 5894
rect 7526 5866 7531 5894
rect 12077 5866 12082 5894
rect 12110 5866 12134 5894
rect 12162 5866 12186 5894
rect 12214 5866 12238 5894
rect 12266 5866 12290 5894
rect 12318 5866 12342 5894
rect 12370 5866 12394 5894
rect 12422 5866 12446 5894
rect 12474 5866 12498 5894
rect 12526 5866 12531 5894
rect 17077 5866 17082 5894
rect 17110 5866 17134 5894
rect 17162 5866 17186 5894
rect 17214 5866 17238 5894
rect 17266 5866 17290 5894
rect 17318 5866 17342 5894
rect 17370 5866 17394 5894
rect 17422 5866 17446 5894
rect 17474 5866 17498 5894
rect 17526 5866 17531 5894
rect 22077 5866 22082 5894
rect 22110 5866 22134 5894
rect 22162 5866 22186 5894
rect 22214 5866 22238 5894
rect 22266 5866 22290 5894
rect 22318 5866 22342 5894
rect 22370 5866 22394 5894
rect 22422 5866 22446 5894
rect 22474 5866 22498 5894
rect 22526 5866 22531 5894
rect 27077 5866 27082 5894
rect 27110 5866 27134 5894
rect 27162 5866 27186 5894
rect 27214 5866 27238 5894
rect 27266 5866 27290 5894
rect 27318 5866 27342 5894
rect 27370 5866 27394 5894
rect 27422 5866 27446 5894
rect 27474 5866 27498 5894
rect 27526 5866 27531 5894
rect 27706 5866 27734 5950
rect 33329 5894 33334 5922
rect 33362 5894 33670 5922
rect 33698 5894 35126 5922
rect 35154 5894 35159 5922
rect 32077 5866 32082 5894
rect 32110 5866 32134 5894
rect 32162 5866 32186 5894
rect 32214 5866 32238 5894
rect 32266 5866 32290 5894
rect 32318 5866 32342 5894
rect 32370 5866 32394 5894
rect 32422 5866 32446 5894
rect 32474 5866 32498 5894
rect 32526 5866 32531 5894
rect 37077 5866 37082 5894
rect 37110 5866 37134 5894
rect 37162 5866 37186 5894
rect 37214 5866 37238 5894
rect 37266 5866 37290 5894
rect 37318 5866 37342 5894
rect 37370 5866 37394 5894
rect 37422 5866 37446 5894
rect 37474 5866 37498 5894
rect 37526 5866 37531 5894
rect 7569 5838 7574 5866
rect 7602 5838 8078 5866
rect 8106 5838 8111 5866
rect 16417 5838 16422 5866
rect 16450 5838 16814 5866
rect 16842 5838 16847 5866
rect 27706 5838 28742 5866
rect 28770 5838 28775 5866
rect 33273 5838 33278 5866
rect 33306 5838 33614 5866
rect 33642 5838 33782 5866
rect 33810 5838 33815 5866
rect 28065 5782 28070 5810
rect 28098 5782 30142 5810
rect 30170 5782 31934 5810
rect 31962 5782 33054 5810
rect 33082 5782 33087 5810
rect 4993 5670 4998 5698
rect 5026 5670 5838 5698
rect 5866 5670 5871 5698
rect 30921 5670 30926 5698
rect 30954 5670 32158 5698
rect 32186 5670 32662 5698
rect 32690 5670 32695 5698
rect 35961 5670 35966 5698
rect 35994 5670 37142 5698
rect 37170 5670 37175 5698
rect 31985 5614 31990 5642
rect 32018 5614 33726 5642
rect 33754 5614 33894 5642
rect 33922 5614 33927 5642
rect 4577 5474 4582 5502
rect 4610 5474 4634 5502
rect 4662 5474 4686 5502
rect 4714 5474 4738 5502
rect 4766 5474 4790 5502
rect 4818 5474 4842 5502
rect 4870 5474 4894 5502
rect 4922 5474 4946 5502
rect 4974 5474 4998 5502
rect 5026 5474 5031 5502
rect 9577 5474 9582 5502
rect 9610 5474 9634 5502
rect 9662 5474 9686 5502
rect 9714 5474 9738 5502
rect 9766 5474 9790 5502
rect 9818 5474 9842 5502
rect 9870 5474 9894 5502
rect 9922 5474 9946 5502
rect 9974 5474 9998 5502
rect 10026 5474 10031 5502
rect 14577 5474 14582 5502
rect 14610 5474 14634 5502
rect 14662 5474 14686 5502
rect 14714 5474 14738 5502
rect 14766 5474 14790 5502
rect 14818 5474 14842 5502
rect 14870 5474 14894 5502
rect 14922 5474 14946 5502
rect 14974 5474 14998 5502
rect 15026 5474 15031 5502
rect 19577 5474 19582 5502
rect 19610 5474 19634 5502
rect 19662 5474 19686 5502
rect 19714 5474 19738 5502
rect 19766 5474 19790 5502
rect 19818 5474 19842 5502
rect 19870 5474 19894 5502
rect 19922 5474 19946 5502
rect 19974 5474 19998 5502
rect 20026 5474 20031 5502
rect 24577 5474 24582 5502
rect 24610 5474 24634 5502
rect 24662 5474 24686 5502
rect 24714 5474 24738 5502
rect 24766 5474 24790 5502
rect 24818 5474 24842 5502
rect 24870 5474 24894 5502
rect 24922 5474 24946 5502
rect 24974 5474 24998 5502
rect 25026 5474 25031 5502
rect 29577 5474 29582 5502
rect 29610 5474 29634 5502
rect 29662 5474 29686 5502
rect 29714 5474 29738 5502
rect 29766 5474 29790 5502
rect 29818 5474 29842 5502
rect 29870 5474 29894 5502
rect 29922 5474 29946 5502
rect 29974 5474 29998 5502
rect 30026 5474 30031 5502
rect 34577 5474 34582 5502
rect 34610 5474 34634 5502
rect 34662 5474 34686 5502
rect 34714 5474 34738 5502
rect 34766 5474 34790 5502
rect 34818 5474 34842 5502
rect 34870 5474 34894 5502
rect 34922 5474 34946 5502
rect 34974 5474 34998 5502
rect 35026 5474 35031 5502
rect 16977 5334 16982 5362
rect 17010 5334 21854 5362
rect 24425 5334 24430 5362
rect 24458 5334 28070 5362
rect 28098 5334 28103 5362
rect 33329 5334 33334 5362
rect 33362 5334 33614 5362
rect 33642 5334 35266 5362
rect 21826 5306 21854 5334
rect 35238 5306 35266 5334
rect 6113 5278 6118 5306
rect 6146 5278 7294 5306
rect 7322 5278 8078 5306
rect 8106 5278 8111 5306
rect 12441 5278 12446 5306
rect 12474 5278 12950 5306
rect 12978 5278 12983 5306
rect 14177 5278 14182 5306
rect 14210 5278 14462 5306
rect 14490 5278 14495 5306
rect 20225 5278 20230 5306
rect 20258 5278 20790 5306
rect 20818 5278 20823 5306
rect 21826 5278 26054 5306
rect 26082 5278 26087 5306
rect 28009 5278 28014 5306
rect 28042 5278 28182 5306
rect 28210 5278 28406 5306
rect 28434 5278 30142 5306
rect 30170 5278 30254 5306
rect 30282 5278 31934 5306
rect 31962 5278 31990 5306
rect 32018 5278 32158 5306
rect 32186 5278 32326 5306
rect 32354 5278 32359 5306
rect 32769 5278 32774 5306
rect 32802 5278 34174 5306
rect 34202 5278 34207 5306
rect 35233 5278 35238 5306
rect 35266 5278 35966 5306
rect 35994 5278 35999 5306
rect 25937 5222 25942 5250
rect 25970 5222 26782 5250
rect 26810 5222 26815 5250
rect 33889 5222 33894 5250
rect 33922 5222 35742 5250
rect 35770 5222 35910 5250
rect 35938 5222 37702 5250
rect 37730 5222 38262 5250
rect 38290 5222 38430 5250
rect 38458 5222 38598 5250
rect 38626 5222 38631 5250
rect 26049 5166 26054 5194
rect 26082 5166 28014 5194
rect 28042 5166 28047 5194
rect 2077 5082 2082 5110
rect 2110 5082 2134 5110
rect 2162 5082 2186 5110
rect 2214 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2394 5110
rect 2422 5082 2446 5110
rect 2474 5082 2498 5110
rect 2526 5082 2531 5110
rect 7077 5082 7082 5110
rect 7110 5082 7134 5110
rect 7162 5082 7186 5110
rect 7214 5082 7238 5110
rect 7266 5082 7290 5110
rect 7318 5082 7342 5110
rect 7370 5082 7394 5110
rect 7422 5082 7446 5110
rect 7474 5082 7498 5110
rect 7526 5082 7531 5110
rect 12077 5082 12082 5110
rect 12110 5082 12134 5110
rect 12162 5082 12186 5110
rect 12214 5082 12238 5110
rect 12266 5082 12290 5110
rect 12318 5082 12342 5110
rect 12370 5082 12394 5110
rect 12422 5082 12446 5110
rect 12474 5082 12498 5110
rect 12526 5082 12531 5110
rect 17077 5082 17082 5110
rect 17110 5082 17134 5110
rect 17162 5082 17186 5110
rect 17214 5082 17238 5110
rect 17266 5082 17290 5110
rect 17318 5082 17342 5110
rect 17370 5082 17394 5110
rect 17422 5082 17446 5110
rect 17474 5082 17498 5110
rect 17526 5082 17531 5110
rect 22077 5082 22082 5110
rect 22110 5082 22134 5110
rect 22162 5082 22186 5110
rect 22214 5082 22238 5110
rect 22266 5082 22290 5110
rect 22318 5082 22342 5110
rect 22370 5082 22394 5110
rect 22422 5082 22446 5110
rect 22474 5082 22498 5110
rect 22526 5082 22531 5110
rect 27077 5082 27082 5110
rect 27110 5082 27134 5110
rect 27162 5082 27186 5110
rect 27214 5082 27238 5110
rect 27266 5082 27290 5110
rect 27318 5082 27342 5110
rect 27370 5082 27394 5110
rect 27422 5082 27446 5110
rect 27474 5082 27498 5110
rect 27526 5082 27531 5110
rect 32077 5082 32082 5110
rect 32110 5082 32134 5110
rect 32162 5082 32186 5110
rect 32214 5082 32238 5110
rect 32266 5082 32290 5110
rect 32318 5082 32342 5110
rect 32370 5082 32394 5110
rect 32422 5082 32446 5110
rect 32474 5082 32498 5110
rect 32526 5082 32531 5110
rect 37077 5082 37082 5110
rect 37110 5082 37134 5110
rect 37162 5082 37186 5110
rect 37214 5082 37238 5110
rect 37266 5082 37290 5110
rect 37318 5082 37342 5110
rect 37370 5082 37394 5110
rect 37422 5082 37446 5110
rect 37474 5082 37498 5110
rect 37526 5082 37531 5110
rect 4489 5054 4494 5082
rect 4522 5054 4998 5082
rect 5026 5054 5950 5082
rect 5978 5054 5983 5082
rect 18769 5054 18774 5082
rect 18802 5054 20230 5082
rect 20258 5054 20263 5082
rect 33833 5054 33838 5082
rect 33866 5054 34510 5082
rect 34538 5054 34543 5082
rect 27706 4942 32942 4970
rect 32970 4942 36134 4970
rect 36162 4942 36694 4970
rect 36722 4942 36727 4970
rect 36857 4942 36862 4970
rect 36890 4942 37310 4970
rect 37338 4942 37646 4970
rect 37674 4942 37679 4970
rect 6449 4886 6454 4914
rect 6482 4886 6790 4914
rect 6818 4886 6823 4914
rect 12945 4830 12950 4858
rect 12978 4830 14182 4858
rect 14210 4830 14215 4858
rect 4577 4690 4582 4718
rect 4610 4690 4634 4718
rect 4662 4690 4686 4718
rect 4714 4690 4738 4718
rect 4766 4690 4790 4718
rect 4818 4690 4842 4718
rect 4870 4690 4894 4718
rect 4922 4690 4946 4718
rect 4974 4690 4998 4718
rect 5026 4690 5031 4718
rect 9577 4690 9582 4718
rect 9610 4690 9634 4718
rect 9662 4690 9686 4718
rect 9714 4690 9738 4718
rect 9766 4690 9790 4718
rect 9818 4690 9842 4718
rect 9870 4690 9894 4718
rect 9922 4690 9946 4718
rect 9974 4690 9998 4718
rect 10026 4690 10031 4718
rect 14577 4690 14582 4718
rect 14610 4690 14634 4718
rect 14662 4690 14686 4718
rect 14714 4690 14738 4718
rect 14766 4690 14790 4718
rect 14818 4690 14842 4718
rect 14870 4690 14894 4718
rect 14922 4690 14946 4718
rect 14974 4690 14998 4718
rect 15026 4690 15031 4718
rect 19577 4690 19582 4718
rect 19610 4690 19634 4718
rect 19662 4690 19686 4718
rect 19714 4690 19738 4718
rect 19766 4690 19790 4718
rect 19818 4690 19842 4718
rect 19870 4690 19894 4718
rect 19922 4690 19946 4718
rect 19974 4690 19998 4718
rect 20026 4690 20031 4718
rect 24577 4690 24582 4718
rect 24610 4690 24634 4718
rect 24662 4690 24686 4718
rect 24714 4690 24738 4718
rect 24766 4690 24790 4718
rect 24818 4690 24842 4718
rect 24870 4690 24894 4718
rect 24922 4690 24946 4718
rect 24974 4690 24998 4718
rect 25026 4690 25031 4718
rect 15806 4662 18214 4690
rect 18242 4662 18247 4690
rect 15806 4634 15834 4662
rect 27706 4634 27734 4942
rect 30193 4886 30198 4914
rect 30226 4886 30310 4914
rect 30338 4886 30343 4914
rect 31985 4886 31990 4914
rect 32018 4886 32158 4914
rect 32186 4886 32191 4914
rect 34169 4886 34174 4914
rect 34202 4886 34678 4914
rect 34706 4886 34711 4914
rect 35681 4886 35686 4914
rect 35714 4886 36078 4914
rect 36106 4886 37590 4914
rect 37618 4886 38150 4914
rect 38178 4886 38878 4914
rect 38906 4886 38911 4914
rect 29577 4690 29582 4718
rect 29610 4690 29634 4718
rect 29662 4690 29686 4718
rect 29714 4690 29738 4718
rect 29766 4690 29790 4718
rect 29818 4690 29842 4718
rect 29870 4690 29894 4718
rect 29922 4690 29946 4718
rect 29974 4690 29998 4718
rect 30026 4690 30031 4718
rect 34577 4690 34582 4718
rect 34610 4690 34634 4718
rect 34662 4690 34686 4718
rect 34714 4690 34738 4718
rect 34766 4690 34790 4718
rect 34818 4690 34842 4718
rect 34870 4690 34894 4718
rect 34922 4690 34946 4718
rect 34974 4690 34998 4718
rect 35026 4690 35031 4718
rect 12665 4606 12670 4634
rect 12698 4606 15834 4634
rect 17985 4606 17990 4634
rect 18018 4606 27734 4634
rect 30086 4662 32606 4690
rect 32634 4662 32639 4690
rect 30086 4522 30114 4662
rect 37865 4550 37870 4578
rect 37898 4550 38262 4578
rect 38290 4550 38430 4578
rect 38458 4550 38463 4578
rect 4489 4494 4494 4522
rect 4522 4494 4774 4522
rect 4802 4494 6790 4522
rect 6818 4494 7014 4522
rect 7042 4494 7047 4522
rect 8465 4494 8470 4522
rect 8498 4494 8974 4522
rect 9002 4494 9007 4522
rect 12441 4494 12446 4522
rect 12474 4494 12726 4522
rect 12754 4494 12759 4522
rect 15465 4494 15470 4522
rect 15498 4494 15694 4522
rect 15722 4494 15727 4522
rect 21401 4494 21406 4522
rect 21434 4494 21798 4522
rect 21826 4494 22694 4522
rect 22722 4494 22918 4522
rect 22946 4494 23198 4522
rect 23226 4494 23231 4522
rect 26329 4494 26334 4522
rect 26362 4494 28126 4522
rect 28154 4494 30114 4522
rect 34169 4494 34174 4522
rect 34202 4494 34678 4522
rect 34706 4494 34711 4522
rect 35681 4438 35686 4466
rect 35714 4438 37590 4466
rect 37618 4438 37623 4466
rect 35065 4382 35070 4410
rect 35098 4382 37646 4410
rect 37674 4382 37679 4410
rect 2077 4298 2082 4326
rect 2110 4298 2134 4326
rect 2162 4298 2186 4326
rect 2214 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2394 4326
rect 2422 4298 2446 4326
rect 2474 4298 2498 4326
rect 2526 4298 2531 4326
rect 7077 4298 7082 4326
rect 7110 4298 7134 4326
rect 7162 4298 7186 4326
rect 7214 4298 7238 4326
rect 7266 4298 7290 4326
rect 7318 4298 7342 4326
rect 7370 4298 7394 4326
rect 7422 4298 7446 4326
rect 7474 4298 7498 4326
rect 7526 4298 7531 4326
rect 12077 4298 12082 4326
rect 12110 4298 12134 4326
rect 12162 4298 12186 4326
rect 12214 4298 12238 4326
rect 12266 4298 12290 4326
rect 12318 4298 12342 4326
rect 12370 4298 12394 4326
rect 12422 4298 12446 4326
rect 12474 4298 12498 4326
rect 12526 4298 12531 4326
rect 17077 4298 17082 4326
rect 17110 4298 17134 4326
rect 17162 4298 17186 4326
rect 17214 4298 17238 4326
rect 17266 4298 17290 4326
rect 17318 4298 17342 4326
rect 17370 4298 17394 4326
rect 17422 4298 17446 4326
rect 17474 4298 17498 4326
rect 17526 4298 17531 4326
rect 22077 4298 22082 4326
rect 22110 4298 22134 4326
rect 22162 4298 22186 4326
rect 22214 4298 22238 4326
rect 22266 4298 22290 4326
rect 22318 4298 22342 4326
rect 22370 4298 22394 4326
rect 22422 4298 22446 4326
rect 22474 4298 22498 4326
rect 22526 4298 22531 4326
rect 27077 4298 27082 4326
rect 27110 4298 27134 4326
rect 27162 4298 27186 4326
rect 27214 4298 27238 4326
rect 27266 4298 27290 4326
rect 27318 4298 27342 4326
rect 27370 4298 27394 4326
rect 27422 4298 27446 4326
rect 27474 4298 27498 4326
rect 27526 4298 27531 4326
rect 32077 4298 32082 4326
rect 32110 4298 32134 4326
rect 32162 4298 32186 4326
rect 32214 4298 32238 4326
rect 32266 4298 32290 4326
rect 32318 4298 32342 4326
rect 32370 4298 32394 4326
rect 32422 4298 32446 4326
rect 32474 4298 32498 4326
rect 32526 4298 32531 4326
rect 37077 4298 37082 4326
rect 37110 4298 37134 4326
rect 37162 4298 37186 4326
rect 37214 4298 37238 4326
rect 37266 4298 37290 4326
rect 37318 4298 37342 4326
rect 37370 4298 37394 4326
rect 37422 4298 37446 4326
rect 37474 4298 37498 4326
rect 37526 4298 37531 4326
rect 3537 4214 3542 4242
rect 3570 4214 3710 4242
rect 3738 4214 3743 4242
rect 2585 4158 2590 4186
rect 2618 4158 3038 4186
rect 3066 4158 3071 4186
rect 7009 4158 7014 4186
rect 7042 4158 8470 4186
rect 8498 4158 8503 4186
rect 20113 4158 20118 4186
rect 20146 4158 21350 4186
rect 21378 4158 21686 4186
rect 21714 4158 21719 4186
rect 3593 4102 3598 4130
rect 3626 4102 4102 4130
rect 4130 4102 5278 4130
rect 5306 4102 5311 4130
rect 5945 4102 5950 4130
rect 5978 4102 6454 4130
rect 6482 4102 6487 4130
rect 9417 4102 9422 4130
rect 9450 4102 9534 4130
rect 9562 4102 10038 4130
rect 10066 4102 10071 4130
rect 22745 4102 22750 4130
rect 22778 4102 24374 4130
rect 24402 4102 24766 4130
rect 24794 4102 24799 4130
rect 27393 4102 27398 4130
rect 27426 4102 27678 4130
rect 27706 4102 27711 4130
rect 31313 4102 31318 4130
rect 31346 4102 34846 4130
rect 34874 4102 35182 4130
rect 35210 4102 35350 4130
rect 35378 4102 35383 4130
rect 37697 4102 37702 4130
rect 37730 4102 37870 4130
rect 37898 4102 38262 4130
rect 38290 4102 38654 4130
rect 38682 4102 38687 4130
rect 23417 4046 23422 4074
rect 23450 4046 24654 4074
rect 24682 4046 24878 4074
rect 24906 4046 25214 4074
rect 25242 4046 25247 4074
rect 31985 4046 31990 4074
rect 32018 4046 32158 4074
rect 32186 4046 32191 4074
rect 30025 3990 30030 4018
rect 30058 3990 30114 4018
rect 4577 3906 4582 3934
rect 4610 3906 4634 3934
rect 4662 3906 4686 3934
rect 4714 3906 4738 3934
rect 4766 3906 4790 3934
rect 4818 3906 4842 3934
rect 4870 3906 4894 3934
rect 4922 3906 4946 3934
rect 4974 3906 4998 3934
rect 5026 3906 5031 3934
rect 9577 3906 9582 3934
rect 9610 3906 9634 3934
rect 9662 3906 9686 3934
rect 9714 3906 9738 3934
rect 9766 3906 9790 3934
rect 9818 3906 9842 3934
rect 9870 3906 9894 3934
rect 9922 3906 9946 3934
rect 9974 3906 9998 3934
rect 10026 3906 10031 3934
rect 14577 3906 14582 3934
rect 14610 3906 14634 3934
rect 14662 3906 14686 3934
rect 14714 3906 14738 3934
rect 14766 3906 14790 3934
rect 14818 3906 14842 3934
rect 14870 3906 14894 3934
rect 14922 3906 14946 3934
rect 14974 3906 14998 3934
rect 15026 3906 15031 3934
rect 19577 3906 19582 3934
rect 19610 3906 19634 3934
rect 19662 3906 19686 3934
rect 19714 3906 19738 3934
rect 19766 3906 19790 3934
rect 19818 3906 19842 3934
rect 19870 3906 19894 3934
rect 19922 3906 19946 3934
rect 19974 3906 19998 3934
rect 20026 3906 20031 3934
rect 24577 3906 24582 3934
rect 24610 3906 24634 3934
rect 24662 3906 24686 3934
rect 24714 3906 24738 3934
rect 24766 3906 24790 3934
rect 24818 3906 24842 3934
rect 24870 3906 24894 3934
rect 24922 3906 24946 3934
rect 24974 3906 24998 3934
rect 25026 3906 25031 3934
rect 29577 3906 29582 3934
rect 29610 3906 29634 3934
rect 29662 3906 29686 3934
rect 29714 3906 29738 3934
rect 29766 3906 29790 3934
rect 29818 3906 29842 3934
rect 29870 3906 29894 3934
rect 29922 3906 29946 3934
rect 29974 3906 29998 3934
rect 30026 3906 30031 3934
rect 30086 3850 30114 3990
rect 34577 3906 34582 3934
rect 34610 3906 34634 3934
rect 34662 3906 34686 3934
rect 34714 3906 34738 3934
rect 34766 3906 34790 3934
rect 34818 3906 34842 3934
rect 34870 3906 34894 3934
rect 34922 3906 34946 3934
rect 34974 3906 34998 3934
rect 35026 3906 35031 3934
rect 30025 3822 30030 3850
rect 30058 3822 30114 3850
rect 28345 3766 28350 3794
rect 28378 3766 30086 3794
rect 30114 3766 30119 3794
rect 35737 3766 35742 3794
rect 35770 3766 35910 3794
rect 35938 3766 35943 3794
rect 5273 3710 5278 3738
rect 5306 3710 5838 3738
rect 5866 3710 5871 3738
rect 6449 3710 6454 3738
rect 6482 3710 6958 3738
rect 6986 3710 8358 3738
rect 8386 3710 8391 3738
rect 10257 3710 10262 3738
rect 10290 3710 10486 3738
rect 10514 3710 10519 3738
rect 12441 3710 12446 3738
rect 12474 3710 12950 3738
rect 12978 3710 12983 3738
rect 13337 3710 13342 3738
rect 13370 3710 13566 3738
rect 13594 3710 13599 3738
rect 14121 3710 14126 3738
rect 14154 3710 14350 3738
rect 14378 3710 14383 3738
rect 15465 3710 15470 3738
rect 15498 3710 15582 3738
rect 15610 3710 15806 3738
rect 15834 3710 15974 3738
rect 16002 3710 16007 3738
rect 24369 3710 24374 3738
rect 24402 3710 24766 3738
rect 24794 3710 24799 3738
rect 25209 3710 25214 3738
rect 25242 3710 25438 3738
rect 25466 3710 26894 3738
rect 26922 3710 27174 3738
rect 27202 3710 27207 3738
rect 29465 3710 29470 3738
rect 29498 3710 29918 3738
rect 29946 3710 31318 3738
rect 31346 3710 31351 3738
rect 32769 3710 32774 3738
rect 32802 3710 34174 3738
rect 34202 3710 34207 3738
rect 2077 3514 2082 3542
rect 2110 3514 2134 3542
rect 2162 3514 2186 3542
rect 2214 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2394 3542
rect 2422 3514 2446 3542
rect 2474 3514 2498 3542
rect 2526 3514 2531 3542
rect 7077 3514 7082 3542
rect 7110 3514 7134 3542
rect 7162 3514 7186 3542
rect 7214 3514 7238 3542
rect 7266 3514 7290 3542
rect 7318 3514 7342 3542
rect 7370 3514 7394 3542
rect 7422 3514 7446 3542
rect 7474 3514 7498 3542
rect 7526 3514 7531 3542
rect 12077 3514 12082 3542
rect 12110 3514 12134 3542
rect 12162 3514 12186 3542
rect 12214 3514 12238 3542
rect 12266 3514 12290 3542
rect 12318 3514 12342 3542
rect 12370 3514 12394 3542
rect 12422 3514 12446 3542
rect 12474 3514 12498 3542
rect 12526 3514 12531 3542
rect 17077 3514 17082 3542
rect 17110 3514 17134 3542
rect 17162 3514 17186 3542
rect 17214 3514 17238 3542
rect 17266 3514 17290 3542
rect 17318 3514 17342 3542
rect 17370 3514 17394 3542
rect 17422 3514 17446 3542
rect 17474 3514 17498 3542
rect 17526 3514 17531 3542
rect 22077 3514 22082 3542
rect 22110 3514 22134 3542
rect 22162 3514 22186 3542
rect 22214 3514 22238 3542
rect 22266 3514 22290 3542
rect 22318 3514 22342 3542
rect 22370 3514 22394 3542
rect 22422 3514 22446 3542
rect 22474 3514 22498 3542
rect 22526 3514 22531 3542
rect 27077 3514 27082 3542
rect 27110 3514 27134 3542
rect 27162 3514 27186 3542
rect 27214 3514 27238 3542
rect 27266 3514 27290 3542
rect 27318 3514 27342 3542
rect 27370 3514 27394 3542
rect 27422 3514 27446 3542
rect 27474 3514 27498 3542
rect 27526 3514 27531 3542
rect 32077 3514 32082 3542
rect 32110 3514 32134 3542
rect 32162 3514 32186 3542
rect 32214 3514 32238 3542
rect 32266 3514 32290 3542
rect 32318 3514 32342 3542
rect 32370 3514 32394 3542
rect 32422 3514 32446 3542
rect 32474 3514 32498 3542
rect 32526 3514 32531 3542
rect 37077 3514 37082 3542
rect 37110 3514 37134 3542
rect 37162 3514 37186 3542
rect 37214 3514 37238 3542
rect 37266 3514 37290 3542
rect 37318 3514 37342 3542
rect 37370 3514 37394 3542
rect 37422 3514 37446 3542
rect 37474 3514 37498 3542
rect 37526 3514 37531 3542
rect 5385 3430 5390 3458
rect 5418 3430 8862 3458
rect 8890 3430 8895 3458
rect 8073 3374 8078 3402
rect 8106 3374 9534 3402
rect 9562 3374 10038 3402
rect 10066 3374 10071 3402
rect 12049 3374 12054 3402
rect 12082 3374 13342 3402
rect 13370 3374 13375 3402
rect 18489 3374 18494 3402
rect 18522 3374 20566 3402
rect 20594 3374 20599 3402
rect 21737 3374 21742 3402
rect 21770 3374 22806 3402
rect 22834 3374 23198 3402
rect 23226 3374 23422 3402
rect 23450 3374 23455 3402
rect 26889 3374 26894 3402
rect 26922 3374 27174 3402
rect 27202 3374 27398 3402
rect 27426 3374 29358 3402
rect 29386 3374 29391 3402
rect 31873 3374 31878 3402
rect 31906 3374 33334 3402
rect 33362 3374 33367 3402
rect 35289 3374 35294 3402
rect 35322 3374 35742 3402
rect 35770 3374 36694 3402
rect 36722 3374 36727 3402
rect 2473 3318 2478 3346
rect 2506 3318 3038 3346
rect 3066 3318 3071 3346
rect 8969 3318 8974 3346
rect 9002 3318 10318 3346
rect 10346 3318 10351 3346
rect 12721 3318 12726 3346
rect 12754 3318 13678 3346
rect 13706 3318 13902 3346
rect 13930 3318 14126 3346
rect 14154 3318 14159 3346
rect 15129 3318 15134 3346
rect 15162 3318 15526 3346
rect 15554 3318 15559 3346
rect 17929 3318 17934 3346
rect 17962 3318 19166 3346
rect 19194 3318 19199 3346
rect 19441 3318 19446 3346
rect 19474 3318 21014 3346
rect 21042 3318 21182 3346
rect 21210 3318 21215 3346
rect 30697 3318 30702 3346
rect 30730 3318 31990 3346
rect 32018 3318 32158 3346
rect 32186 3318 32191 3346
rect 33777 3318 33782 3346
rect 33810 3318 33950 3346
rect 33978 3318 35854 3346
rect 35882 3318 35887 3346
rect 37585 3318 37590 3346
rect 37618 3318 38150 3346
rect 38178 3318 38183 3346
rect 14126 3290 14154 3318
rect 6449 3262 6454 3290
rect 6482 3262 7014 3290
rect 7042 3262 7047 3290
rect 14126 3262 15246 3290
rect 15274 3262 15279 3290
rect 28345 3262 28350 3290
rect 28378 3262 30030 3290
rect 30058 3262 31990 3290
rect 32018 3262 32023 3290
rect 33889 3262 33894 3290
rect 33922 3262 37030 3290
rect 37058 3262 37063 3290
rect 37697 3262 37702 3290
rect 37730 3262 37926 3290
rect 37954 3262 38262 3290
rect 38290 3262 38295 3290
rect 4577 3122 4582 3150
rect 4610 3122 4634 3150
rect 4662 3122 4686 3150
rect 4714 3122 4738 3150
rect 4766 3122 4790 3150
rect 4818 3122 4842 3150
rect 4870 3122 4894 3150
rect 4922 3122 4946 3150
rect 4974 3122 4998 3150
rect 5026 3122 5031 3150
rect 9577 3122 9582 3150
rect 9610 3122 9634 3150
rect 9662 3122 9686 3150
rect 9714 3122 9738 3150
rect 9766 3122 9790 3150
rect 9818 3122 9842 3150
rect 9870 3122 9894 3150
rect 9922 3122 9946 3150
rect 9974 3122 9998 3150
rect 10026 3122 10031 3150
rect 14577 3122 14582 3150
rect 14610 3122 14634 3150
rect 14662 3122 14686 3150
rect 14714 3122 14738 3150
rect 14766 3122 14790 3150
rect 14818 3122 14842 3150
rect 14870 3122 14894 3150
rect 14922 3122 14946 3150
rect 14974 3122 14998 3150
rect 15026 3122 15031 3150
rect 19577 3122 19582 3150
rect 19610 3122 19634 3150
rect 19662 3122 19686 3150
rect 19714 3122 19738 3150
rect 19766 3122 19790 3150
rect 19818 3122 19842 3150
rect 19870 3122 19894 3150
rect 19922 3122 19946 3150
rect 19974 3122 19998 3150
rect 20026 3122 20031 3150
rect 24577 3122 24582 3150
rect 24610 3122 24634 3150
rect 24662 3122 24686 3150
rect 24714 3122 24738 3150
rect 24766 3122 24790 3150
rect 24818 3122 24842 3150
rect 24870 3122 24894 3150
rect 24922 3122 24946 3150
rect 24974 3122 24998 3150
rect 25026 3122 25031 3150
rect 29577 3122 29582 3150
rect 29610 3122 29634 3150
rect 29662 3122 29686 3150
rect 29714 3122 29738 3150
rect 29766 3122 29790 3150
rect 29818 3122 29842 3150
rect 29870 3122 29894 3150
rect 29922 3122 29946 3150
rect 29974 3122 29998 3150
rect 30026 3122 30031 3150
rect 34577 3122 34582 3150
rect 34610 3122 34634 3150
rect 34662 3122 34686 3150
rect 34714 3122 34738 3150
rect 34766 3122 34790 3150
rect 34818 3122 34842 3150
rect 34870 3122 34894 3150
rect 34922 3122 34946 3150
rect 34974 3122 34998 3150
rect 35026 3122 35031 3150
rect 21401 3038 21406 3066
rect 21434 3038 28630 3066
rect 28658 3038 28663 3066
rect 12441 2982 12446 3010
rect 12474 2982 12726 3010
rect 12754 2982 12759 3010
rect 30305 2982 30310 3010
rect 30338 2982 31094 3010
rect 32041 2982 32046 3010
rect 32074 2982 33670 3010
rect 33698 2982 33703 3010
rect 35737 2982 35742 3010
rect 35770 2982 35910 3010
rect 35938 2982 37702 3010
rect 37730 2982 37735 3010
rect 31066 2954 31094 2982
rect 14121 2926 14126 2954
rect 14154 2926 18886 2954
rect 18914 2926 18919 2954
rect 20785 2926 20790 2954
rect 20818 2926 22246 2954
rect 22274 2926 22582 2954
rect 22610 2926 22615 2954
rect 31066 2926 32214 2954
rect 32242 2926 32382 2954
rect 32410 2926 32606 2954
rect 32634 2926 33782 2954
rect 33810 2926 33815 2954
rect 36129 2926 36134 2954
rect 36162 2926 36694 2954
rect 36722 2926 36727 2954
rect 36857 2926 36862 2954
rect 36890 2926 37142 2954
rect 37170 2926 37366 2954
rect 37394 2926 37399 2954
rect 15297 2870 15302 2898
rect 15330 2870 15470 2898
rect 15498 2870 15503 2898
rect 33329 2870 33334 2898
rect 33362 2870 33894 2898
rect 33922 2870 33927 2898
rect 2077 2730 2082 2758
rect 2110 2730 2134 2758
rect 2162 2730 2186 2758
rect 2214 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2394 2758
rect 2422 2730 2446 2758
rect 2474 2730 2498 2758
rect 2526 2730 2531 2758
rect 7077 2730 7082 2758
rect 7110 2730 7134 2758
rect 7162 2730 7186 2758
rect 7214 2730 7238 2758
rect 7266 2730 7290 2758
rect 7318 2730 7342 2758
rect 7370 2730 7394 2758
rect 7422 2730 7446 2758
rect 7474 2730 7498 2758
rect 7526 2730 7531 2758
rect 12077 2730 12082 2758
rect 12110 2730 12134 2758
rect 12162 2730 12186 2758
rect 12214 2730 12238 2758
rect 12266 2730 12290 2758
rect 12318 2730 12342 2758
rect 12370 2730 12394 2758
rect 12422 2730 12446 2758
rect 12474 2730 12498 2758
rect 12526 2730 12531 2758
rect 17077 2730 17082 2758
rect 17110 2730 17134 2758
rect 17162 2730 17186 2758
rect 17214 2730 17238 2758
rect 17266 2730 17290 2758
rect 17318 2730 17342 2758
rect 17370 2730 17394 2758
rect 17422 2730 17446 2758
rect 17474 2730 17498 2758
rect 17526 2730 17531 2758
rect 22077 2730 22082 2758
rect 22110 2730 22134 2758
rect 22162 2730 22186 2758
rect 22214 2730 22238 2758
rect 22266 2730 22290 2758
rect 22318 2730 22342 2758
rect 22370 2730 22394 2758
rect 22422 2730 22446 2758
rect 22474 2730 22498 2758
rect 22526 2730 22531 2758
rect 27077 2730 27082 2758
rect 27110 2730 27134 2758
rect 27162 2730 27186 2758
rect 27214 2730 27238 2758
rect 27266 2730 27290 2758
rect 27318 2730 27342 2758
rect 27370 2730 27394 2758
rect 27422 2730 27446 2758
rect 27474 2730 27498 2758
rect 27526 2730 27531 2758
rect 32077 2730 32082 2758
rect 32110 2730 32134 2758
rect 32162 2730 32186 2758
rect 32214 2730 32238 2758
rect 32266 2730 32290 2758
rect 32318 2730 32342 2758
rect 32370 2730 32394 2758
rect 32422 2730 32446 2758
rect 32474 2730 32498 2758
rect 32526 2730 32531 2758
rect 37077 2730 37082 2758
rect 37110 2730 37134 2758
rect 37162 2730 37186 2758
rect 37214 2730 37238 2758
rect 37266 2730 37290 2758
rect 37318 2730 37342 2758
rect 37370 2730 37394 2758
rect 37422 2730 37446 2758
rect 37474 2730 37498 2758
rect 37526 2730 37531 2758
rect 26889 2646 26894 2674
rect 26922 2646 27174 2674
rect 27202 2646 27207 2674
rect 28681 2646 28686 2674
rect 28714 2646 32438 2674
rect 32466 2646 32471 2674
rect 14233 2590 14238 2618
rect 14266 2590 17598 2618
rect 17626 2590 19222 2618
rect 19250 2590 19255 2618
rect 20953 2590 20958 2618
rect 20986 2590 33334 2618
rect 33362 2590 33367 2618
rect 34673 2590 34678 2618
rect 34706 2590 36134 2618
rect 36162 2590 36167 2618
rect 38425 2590 38430 2618
rect 38458 2590 38822 2618
rect 38850 2590 38855 2618
rect 2473 2534 2478 2562
rect 2506 2534 3038 2562
rect 3066 2534 3071 2562
rect 15913 2534 15918 2562
rect 15946 2534 17150 2562
rect 17178 2534 17374 2562
rect 17402 2534 17654 2562
rect 17682 2534 17687 2562
rect 20113 2534 20118 2562
rect 20146 2534 21406 2562
rect 21434 2534 21439 2562
rect 23193 2534 23198 2562
rect 23226 2534 23534 2562
rect 23562 2534 24654 2562
rect 24682 2534 24878 2562
rect 24906 2534 25214 2562
rect 25242 2534 25438 2562
rect 25466 2534 25471 2562
rect 26273 2534 26278 2562
rect 26306 2534 26726 2562
rect 26754 2534 28462 2562
rect 28490 2534 28630 2562
rect 28658 2534 29022 2562
rect 29050 2534 30366 2562
rect 30394 2534 30702 2562
rect 30730 2534 30735 2562
rect 33665 2534 33670 2562
rect 33698 2534 35686 2562
rect 35714 2534 35719 2562
rect 38145 2534 38150 2562
rect 38178 2534 38878 2562
rect 38906 2534 38911 2562
rect 1633 2478 1638 2506
rect 1666 2478 4494 2506
rect 4522 2478 4998 2506
rect 5026 2478 6342 2506
rect 6370 2478 6375 2506
rect 8465 2478 8470 2506
rect 8498 2478 8974 2506
rect 9002 2478 10262 2506
rect 10290 2478 10295 2506
rect 15241 2478 15246 2506
rect 15274 2478 16814 2506
rect 16842 2478 16847 2506
rect 18769 2478 18774 2506
rect 18802 2478 20230 2506
rect 20258 2478 20790 2506
rect 20818 2478 20823 2506
rect 24089 2478 24094 2506
rect 24122 2478 26054 2506
rect 26082 2478 26222 2506
rect 26250 2478 28238 2506
rect 28266 2478 30030 2506
rect 30058 2478 30063 2506
rect 34510 2478 35518 2506
rect 35546 2478 38990 2506
rect 39018 2478 39023 2506
rect 34510 2450 34538 2478
rect 22745 2422 22750 2450
rect 22778 2422 24374 2450
rect 24402 2422 24486 2450
rect 24514 2422 24766 2450
rect 24794 2422 24799 2450
rect 26329 2422 26334 2450
rect 26362 2422 31598 2450
rect 31626 2422 31631 2450
rect 34505 2422 34510 2450
rect 34538 2422 34543 2450
rect 4577 2338 4582 2366
rect 4610 2338 4634 2366
rect 4662 2338 4686 2366
rect 4714 2338 4738 2366
rect 4766 2338 4790 2366
rect 4818 2338 4842 2366
rect 4870 2338 4894 2366
rect 4922 2338 4946 2366
rect 4974 2338 4998 2366
rect 5026 2338 5031 2366
rect 9577 2338 9582 2366
rect 9610 2338 9634 2366
rect 9662 2338 9686 2366
rect 9714 2338 9738 2366
rect 9766 2338 9790 2366
rect 9818 2338 9842 2366
rect 9870 2338 9894 2366
rect 9922 2338 9946 2366
rect 9974 2338 9998 2366
rect 10026 2338 10031 2366
rect 14577 2338 14582 2366
rect 14610 2338 14634 2366
rect 14662 2338 14686 2366
rect 14714 2338 14738 2366
rect 14766 2338 14790 2366
rect 14818 2338 14842 2366
rect 14870 2338 14894 2366
rect 14922 2338 14946 2366
rect 14974 2338 14998 2366
rect 15026 2338 15031 2366
rect 19577 2338 19582 2366
rect 19610 2338 19634 2366
rect 19662 2338 19686 2366
rect 19714 2338 19738 2366
rect 19766 2338 19790 2366
rect 19818 2338 19842 2366
rect 19870 2338 19894 2366
rect 19922 2338 19946 2366
rect 19974 2338 19998 2366
rect 20026 2338 20031 2366
rect 24577 2338 24582 2366
rect 24610 2338 24634 2366
rect 24662 2338 24686 2366
rect 24714 2338 24738 2366
rect 24766 2338 24790 2366
rect 24818 2338 24842 2366
rect 24870 2338 24894 2366
rect 24922 2338 24946 2366
rect 24974 2338 24998 2366
rect 25026 2338 25031 2366
rect 29577 2338 29582 2366
rect 29610 2338 29634 2366
rect 29662 2338 29686 2366
rect 29714 2338 29738 2366
rect 29766 2338 29790 2366
rect 29818 2338 29842 2366
rect 29870 2338 29894 2366
rect 29922 2338 29946 2366
rect 29974 2338 29998 2366
rect 30026 2338 30031 2366
rect 34577 2338 34582 2366
rect 34610 2338 34634 2366
rect 34662 2338 34686 2366
rect 34714 2338 34738 2366
rect 34766 2338 34790 2366
rect 34818 2338 34842 2366
rect 34870 2338 34894 2366
rect 34922 2338 34946 2366
rect 34974 2338 34998 2366
rect 35026 2338 35031 2366
rect 2025 2198 2030 2226
rect 2058 2198 2478 2226
rect 2506 2198 4438 2226
rect 4466 2198 4471 2226
rect 11993 2198 11998 2226
rect 12026 2198 12446 2226
rect 12474 2198 12726 2226
rect 12754 2198 13510 2226
rect 13538 2198 14070 2226
rect 14098 2198 14294 2226
rect 14322 2198 14327 2226
rect 29409 2198 29414 2226
rect 29442 2198 31262 2226
rect 31290 2198 31295 2226
rect 3033 2142 3038 2170
rect 3066 2142 3486 2170
rect 3514 2142 3519 2170
rect 5889 2142 5894 2170
rect 5922 2142 7294 2170
rect 7322 2142 7574 2170
rect 7602 2142 7798 2170
rect 7826 2142 7831 2170
rect 10033 2142 10038 2170
rect 10066 2142 11214 2170
rect 11242 2142 11247 2170
rect 13337 2142 13342 2170
rect 13370 2142 13622 2170
rect 13650 2142 15134 2170
rect 15162 2142 15167 2170
rect 16585 2142 16590 2170
rect 16618 2142 18270 2170
rect 18298 2142 18550 2170
rect 18578 2142 18774 2170
rect 18802 2142 18807 2170
rect 24481 2142 24486 2170
rect 24514 2142 24766 2170
rect 24794 2142 26222 2170
rect 26250 2142 26255 2170
rect 30249 2142 30254 2170
rect 30282 2142 31654 2170
rect 31682 2142 31687 2170
rect 2077 1946 2082 1974
rect 2110 1946 2134 1974
rect 2162 1946 2186 1974
rect 2214 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2394 1974
rect 2422 1946 2446 1974
rect 2474 1946 2498 1974
rect 2526 1946 2531 1974
rect 7077 1946 7082 1974
rect 7110 1946 7134 1974
rect 7162 1946 7186 1974
rect 7214 1946 7238 1974
rect 7266 1946 7290 1974
rect 7318 1946 7342 1974
rect 7370 1946 7394 1974
rect 7422 1946 7446 1974
rect 7474 1946 7498 1974
rect 7526 1946 7531 1974
rect 12077 1946 12082 1974
rect 12110 1946 12134 1974
rect 12162 1946 12186 1974
rect 12214 1946 12238 1974
rect 12266 1946 12290 1974
rect 12318 1946 12342 1974
rect 12370 1946 12394 1974
rect 12422 1946 12446 1974
rect 12474 1946 12498 1974
rect 12526 1946 12531 1974
rect 17077 1946 17082 1974
rect 17110 1946 17134 1974
rect 17162 1946 17186 1974
rect 17214 1946 17238 1974
rect 17266 1946 17290 1974
rect 17318 1946 17342 1974
rect 17370 1946 17394 1974
rect 17422 1946 17446 1974
rect 17474 1946 17498 1974
rect 17526 1946 17531 1974
rect 22077 1946 22082 1974
rect 22110 1946 22134 1974
rect 22162 1946 22186 1974
rect 22214 1946 22238 1974
rect 22266 1946 22290 1974
rect 22318 1946 22342 1974
rect 22370 1946 22394 1974
rect 22422 1946 22446 1974
rect 22474 1946 22498 1974
rect 22526 1946 22531 1974
rect 27077 1946 27082 1974
rect 27110 1946 27134 1974
rect 27162 1946 27186 1974
rect 27214 1946 27238 1974
rect 27266 1946 27290 1974
rect 27318 1946 27342 1974
rect 27370 1946 27394 1974
rect 27422 1946 27446 1974
rect 27474 1946 27498 1974
rect 27526 1946 27531 1974
rect 32077 1946 32082 1974
rect 32110 1946 32134 1974
rect 32162 1946 32186 1974
rect 32214 1946 32238 1974
rect 32266 1946 32290 1974
rect 32318 1946 32342 1974
rect 32370 1946 32394 1974
rect 32422 1946 32446 1974
rect 32474 1946 32498 1974
rect 32526 1946 32531 1974
rect 37077 1946 37082 1974
rect 37110 1946 37134 1974
rect 37162 1946 37186 1974
rect 37214 1946 37238 1974
rect 37266 1946 37290 1974
rect 37318 1946 37342 1974
rect 37370 1946 37394 1974
rect 37422 1946 37446 1974
rect 37474 1946 37498 1974
rect 37526 1946 37531 1974
rect 7569 1862 7574 1890
rect 7602 1862 8302 1890
rect 8330 1862 9422 1890
rect 9450 1862 16590 1890
rect 16618 1862 16623 1890
rect 17033 1862 17038 1890
rect 17066 1862 17990 1890
rect 18018 1862 18023 1890
rect 24313 1862 24318 1890
rect 24346 1862 36190 1890
rect 36218 1862 37590 1890
rect 37618 1862 37623 1890
rect 3481 1806 3486 1834
rect 3514 1806 3822 1834
rect 3850 1806 5502 1834
rect 5530 1806 13454 1834
rect 15297 1806 15302 1834
rect 15330 1806 15526 1834
rect 15554 1806 15559 1834
rect 20118 1806 22470 1834
rect 22498 1806 22503 1834
rect 31593 1806 31598 1834
rect 31626 1806 38150 1834
rect 38178 1806 38934 1834
rect 38962 1806 38967 1834
rect 13426 1778 13454 1806
rect 20118 1778 20146 1806
rect 6505 1750 6510 1778
rect 6538 1750 8134 1778
rect 8162 1750 8167 1778
rect 13426 1750 20118 1778
rect 20146 1750 20151 1778
rect 21177 1750 21182 1778
rect 21210 1750 22862 1778
rect 22890 1750 23086 1778
rect 23114 1750 23119 1778
rect 35681 1750 35686 1778
rect 35714 1750 37422 1778
rect 37450 1750 37455 1778
rect 38649 1750 38654 1778
rect 38682 1750 38822 1778
rect 38850 1750 38855 1778
rect 2478 1694 2926 1722
rect 2954 1694 2959 1722
rect 4433 1694 4438 1722
rect 4466 1694 5082 1722
rect 21793 1694 21798 1722
rect 21826 1694 33446 1722
rect 33474 1694 35070 1722
rect 35098 1694 37142 1722
rect 37170 1694 37175 1722
rect 2478 1666 2506 1694
rect 5054 1666 5082 1694
rect 2473 1638 2478 1666
rect 2506 1638 2511 1666
rect 5054 1638 28798 1666
rect 28826 1638 29022 1666
rect 29050 1638 29055 1666
rect 4577 1554 4582 1582
rect 4610 1554 4634 1582
rect 4662 1554 4686 1582
rect 4714 1554 4738 1582
rect 4766 1554 4790 1582
rect 4818 1554 4842 1582
rect 4870 1554 4894 1582
rect 4922 1554 4946 1582
rect 4974 1554 4998 1582
rect 5026 1554 5031 1582
rect 9577 1554 9582 1582
rect 9610 1554 9634 1582
rect 9662 1554 9686 1582
rect 9714 1554 9738 1582
rect 9766 1554 9790 1582
rect 9818 1554 9842 1582
rect 9870 1554 9894 1582
rect 9922 1554 9946 1582
rect 9974 1554 9998 1582
rect 10026 1554 10031 1582
rect 14577 1554 14582 1582
rect 14610 1554 14634 1582
rect 14662 1554 14686 1582
rect 14714 1554 14738 1582
rect 14766 1554 14790 1582
rect 14818 1554 14842 1582
rect 14870 1554 14894 1582
rect 14922 1554 14946 1582
rect 14974 1554 14998 1582
rect 15026 1554 15031 1582
rect 19577 1554 19582 1582
rect 19610 1554 19634 1582
rect 19662 1554 19686 1582
rect 19714 1554 19738 1582
rect 19766 1554 19790 1582
rect 19818 1554 19842 1582
rect 19870 1554 19894 1582
rect 19922 1554 19946 1582
rect 19974 1554 19998 1582
rect 20026 1554 20031 1582
rect 24577 1554 24582 1582
rect 24610 1554 24634 1582
rect 24662 1554 24686 1582
rect 24714 1554 24738 1582
rect 24766 1554 24790 1582
rect 24818 1554 24842 1582
rect 24870 1554 24894 1582
rect 24922 1554 24946 1582
rect 24974 1554 24998 1582
rect 25026 1554 25031 1582
rect 29577 1554 29582 1582
rect 29610 1554 29634 1582
rect 29662 1554 29686 1582
rect 29714 1554 29738 1582
rect 29766 1554 29790 1582
rect 29818 1554 29842 1582
rect 29870 1554 29894 1582
rect 29922 1554 29946 1582
rect 29974 1554 29998 1582
rect 30026 1554 30031 1582
rect 34577 1554 34582 1582
rect 34610 1554 34634 1582
rect 34662 1554 34686 1582
rect 34714 1554 34738 1582
rect 34766 1554 34790 1582
rect 34818 1554 34842 1582
rect 34870 1554 34894 1582
rect 34922 1554 34946 1582
rect 34974 1554 34998 1582
rect 35026 1554 35031 1582
rect 2529 1470 2534 1498
rect 2562 1470 18494 1498
rect 18522 1470 18527 1498
rect 6393 1414 6398 1442
rect 6426 1414 22918 1442
rect 22946 1414 22951 1442
<< via3 >>
rect 2082 18410 2110 18438
rect 2134 18410 2162 18438
rect 2186 18410 2214 18438
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 2394 18410 2422 18438
rect 2446 18410 2474 18438
rect 2498 18410 2526 18438
rect 7082 18410 7110 18438
rect 7134 18410 7162 18438
rect 7186 18410 7214 18438
rect 7238 18410 7266 18438
rect 7290 18410 7318 18438
rect 7342 18410 7370 18438
rect 7394 18410 7422 18438
rect 7446 18410 7474 18438
rect 7498 18410 7526 18438
rect 12082 18410 12110 18438
rect 12134 18410 12162 18438
rect 12186 18410 12214 18438
rect 12238 18410 12266 18438
rect 12290 18410 12318 18438
rect 12342 18410 12370 18438
rect 12394 18410 12422 18438
rect 12446 18410 12474 18438
rect 12498 18410 12526 18438
rect 17082 18410 17110 18438
rect 17134 18410 17162 18438
rect 17186 18410 17214 18438
rect 17238 18410 17266 18438
rect 17290 18410 17318 18438
rect 17342 18410 17370 18438
rect 17394 18410 17422 18438
rect 17446 18410 17474 18438
rect 17498 18410 17526 18438
rect 22082 18410 22110 18438
rect 22134 18410 22162 18438
rect 22186 18410 22214 18438
rect 22238 18410 22266 18438
rect 22290 18410 22318 18438
rect 22342 18410 22370 18438
rect 22394 18410 22422 18438
rect 22446 18410 22474 18438
rect 22498 18410 22526 18438
rect 27082 18410 27110 18438
rect 27134 18410 27162 18438
rect 27186 18410 27214 18438
rect 27238 18410 27266 18438
rect 27290 18410 27318 18438
rect 27342 18410 27370 18438
rect 27394 18410 27422 18438
rect 27446 18410 27474 18438
rect 27498 18410 27526 18438
rect 32082 18410 32110 18438
rect 32134 18410 32162 18438
rect 32186 18410 32214 18438
rect 32238 18410 32266 18438
rect 32290 18410 32318 18438
rect 32342 18410 32370 18438
rect 32394 18410 32422 18438
rect 32446 18410 32474 18438
rect 32498 18410 32526 18438
rect 37082 18410 37110 18438
rect 37134 18410 37162 18438
rect 37186 18410 37214 18438
rect 37238 18410 37266 18438
rect 37290 18410 37318 18438
rect 37342 18410 37370 18438
rect 37394 18410 37422 18438
rect 37446 18410 37474 18438
rect 37498 18410 37526 18438
rect 4582 18018 4610 18046
rect 4634 18018 4662 18046
rect 4686 18018 4714 18046
rect 4738 18018 4766 18046
rect 4790 18018 4818 18046
rect 4842 18018 4870 18046
rect 4894 18018 4922 18046
rect 4946 18018 4974 18046
rect 4998 18018 5026 18046
rect 9582 18018 9610 18046
rect 9634 18018 9662 18046
rect 9686 18018 9714 18046
rect 9738 18018 9766 18046
rect 9790 18018 9818 18046
rect 9842 18018 9870 18046
rect 9894 18018 9922 18046
rect 9946 18018 9974 18046
rect 9998 18018 10026 18046
rect 14582 18018 14610 18046
rect 14634 18018 14662 18046
rect 14686 18018 14714 18046
rect 14738 18018 14766 18046
rect 14790 18018 14818 18046
rect 14842 18018 14870 18046
rect 14894 18018 14922 18046
rect 14946 18018 14974 18046
rect 14998 18018 15026 18046
rect 19582 18018 19610 18046
rect 19634 18018 19662 18046
rect 19686 18018 19714 18046
rect 19738 18018 19766 18046
rect 19790 18018 19818 18046
rect 19842 18018 19870 18046
rect 19894 18018 19922 18046
rect 19946 18018 19974 18046
rect 19998 18018 20026 18046
rect 24582 18018 24610 18046
rect 24634 18018 24662 18046
rect 24686 18018 24714 18046
rect 24738 18018 24766 18046
rect 24790 18018 24818 18046
rect 24842 18018 24870 18046
rect 24894 18018 24922 18046
rect 24946 18018 24974 18046
rect 24998 18018 25026 18046
rect 29582 18018 29610 18046
rect 29634 18018 29662 18046
rect 29686 18018 29714 18046
rect 29738 18018 29766 18046
rect 29790 18018 29818 18046
rect 29842 18018 29870 18046
rect 29894 18018 29922 18046
rect 29946 18018 29974 18046
rect 29998 18018 30026 18046
rect 34582 18018 34610 18046
rect 34634 18018 34662 18046
rect 34686 18018 34714 18046
rect 34738 18018 34766 18046
rect 34790 18018 34818 18046
rect 34842 18018 34870 18046
rect 34894 18018 34922 18046
rect 34946 18018 34974 18046
rect 34998 18018 35026 18046
rect 2082 17626 2110 17654
rect 2134 17626 2162 17654
rect 2186 17626 2214 17654
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 2394 17626 2422 17654
rect 2446 17626 2474 17654
rect 2498 17626 2526 17654
rect 7082 17626 7110 17654
rect 7134 17626 7162 17654
rect 7186 17626 7214 17654
rect 7238 17626 7266 17654
rect 7290 17626 7318 17654
rect 7342 17626 7370 17654
rect 7394 17626 7422 17654
rect 7446 17626 7474 17654
rect 7498 17626 7526 17654
rect 12082 17626 12110 17654
rect 12134 17626 12162 17654
rect 12186 17626 12214 17654
rect 12238 17626 12266 17654
rect 12290 17626 12318 17654
rect 12342 17626 12370 17654
rect 12394 17626 12422 17654
rect 12446 17626 12474 17654
rect 12498 17626 12526 17654
rect 17082 17626 17110 17654
rect 17134 17626 17162 17654
rect 17186 17626 17214 17654
rect 17238 17626 17266 17654
rect 17290 17626 17318 17654
rect 17342 17626 17370 17654
rect 17394 17626 17422 17654
rect 17446 17626 17474 17654
rect 17498 17626 17526 17654
rect 22082 17626 22110 17654
rect 22134 17626 22162 17654
rect 22186 17626 22214 17654
rect 22238 17626 22266 17654
rect 22290 17626 22318 17654
rect 22342 17626 22370 17654
rect 22394 17626 22422 17654
rect 22446 17626 22474 17654
rect 22498 17626 22526 17654
rect 27082 17626 27110 17654
rect 27134 17626 27162 17654
rect 27186 17626 27214 17654
rect 27238 17626 27266 17654
rect 27290 17626 27318 17654
rect 27342 17626 27370 17654
rect 27394 17626 27422 17654
rect 27446 17626 27474 17654
rect 27498 17626 27526 17654
rect 32082 17626 32110 17654
rect 32134 17626 32162 17654
rect 32186 17626 32214 17654
rect 32238 17626 32266 17654
rect 32290 17626 32318 17654
rect 32342 17626 32370 17654
rect 32394 17626 32422 17654
rect 32446 17626 32474 17654
rect 32498 17626 32526 17654
rect 37082 17626 37110 17654
rect 37134 17626 37162 17654
rect 37186 17626 37214 17654
rect 37238 17626 37266 17654
rect 37290 17626 37318 17654
rect 37342 17626 37370 17654
rect 37394 17626 37422 17654
rect 37446 17626 37474 17654
rect 37498 17626 37526 17654
rect 4582 17234 4610 17262
rect 4634 17234 4662 17262
rect 4686 17234 4714 17262
rect 4738 17234 4766 17262
rect 4790 17234 4818 17262
rect 4842 17234 4870 17262
rect 4894 17234 4922 17262
rect 4946 17234 4974 17262
rect 4998 17234 5026 17262
rect 9582 17234 9610 17262
rect 9634 17234 9662 17262
rect 9686 17234 9714 17262
rect 9738 17234 9766 17262
rect 9790 17234 9818 17262
rect 9842 17234 9870 17262
rect 9894 17234 9922 17262
rect 9946 17234 9974 17262
rect 9998 17234 10026 17262
rect 14582 17234 14610 17262
rect 14634 17234 14662 17262
rect 14686 17234 14714 17262
rect 14738 17234 14766 17262
rect 14790 17234 14818 17262
rect 14842 17234 14870 17262
rect 14894 17234 14922 17262
rect 14946 17234 14974 17262
rect 14998 17234 15026 17262
rect 19582 17234 19610 17262
rect 19634 17234 19662 17262
rect 19686 17234 19714 17262
rect 19738 17234 19766 17262
rect 19790 17234 19818 17262
rect 19842 17234 19870 17262
rect 19894 17234 19922 17262
rect 19946 17234 19974 17262
rect 19998 17234 20026 17262
rect 24582 17234 24610 17262
rect 24634 17234 24662 17262
rect 24686 17234 24714 17262
rect 24738 17234 24766 17262
rect 24790 17234 24818 17262
rect 24842 17234 24870 17262
rect 24894 17234 24922 17262
rect 24946 17234 24974 17262
rect 24998 17234 25026 17262
rect 29582 17234 29610 17262
rect 29634 17234 29662 17262
rect 29686 17234 29714 17262
rect 29738 17234 29766 17262
rect 29790 17234 29818 17262
rect 29842 17234 29870 17262
rect 29894 17234 29922 17262
rect 29946 17234 29974 17262
rect 29998 17234 30026 17262
rect 34582 17234 34610 17262
rect 34634 17234 34662 17262
rect 34686 17234 34714 17262
rect 34738 17234 34766 17262
rect 34790 17234 34818 17262
rect 34842 17234 34870 17262
rect 34894 17234 34922 17262
rect 34946 17234 34974 17262
rect 34998 17234 35026 17262
rect 2082 16842 2110 16870
rect 2134 16842 2162 16870
rect 2186 16842 2214 16870
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 2394 16842 2422 16870
rect 2446 16842 2474 16870
rect 2498 16842 2526 16870
rect 7082 16842 7110 16870
rect 7134 16842 7162 16870
rect 7186 16842 7214 16870
rect 7238 16842 7266 16870
rect 7290 16842 7318 16870
rect 7342 16842 7370 16870
rect 7394 16842 7422 16870
rect 7446 16842 7474 16870
rect 7498 16842 7526 16870
rect 12082 16842 12110 16870
rect 12134 16842 12162 16870
rect 12186 16842 12214 16870
rect 12238 16842 12266 16870
rect 12290 16842 12318 16870
rect 12342 16842 12370 16870
rect 12394 16842 12422 16870
rect 12446 16842 12474 16870
rect 12498 16842 12526 16870
rect 17082 16842 17110 16870
rect 17134 16842 17162 16870
rect 17186 16842 17214 16870
rect 17238 16842 17266 16870
rect 17290 16842 17318 16870
rect 17342 16842 17370 16870
rect 17394 16842 17422 16870
rect 17446 16842 17474 16870
rect 17498 16842 17526 16870
rect 22082 16842 22110 16870
rect 22134 16842 22162 16870
rect 22186 16842 22214 16870
rect 22238 16842 22266 16870
rect 22290 16842 22318 16870
rect 22342 16842 22370 16870
rect 22394 16842 22422 16870
rect 22446 16842 22474 16870
rect 22498 16842 22526 16870
rect 27082 16842 27110 16870
rect 27134 16842 27162 16870
rect 27186 16842 27214 16870
rect 27238 16842 27266 16870
rect 27290 16842 27318 16870
rect 27342 16842 27370 16870
rect 27394 16842 27422 16870
rect 27446 16842 27474 16870
rect 27498 16842 27526 16870
rect 32082 16842 32110 16870
rect 32134 16842 32162 16870
rect 32186 16842 32214 16870
rect 32238 16842 32266 16870
rect 32290 16842 32318 16870
rect 32342 16842 32370 16870
rect 32394 16842 32422 16870
rect 32446 16842 32474 16870
rect 32498 16842 32526 16870
rect 37082 16842 37110 16870
rect 37134 16842 37162 16870
rect 37186 16842 37214 16870
rect 37238 16842 37266 16870
rect 37290 16842 37318 16870
rect 37342 16842 37370 16870
rect 37394 16842 37422 16870
rect 37446 16842 37474 16870
rect 37498 16842 37526 16870
rect 4582 16450 4610 16478
rect 4634 16450 4662 16478
rect 4686 16450 4714 16478
rect 4738 16450 4766 16478
rect 4790 16450 4818 16478
rect 4842 16450 4870 16478
rect 4894 16450 4922 16478
rect 4946 16450 4974 16478
rect 4998 16450 5026 16478
rect 9582 16450 9610 16478
rect 9634 16450 9662 16478
rect 9686 16450 9714 16478
rect 9738 16450 9766 16478
rect 9790 16450 9818 16478
rect 9842 16450 9870 16478
rect 9894 16450 9922 16478
rect 9946 16450 9974 16478
rect 9998 16450 10026 16478
rect 14582 16450 14610 16478
rect 14634 16450 14662 16478
rect 14686 16450 14714 16478
rect 14738 16450 14766 16478
rect 14790 16450 14818 16478
rect 14842 16450 14870 16478
rect 14894 16450 14922 16478
rect 14946 16450 14974 16478
rect 14998 16450 15026 16478
rect 19582 16450 19610 16478
rect 19634 16450 19662 16478
rect 19686 16450 19714 16478
rect 19738 16450 19766 16478
rect 19790 16450 19818 16478
rect 19842 16450 19870 16478
rect 19894 16450 19922 16478
rect 19946 16450 19974 16478
rect 19998 16450 20026 16478
rect 24582 16450 24610 16478
rect 24634 16450 24662 16478
rect 24686 16450 24714 16478
rect 24738 16450 24766 16478
rect 24790 16450 24818 16478
rect 24842 16450 24870 16478
rect 24894 16450 24922 16478
rect 24946 16450 24974 16478
rect 24998 16450 25026 16478
rect 29582 16450 29610 16478
rect 29634 16450 29662 16478
rect 29686 16450 29714 16478
rect 29738 16450 29766 16478
rect 29790 16450 29818 16478
rect 29842 16450 29870 16478
rect 29894 16450 29922 16478
rect 29946 16450 29974 16478
rect 29998 16450 30026 16478
rect 34582 16450 34610 16478
rect 34634 16450 34662 16478
rect 34686 16450 34714 16478
rect 34738 16450 34766 16478
rect 34790 16450 34818 16478
rect 34842 16450 34870 16478
rect 34894 16450 34922 16478
rect 34946 16450 34974 16478
rect 34998 16450 35026 16478
rect 10094 16254 10122 16282
rect 2082 16058 2110 16086
rect 2134 16058 2162 16086
rect 2186 16058 2214 16086
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 2394 16058 2422 16086
rect 2446 16058 2474 16086
rect 2498 16058 2526 16086
rect 7082 16058 7110 16086
rect 7134 16058 7162 16086
rect 7186 16058 7214 16086
rect 7238 16058 7266 16086
rect 7290 16058 7318 16086
rect 7342 16058 7370 16086
rect 7394 16058 7422 16086
rect 7446 16058 7474 16086
rect 7498 16058 7526 16086
rect 12082 16058 12110 16086
rect 12134 16058 12162 16086
rect 12186 16058 12214 16086
rect 12238 16058 12266 16086
rect 12290 16058 12318 16086
rect 12342 16058 12370 16086
rect 12394 16058 12422 16086
rect 12446 16058 12474 16086
rect 12498 16058 12526 16086
rect 17082 16058 17110 16086
rect 17134 16058 17162 16086
rect 17186 16058 17214 16086
rect 17238 16058 17266 16086
rect 17290 16058 17318 16086
rect 17342 16058 17370 16086
rect 17394 16058 17422 16086
rect 17446 16058 17474 16086
rect 17498 16058 17526 16086
rect 22082 16058 22110 16086
rect 22134 16058 22162 16086
rect 22186 16058 22214 16086
rect 22238 16058 22266 16086
rect 22290 16058 22318 16086
rect 22342 16058 22370 16086
rect 22394 16058 22422 16086
rect 22446 16058 22474 16086
rect 22498 16058 22526 16086
rect 27082 16058 27110 16086
rect 27134 16058 27162 16086
rect 27186 16058 27214 16086
rect 27238 16058 27266 16086
rect 27290 16058 27318 16086
rect 27342 16058 27370 16086
rect 27394 16058 27422 16086
rect 27446 16058 27474 16086
rect 27498 16058 27526 16086
rect 32082 16058 32110 16086
rect 32134 16058 32162 16086
rect 32186 16058 32214 16086
rect 32238 16058 32266 16086
rect 32290 16058 32318 16086
rect 32342 16058 32370 16086
rect 32394 16058 32422 16086
rect 32446 16058 32474 16086
rect 32498 16058 32526 16086
rect 37082 16058 37110 16086
rect 37134 16058 37162 16086
rect 37186 16058 37214 16086
rect 37238 16058 37266 16086
rect 37290 16058 37318 16086
rect 37342 16058 37370 16086
rect 37394 16058 37422 16086
rect 37446 16058 37474 16086
rect 37498 16058 37526 16086
rect 4582 15666 4610 15694
rect 4634 15666 4662 15694
rect 4686 15666 4714 15694
rect 4738 15666 4766 15694
rect 4790 15666 4818 15694
rect 4842 15666 4870 15694
rect 4894 15666 4922 15694
rect 4946 15666 4974 15694
rect 4998 15666 5026 15694
rect 9582 15666 9610 15694
rect 9634 15666 9662 15694
rect 9686 15666 9714 15694
rect 9738 15666 9766 15694
rect 9790 15666 9818 15694
rect 9842 15666 9870 15694
rect 9894 15666 9922 15694
rect 9946 15666 9974 15694
rect 9998 15666 10026 15694
rect 14582 15666 14610 15694
rect 14634 15666 14662 15694
rect 14686 15666 14714 15694
rect 14738 15666 14766 15694
rect 14790 15666 14818 15694
rect 14842 15666 14870 15694
rect 14894 15666 14922 15694
rect 14946 15666 14974 15694
rect 14998 15666 15026 15694
rect 19582 15666 19610 15694
rect 19634 15666 19662 15694
rect 19686 15666 19714 15694
rect 19738 15666 19766 15694
rect 19790 15666 19818 15694
rect 19842 15666 19870 15694
rect 19894 15666 19922 15694
rect 19946 15666 19974 15694
rect 19998 15666 20026 15694
rect 24582 15666 24610 15694
rect 24634 15666 24662 15694
rect 24686 15666 24714 15694
rect 24738 15666 24766 15694
rect 24790 15666 24818 15694
rect 24842 15666 24870 15694
rect 24894 15666 24922 15694
rect 24946 15666 24974 15694
rect 24998 15666 25026 15694
rect 29582 15666 29610 15694
rect 29634 15666 29662 15694
rect 29686 15666 29714 15694
rect 29738 15666 29766 15694
rect 29790 15666 29818 15694
rect 29842 15666 29870 15694
rect 29894 15666 29922 15694
rect 29946 15666 29974 15694
rect 29998 15666 30026 15694
rect 34582 15666 34610 15694
rect 34634 15666 34662 15694
rect 34686 15666 34714 15694
rect 34738 15666 34766 15694
rect 34790 15666 34818 15694
rect 34842 15666 34870 15694
rect 34894 15666 34922 15694
rect 34946 15666 34974 15694
rect 34998 15666 35026 15694
rect 10094 15470 10122 15498
rect 2082 15274 2110 15302
rect 2134 15274 2162 15302
rect 2186 15274 2214 15302
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 2394 15274 2422 15302
rect 2446 15274 2474 15302
rect 2498 15274 2526 15302
rect 7082 15274 7110 15302
rect 7134 15274 7162 15302
rect 7186 15274 7214 15302
rect 7238 15274 7266 15302
rect 7290 15274 7318 15302
rect 7342 15274 7370 15302
rect 7394 15274 7422 15302
rect 7446 15274 7474 15302
rect 7498 15274 7526 15302
rect 12082 15274 12110 15302
rect 12134 15274 12162 15302
rect 12186 15274 12214 15302
rect 12238 15274 12266 15302
rect 12290 15274 12318 15302
rect 12342 15274 12370 15302
rect 12394 15274 12422 15302
rect 12446 15274 12474 15302
rect 12498 15274 12526 15302
rect 17082 15274 17110 15302
rect 17134 15274 17162 15302
rect 17186 15274 17214 15302
rect 17238 15274 17266 15302
rect 17290 15274 17318 15302
rect 17342 15274 17370 15302
rect 17394 15274 17422 15302
rect 17446 15274 17474 15302
rect 17498 15274 17526 15302
rect 22082 15274 22110 15302
rect 22134 15274 22162 15302
rect 22186 15274 22214 15302
rect 22238 15274 22266 15302
rect 22290 15274 22318 15302
rect 22342 15274 22370 15302
rect 22394 15274 22422 15302
rect 22446 15274 22474 15302
rect 22498 15274 22526 15302
rect 27082 15274 27110 15302
rect 27134 15274 27162 15302
rect 27186 15274 27214 15302
rect 27238 15274 27266 15302
rect 27290 15274 27318 15302
rect 27342 15274 27370 15302
rect 27394 15274 27422 15302
rect 27446 15274 27474 15302
rect 27498 15274 27526 15302
rect 32082 15274 32110 15302
rect 32134 15274 32162 15302
rect 32186 15274 32214 15302
rect 32238 15274 32266 15302
rect 32290 15274 32318 15302
rect 32342 15274 32370 15302
rect 32394 15274 32422 15302
rect 32446 15274 32474 15302
rect 32498 15274 32526 15302
rect 37082 15274 37110 15302
rect 37134 15274 37162 15302
rect 37186 15274 37214 15302
rect 37238 15274 37266 15302
rect 37290 15274 37318 15302
rect 37342 15274 37370 15302
rect 37394 15274 37422 15302
rect 37446 15274 37474 15302
rect 37498 15274 37526 15302
rect 4582 14882 4610 14910
rect 4634 14882 4662 14910
rect 4686 14882 4714 14910
rect 4738 14882 4766 14910
rect 4790 14882 4818 14910
rect 4842 14882 4870 14910
rect 4894 14882 4922 14910
rect 4946 14882 4974 14910
rect 4998 14882 5026 14910
rect 9582 14882 9610 14910
rect 9634 14882 9662 14910
rect 9686 14882 9714 14910
rect 9738 14882 9766 14910
rect 9790 14882 9818 14910
rect 9842 14882 9870 14910
rect 9894 14882 9922 14910
rect 9946 14882 9974 14910
rect 9998 14882 10026 14910
rect 14582 14882 14610 14910
rect 14634 14882 14662 14910
rect 14686 14882 14714 14910
rect 14738 14882 14766 14910
rect 14790 14882 14818 14910
rect 14842 14882 14870 14910
rect 14894 14882 14922 14910
rect 14946 14882 14974 14910
rect 14998 14882 15026 14910
rect 19582 14882 19610 14910
rect 19634 14882 19662 14910
rect 19686 14882 19714 14910
rect 19738 14882 19766 14910
rect 19790 14882 19818 14910
rect 19842 14882 19870 14910
rect 19894 14882 19922 14910
rect 19946 14882 19974 14910
rect 19998 14882 20026 14910
rect 24582 14882 24610 14910
rect 24634 14882 24662 14910
rect 24686 14882 24714 14910
rect 24738 14882 24766 14910
rect 24790 14882 24818 14910
rect 24842 14882 24870 14910
rect 24894 14882 24922 14910
rect 24946 14882 24974 14910
rect 24998 14882 25026 14910
rect 29582 14882 29610 14910
rect 29634 14882 29662 14910
rect 29686 14882 29714 14910
rect 29738 14882 29766 14910
rect 29790 14882 29818 14910
rect 29842 14882 29870 14910
rect 29894 14882 29922 14910
rect 29946 14882 29974 14910
rect 29998 14882 30026 14910
rect 34582 14882 34610 14910
rect 34634 14882 34662 14910
rect 34686 14882 34714 14910
rect 34738 14882 34766 14910
rect 34790 14882 34818 14910
rect 34842 14882 34870 14910
rect 34894 14882 34922 14910
rect 34946 14882 34974 14910
rect 34998 14882 35026 14910
rect 2082 14490 2110 14518
rect 2134 14490 2162 14518
rect 2186 14490 2214 14518
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 2394 14490 2422 14518
rect 2446 14490 2474 14518
rect 2498 14490 2526 14518
rect 7082 14490 7110 14518
rect 7134 14490 7162 14518
rect 7186 14490 7214 14518
rect 7238 14490 7266 14518
rect 7290 14490 7318 14518
rect 7342 14490 7370 14518
rect 7394 14490 7422 14518
rect 7446 14490 7474 14518
rect 7498 14490 7526 14518
rect 12082 14490 12110 14518
rect 12134 14490 12162 14518
rect 12186 14490 12214 14518
rect 12238 14490 12266 14518
rect 12290 14490 12318 14518
rect 12342 14490 12370 14518
rect 12394 14490 12422 14518
rect 12446 14490 12474 14518
rect 12498 14490 12526 14518
rect 17082 14490 17110 14518
rect 17134 14490 17162 14518
rect 17186 14490 17214 14518
rect 17238 14490 17266 14518
rect 17290 14490 17318 14518
rect 17342 14490 17370 14518
rect 17394 14490 17422 14518
rect 17446 14490 17474 14518
rect 17498 14490 17526 14518
rect 22082 14490 22110 14518
rect 22134 14490 22162 14518
rect 22186 14490 22214 14518
rect 22238 14490 22266 14518
rect 22290 14490 22318 14518
rect 22342 14490 22370 14518
rect 22394 14490 22422 14518
rect 22446 14490 22474 14518
rect 22498 14490 22526 14518
rect 27082 14490 27110 14518
rect 27134 14490 27162 14518
rect 27186 14490 27214 14518
rect 27238 14490 27266 14518
rect 27290 14490 27318 14518
rect 27342 14490 27370 14518
rect 27394 14490 27422 14518
rect 27446 14490 27474 14518
rect 27498 14490 27526 14518
rect 32082 14490 32110 14518
rect 32134 14490 32162 14518
rect 32186 14490 32214 14518
rect 32238 14490 32266 14518
rect 32290 14490 32318 14518
rect 32342 14490 32370 14518
rect 32394 14490 32422 14518
rect 32446 14490 32474 14518
rect 32498 14490 32526 14518
rect 37082 14490 37110 14518
rect 37134 14490 37162 14518
rect 37186 14490 37214 14518
rect 37238 14490 37266 14518
rect 37290 14490 37318 14518
rect 37342 14490 37370 14518
rect 37394 14490 37422 14518
rect 37446 14490 37474 14518
rect 37498 14490 37526 14518
rect 4582 14098 4610 14126
rect 4634 14098 4662 14126
rect 4686 14098 4714 14126
rect 4738 14098 4766 14126
rect 4790 14098 4818 14126
rect 4842 14098 4870 14126
rect 4894 14098 4922 14126
rect 4946 14098 4974 14126
rect 4998 14098 5026 14126
rect 9582 14098 9610 14126
rect 9634 14098 9662 14126
rect 9686 14098 9714 14126
rect 9738 14098 9766 14126
rect 9790 14098 9818 14126
rect 9842 14098 9870 14126
rect 9894 14098 9922 14126
rect 9946 14098 9974 14126
rect 9998 14098 10026 14126
rect 14582 14098 14610 14126
rect 14634 14098 14662 14126
rect 14686 14098 14714 14126
rect 14738 14098 14766 14126
rect 14790 14098 14818 14126
rect 14842 14098 14870 14126
rect 14894 14098 14922 14126
rect 14946 14098 14974 14126
rect 14998 14098 15026 14126
rect 19582 14098 19610 14126
rect 19634 14098 19662 14126
rect 19686 14098 19714 14126
rect 19738 14098 19766 14126
rect 19790 14098 19818 14126
rect 19842 14098 19870 14126
rect 19894 14098 19922 14126
rect 19946 14098 19974 14126
rect 19998 14098 20026 14126
rect 24582 14098 24610 14126
rect 24634 14098 24662 14126
rect 24686 14098 24714 14126
rect 24738 14098 24766 14126
rect 24790 14098 24818 14126
rect 24842 14098 24870 14126
rect 24894 14098 24922 14126
rect 24946 14098 24974 14126
rect 24998 14098 25026 14126
rect 29582 14098 29610 14126
rect 29634 14098 29662 14126
rect 29686 14098 29714 14126
rect 29738 14098 29766 14126
rect 29790 14098 29818 14126
rect 29842 14098 29870 14126
rect 29894 14098 29922 14126
rect 29946 14098 29974 14126
rect 29998 14098 30026 14126
rect 34582 14098 34610 14126
rect 34634 14098 34662 14126
rect 34686 14098 34714 14126
rect 34738 14098 34766 14126
rect 34790 14098 34818 14126
rect 34842 14098 34870 14126
rect 34894 14098 34922 14126
rect 34946 14098 34974 14126
rect 34998 14098 35026 14126
rect 2082 13706 2110 13734
rect 2134 13706 2162 13734
rect 2186 13706 2214 13734
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 2394 13706 2422 13734
rect 2446 13706 2474 13734
rect 2498 13706 2526 13734
rect 7082 13706 7110 13734
rect 7134 13706 7162 13734
rect 7186 13706 7214 13734
rect 7238 13706 7266 13734
rect 7290 13706 7318 13734
rect 7342 13706 7370 13734
rect 7394 13706 7422 13734
rect 7446 13706 7474 13734
rect 7498 13706 7526 13734
rect 12082 13706 12110 13734
rect 12134 13706 12162 13734
rect 12186 13706 12214 13734
rect 12238 13706 12266 13734
rect 12290 13706 12318 13734
rect 12342 13706 12370 13734
rect 12394 13706 12422 13734
rect 12446 13706 12474 13734
rect 12498 13706 12526 13734
rect 17082 13706 17110 13734
rect 17134 13706 17162 13734
rect 17186 13706 17214 13734
rect 17238 13706 17266 13734
rect 17290 13706 17318 13734
rect 17342 13706 17370 13734
rect 17394 13706 17422 13734
rect 17446 13706 17474 13734
rect 17498 13706 17526 13734
rect 22082 13706 22110 13734
rect 22134 13706 22162 13734
rect 22186 13706 22214 13734
rect 22238 13706 22266 13734
rect 22290 13706 22318 13734
rect 22342 13706 22370 13734
rect 22394 13706 22422 13734
rect 22446 13706 22474 13734
rect 22498 13706 22526 13734
rect 27082 13706 27110 13734
rect 27134 13706 27162 13734
rect 27186 13706 27214 13734
rect 27238 13706 27266 13734
rect 27290 13706 27318 13734
rect 27342 13706 27370 13734
rect 27394 13706 27422 13734
rect 27446 13706 27474 13734
rect 27498 13706 27526 13734
rect 32082 13706 32110 13734
rect 32134 13706 32162 13734
rect 32186 13706 32214 13734
rect 32238 13706 32266 13734
rect 32290 13706 32318 13734
rect 32342 13706 32370 13734
rect 32394 13706 32422 13734
rect 32446 13706 32474 13734
rect 32498 13706 32526 13734
rect 37082 13706 37110 13734
rect 37134 13706 37162 13734
rect 37186 13706 37214 13734
rect 37238 13706 37266 13734
rect 37290 13706 37318 13734
rect 37342 13706 37370 13734
rect 37394 13706 37422 13734
rect 37446 13706 37474 13734
rect 37498 13706 37526 13734
rect 4582 13314 4610 13342
rect 4634 13314 4662 13342
rect 4686 13314 4714 13342
rect 4738 13314 4766 13342
rect 4790 13314 4818 13342
rect 4842 13314 4870 13342
rect 4894 13314 4922 13342
rect 4946 13314 4974 13342
rect 4998 13314 5026 13342
rect 9582 13314 9610 13342
rect 9634 13314 9662 13342
rect 9686 13314 9714 13342
rect 9738 13314 9766 13342
rect 9790 13314 9818 13342
rect 9842 13314 9870 13342
rect 9894 13314 9922 13342
rect 9946 13314 9974 13342
rect 9998 13314 10026 13342
rect 14582 13314 14610 13342
rect 14634 13314 14662 13342
rect 14686 13314 14714 13342
rect 14738 13314 14766 13342
rect 14790 13314 14818 13342
rect 14842 13314 14870 13342
rect 14894 13314 14922 13342
rect 14946 13314 14974 13342
rect 14998 13314 15026 13342
rect 19582 13314 19610 13342
rect 19634 13314 19662 13342
rect 19686 13314 19714 13342
rect 19738 13314 19766 13342
rect 19790 13314 19818 13342
rect 19842 13314 19870 13342
rect 19894 13314 19922 13342
rect 19946 13314 19974 13342
rect 19998 13314 20026 13342
rect 24582 13314 24610 13342
rect 24634 13314 24662 13342
rect 24686 13314 24714 13342
rect 24738 13314 24766 13342
rect 24790 13314 24818 13342
rect 24842 13314 24870 13342
rect 24894 13314 24922 13342
rect 24946 13314 24974 13342
rect 24998 13314 25026 13342
rect 29582 13314 29610 13342
rect 29634 13314 29662 13342
rect 29686 13314 29714 13342
rect 29738 13314 29766 13342
rect 29790 13314 29818 13342
rect 29842 13314 29870 13342
rect 29894 13314 29922 13342
rect 29946 13314 29974 13342
rect 29998 13314 30026 13342
rect 34582 13314 34610 13342
rect 34634 13314 34662 13342
rect 34686 13314 34714 13342
rect 34738 13314 34766 13342
rect 34790 13314 34818 13342
rect 34842 13314 34870 13342
rect 34894 13314 34922 13342
rect 34946 13314 34974 13342
rect 34998 13314 35026 13342
rect 2082 12922 2110 12950
rect 2134 12922 2162 12950
rect 2186 12922 2214 12950
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 2394 12922 2422 12950
rect 2446 12922 2474 12950
rect 2498 12922 2526 12950
rect 7082 12922 7110 12950
rect 7134 12922 7162 12950
rect 7186 12922 7214 12950
rect 7238 12922 7266 12950
rect 7290 12922 7318 12950
rect 7342 12922 7370 12950
rect 7394 12922 7422 12950
rect 7446 12922 7474 12950
rect 7498 12922 7526 12950
rect 12082 12922 12110 12950
rect 12134 12922 12162 12950
rect 12186 12922 12214 12950
rect 12238 12922 12266 12950
rect 12290 12922 12318 12950
rect 12342 12922 12370 12950
rect 12394 12922 12422 12950
rect 12446 12922 12474 12950
rect 12498 12922 12526 12950
rect 17082 12922 17110 12950
rect 17134 12922 17162 12950
rect 17186 12922 17214 12950
rect 17238 12922 17266 12950
rect 17290 12922 17318 12950
rect 17342 12922 17370 12950
rect 17394 12922 17422 12950
rect 17446 12922 17474 12950
rect 17498 12922 17526 12950
rect 22082 12922 22110 12950
rect 22134 12922 22162 12950
rect 22186 12922 22214 12950
rect 22238 12922 22266 12950
rect 22290 12922 22318 12950
rect 22342 12922 22370 12950
rect 22394 12922 22422 12950
rect 22446 12922 22474 12950
rect 22498 12922 22526 12950
rect 27082 12922 27110 12950
rect 27134 12922 27162 12950
rect 27186 12922 27214 12950
rect 27238 12922 27266 12950
rect 27290 12922 27318 12950
rect 27342 12922 27370 12950
rect 27394 12922 27422 12950
rect 27446 12922 27474 12950
rect 27498 12922 27526 12950
rect 32082 12922 32110 12950
rect 32134 12922 32162 12950
rect 32186 12922 32214 12950
rect 32238 12922 32266 12950
rect 32290 12922 32318 12950
rect 32342 12922 32370 12950
rect 32394 12922 32422 12950
rect 32446 12922 32474 12950
rect 32498 12922 32526 12950
rect 37082 12922 37110 12950
rect 37134 12922 37162 12950
rect 37186 12922 37214 12950
rect 37238 12922 37266 12950
rect 37290 12922 37318 12950
rect 37342 12922 37370 12950
rect 37394 12922 37422 12950
rect 37446 12922 37474 12950
rect 37498 12922 37526 12950
rect 4582 12530 4610 12558
rect 4634 12530 4662 12558
rect 4686 12530 4714 12558
rect 4738 12530 4766 12558
rect 4790 12530 4818 12558
rect 4842 12530 4870 12558
rect 4894 12530 4922 12558
rect 4946 12530 4974 12558
rect 4998 12530 5026 12558
rect 9582 12530 9610 12558
rect 9634 12530 9662 12558
rect 9686 12530 9714 12558
rect 9738 12530 9766 12558
rect 9790 12530 9818 12558
rect 9842 12530 9870 12558
rect 9894 12530 9922 12558
rect 9946 12530 9974 12558
rect 9998 12530 10026 12558
rect 14582 12530 14610 12558
rect 14634 12530 14662 12558
rect 14686 12530 14714 12558
rect 14738 12530 14766 12558
rect 14790 12530 14818 12558
rect 14842 12530 14870 12558
rect 14894 12530 14922 12558
rect 14946 12530 14974 12558
rect 14998 12530 15026 12558
rect 19582 12530 19610 12558
rect 19634 12530 19662 12558
rect 19686 12530 19714 12558
rect 19738 12530 19766 12558
rect 19790 12530 19818 12558
rect 19842 12530 19870 12558
rect 19894 12530 19922 12558
rect 19946 12530 19974 12558
rect 19998 12530 20026 12558
rect 24582 12530 24610 12558
rect 24634 12530 24662 12558
rect 24686 12530 24714 12558
rect 24738 12530 24766 12558
rect 24790 12530 24818 12558
rect 24842 12530 24870 12558
rect 24894 12530 24922 12558
rect 24946 12530 24974 12558
rect 24998 12530 25026 12558
rect 29582 12530 29610 12558
rect 29634 12530 29662 12558
rect 29686 12530 29714 12558
rect 29738 12530 29766 12558
rect 29790 12530 29818 12558
rect 29842 12530 29870 12558
rect 29894 12530 29922 12558
rect 29946 12530 29974 12558
rect 29998 12530 30026 12558
rect 34582 12530 34610 12558
rect 34634 12530 34662 12558
rect 34686 12530 34714 12558
rect 34738 12530 34766 12558
rect 34790 12530 34818 12558
rect 34842 12530 34870 12558
rect 34894 12530 34922 12558
rect 34946 12530 34974 12558
rect 34998 12530 35026 12558
rect 2082 12138 2110 12166
rect 2134 12138 2162 12166
rect 2186 12138 2214 12166
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 2394 12138 2422 12166
rect 2446 12138 2474 12166
rect 2498 12138 2526 12166
rect 7082 12138 7110 12166
rect 7134 12138 7162 12166
rect 7186 12138 7214 12166
rect 7238 12138 7266 12166
rect 7290 12138 7318 12166
rect 7342 12138 7370 12166
rect 7394 12138 7422 12166
rect 7446 12138 7474 12166
rect 7498 12138 7526 12166
rect 12082 12138 12110 12166
rect 12134 12138 12162 12166
rect 12186 12138 12214 12166
rect 12238 12138 12266 12166
rect 12290 12138 12318 12166
rect 12342 12138 12370 12166
rect 12394 12138 12422 12166
rect 12446 12138 12474 12166
rect 12498 12138 12526 12166
rect 17082 12138 17110 12166
rect 17134 12138 17162 12166
rect 17186 12138 17214 12166
rect 17238 12138 17266 12166
rect 17290 12138 17318 12166
rect 17342 12138 17370 12166
rect 17394 12138 17422 12166
rect 17446 12138 17474 12166
rect 17498 12138 17526 12166
rect 22082 12138 22110 12166
rect 22134 12138 22162 12166
rect 22186 12138 22214 12166
rect 22238 12138 22266 12166
rect 22290 12138 22318 12166
rect 22342 12138 22370 12166
rect 22394 12138 22422 12166
rect 22446 12138 22474 12166
rect 22498 12138 22526 12166
rect 27082 12138 27110 12166
rect 27134 12138 27162 12166
rect 27186 12138 27214 12166
rect 27238 12138 27266 12166
rect 27290 12138 27318 12166
rect 27342 12138 27370 12166
rect 27394 12138 27422 12166
rect 27446 12138 27474 12166
rect 27498 12138 27526 12166
rect 32082 12138 32110 12166
rect 32134 12138 32162 12166
rect 32186 12138 32214 12166
rect 32238 12138 32266 12166
rect 32290 12138 32318 12166
rect 32342 12138 32370 12166
rect 32394 12138 32422 12166
rect 32446 12138 32474 12166
rect 32498 12138 32526 12166
rect 37082 12138 37110 12166
rect 37134 12138 37162 12166
rect 37186 12138 37214 12166
rect 37238 12138 37266 12166
rect 37290 12138 37318 12166
rect 37342 12138 37370 12166
rect 37394 12138 37422 12166
rect 37446 12138 37474 12166
rect 37498 12138 37526 12166
rect 4582 11746 4610 11774
rect 4634 11746 4662 11774
rect 4686 11746 4714 11774
rect 4738 11746 4766 11774
rect 4790 11746 4818 11774
rect 4842 11746 4870 11774
rect 4894 11746 4922 11774
rect 4946 11746 4974 11774
rect 4998 11746 5026 11774
rect 9582 11746 9610 11774
rect 9634 11746 9662 11774
rect 9686 11746 9714 11774
rect 9738 11746 9766 11774
rect 9790 11746 9818 11774
rect 9842 11746 9870 11774
rect 9894 11746 9922 11774
rect 9946 11746 9974 11774
rect 9998 11746 10026 11774
rect 14582 11746 14610 11774
rect 14634 11746 14662 11774
rect 14686 11746 14714 11774
rect 14738 11746 14766 11774
rect 14790 11746 14818 11774
rect 14842 11746 14870 11774
rect 14894 11746 14922 11774
rect 14946 11746 14974 11774
rect 14998 11746 15026 11774
rect 19582 11746 19610 11774
rect 19634 11746 19662 11774
rect 19686 11746 19714 11774
rect 19738 11746 19766 11774
rect 19790 11746 19818 11774
rect 19842 11746 19870 11774
rect 19894 11746 19922 11774
rect 19946 11746 19974 11774
rect 19998 11746 20026 11774
rect 24582 11746 24610 11774
rect 24634 11746 24662 11774
rect 24686 11746 24714 11774
rect 24738 11746 24766 11774
rect 24790 11746 24818 11774
rect 24842 11746 24870 11774
rect 24894 11746 24922 11774
rect 24946 11746 24974 11774
rect 24998 11746 25026 11774
rect 29582 11746 29610 11774
rect 29634 11746 29662 11774
rect 29686 11746 29714 11774
rect 29738 11746 29766 11774
rect 29790 11746 29818 11774
rect 29842 11746 29870 11774
rect 29894 11746 29922 11774
rect 29946 11746 29974 11774
rect 29998 11746 30026 11774
rect 34582 11746 34610 11774
rect 34634 11746 34662 11774
rect 34686 11746 34714 11774
rect 34738 11746 34766 11774
rect 34790 11746 34818 11774
rect 34842 11746 34870 11774
rect 34894 11746 34922 11774
rect 34946 11746 34974 11774
rect 34998 11746 35026 11774
rect 2082 11354 2110 11382
rect 2134 11354 2162 11382
rect 2186 11354 2214 11382
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 2394 11354 2422 11382
rect 2446 11354 2474 11382
rect 2498 11354 2526 11382
rect 7082 11354 7110 11382
rect 7134 11354 7162 11382
rect 7186 11354 7214 11382
rect 7238 11354 7266 11382
rect 7290 11354 7318 11382
rect 7342 11354 7370 11382
rect 7394 11354 7422 11382
rect 7446 11354 7474 11382
rect 7498 11354 7526 11382
rect 12082 11354 12110 11382
rect 12134 11354 12162 11382
rect 12186 11354 12214 11382
rect 12238 11354 12266 11382
rect 12290 11354 12318 11382
rect 12342 11354 12370 11382
rect 12394 11354 12422 11382
rect 12446 11354 12474 11382
rect 12498 11354 12526 11382
rect 17082 11354 17110 11382
rect 17134 11354 17162 11382
rect 17186 11354 17214 11382
rect 17238 11354 17266 11382
rect 17290 11354 17318 11382
rect 17342 11354 17370 11382
rect 17394 11354 17422 11382
rect 17446 11354 17474 11382
rect 17498 11354 17526 11382
rect 22082 11354 22110 11382
rect 22134 11354 22162 11382
rect 22186 11354 22214 11382
rect 22238 11354 22266 11382
rect 22290 11354 22318 11382
rect 22342 11354 22370 11382
rect 22394 11354 22422 11382
rect 22446 11354 22474 11382
rect 22498 11354 22526 11382
rect 27082 11354 27110 11382
rect 27134 11354 27162 11382
rect 27186 11354 27214 11382
rect 27238 11354 27266 11382
rect 27290 11354 27318 11382
rect 27342 11354 27370 11382
rect 27394 11354 27422 11382
rect 27446 11354 27474 11382
rect 27498 11354 27526 11382
rect 32082 11354 32110 11382
rect 32134 11354 32162 11382
rect 32186 11354 32214 11382
rect 32238 11354 32266 11382
rect 32290 11354 32318 11382
rect 32342 11354 32370 11382
rect 32394 11354 32422 11382
rect 32446 11354 32474 11382
rect 32498 11354 32526 11382
rect 37082 11354 37110 11382
rect 37134 11354 37162 11382
rect 37186 11354 37214 11382
rect 37238 11354 37266 11382
rect 37290 11354 37318 11382
rect 37342 11354 37370 11382
rect 37394 11354 37422 11382
rect 37446 11354 37474 11382
rect 37498 11354 37526 11382
rect 4582 10962 4610 10990
rect 4634 10962 4662 10990
rect 4686 10962 4714 10990
rect 4738 10962 4766 10990
rect 4790 10962 4818 10990
rect 4842 10962 4870 10990
rect 4894 10962 4922 10990
rect 4946 10962 4974 10990
rect 4998 10962 5026 10990
rect 9582 10962 9610 10990
rect 9634 10962 9662 10990
rect 9686 10962 9714 10990
rect 9738 10962 9766 10990
rect 9790 10962 9818 10990
rect 9842 10962 9870 10990
rect 9894 10962 9922 10990
rect 9946 10962 9974 10990
rect 9998 10962 10026 10990
rect 14582 10962 14610 10990
rect 14634 10962 14662 10990
rect 14686 10962 14714 10990
rect 14738 10962 14766 10990
rect 14790 10962 14818 10990
rect 14842 10962 14870 10990
rect 14894 10962 14922 10990
rect 14946 10962 14974 10990
rect 14998 10962 15026 10990
rect 19582 10962 19610 10990
rect 19634 10962 19662 10990
rect 19686 10962 19714 10990
rect 19738 10962 19766 10990
rect 19790 10962 19818 10990
rect 19842 10962 19870 10990
rect 19894 10962 19922 10990
rect 19946 10962 19974 10990
rect 19998 10962 20026 10990
rect 24582 10962 24610 10990
rect 24634 10962 24662 10990
rect 24686 10962 24714 10990
rect 24738 10962 24766 10990
rect 24790 10962 24818 10990
rect 24842 10962 24870 10990
rect 24894 10962 24922 10990
rect 24946 10962 24974 10990
rect 24998 10962 25026 10990
rect 29582 10962 29610 10990
rect 29634 10962 29662 10990
rect 29686 10962 29714 10990
rect 29738 10962 29766 10990
rect 29790 10962 29818 10990
rect 29842 10962 29870 10990
rect 29894 10962 29922 10990
rect 29946 10962 29974 10990
rect 29998 10962 30026 10990
rect 34582 10962 34610 10990
rect 34634 10962 34662 10990
rect 34686 10962 34714 10990
rect 34738 10962 34766 10990
rect 34790 10962 34818 10990
rect 34842 10962 34870 10990
rect 34894 10962 34922 10990
rect 34946 10962 34974 10990
rect 34998 10962 35026 10990
rect 2082 10570 2110 10598
rect 2134 10570 2162 10598
rect 2186 10570 2214 10598
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 2394 10570 2422 10598
rect 2446 10570 2474 10598
rect 2498 10570 2526 10598
rect 7082 10570 7110 10598
rect 7134 10570 7162 10598
rect 7186 10570 7214 10598
rect 7238 10570 7266 10598
rect 7290 10570 7318 10598
rect 7342 10570 7370 10598
rect 7394 10570 7422 10598
rect 7446 10570 7474 10598
rect 7498 10570 7526 10598
rect 12082 10570 12110 10598
rect 12134 10570 12162 10598
rect 12186 10570 12214 10598
rect 12238 10570 12266 10598
rect 12290 10570 12318 10598
rect 12342 10570 12370 10598
rect 12394 10570 12422 10598
rect 12446 10570 12474 10598
rect 12498 10570 12526 10598
rect 17082 10570 17110 10598
rect 17134 10570 17162 10598
rect 17186 10570 17214 10598
rect 17238 10570 17266 10598
rect 17290 10570 17318 10598
rect 17342 10570 17370 10598
rect 17394 10570 17422 10598
rect 17446 10570 17474 10598
rect 17498 10570 17526 10598
rect 22082 10570 22110 10598
rect 22134 10570 22162 10598
rect 22186 10570 22214 10598
rect 22238 10570 22266 10598
rect 22290 10570 22318 10598
rect 22342 10570 22370 10598
rect 22394 10570 22422 10598
rect 22446 10570 22474 10598
rect 22498 10570 22526 10598
rect 27082 10570 27110 10598
rect 27134 10570 27162 10598
rect 27186 10570 27214 10598
rect 27238 10570 27266 10598
rect 27290 10570 27318 10598
rect 27342 10570 27370 10598
rect 27394 10570 27422 10598
rect 27446 10570 27474 10598
rect 27498 10570 27526 10598
rect 32082 10570 32110 10598
rect 32134 10570 32162 10598
rect 32186 10570 32214 10598
rect 32238 10570 32266 10598
rect 32290 10570 32318 10598
rect 32342 10570 32370 10598
rect 32394 10570 32422 10598
rect 32446 10570 32474 10598
rect 32498 10570 32526 10598
rect 37082 10570 37110 10598
rect 37134 10570 37162 10598
rect 37186 10570 37214 10598
rect 37238 10570 37266 10598
rect 37290 10570 37318 10598
rect 37342 10570 37370 10598
rect 37394 10570 37422 10598
rect 37446 10570 37474 10598
rect 37498 10570 37526 10598
rect 4582 10178 4610 10206
rect 4634 10178 4662 10206
rect 4686 10178 4714 10206
rect 4738 10178 4766 10206
rect 4790 10178 4818 10206
rect 4842 10178 4870 10206
rect 4894 10178 4922 10206
rect 4946 10178 4974 10206
rect 4998 10178 5026 10206
rect 9582 10178 9610 10206
rect 9634 10178 9662 10206
rect 9686 10178 9714 10206
rect 9738 10178 9766 10206
rect 9790 10178 9818 10206
rect 9842 10178 9870 10206
rect 9894 10178 9922 10206
rect 9946 10178 9974 10206
rect 9998 10178 10026 10206
rect 14582 10178 14610 10206
rect 14634 10178 14662 10206
rect 14686 10178 14714 10206
rect 14738 10178 14766 10206
rect 14790 10178 14818 10206
rect 14842 10178 14870 10206
rect 14894 10178 14922 10206
rect 14946 10178 14974 10206
rect 14998 10178 15026 10206
rect 19582 10178 19610 10206
rect 19634 10178 19662 10206
rect 19686 10178 19714 10206
rect 19738 10178 19766 10206
rect 19790 10178 19818 10206
rect 19842 10178 19870 10206
rect 19894 10178 19922 10206
rect 19946 10178 19974 10206
rect 19998 10178 20026 10206
rect 24582 10178 24610 10206
rect 24634 10178 24662 10206
rect 24686 10178 24714 10206
rect 24738 10178 24766 10206
rect 24790 10178 24818 10206
rect 24842 10178 24870 10206
rect 24894 10178 24922 10206
rect 24946 10178 24974 10206
rect 24998 10178 25026 10206
rect 29582 10178 29610 10206
rect 29634 10178 29662 10206
rect 29686 10178 29714 10206
rect 29738 10178 29766 10206
rect 29790 10178 29818 10206
rect 29842 10178 29870 10206
rect 29894 10178 29922 10206
rect 29946 10178 29974 10206
rect 29998 10178 30026 10206
rect 34582 10178 34610 10206
rect 34634 10178 34662 10206
rect 34686 10178 34714 10206
rect 34738 10178 34766 10206
rect 34790 10178 34818 10206
rect 34842 10178 34870 10206
rect 34894 10178 34922 10206
rect 34946 10178 34974 10206
rect 34998 10178 35026 10206
rect 2082 9786 2110 9814
rect 2134 9786 2162 9814
rect 2186 9786 2214 9814
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 2394 9786 2422 9814
rect 2446 9786 2474 9814
rect 2498 9786 2526 9814
rect 7082 9786 7110 9814
rect 7134 9786 7162 9814
rect 7186 9786 7214 9814
rect 7238 9786 7266 9814
rect 7290 9786 7318 9814
rect 7342 9786 7370 9814
rect 7394 9786 7422 9814
rect 7446 9786 7474 9814
rect 7498 9786 7526 9814
rect 12082 9786 12110 9814
rect 12134 9786 12162 9814
rect 12186 9786 12214 9814
rect 12238 9786 12266 9814
rect 12290 9786 12318 9814
rect 12342 9786 12370 9814
rect 12394 9786 12422 9814
rect 12446 9786 12474 9814
rect 12498 9786 12526 9814
rect 17082 9786 17110 9814
rect 17134 9786 17162 9814
rect 17186 9786 17214 9814
rect 17238 9786 17266 9814
rect 17290 9786 17318 9814
rect 17342 9786 17370 9814
rect 17394 9786 17422 9814
rect 17446 9786 17474 9814
rect 17498 9786 17526 9814
rect 22082 9786 22110 9814
rect 22134 9786 22162 9814
rect 22186 9786 22214 9814
rect 22238 9786 22266 9814
rect 22290 9786 22318 9814
rect 22342 9786 22370 9814
rect 22394 9786 22422 9814
rect 22446 9786 22474 9814
rect 22498 9786 22526 9814
rect 27082 9786 27110 9814
rect 27134 9786 27162 9814
rect 27186 9786 27214 9814
rect 27238 9786 27266 9814
rect 27290 9786 27318 9814
rect 27342 9786 27370 9814
rect 27394 9786 27422 9814
rect 27446 9786 27474 9814
rect 27498 9786 27526 9814
rect 32082 9786 32110 9814
rect 32134 9786 32162 9814
rect 32186 9786 32214 9814
rect 32238 9786 32266 9814
rect 32290 9786 32318 9814
rect 32342 9786 32370 9814
rect 32394 9786 32422 9814
rect 32446 9786 32474 9814
rect 32498 9786 32526 9814
rect 37082 9786 37110 9814
rect 37134 9786 37162 9814
rect 37186 9786 37214 9814
rect 37238 9786 37266 9814
rect 37290 9786 37318 9814
rect 37342 9786 37370 9814
rect 37394 9786 37422 9814
rect 37446 9786 37474 9814
rect 37498 9786 37526 9814
rect 4582 9394 4610 9422
rect 4634 9394 4662 9422
rect 4686 9394 4714 9422
rect 4738 9394 4766 9422
rect 4790 9394 4818 9422
rect 4842 9394 4870 9422
rect 4894 9394 4922 9422
rect 4946 9394 4974 9422
rect 4998 9394 5026 9422
rect 9582 9394 9610 9422
rect 9634 9394 9662 9422
rect 9686 9394 9714 9422
rect 9738 9394 9766 9422
rect 9790 9394 9818 9422
rect 9842 9394 9870 9422
rect 9894 9394 9922 9422
rect 9946 9394 9974 9422
rect 9998 9394 10026 9422
rect 14582 9394 14610 9422
rect 14634 9394 14662 9422
rect 14686 9394 14714 9422
rect 14738 9394 14766 9422
rect 14790 9394 14818 9422
rect 14842 9394 14870 9422
rect 14894 9394 14922 9422
rect 14946 9394 14974 9422
rect 14998 9394 15026 9422
rect 19582 9394 19610 9422
rect 19634 9394 19662 9422
rect 19686 9394 19714 9422
rect 19738 9394 19766 9422
rect 19790 9394 19818 9422
rect 19842 9394 19870 9422
rect 19894 9394 19922 9422
rect 19946 9394 19974 9422
rect 19998 9394 20026 9422
rect 24582 9394 24610 9422
rect 24634 9394 24662 9422
rect 24686 9394 24714 9422
rect 24738 9394 24766 9422
rect 24790 9394 24818 9422
rect 24842 9394 24870 9422
rect 24894 9394 24922 9422
rect 24946 9394 24974 9422
rect 24998 9394 25026 9422
rect 29582 9394 29610 9422
rect 29634 9394 29662 9422
rect 29686 9394 29714 9422
rect 29738 9394 29766 9422
rect 29790 9394 29818 9422
rect 29842 9394 29870 9422
rect 29894 9394 29922 9422
rect 29946 9394 29974 9422
rect 29998 9394 30026 9422
rect 34582 9394 34610 9422
rect 34634 9394 34662 9422
rect 34686 9394 34714 9422
rect 34738 9394 34766 9422
rect 34790 9394 34818 9422
rect 34842 9394 34870 9422
rect 34894 9394 34922 9422
rect 34946 9394 34974 9422
rect 34998 9394 35026 9422
rect 2082 9002 2110 9030
rect 2134 9002 2162 9030
rect 2186 9002 2214 9030
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 2394 9002 2422 9030
rect 2446 9002 2474 9030
rect 2498 9002 2526 9030
rect 7082 9002 7110 9030
rect 7134 9002 7162 9030
rect 7186 9002 7214 9030
rect 7238 9002 7266 9030
rect 7290 9002 7318 9030
rect 7342 9002 7370 9030
rect 7394 9002 7422 9030
rect 7446 9002 7474 9030
rect 7498 9002 7526 9030
rect 12082 9002 12110 9030
rect 12134 9002 12162 9030
rect 12186 9002 12214 9030
rect 12238 9002 12266 9030
rect 12290 9002 12318 9030
rect 12342 9002 12370 9030
rect 12394 9002 12422 9030
rect 12446 9002 12474 9030
rect 12498 9002 12526 9030
rect 17082 9002 17110 9030
rect 17134 9002 17162 9030
rect 17186 9002 17214 9030
rect 17238 9002 17266 9030
rect 17290 9002 17318 9030
rect 17342 9002 17370 9030
rect 17394 9002 17422 9030
rect 17446 9002 17474 9030
rect 17498 9002 17526 9030
rect 22082 9002 22110 9030
rect 22134 9002 22162 9030
rect 22186 9002 22214 9030
rect 22238 9002 22266 9030
rect 22290 9002 22318 9030
rect 22342 9002 22370 9030
rect 22394 9002 22422 9030
rect 22446 9002 22474 9030
rect 22498 9002 22526 9030
rect 27082 9002 27110 9030
rect 27134 9002 27162 9030
rect 27186 9002 27214 9030
rect 27238 9002 27266 9030
rect 27290 9002 27318 9030
rect 27342 9002 27370 9030
rect 27394 9002 27422 9030
rect 27446 9002 27474 9030
rect 27498 9002 27526 9030
rect 32082 9002 32110 9030
rect 32134 9002 32162 9030
rect 32186 9002 32214 9030
rect 32238 9002 32266 9030
rect 32290 9002 32318 9030
rect 32342 9002 32370 9030
rect 32394 9002 32422 9030
rect 32446 9002 32474 9030
rect 32498 9002 32526 9030
rect 37082 9002 37110 9030
rect 37134 9002 37162 9030
rect 37186 9002 37214 9030
rect 37238 9002 37266 9030
rect 37290 9002 37318 9030
rect 37342 9002 37370 9030
rect 37394 9002 37422 9030
rect 37446 9002 37474 9030
rect 37498 9002 37526 9030
rect 4582 8610 4610 8638
rect 4634 8610 4662 8638
rect 4686 8610 4714 8638
rect 4738 8610 4766 8638
rect 4790 8610 4818 8638
rect 4842 8610 4870 8638
rect 4894 8610 4922 8638
rect 4946 8610 4974 8638
rect 4998 8610 5026 8638
rect 9582 8610 9610 8638
rect 9634 8610 9662 8638
rect 9686 8610 9714 8638
rect 9738 8610 9766 8638
rect 9790 8610 9818 8638
rect 9842 8610 9870 8638
rect 9894 8610 9922 8638
rect 9946 8610 9974 8638
rect 9998 8610 10026 8638
rect 14582 8610 14610 8638
rect 14634 8610 14662 8638
rect 14686 8610 14714 8638
rect 14738 8610 14766 8638
rect 14790 8610 14818 8638
rect 14842 8610 14870 8638
rect 14894 8610 14922 8638
rect 14946 8610 14974 8638
rect 14998 8610 15026 8638
rect 19582 8610 19610 8638
rect 19634 8610 19662 8638
rect 19686 8610 19714 8638
rect 19738 8610 19766 8638
rect 19790 8610 19818 8638
rect 19842 8610 19870 8638
rect 19894 8610 19922 8638
rect 19946 8610 19974 8638
rect 19998 8610 20026 8638
rect 24582 8610 24610 8638
rect 24634 8610 24662 8638
rect 24686 8610 24714 8638
rect 24738 8610 24766 8638
rect 24790 8610 24818 8638
rect 24842 8610 24870 8638
rect 24894 8610 24922 8638
rect 24946 8610 24974 8638
rect 24998 8610 25026 8638
rect 29582 8610 29610 8638
rect 29634 8610 29662 8638
rect 29686 8610 29714 8638
rect 29738 8610 29766 8638
rect 29790 8610 29818 8638
rect 29842 8610 29870 8638
rect 29894 8610 29922 8638
rect 29946 8610 29974 8638
rect 29998 8610 30026 8638
rect 34582 8610 34610 8638
rect 34634 8610 34662 8638
rect 34686 8610 34714 8638
rect 34738 8610 34766 8638
rect 34790 8610 34818 8638
rect 34842 8610 34870 8638
rect 34894 8610 34922 8638
rect 34946 8610 34974 8638
rect 34998 8610 35026 8638
rect 31934 8526 31962 8554
rect 2082 8218 2110 8246
rect 2134 8218 2162 8246
rect 2186 8218 2214 8246
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 2394 8218 2422 8246
rect 2446 8218 2474 8246
rect 2498 8218 2526 8246
rect 7082 8218 7110 8246
rect 7134 8218 7162 8246
rect 7186 8218 7214 8246
rect 7238 8218 7266 8246
rect 7290 8218 7318 8246
rect 7342 8218 7370 8246
rect 7394 8218 7422 8246
rect 7446 8218 7474 8246
rect 7498 8218 7526 8246
rect 12082 8218 12110 8246
rect 12134 8218 12162 8246
rect 12186 8218 12214 8246
rect 12238 8218 12266 8246
rect 12290 8218 12318 8246
rect 12342 8218 12370 8246
rect 12394 8218 12422 8246
rect 12446 8218 12474 8246
rect 12498 8218 12526 8246
rect 17082 8218 17110 8246
rect 17134 8218 17162 8246
rect 17186 8218 17214 8246
rect 17238 8218 17266 8246
rect 17290 8218 17318 8246
rect 17342 8218 17370 8246
rect 17394 8218 17422 8246
rect 17446 8218 17474 8246
rect 17498 8218 17526 8246
rect 22082 8218 22110 8246
rect 22134 8218 22162 8246
rect 22186 8218 22214 8246
rect 22238 8218 22266 8246
rect 22290 8218 22318 8246
rect 22342 8218 22370 8246
rect 22394 8218 22422 8246
rect 22446 8218 22474 8246
rect 22498 8218 22526 8246
rect 27082 8218 27110 8246
rect 27134 8218 27162 8246
rect 27186 8218 27214 8246
rect 27238 8218 27266 8246
rect 27290 8218 27318 8246
rect 27342 8218 27370 8246
rect 27394 8218 27422 8246
rect 27446 8218 27474 8246
rect 27498 8218 27526 8246
rect 32082 8218 32110 8246
rect 32134 8218 32162 8246
rect 32186 8218 32214 8246
rect 32238 8218 32266 8246
rect 32290 8218 32318 8246
rect 32342 8218 32370 8246
rect 32394 8218 32422 8246
rect 32446 8218 32474 8246
rect 32498 8218 32526 8246
rect 37082 8218 37110 8246
rect 37134 8218 37162 8246
rect 37186 8218 37214 8246
rect 37238 8218 37266 8246
rect 37290 8218 37318 8246
rect 37342 8218 37370 8246
rect 37394 8218 37422 8246
rect 37446 8218 37474 8246
rect 37498 8218 37526 8246
rect 4582 7826 4610 7854
rect 4634 7826 4662 7854
rect 4686 7826 4714 7854
rect 4738 7826 4766 7854
rect 4790 7826 4818 7854
rect 4842 7826 4870 7854
rect 4894 7826 4922 7854
rect 4946 7826 4974 7854
rect 4998 7826 5026 7854
rect 9582 7826 9610 7854
rect 9634 7826 9662 7854
rect 9686 7826 9714 7854
rect 9738 7826 9766 7854
rect 9790 7826 9818 7854
rect 9842 7826 9870 7854
rect 9894 7826 9922 7854
rect 9946 7826 9974 7854
rect 9998 7826 10026 7854
rect 14582 7826 14610 7854
rect 14634 7826 14662 7854
rect 14686 7826 14714 7854
rect 14738 7826 14766 7854
rect 14790 7826 14818 7854
rect 14842 7826 14870 7854
rect 14894 7826 14922 7854
rect 14946 7826 14974 7854
rect 14998 7826 15026 7854
rect 19582 7826 19610 7854
rect 19634 7826 19662 7854
rect 19686 7826 19714 7854
rect 19738 7826 19766 7854
rect 19790 7826 19818 7854
rect 19842 7826 19870 7854
rect 19894 7826 19922 7854
rect 19946 7826 19974 7854
rect 19998 7826 20026 7854
rect 24582 7826 24610 7854
rect 24634 7826 24662 7854
rect 24686 7826 24714 7854
rect 24738 7826 24766 7854
rect 24790 7826 24818 7854
rect 24842 7826 24870 7854
rect 24894 7826 24922 7854
rect 24946 7826 24974 7854
rect 24998 7826 25026 7854
rect 29582 7826 29610 7854
rect 29634 7826 29662 7854
rect 29686 7826 29714 7854
rect 29738 7826 29766 7854
rect 29790 7826 29818 7854
rect 29842 7826 29870 7854
rect 29894 7826 29922 7854
rect 29946 7826 29974 7854
rect 29998 7826 30026 7854
rect 34582 7826 34610 7854
rect 34634 7826 34662 7854
rect 34686 7826 34714 7854
rect 34738 7826 34766 7854
rect 34790 7826 34818 7854
rect 34842 7826 34870 7854
rect 34894 7826 34922 7854
rect 34946 7826 34974 7854
rect 34998 7826 35026 7854
rect 31990 7630 32018 7658
rect 2082 7434 2110 7462
rect 2134 7434 2162 7462
rect 2186 7434 2214 7462
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 2394 7434 2422 7462
rect 2446 7434 2474 7462
rect 2498 7434 2526 7462
rect 7082 7434 7110 7462
rect 7134 7434 7162 7462
rect 7186 7434 7214 7462
rect 7238 7434 7266 7462
rect 7290 7434 7318 7462
rect 7342 7434 7370 7462
rect 7394 7434 7422 7462
rect 7446 7434 7474 7462
rect 7498 7434 7526 7462
rect 12082 7434 12110 7462
rect 12134 7434 12162 7462
rect 12186 7434 12214 7462
rect 12238 7434 12266 7462
rect 12290 7434 12318 7462
rect 12342 7434 12370 7462
rect 12394 7434 12422 7462
rect 12446 7434 12474 7462
rect 12498 7434 12526 7462
rect 17082 7434 17110 7462
rect 17134 7434 17162 7462
rect 17186 7434 17214 7462
rect 17238 7434 17266 7462
rect 17290 7434 17318 7462
rect 17342 7434 17370 7462
rect 17394 7434 17422 7462
rect 17446 7434 17474 7462
rect 17498 7434 17526 7462
rect 22082 7434 22110 7462
rect 22134 7434 22162 7462
rect 22186 7434 22214 7462
rect 22238 7434 22266 7462
rect 22290 7434 22318 7462
rect 22342 7434 22370 7462
rect 22394 7434 22422 7462
rect 22446 7434 22474 7462
rect 22498 7434 22526 7462
rect 27082 7434 27110 7462
rect 27134 7434 27162 7462
rect 27186 7434 27214 7462
rect 27238 7434 27266 7462
rect 27290 7434 27318 7462
rect 27342 7434 27370 7462
rect 27394 7434 27422 7462
rect 27446 7434 27474 7462
rect 27498 7434 27526 7462
rect 32082 7434 32110 7462
rect 32134 7434 32162 7462
rect 32186 7434 32214 7462
rect 32238 7434 32266 7462
rect 32290 7434 32318 7462
rect 32342 7434 32370 7462
rect 32394 7434 32422 7462
rect 32446 7434 32474 7462
rect 32498 7434 32526 7462
rect 37082 7434 37110 7462
rect 37134 7434 37162 7462
rect 37186 7434 37214 7462
rect 37238 7434 37266 7462
rect 37290 7434 37318 7462
rect 37342 7434 37370 7462
rect 37394 7434 37422 7462
rect 37446 7434 37474 7462
rect 37498 7434 37526 7462
rect 4582 7042 4610 7070
rect 4634 7042 4662 7070
rect 4686 7042 4714 7070
rect 4738 7042 4766 7070
rect 4790 7042 4818 7070
rect 4842 7042 4870 7070
rect 4894 7042 4922 7070
rect 4946 7042 4974 7070
rect 4998 7042 5026 7070
rect 9582 7042 9610 7070
rect 9634 7042 9662 7070
rect 9686 7042 9714 7070
rect 9738 7042 9766 7070
rect 9790 7042 9818 7070
rect 9842 7042 9870 7070
rect 9894 7042 9922 7070
rect 9946 7042 9974 7070
rect 9998 7042 10026 7070
rect 14582 7042 14610 7070
rect 14634 7042 14662 7070
rect 14686 7042 14714 7070
rect 14738 7042 14766 7070
rect 14790 7042 14818 7070
rect 14842 7042 14870 7070
rect 14894 7042 14922 7070
rect 14946 7042 14974 7070
rect 14998 7042 15026 7070
rect 19582 7042 19610 7070
rect 19634 7042 19662 7070
rect 19686 7042 19714 7070
rect 19738 7042 19766 7070
rect 19790 7042 19818 7070
rect 19842 7042 19870 7070
rect 19894 7042 19922 7070
rect 19946 7042 19974 7070
rect 19998 7042 20026 7070
rect 24582 7042 24610 7070
rect 24634 7042 24662 7070
rect 24686 7042 24714 7070
rect 24738 7042 24766 7070
rect 24790 7042 24818 7070
rect 24842 7042 24870 7070
rect 24894 7042 24922 7070
rect 24946 7042 24974 7070
rect 24998 7042 25026 7070
rect 29582 7042 29610 7070
rect 29634 7042 29662 7070
rect 29686 7042 29714 7070
rect 29738 7042 29766 7070
rect 29790 7042 29818 7070
rect 29842 7042 29870 7070
rect 29894 7042 29922 7070
rect 29946 7042 29974 7070
rect 29998 7042 30026 7070
rect 34582 7042 34610 7070
rect 34634 7042 34662 7070
rect 34686 7042 34714 7070
rect 34738 7042 34766 7070
rect 34790 7042 34818 7070
rect 34842 7042 34870 7070
rect 34894 7042 34922 7070
rect 34946 7042 34974 7070
rect 34998 7042 35026 7070
rect 31990 6734 32018 6762
rect 2082 6650 2110 6678
rect 2134 6650 2162 6678
rect 2186 6650 2214 6678
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 2394 6650 2422 6678
rect 2446 6650 2474 6678
rect 2498 6650 2526 6678
rect 7082 6650 7110 6678
rect 7134 6650 7162 6678
rect 7186 6650 7214 6678
rect 7238 6650 7266 6678
rect 7290 6650 7318 6678
rect 7342 6650 7370 6678
rect 7394 6650 7422 6678
rect 7446 6650 7474 6678
rect 7498 6650 7526 6678
rect 12082 6650 12110 6678
rect 12134 6650 12162 6678
rect 12186 6650 12214 6678
rect 12238 6650 12266 6678
rect 12290 6650 12318 6678
rect 12342 6650 12370 6678
rect 12394 6650 12422 6678
rect 12446 6650 12474 6678
rect 12498 6650 12526 6678
rect 17082 6650 17110 6678
rect 17134 6650 17162 6678
rect 17186 6650 17214 6678
rect 17238 6650 17266 6678
rect 17290 6650 17318 6678
rect 17342 6650 17370 6678
rect 17394 6650 17422 6678
rect 17446 6650 17474 6678
rect 17498 6650 17526 6678
rect 22082 6650 22110 6678
rect 22134 6650 22162 6678
rect 22186 6650 22214 6678
rect 22238 6650 22266 6678
rect 22290 6650 22318 6678
rect 22342 6650 22370 6678
rect 22394 6650 22422 6678
rect 22446 6650 22474 6678
rect 22498 6650 22526 6678
rect 27082 6650 27110 6678
rect 27134 6650 27162 6678
rect 27186 6650 27214 6678
rect 27238 6650 27266 6678
rect 27290 6650 27318 6678
rect 27342 6650 27370 6678
rect 27394 6650 27422 6678
rect 27446 6650 27474 6678
rect 27498 6650 27526 6678
rect 32082 6650 32110 6678
rect 32134 6650 32162 6678
rect 32186 6650 32214 6678
rect 32238 6650 32266 6678
rect 32290 6650 32318 6678
rect 32342 6650 32370 6678
rect 32394 6650 32422 6678
rect 32446 6650 32474 6678
rect 32498 6650 32526 6678
rect 37082 6650 37110 6678
rect 37134 6650 37162 6678
rect 37186 6650 37214 6678
rect 37238 6650 37266 6678
rect 37290 6650 37318 6678
rect 37342 6650 37370 6678
rect 37394 6650 37422 6678
rect 37446 6650 37474 6678
rect 37498 6650 37526 6678
rect 4582 6258 4610 6286
rect 4634 6258 4662 6286
rect 4686 6258 4714 6286
rect 4738 6258 4766 6286
rect 4790 6258 4818 6286
rect 4842 6258 4870 6286
rect 4894 6258 4922 6286
rect 4946 6258 4974 6286
rect 4998 6258 5026 6286
rect 9582 6258 9610 6286
rect 9634 6258 9662 6286
rect 9686 6258 9714 6286
rect 9738 6258 9766 6286
rect 9790 6258 9818 6286
rect 9842 6258 9870 6286
rect 9894 6258 9922 6286
rect 9946 6258 9974 6286
rect 9998 6258 10026 6286
rect 14582 6258 14610 6286
rect 14634 6258 14662 6286
rect 14686 6258 14714 6286
rect 14738 6258 14766 6286
rect 14790 6258 14818 6286
rect 14842 6258 14870 6286
rect 14894 6258 14922 6286
rect 14946 6258 14974 6286
rect 14998 6258 15026 6286
rect 19582 6258 19610 6286
rect 19634 6258 19662 6286
rect 19686 6258 19714 6286
rect 19738 6258 19766 6286
rect 19790 6258 19818 6286
rect 19842 6258 19870 6286
rect 19894 6258 19922 6286
rect 19946 6258 19974 6286
rect 19998 6258 20026 6286
rect 24582 6258 24610 6286
rect 24634 6258 24662 6286
rect 24686 6258 24714 6286
rect 24738 6258 24766 6286
rect 24790 6258 24818 6286
rect 24842 6258 24870 6286
rect 24894 6258 24922 6286
rect 24946 6258 24974 6286
rect 24998 6258 25026 6286
rect 29582 6258 29610 6286
rect 29634 6258 29662 6286
rect 29686 6258 29714 6286
rect 29738 6258 29766 6286
rect 29790 6258 29818 6286
rect 29842 6258 29870 6286
rect 29894 6258 29922 6286
rect 29946 6258 29974 6286
rect 29998 6258 30026 6286
rect 34582 6258 34610 6286
rect 34634 6258 34662 6286
rect 34686 6258 34714 6286
rect 34738 6258 34766 6286
rect 34790 6258 34818 6286
rect 34842 6258 34870 6286
rect 34894 6258 34922 6286
rect 34946 6258 34974 6286
rect 34998 6258 35026 6286
rect 31990 6062 32018 6090
rect 2082 5866 2110 5894
rect 2134 5866 2162 5894
rect 2186 5866 2214 5894
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 2394 5866 2422 5894
rect 2446 5866 2474 5894
rect 2498 5866 2526 5894
rect 7082 5866 7110 5894
rect 7134 5866 7162 5894
rect 7186 5866 7214 5894
rect 7238 5866 7266 5894
rect 7290 5866 7318 5894
rect 7342 5866 7370 5894
rect 7394 5866 7422 5894
rect 7446 5866 7474 5894
rect 7498 5866 7526 5894
rect 12082 5866 12110 5894
rect 12134 5866 12162 5894
rect 12186 5866 12214 5894
rect 12238 5866 12266 5894
rect 12290 5866 12318 5894
rect 12342 5866 12370 5894
rect 12394 5866 12422 5894
rect 12446 5866 12474 5894
rect 12498 5866 12526 5894
rect 17082 5866 17110 5894
rect 17134 5866 17162 5894
rect 17186 5866 17214 5894
rect 17238 5866 17266 5894
rect 17290 5866 17318 5894
rect 17342 5866 17370 5894
rect 17394 5866 17422 5894
rect 17446 5866 17474 5894
rect 17498 5866 17526 5894
rect 22082 5866 22110 5894
rect 22134 5866 22162 5894
rect 22186 5866 22214 5894
rect 22238 5866 22266 5894
rect 22290 5866 22318 5894
rect 22342 5866 22370 5894
rect 22394 5866 22422 5894
rect 22446 5866 22474 5894
rect 22498 5866 22526 5894
rect 27082 5866 27110 5894
rect 27134 5866 27162 5894
rect 27186 5866 27214 5894
rect 27238 5866 27266 5894
rect 27290 5866 27318 5894
rect 27342 5866 27370 5894
rect 27394 5866 27422 5894
rect 27446 5866 27474 5894
rect 27498 5866 27526 5894
rect 32082 5866 32110 5894
rect 32134 5866 32162 5894
rect 32186 5866 32214 5894
rect 32238 5866 32266 5894
rect 32290 5866 32318 5894
rect 32342 5866 32370 5894
rect 32394 5866 32422 5894
rect 32446 5866 32474 5894
rect 32498 5866 32526 5894
rect 37082 5866 37110 5894
rect 37134 5866 37162 5894
rect 37186 5866 37214 5894
rect 37238 5866 37266 5894
rect 37290 5866 37318 5894
rect 37342 5866 37370 5894
rect 37394 5866 37422 5894
rect 37446 5866 37474 5894
rect 37498 5866 37526 5894
rect 31990 5614 32018 5642
rect 4582 5474 4610 5502
rect 4634 5474 4662 5502
rect 4686 5474 4714 5502
rect 4738 5474 4766 5502
rect 4790 5474 4818 5502
rect 4842 5474 4870 5502
rect 4894 5474 4922 5502
rect 4946 5474 4974 5502
rect 4998 5474 5026 5502
rect 9582 5474 9610 5502
rect 9634 5474 9662 5502
rect 9686 5474 9714 5502
rect 9738 5474 9766 5502
rect 9790 5474 9818 5502
rect 9842 5474 9870 5502
rect 9894 5474 9922 5502
rect 9946 5474 9974 5502
rect 9998 5474 10026 5502
rect 14582 5474 14610 5502
rect 14634 5474 14662 5502
rect 14686 5474 14714 5502
rect 14738 5474 14766 5502
rect 14790 5474 14818 5502
rect 14842 5474 14870 5502
rect 14894 5474 14922 5502
rect 14946 5474 14974 5502
rect 14998 5474 15026 5502
rect 19582 5474 19610 5502
rect 19634 5474 19662 5502
rect 19686 5474 19714 5502
rect 19738 5474 19766 5502
rect 19790 5474 19818 5502
rect 19842 5474 19870 5502
rect 19894 5474 19922 5502
rect 19946 5474 19974 5502
rect 19998 5474 20026 5502
rect 24582 5474 24610 5502
rect 24634 5474 24662 5502
rect 24686 5474 24714 5502
rect 24738 5474 24766 5502
rect 24790 5474 24818 5502
rect 24842 5474 24870 5502
rect 24894 5474 24922 5502
rect 24946 5474 24974 5502
rect 24998 5474 25026 5502
rect 29582 5474 29610 5502
rect 29634 5474 29662 5502
rect 29686 5474 29714 5502
rect 29738 5474 29766 5502
rect 29790 5474 29818 5502
rect 29842 5474 29870 5502
rect 29894 5474 29922 5502
rect 29946 5474 29974 5502
rect 29998 5474 30026 5502
rect 34582 5474 34610 5502
rect 34634 5474 34662 5502
rect 34686 5474 34714 5502
rect 34738 5474 34766 5502
rect 34790 5474 34818 5502
rect 34842 5474 34870 5502
rect 34894 5474 34922 5502
rect 34946 5474 34974 5502
rect 34998 5474 35026 5502
rect 31990 5278 32018 5306
rect 2082 5082 2110 5110
rect 2134 5082 2162 5110
rect 2186 5082 2214 5110
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 2394 5082 2422 5110
rect 2446 5082 2474 5110
rect 2498 5082 2526 5110
rect 7082 5082 7110 5110
rect 7134 5082 7162 5110
rect 7186 5082 7214 5110
rect 7238 5082 7266 5110
rect 7290 5082 7318 5110
rect 7342 5082 7370 5110
rect 7394 5082 7422 5110
rect 7446 5082 7474 5110
rect 7498 5082 7526 5110
rect 12082 5082 12110 5110
rect 12134 5082 12162 5110
rect 12186 5082 12214 5110
rect 12238 5082 12266 5110
rect 12290 5082 12318 5110
rect 12342 5082 12370 5110
rect 12394 5082 12422 5110
rect 12446 5082 12474 5110
rect 12498 5082 12526 5110
rect 17082 5082 17110 5110
rect 17134 5082 17162 5110
rect 17186 5082 17214 5110
rect 17238 5082 17266 5110
rect 17290 5082 17318 5110
rect 17342 5082 17370 5110
rect 17394 5082 17422 5110
rect 17446 5082 17474 5110
rect 17498 5082 17526 5110
rect 22082 5082 22110 5110
rect 22134 5082 22162 5110
rect 22186 5082 22214 5110
rect 22238 5082 22266 5110
rect 22290 5082 22318 5110
rect 22342 5082 22370 5110
rect 22394 5082 22422 5110
rect 22446 5082 22474 5110
rect 22498 5082 22526 5110
rect 27082 5082 27110 5110
rect 27134 5082 27162 5110
rect 27186 5082 27214 5110
rect 27238 5082 27266 5110
rect 27290 5082 27318 5110
rect 27342 5082 27370 5110
rect 27394 5082 27422 5110
rect 27446 5082 27474 5110
rect 27498 5082 27526 5110
rect 32082 5082 32110 5110
rect 32134 5082 32162 5110
rect 32186 5082 32214 5110
rect 32238 5082 32266 5110
rect 32290 5082 32318 5110
rect 32342 5082 32370 5110
rect 32394 5082 32422 5110
rect 32446 5082 32474 5110
rect 32498 5082 32526 5110
rect 37082 5082 37110 5110
rect 37134 5082 37162 5110
rect 37186 5082 37214 5110
rect 37238 5082 37266 5110
rect 37290 5082 37318 5110
rect 37342 5082 37370 5110
rect 37394 5082 37422 5110
rect 37446 5082 37474 5110
rect 37498 5082 37526 5110
rect 4582 4690 4610 4718
rect 4634 4690 4662 4718
rect 4686 4690 4714 4718
rect 4738 4690 4766 4718
rect 4790 4690 4818 4718
rect 4842 4690 4870 4718
rect 4894 4690 4922 4718
rect 4946 4690 4974 4718
rect 4998 4690 5026 4718
rect 9582 4690 9610 4718
rect 9634 4690 9662 4718
rect 9686 4690 9714 4718
rect 9738 4690 9766 4718
rect 9790 4690 9818 4718
rect 9842 4690 9870 4718
rect 9894 4690 9922 4718
rect 9946 4690 9974 4718
rect 9998 4690 10026 4718
rect 14582 4690 14610 4718
rect 14634 4690 14662 4718
rect 14686 4690 14714 4718
rect 14738 4690 14766 4718
rect 14790 4690 14818 4718
rect 14842 4690 14870 4718
rect 14894 4690 14922 4718
rect 14946 4690 14974 4718
rect 14998 4690 15026 4718
rect 19582 4690 19610 4718
rect 19634 4690 19662 4718
rect 19686 4690 19714 4718
rect 19738 4690 19766 4718
rect 19790 4690 19818 4718
rect 19842 4690 19870 4718
rect 19894 4690 19922 4718
rect 19946 4690 19974 4718
rect 19998 4690 20026 4718
rect 24582 4690 24610 4718
rect 24634 4690 24662 4718
rect 24686 4690 24714 4718
rect 24738 4690 24766 4718
rect 24790 4690 24818 4718
rect 24842 4690 24870 4718
rect 24894 4690 24922 4718
rect 24946 4690 24974 4718
rect 24998 4690 25026 4718
rect 31990 4886 32018 4914
rect 29582 4690 29610 4718
rect 29634 4690 29662 4718
rect 29686 4690 29714 4718
rect 29738 4690 29766 4718
rect 29790 4690 29818 4718
rect 29842 4690 29870 4718
rect 29894 4690 29922 4718
rect 29946 4690 29974 4718
rect 29998 4690 30026 4718
rect 34582 4690 34610 4718
rect 34634 4690 34662 4718
rect 34686 4690 34714 4718
rect 34738 4690 34766 4718
rect 34790 4690 34818 4718
rect 34842 4690 34870 4718
rect 34894 4690 34922 4718
rect 34946 4690 34974 4718
rect 34998 4690 35026 4718
rect 2082 4298 2110 4326
rect 2134 4298 2162 4326
rect 2186 4298 2214 4326
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 2394 4298 2422 4326
rect 2446 4298 2474 4326
rect 2498 4298 2526 4326
rect 7082 4298 7110 4326
rect 7134 4298 7162 4326
rect 7186 4298 7214 4326
rect 7238 4298 7266 4326
rect 7290 4298 7318 4326
rect 7342 4298 7370 4326
rect 7394 4298 7422 4326
rect 7446 4298 7474 4326
rect 7498 4298 7526 4326
rect 12082 4298 12110 4326
rect 12134 4298 12162 4326
rect 12186 4298 12214 4326
rect 12238 4298 12266 4326
rect 12290 4298 12318 4326
rect 12342 4298 12370 4326
rect 12394 4298 12422 4326
rect 12446 4298 12474 4326
rect 12498 4298 12526 4326
rect 17082 4298 17110 4326
rect 17134 4298 17162 4326
rect 17186 4298 17214 4326
rect 17238 4298 17266 4326
rect 17290 4298 17318 4326
rect 17342 4298 17370 4326
rect 17394 4298 17422 4326
rect 17446 4298 17474 4326
rect 17498 4298 17526 4326
rect 22082 4298 22110 4326
rect 22134 4298 22162 4326
rect 22186 4298 22214 4326
rect 22238 4298 22266 4326
rect 22290 4298 22318 4326
rect 22342 4298 22370 4326
rect 22394 4298 22422 4326
rect 22446 4298 22474 4326
rect 22498 4298 22526 4326
rect 27082 4298 27110 4326
rect 27134 4298 27162 4326
rect 27186 4298 27214 4326
rect 27238 4298 27266 4326
rect 27290 4298 27318 4326
rect 27342 4298 27370 4326
rect 27394 4298 27422 4326
rect 27446 4298 27474 4326
rect 27498 4298 27526 4326
rect 32082 4298 32110 4326
rect 32134 4298 32162 4326
rect 32186 4298 32214 4326
rect 32238 4298 32266 4326
rect 32290 4298 32318 4326
rect 32342 4298 32370 4326
rect 32394 4298 32422 4326
rect 32446 4298 32474 4326
rect 32498 4298 32526 4326
rect 37082 4298 37110 4326
rect 37134 4298 37162 4326
rect 37186 4298 37214 4326
rect 37238 4298 37266 4326
rect 37290 4298 37318 4326
rect 37342 4298 37370 4326
rect 37394 4298 37422 4326
rect 37446 4298 37474 4326
rect 37498 4298 37526 4326
rect 31990 4046 32018 4074
rect 4582 3906 4610 3934
rect 4634 3906 4662 3934
rect 4686 3906 4714 3934
rect 4738 3906 4766 3934
rect 4790 3906 4818 3934
rect 4842 3906 4870 3934
rect 4894 3906 4922 3934
rect 4946 3906 4974 3934
rect 4998 3906 5026 3934
rect 9582 3906 9610 3934
rect 9634 3906 9662 3934
rect 9686 3906 9714 3934
rect 9738 3906 9766 3934
rect 9790 3906 9818 3934
rect 9842 3906 9870 3934
rect 9894 3906 9922 3934
rect 9946 3906 9974 3934
rect 9998 3906 10026 3934
rect 14582 3906 14610 3934
rect 14634 3906 14662 3934
rect 14686 3906 14714 3934
rect 14738 3906 14766 3934
rect 14790 3906 14818 3934
rect 14842 3906 14870 3934
rect 14894 3906 14922 3934
rect 14946 3906 14974 3934
rect 14998 3906 15026 3934
rect 19582 3906 19610 3934
rect 19634 3906 19662 3934
rect 19686 3906 19714 3934
rect 19738 3906 19766 3934
rect 19790 3906 19818 3934
rect 19842 3906 19870 3934
rect 19894 3906 19922 3934
rect 19946 3906 19974 3934
rect 19998 3906 20026 3934
rect 24582 3906 24610 3934
rect 24634 3906 24662 3934
rect 24686 3906 24714 3934
rect 24738 3906 24766 3934
rect 24790 3906 24818 3934
rect 24842 3906 24870 3934
rect 24894 3906 24922 3934
rect 24946 3906 24974 3934
rect 24998 3906 25026 3934
rect 29582 3906 29610 3934
rect 29634 3906 29662 3934
rect 29686 3906 29714 3934
rect 29738 3906 29766 3934
rect 29790 3906 29818 3934
rect 29842 3906 29870 3934
rect 29894 3906 29922 3934
rect 29946 3906 29974 3934
rect 29998 3906 30026 3934
rect 34582 3906 34610 3934
rect 34634 3906 34662 3934
rect 34686 3906 34714 3934
rect 34738 3906 34766 3934
rect 34790 3906 34818 3934
rect 34842 3906 34870 3934
rect 34894 3906 34922 3934
rect 34946 3906 34974 3934
rect 34998 3906 35026 3934
rect 2082 3514 2110 3542
rect 2134 3514 2162 3542
rect 2186 3514 2214 3542
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 2394 3514 2422 3542
rect 2446 3514 2474 3542
rect 2498 3514 2526 3542
rect 7082 3514 7110 3542
rect 7134 3514 7162 3542
rect 7186 3514 7214 3542
rect 7238 3514 7266 3542
rect 7290 3514 7318 3542
rect 7342 3514 7370 3542
rect 7394 3514 7422 3542
rect 7446 3514 7474 3542
rect 7498 3514 7526 3542
rect 12082 3514 12110 3542
rect 12134 3514 12162 3542
rect 12186 3514 12214 3542
rect 12238 3514 12266 3542
rect 12290 3514 12318 3542
rect 12342 3514 12370 3542
rect 12394 3514 12422 3542
rect 12446 3514 12474 3542
rect 12498 3514 12526 3542
rect 17082 3514 17110 3542
rect 17134 3514 17162 3542
rect 17186 3514 17214 3542
rect 17238 3514 17266 3542
rect 17290 3514 17318 3542
rect 17342 3514 17370 3542
rect 17394 3514 17422 3542
rect 17446 3514 17474 3542
rect 17498 3514 17526 3542
rect 22082 3514 22110 3542
rect 22134 3514 22162 3542
rect 22186 3514 22214 3542
rect 22238 3514 22266 3542
rect 22290 3514 22318 3542
rect 22342 3514 22370 3542
rect 22394 3514 22422 3542
rect 22446 3514 22474 3542
rect 22498 3514 22526 3542
rect 27082 3514 27110 3542
rect 27134 3514 27162 3542
rect 27186 3514 27214 3542
rect 27238 3514 27266 3542
rect 27290 3514 27318 3542
rect 27342 3514 27370 3542
rect 27394 3514 27422 3542
rect 27446 3514 27474 3542
rect 27498 3514 27526 3542
rect 32082 3514 32110 3542
rect 32134 3514 32162 3542
rect 32186 3514 32214 3542
rect 32238 3514 32266 3542
rect 32290 3514 32318 3542
rect 32342 3514 32370 3542
rect 32394 3514 32422 3542
rect 32446 3514 32474 3542
rect 32498 3514 32526 3542
rect 37082 3514 37110 3542
rect 37134 3514 37162 3542
rect 37186 3514 37214 3542
rect 37238 3514 37266 3542
rect 37290 3514 37318 3542
rect 37342 3514 37370 3542
rect 37394 3514 37422 3542
rect 37446 3514 37474 3542
rect 37498 3514 37526 3542
rect 31990 3318 32018 3346
rect 4582 3122 4610 3150
rect 4634 3122 4662 3150
rect 4686 3122 4714 3150
rect 4738 3122 4766 3150
rect 4790 3122 4818 3150
rect 4842 3122 4870 3150
rect 4894 3122 4922 3150
rect 4946 3122 4974 3150
rect 4998 3122 5026 3150
rect 9582 3122 9610 3150
rect 9634 3122 9662 3150
rect 9686 3122 9714 3150
rect 9738 3122 9766 3150
rect 9790 3122 9818 3150
rect 9842 3122 9870 3150
rect 9894 3122 9922 3150
rect 9946 3122 9974 3150
rect 9998 3122 10026 3150
rect 14582 3122 14610 3150
rect 14634 3122 14662 3150
rect 14686 3122 14714 3150
rect 14738 3122 14766 3150
rect 14790 3122 14818 3150
rect 14842 3122 14870 3150
rect 14894 3122 14922 3150
rect 14946 3122 14974 3150
rect 14998 3122 15026 3150
rect 19582 3122 19610 3150
rect 19634 3122 19662 3150
rect 19686 3122 19714 3150
rect 19738 3122 19766 3150
rect 19790 3122 19818 3150
rect 19842 3122 19870 3150
rect 19894 3122 19922 3150
rect 19946 3122 19974 3150
rect 19998 3122 20026 3150
rect 24582 3122 24610 3150
rect 24634 3122 24662 3150
rect 24686 3122 24714 3150
rect 24738 3122 24766 3150
rect 24790 3122 24818 3150
rect 24842 3122 24870 3150
rect 24894 3122 24922 3150
rect 24946 3122 24974 3150
rect 24998 3122 25026 3150
rect 29582 3122 29610 3150
rect 29634 3122 29662 3150
rect 29686 3122 29714 3150
rect 29738 3122 29766 3150
rect 29790 3122 29818 3150
rect 29842 3122 29870 3150
rect 29894 3122 29922 3150
rect 29946 3122 29974 3150
rect 29998 3122 30026 3150
rect 34582 3122 34610 3150
rect 34634 3122 34662 3150
rect 34686 3122 34714 3150
rect 34738 3122 34766 3150
rect 34790 3122 34818 3150
rect 34842 3122 34870 3150
rect 34894 3122 34922 3150
rect 34946 3122 34974 3150
rect 34998 3122 35026 3150
rect 2082 2730 2110 2758
rect 2134 2730 2162 2758
rect 2186 2730 2214 2758
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 2394 2730 2422 2758
rect 2446 2730 2474 2758
rect 2498 2730 2526 2758
rect 7082 2730 7110 2758
rect 7134 2730 7162 2758
rect 7186 2730 7214 2758
rect 7238 2730 7266 2758
rect 7290 2730 7318 2758
rect 7342 2730 7370 2758
rect 7394 2730 7422 2758
rect 7446 2730 7474 2758
rect 7498 2730 7526 2758
rect 12082 2730 12110 2758
rect 12134 2730 12162 2758
rect 12186 2730 12214 2758
rect 12238 2730 12266 2758
rect 12290 2730 12318 2758
rect 12342 2730 12370 2758
rect 12394 2730 12422 2758
rect 12446 2730 12474 2758
rect 12498 2730 12526 2758
rect 17082 2730 17110 2758
rect 17134 2730 17162 2758
rect 17186 2730 17214 2758
rect 17238 2730 17266 2758
rect 17290 2730 17318 2758
rect 17342 2730 17370 2758
rect 17394 2730 17422 2758
rect 17446 2730 17474 2758
rect 17498 2730 17526 2758
rect 22082 2730 22110 2758
rect 22134 2730 22162 2758
rect 22186 2730 22214 2758
rect 22238 2730 22266 2758
rect 22290 2730 22318 2758
rect 22342 2730 22370 2758
rect 22394 2730 22422 2758
rect 22446 2730 22474 2758
rect 22498 2730 22526 2758
rect 27082 2730 27110 2758
rect 27134 2730 27162 2758
rect 27186 2730 27214 2758
rect 27238 2730 27266 2758
rect 27290 2730 27318 2758
rect 27342 2730 27370 2758
rect 27394 2730 27422 2758
rect 27446 2730 27474 2758
rect 27498 2730 27526 2758
rect 32082 2730 32110 2758
rect 32134 2730 32162 2758
rect 32186 2730 32214 2758
rect 32238 2730 32266 2758
rect 32290 2730 32318 2758
rect 32342 2730 32370 2758
rect 32394 2730 32422 2758
rect 32446 2730 32474 2758
rect 32498 2730 32526 2758
rect 37082 2730 37110 2758
rect 37134 2730 37162 2758
rect 37186 2730 37214 2758
rect 37238 2730 37266 2758
rect 37290 2730 37318 2758
rect 37342 2730 37370 2758
rect 37394 2730 37422 2758
rect 37446 2730 37474 2758
rect 37498 2730 37526 2758
rect 4582 2338 4610 2366
rect 4634 2338 4662 2366
rect 4686 2338 4714 2366
rect 4738 2338 4766 2366
rect 4790 2338 4818 2366
rect 4842 2338 4870 2366
rect 4894 2338 4922 2366
rect 4946 2338 4974 2366
rect 4998 2338 5026 2366
rect 9582 2338 9610 2366
rect 9634 2338 9662 2366
rect 9686 2338 9714 2366
rect 9738 2338 9766 2366
rect 9790 2338 9818 2366
rect 9842 2338 9870 2366
rect 9894 2338 9922 2366
rect 9946 2338 9974 2366
rect 9998 2338 10026 2366
rect 14582 2338 14610 2366
rect 14634 2338 14662 2366
rect 14686 2338 14714 2366
rect 14738 2338 14766 2366
rect 14790 2338 14818 2366
rect 14842 2338 14870 2366
rect 14894 2338 14922 2366
rect 14946 2338 14974 2366
rect 14998 2338 15026 2366
rect 19582 2338 19610 2366
rect 19634 2338 19662 2366
rect 19686 2338 19714 2366
rect 19738 2338 19766 2366
rect 19790 2338 19818 2366
rect 19842 2338 19870 2366
rect 19894 2338 19922 2366
rect 19946 2338 19974 2366
rect 19998 2338 20026 2366
rect 24582 2338 24610 2366
rect 24634 2338 24662 2366
rect 24686 2338 24714 2366
rect 24738 2338 24766 2366
rect 24790 2338 24818 2366
rect 24842 2338 24870 2366
rect 24894 2338 24922 2366
rect 24946 2338 24974 2366
rect 24998 2338 25026 2366
rect 29582 2338 29610 2366
rect 29634 2338 29662 2366
rect 29686 2338 29714 2366
rect 29738 2338 29766 2366
rect 29790 2338 29818 2366
rect 29842 2338 29870 2366
rect 29894 2338 29922 2366
rect 29946 2338 29974 2366
rect 29998 2338 30026 2366
rect 34582 2338 34610 2366
rect 34634 2338 34662 2366
rect 34686 2338 34714 2366
rect 34738 2338 34766 2366
rect 34790 2338 34818 2366
rect 34842 2338 34870 2366
rect 34894 2338 34922 2366
rect 34946 2338 34974 2366
rect 34998 2338 35026 2366
rect 2082 1946 2110 1974
rect 2134 1946 2162 1974
rect 2186 1946 2214 1974
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 2394 1946 2422 1974
rect 2446 1946 2474 1974
rect 2498 1946 2526 1974
rect 7082 1946 7110 1974
rect 7134 1946 7162 1974
rect 7186 1946 7214 1974
rect 7238 1946 7266 1974
rect 7290 1946 7318 1974
rect 7342 1946 7370 1974
rect 7394 1946 7422 1974
rect 7446 1946 7474 1974
rect 7498 1946 7526 1974
rect 12082 1946 12110 1974
rect 12134 1946 12162 1974
rect 12186 1946 12214 1974
rect 12238 1946 12266 1974
rect 12290 1946 12318 1974
rect 12342 1946 12370 1974
rect 12394 1946 12422 1974
rect 12446 1946 12474 1974
rect 12498 1946 12526 1974
rect 17082 1946 17110 1974
rect 17134 1946 17162 1974
rect 17186 1946 17214 1974
rect 17238 1946 17266 1974
rect 17290 1946 17318 1974
rect 17342 1946 17370 1974
rect 17394 1946 17422 1974
rect 17446 1946 17474 1974
rect 17498 1946 17526 1974
rect 22082 1946 22110 1974
rect 22134 1946 22162 1974
rect 22186 1946 22214 1974
rect 22238 1946 22266 1974
rect 22290 1946 22318 1974
rect 22342 1946 22370 1974
rect 22394 1946 22422 1974
rect 22446 1946 22474 1974
rect 22498 1946 22526 1974
rect 27082 1946 27110 1974
rect 27134 1946 27162 1974
rect 27186 1946 27214 1974
rect 27238 1946 27266 1974
rect 27290 1946 27318 1974
rect 27342 1946 27370 1974
rect 27394 1946 27422 1974
rect 27446 1946 27474 1974
rect 27498 1946 27526 1974
rect 32082 1946 32110 1974
rect 32134 1946 32162 1974
rect 32186 1946 32214 1974
rect 32238 1946 32266 1974
rect 32290 1946 32318 1974
rect 32342 1946 32370 1974
rect 32394 1946 32422 1974
rect 32446 1946 32474 1974
rect 32498 1946 32526 1974
rect 37082 1946 37110 1974
rect 37134 1946 37162 1974
rect 37186 1946 37214 1974
rect 37238 1946 37266 1974
rect 37290 1946 37318 1974
rect 37342 1946 37370 1974
rect 37394 1946 37422 1974
rect 37446 1946 37474 1974
rect 37498 1946 37526 1974
rect 4582 1554 4610 1582
rect 4634 1554 4662 1582
rect 4686 1554 4714 1582
rect 4738 1554 4766 1582
rect 4790 1554 4818 1582
rect 4842 1554 4870 1582
rect 4894 1554 4922 1582
rect 4946 1554 4974 1582
rect 4998 1554 5026 1582
rect 9582 1554 9610 1582
rect 9634 1554 9662 1582
rect 9686 1554 9714 1582
rect 9738 1554 9766 1582
rect 9790 1554 9818 1582
rect 9842 1554 9870 1582
rect 9894 1554 9922 1582
rect 9946 1554 9974 1582
rect 9998 1554 10026 1582
rect 14582 1554 14610 1582
rect 14634 1554 14662 1582
rect 14686 1554 14714 1582
rect 14738 1554 14766 1582
rect 14790 1554 14818 1582
rect 14842 1554 14870 1582
rect 14894 1554 14922 1582
rect 14946 1554 14974 1582
rect 14998 1554 15026 1582
rect 19582 1554 19610 1582
rect 19634 1554 19662 1582
rect 19686 1554 19714 1582
rect 19738 1554 19766 1582
rect 19790 1554 19818 1582
rect 19842 1554 19870 1582
rect 19894 1554 19922 1582
rect 19946 1554 19974 1582
rect 19998 1554 20026 1582
rect 24582 1554 24610 1582
rect 24634 1554 24662 1582
rect 24686 1554 24714 1582
rect 24738 1554 24766 1582
rect 24790 1554 24818 1582
rect 24842 1554 24870 1582
rect 24894 1554 24922 1582
rect 24946 1554 24974 1582
rect 24998 1554 25026 1582
rect 29582 1554 29610 1582
rect 29634 1554 29662 1582
rect 29686 1554 29714 1582
rect 29738 1554 29766 1582
rect 29790 1554 29818 1582
rect 29842 1554 29870 1582
rect 29894 1554 29922 1582
rect 29946 1554 29974 1582
rect 29998 1554 30026 1582
rect 34582 1554 34610 1582
rect 34634 1554 34662 1582
rect 34686 1554 34714 1582
rect 34738 1554 34766 1582
rect 34790 1554 34818 1582
rect 34842 1554 34870 1582
rect 34894 1554 34922 1582
rect 34946 1554 34974 1582
rect 34998 1554 35026 1582
<< metal4 >>
rect 2054 18438 2554 18454
rect 2054 18410 2082 18438
rect 2110 18410 2134 18438
rect 2162 18410 2186 18438
rect 2214 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2394 18438
rect 2422 18410 2446 18438
rect 2474 18410 2498 18438
rect 2526 18410 2554 18438
rect 2054 17654 2554 18410
rect 2054 17626 2082 17654
rect 2110 17626 2134 17654
rect 2162 17626 2186 17654
rect 2214 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2394 17654
rect 2422 17626 2446 17654
rect 2474 17626 2498 17654
rect 2526 17626 2554 17654
rect 2054 16870 2554 17626
rect 2054 16842 2082 16870
rect 2110 16842 2134 16870
rect 2162 16842 2186 16870
rect 2214 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2394 16870
rect 2422 16842 2446 16870
rect 2474 16842 2498 16870
rect 2526 16842 2554 16870
rect 2054 16086 2554 16842
rect 2054 16058 2082 16086
rect 2110 16058 2134 16086
rect 2162 16058 2186 16086
rect 2214 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2394 16086
rect 2422 16058 2446 16086
rect 2474 16058 2498 16086
rect 2526 16058 2554 16086
rect 2054 15302 2554 16058
rect 2054 15274 2082 15302
rect 2110 15274 2134 15302
rect 2162 15274 2186 15302
rect 2214 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2394 15302
rect 2422 15274 2446 15302
rect 2474 15274 2498 15302
rect 2526 15274 2554 15302
rect 2054 14518 2554 15274
rect 2054 14490 2082 14518
rect 2110 14490 2134 14518
rect 2162 14490 2186 14518
rect 2214 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2394 14518
rect 2422 14490 2446 14518
rect 2474 14490 2498 14518
rect 2526 14490 2554 14518
rect 2054 13734 2554 14490
rect 2054 13706 2082 13734
rect 2110 13706 2134 13734
rect 2162 13706 2186 13734
rect 2214 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2394 13734
rect 2422 13706 2446 13734
rect 2474 13706 2498 13734
rect 2526 13706 2554 13734
rect 2054 12950 2554 13706
rect 2054 12922 2082 12950
rect 2110 12922 2134 12950
rect 2162 12922 2186 12950
rect 2214 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2394 12950
rect 2422 12922 2446 12950
rect 2474 12922 2498 12950
rect 2526 12922 2554 12950
rect 2054 12166 2554 12922
rect 2054 12138 2082 12166
rect 2110 12138 2134 12166
rect 2162 12138 2186 12166
rect 2214 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2394 12166
rect 2422 12138 2446 12166
rect 2474 12138 2498 12166
rect 2526 12138 2554 12166
rect 2054 11382 2554 12138
rect 2054 11354 2082 11382
rect 2110 11354 2134 11382
rect 2162 11354 2186 11382
rect 2214 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2394 11382
rect 2422 11354 2446 11382
rect 2474 11354 2498 11382
rect 2526 11354 2554 11382
rect 2054 10598 2554 11354
rect 2054 10570 2082 10598
rect 2110 10570 2134 10598
rect 2162 10570 2186 10598
rect 2214 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2394 10598
rect 2422 10570 2446 10598
rect 2474 10570 2498 10598
rect 2526 10570 2554 10598
rect 2054 9814 2554 10570
rect 2054 9786 2082 9814
rect 2110 9786 2134 9814
rect 2162 9786 2186 9814
rect 2214 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2394 9814
rect 2422 9786 2446 9814
rect 2474 9786 2498 9814
rect 2526 9786 2554 9814
rect 2054 9030 2554 9786
rect 2054 9002 2082 9030
rect 2110 9002 2134 9030
rect 2162 9002 2186 9030
rect 2214 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2394 9030
rect 2422 9002 2446 9030
rect 2474 9002 2498 9030
rect 2526 9002 2554 9030
rect 2054 8246 2554 9002
rect 2054 8218 2082 8246
rect 2110 8218 2134 8246
rect 2162 8218 2186 8246
rect 2214 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2394 8246
rect 2422 8218 2446 8246
rect 2474 8218 2498 8246
rect 2526 8218 2554 8246
rect 2054 7462 2554 8218
rect 2054 7434 2082 7462
rect 2110 7434 2134 7462
rect 2162 7434 2186 7462
rect 2214 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2394 7462
rect 2422 7434 2446 7462
rect 2474 7434 2498 7462
rect 2526 7434 2554 7462
rect 2054 6678 2554 7434
rect 2054 6650 2082 6678
rect 2110 6650 2134 6678
rect 2162 6650 2186 6678
rect 2214 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2394 6678
rect 2422 6650 2446 6678
rect 2474 6650 2498 6678
rect 2526 6650 2554 6678
rect 2054 5894 2554 6650
rect 2054 5866 2082 5894
rect 2110 5866 2134 5894
rect 2162 5866 2186 5894
rect 2214 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2394 5894
rect 2422 5866 2446 5894
rect 2474 5866 2498 5894
rect 2526 5866 2554 5894
rect 2054 5110 2554 5866
rect 2054 5082 2082 5110
rect 2110 5082 2134 5110
rect 2162 5082 2186 5110
rect 2214 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2394 5110
rect 2422 5082 2446 5110
rect 2474 5082 2498 5110
rect 2526 5082 2554 5110
rect 2054 4326 2554 5082
rect 2054 4298 2082 4326
rect 2110 4298 2134 4326
rect 2162 4298 2186 4326
rect 2214 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2394 4326
rect 2422 4298 2446 4326
rect 2474 4298 2498 4326
rect 2526 4298 2554 4326
rect 2054 3542 2554 4298
rect 2054 3514 2082 3542
rect 2110 3514 2134 3542
rect 2162 3514 2186 3542
rect 2214 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2394 3542
rect 2422 3514 2446 3542
rect 2474 3514 2498 3542
rect 2526 3514 2554 3542
rect 2054 2758 2554 3514
rect 2054 2730 2082 2758
rect 2110 2730 2134 2758
rect 2162 2730 2186 2758
rect 2214 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2394 2758
rect 2422 2730 2446 2758
rect 2474 2730 2498 2758
rect 2526 2730 2554 2758
rect 2054 1974 2554 2730
rect 2054 1946 2082 1974
rect 2110 1946 2134 1974
rect 2162 1946 2186 1974
rect 2214 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2394 1974
rect 2422 1946 2446 1974
rect 2474 1946 2498 1974
rect 2526 1946 2554 1974
rect 2054 1538 2554 1946
rect 4554 18046 5054 18454
rect 4554 18018 4582 18046
rect 4610 18018 4634 18046
rect 4662 18018 4686 18046
rect 4714 18018 4738 18046
rect 4766 18018 4790 18046
rect 4818 18018 4842 18046
rect 4870 18018 4894 18046
rect 4922 18018 4946 18046
rect 4974 18018 4998 18046
rect 5026 18018 5054 18046
rect 4554 17262 5054 18018
rect 4554 17234 4582 17262
rect 4610 17234 4634 17262
rect 4662 17234 4686 17262
rect 4714 17234 4738 17262
rect 4766 17234 4790 17262
rect 4818 17234 4842 17262
rect 4870 17234 4894 17262
rect 4922 17234 4946 17262
rect 4974 17234 4998 17262
rect 5026 17234 5054 17262
rect 4554 16478 5054 17234
rect 4554 16450 4582 16478
rect 4610 16450 4634 16478
rect 4662 16450 4686 16478
rect 4714 16450 4738 16478
rect 4766 16450 4790 16478
rect 4818 16450 4842 16478
rect 4870 16450 4894 16478
rect 4922 16450 4946 16478
rect 4974 16450 4998 16478
rect 5026 16450 5054 16478
rect 4554 15694 5054 16450
rect 4554 15666 4582 15694
rect 4610 15666 4634 15694
rect 4662 15666 4686 15694
rect 4714 15666 4738 15694
rect 4766 15666 4790 15694
rect 4818 15666 4842 15694
rect 4870 15666 4894 15694
rect 4922 15666 4946 15694
rect 4974 15666 4998 15694
rect 5026 15666 5054 15694
rect 4554 14910 5054 15666
rect 4554 14882 4582 14910
rect 4610 14882 4634 14910
rect 4662 14882 4686 14910
rect 4714 14882 4738 14910
rect 4766 14882 4790 14910
rect 4818 14882 4842 14910
rect 4870 14882 4894 14910
rect 4922 14882 4946 14910
rect 4974 14882 4998 14910
rect 5026 14882 5054 14910
rect 4554 14126 5054 14882
rect 4554 14098 4582 14126
rect 4610 14098 4634 14126
rect 4662 14098 4686 14126
rect 4714 14098 4738 14126
rect 4766 14098 4790 14126
rect 4818 14098 4842 14126
rect 4870 14098 4894 14126
rect 4922 14098 4946 14126
rect 4974 14098 4998 14126
rect 5026 14098 5054 14126
rect 4554 13342 5054 14098
rect 4554 13314 4582 13342
rect 4610 13314 4634 13342
rect 4662 13314 4686 13342
rect 4714 13314 4738 13342
rect 4766 13314 4790 13342
rect 4818 13314 4842 13342
rect 4870 13314 4894 13342
rect 4922 13314 4946 13342
rect 4974 13314 4998 13342
rect 5026 13314 5054 13342
rect 4554 12558 5054 13314
rect 4554 12530 4582 12558
rect 4610 12530 4634 12558
rect 4662 12530 4686 12558
rect 4714 12530 4738 12558
rect 4766 12530 4790 12558
rect 4818 12530 4842 12558
rect 4870 12530 4894 12558
rect 4922 12530 4946 12558
rect 4974 12530 4998 12558
rect 5026 12530 5054 12558
rect 4554 11774 5054 12530
rect 4554 11746 4582 11774
rect 4610 11746 4634 11774
rect 4662 11746 4686 11774
rect 4714 11746 4738 11774
rect 4766 11746 4790 11774
rect 4818 11746 4842 11774
rect 4870 11746 4894 11774
rect 4922 11746 4946 11774
rect 4974 11746 4998 11774
rect 5026 11746 5054 11774
rect 4554 10990 5054 11746
rect 4554 10962 4582 10990
rect 4610 10962 4634 10990
rect 4662 10962 4686 10990
rect 4714 10962 4738 10990
rect 4766 10962 4790 10990
rect 4818 10962 4842 10990
rect 4870 10962 4894 10990
rect 4922 10962 4946 10990
rect 4974 10962 4998 10990
rect 5026 10962 5054 10990
rect 4554 10206 5054 10962
rect 4554 10178 4582 10206
rect 4610 10178 4634 10206
rect 4662 10178 4686 10206
rect 4714 10178 4738 10206
rect 4766 10178 4790 10206
rect 4818 10178 4842 10206
rect 4870 10178 4894 10206
rect 4922 10178 4946 10206
rect 4974 10178 4998 10206
rect 5026 10178 5054 10206
rect 4554 9422 5054 10178
rect 4554 9394 4582 9422
rect 4610 9394 4634 9422
rect 4662 9394 4686 9422
rect 4714 9394 4738 9422
rect 4766 9394 4790 9422
rect 4818 9394 4842 9422
rect 4870 9394 4894 9422
rect 4922 9394 4946 9422
rect 4974 9394 4998 9422
rect 5026 9394 5054 9422
rect 4554 8638 5054 9394
rect 4554 8610 4582 8638
rect 4610 8610 4634 8638
rect 4662 8610 4686 8638
rect 4714 8610 4738 8638
rect 4766 8610 4790 8638
rect 4818 8610 4842 8638
rect 4870 8610 4894 8638
rect 4922 8610 4946 8638
rect 4974 8610 4998 8638
rect 5026 8610 5054 8638
rect 4554 7854 5054 8610
rect 4554 7826 4582 7854
rect 4610 7826 4634 7854
rect 4662 7826 4686 7854
rect 4714 7826 4738 7854
rect 4766 7826 4790 7854
rect 4818 7826 4842 7854
rect 4870 7826 4894 7854
rect 4922 7826 4946 7854
rect 4974 7826 4998 7854
rect 5026 7826 5054 7854
rect 4554 7070 5054 7826
rect 4554 7042 4582 7070
rect 4610 7042 4634 7070
rect 4662 7042 4686 7070
rect 4714 7042 4738 7070
rect 4766 7042 4790 7070
rect 4818 7042 4842 7070
rect 4870 7042 4894 7070
rect 4922 7042 4946 7070
rect 4974 7042 4998 7070
rect 5026 7042 5054 7070
rect 4554 6286 5054 7042
rect 4554 6258 4582 6286
rect 4610 6258 4634 6286
rect 4662 6258 4686 6286
rect 4714 6258 4738 6286
rect 4766 6258 4790 6286
rect 4818 6258 4842 6286
rect 4870 6258 4894 6286
rect 4922 6258 4946 6286
rect 4974 6258 4998 6286
rect 5026 6258 5054 6286
rect 4554 5502 5054 6258
rect 4554 5474 4582 5502
rect 4610 5474 4634 5502
rect 4662 5474 4686 5502
rect 4714 5474 4738 5502
rect 4766 5474 4790 5502
rect 4818 5474 4842 5502
rect 4870 5474 4894 5502
rect 4922 5474 4946 5502
rect 4974 5474 4998 5502
rect 5026 5474 5054 5502
rect 4554 4718 5054 5474
rect 4554 4690 4582 4718
rect 4610 4690 4634 4718
rect 4662 4690 4686 4718
rect 4714 4690 4738 4718
rect 4766 4690 4790 4718
rect 4818 4690 4842 4718
rect 4870 4690 4894 4718
rect 4922 4690 4946 4718
rect 4974 4690 4998 4718
rect 5026 4690 5054 4718
rect 4554 3934 5054 4690
rect 4554 3906 4582 3934
rect 4610 3906 4634 3934
rect 4662 3906 4686 3934
rect 4714 3906 4738 3934
rect 4766 3906 4790 3934
rect 4818 3906 4842 3934
rect 4870 3906 4894 3934
rect 4922 3906 4946 3934
rect 4974 3906 4998 3934
rect 5026 3906 5054 3934
rect 4554 3150 5054 3906
rect 4554 3122 4582 3150
rect 4610 3122 4634 3150
rect 4662 3122 4686 3150
rect 4714 3122 4738 3150
rect 4766 3122 4790 3150
rect 4818 3122 4842 3150
rect 4870 3122 4894 3150
rect 4922 3122 4946 3150
rect 4974 3122 4998 3150
rect 5026 3122 5054 3150
rect 4554 2366 5054 3122
rect 4554 2338 4582 2366
rect 4610 2338 4634 2366
rect 4662 2338 4686 2366
rect 4714 2338 4738 2366
rect 4766 2338 4790 2366
rect 4818 2338 4842 2366
rect 4870 2338 4894 2366
rect 4922 2338 4946 2366
rect 4974 2338 4998 2366
rect 5026 2338 5054 2366
rect 4554 1582 5054 2338
rect 4554 1554 4582 1582
rect 4610 1554 4634 1582
rect 4662 1554 4686 1582
rect 4714 1554 4738 1582
rect 4766 1554 4790 1582
rect 4818 1554 4842 1582
rect 4870 1554 4894 1582
rect 4922 1554 4946 1582
rect 4974 1554 4998 1582
rect 5026 1554 5054 1582
rect 4554 1538 5054 1554
rect 7054 18438 7554 18454
rect 7054 18410 7082 18438
rect 7110 18410 7134 18438
rect 7162 18410 7186 18438
rect 7214 18410 7238 18438
rect 7266 18410 7290 18438
rect 7318 18410 7342 18438
rect 7370 18410 7394 18438
rect 7422 18410 7446 18438
rect 7474 18410 7498 18438
rect 7526 18410 7554 18438
rect 7054 17654 7554 18410
rect 7054 17626 7082 17654
rect 7110 17626 7134 17654
rect 7162 17626 7186 17654
rect 7214 17626 7238 17654
rect 7266 17626 7290 17654
rect 7318 17626 7342 17654
rect 7370 17626 7394 17654
rect 7422 17626 7446 17654
rect 7474 17626 7498 17654
rect 7526 17626 7554 17654
rect 7054 16870 7554 17626
rect 7054 16842 7082 16870
rect 7110 16842 7134 16870
rect 7162 16842 7186 16870
rect 7214 16842 7238 16870
rect 7266 16842 7290 16870
rect 7318 16842 7342 16870
rect 7370 16842 7394 16870
rect 7422 16842 7446 16870
rect 7474 16842 7498 16870
rect 7526 16842 7554 16870
rect 7054 16086 7554 16842
rect 7054 16058 7082 16086
rect 7110 16058 7134 16086
rect 7162 16058 7186 16086
rect 7214 16058 7238 16086
rect 7266 16058 7290 16086
rect 7318 16058 7342 16086
rect 7370 16058 7394 16086
rect 7422 16058 7446 16086
rect 7474 16058 7498 16086
rect 7526 16058 7554 16086
rect 7054 15302 7554 16058
rect 7054 15274 7082 15302
rect 7110 15274 7134 15302
rect 7162 15274 7186 15302
rect 7214 15274 7238 15302
rect 7266 15274 7290 15302
rect 7318 15274 7342 15302
rect 7370 15274 7394 15302
rect 7422 15274 7446 15302
rect 7474 15274 7498 15302
rect 7526 15274 7554 15302
rect 7054 14518 7554 15274
rect 7054 14490 7082 14518
rect 7110 14490 7134 14518
rect 7162 14490 7186 14518
rect 7214 14490 7238 14518
rect 7266 14490 7290 14518
rect 7318 14490 7342 14518
rect 7370 14490 7394 14518
rect 7422 14490 7446 14518
rect 7474 14490 7498 14518
rect 7526 14490 7554 14518
rect 7054 13734 7554 14490
rect 7054 13706 7082 13734
rect 7110 13706 7134 13734
rect 7162 13706 7186 13734
rect 7214 13706 7238 13734
rect 7266 13706 7290 13734
rect 7318 13706 7342 13734
rect 7370 13706 7394 13734
rect 7422 13706 7446 13734
rect 7474 13706 7498 13734
rect 7526 13706 7554 13734
rect 7054 12950 7554 13706
rect 7054 12922 7082 12950
rect 7110 12922 7134 12950
rect 7162 12922 7186 12950
rect 7214 12922 7238 12950
rect 7266 12922 7290 12950
rect 7318 12922 7342 12950
rect 7370 12922 7394 12950
rect 7422 12922 7446 12950
rect 7474 12922 7498 12950
rect 7526 12922 7554 12950
rect 7054 12166 7554 12922
rect 7054 12138 7082 12166
rect 7110 12138 7134 12166
rect 7162 12138 7186 12166
rect 7214 12138 7238 12166
rect 7266 12138 7290 12166
rect 7318 12138 7342 12166
rect 7370 12138 7394 12166
rect 7422 12138 7446 12166
rect 7474 12138 7498 12166
rect 7526 12138 7554 12166
rect 7054 11382 7554 12138
rect 7054 11354 7082 11382
rect 7110 11354 7134 11382
rect 7162 11354 7186 11382
rect 7214 11354 7238 11382
rect 7266 11354 7290 11382
rect 7318 11354 7342 11382
rect 7370 11354 7394 11382
rect 7422 11354 7446 11382
rect 7474 11354 7498 11382
rect 7526 11354 7554 11382
rect 7054 10598 7554 11354
rect 7054 10570 7082 10598
rect 7110 10570 7134 10598
rect 7162 10570 7186 10598
rect 7214 10570 7238 10598
rect 7266 10570 7290 10598
rect 7318 10570 7342 10598
rect 7370 10570 7394 10598
rect 7422 10570 7446 10598
rect 7474 10570 7498 10598
rect 7526 10570 7554 10598
rect 7054 9814 7554 10570
rect 7054 9786 7082 9814
rect 7110 9786 7134 9814
rect 7162 9786 7186 9814
rect 7214 9786 7238 9814
rect 7266 9786 7290 9814
rect 7318 9786 7342 9814
rect 7370 9786 7394 9814
rect 7422 9786 7446 9814
rect 7474 9786 7498 9814
rect 7526 9786 7554 9814
rect 7054 9030 7554 9786
rect 7054 9002 7082 9030
rect 7110 9002 7134 9030
rect 7162 9002 7186 9030
rect 7214 9002 7238 9030
rect 7266 9002 7290 9030
rect 7318 9002 7342 9030
rect 7370 9002 7394 9030
rect 7422 9002 7446 9030
rect 7474 9002 7498 9030
rect 7526 9002 7554 9030
rect 7054 8246 7554 9002
rect 7054 8218 7082 8246
rect 7110 8218 7134 8246
rect 7162 8218 7186 8246
rect 7214 8218 7238 8246
rect 7266 8218 7290 8246
rect 7318 8218 7342 8246
rect 7370 8218 7394 8246
rect 7422 8218 7446 8246
rect 7474 8218 7498 8246
rect 7526 8218 7554 8246
rect 7054 7462 7554 8218
rect 7054 7434 7082 7462
rect 7110 7434 7134 7462
rect 7162 7434 7186 7462
rect 7214 7434 7238 7462
rect 7266 7434 7290 7462
rect 7318 7434 7342 7462
rect 7370 7434 7394 7462
rect 7422 7434 7446 7462
rect 7474 7434 7498 7462
rect 7526 7434 7554 7462
rect 7054 6678 7554 7434
rect 7054 6650 7082 6678
rect 7110 6650 7134 6678
rect 7162 6650 7186 6678
rect 7214 6650 7238 6678
rect 7266 6650 7290 6678
rect 7318 6650 7342 6678
rect 7370 6650 7394 6678
rect 7422 6650 7446 6678
rect 7474 6650 7498 6678
rect 7526 6650 7554 6678
rect 7054 5894 7554 6650
rect 7054 5866 7082 5894
rect 7110 5866 7134 5894
rect 7162 5866 7186 5894
rect 7214 5866 7238 5894
rect 7266 5866 7290 5894
rect 7318 5866 7342 5894
rect 7370 5866 7394 5894
rect 7422 5866 7446 5894
rect 7474 5866 7498 5894
rect 7526 5866 7554 5894
rect 7054 5110 7554 5866
rect 7054 5082 7082 5110
rect 7110 5082 7134 5110
rect 7162 5082 7186 5110
rect 7214 5082 7238 5110
rect 7266 5082 7290 5110
rect 7318 5082 7342 5110
rect 7370 5082 7394 5110
rect 7422 5082 7446 5110
rect 7474 5082 7498 5110
rect 7526 5082 7554 5110
rect 7054 4326 7554 5082
rect 7054 4298 7082 4326
rect 7110 4298 7134 4326
rect 7162 4298 7186 4326
rect 7214 4298 7238 4326
rect 7266 4298 7290 4326
rect 7318 4298 7342 4326
rect 7370 4298 7394 4326
rect 7422 4298 7446 4326
rect 7474 4298 7498 4326
rect 7526 4298 7554 4326
rect 7054 3542 7554 4298
rect 7054 3514 7082 3542
rect 7110 3514 7134 3542
rect 7162 3514 7186 3542
rect 7214 3514 7238 3542
rect 7266 3514 7290 3542
rect 7318 3514 7342 3542
rect 7370 3514 7394 3542
rect 7422 3514 7446 3542
rect 7474 3514 7498 3542
rect 7526 3514 7554 3542
rect 7054 2758 7554 3514
rect 7054 2730 7082 2758
rect 7110 2730 7134 2758
rect 7162 2730 7186 2758
rect 7214 2730 7238 2758
rect 7266 2730 7290 2758
rect 7318 2730 7342 2758
rect 7370 2730 7394 2758
rect 7422 2730 7446 2758
rect 7474 2730 7498 2758
rect 7526 2730 7554 2758
rect 7054 1974 7554 2730
rect 7054 1946 7082 1974
rect 7110 1946 7134 1974
rect 7162 1946 7186 1974
rect 7214 1946 7238 1974
rect 7266 1946 7290 1974
rect 7318 1946 7342 1974
rect 7370 1946 7394 1974
rect 7422 1946 7446 1974
rect 7474 1946 7498 1974
rect 7526 1946 7554 1974
rect 7054 1538 7554 1946
rect 9554 18046 10054 18454
rect 9554 18018 9582 18046
rect 9610 18018 9634 18046
rect 9662 18018 9686 18046
rect 9714 18018 9738 18046
rect 9766 18018 9790 18046
rect 9818 18018 9842 18046
rect 9870 18018 9894 18046
rect 9922 18018 9946 18046
rect 9974 18018 9998 18046
rect 10026 18018 10054 18046
rect 9554 17262 10054 18018
rect 9554 17234 9582 17262
rect 9610 17234 9634 17262
rect 9662 17234 9686 17262
rect 9714 17234 9738 17262
rect 9766 17234 9790 17262
rect 9818 17234 9842 17262
rect 9870 17234 9894 17262
rect 9922 17234 9946 17262
rect 9974 17234 9998 17262
rect 10026 17234 10054 17262
rect 9554 16478 10054 17234
rect 9554 16450 9582 16478
rect 9610 16450 9634 16478
rect 9662 16450 9686 16478
rect 9714 16450 9738 16478
rect 9766 16450 9790 16478
rect 9818 16450 9842 16478
rect 9870 16450 9894 16478
rect 9922 16450 9946 16478
rect 9974 16450 9998 16478
rect 10026 16450 10054 16478
rect 9554 15694 10054 16450
rect 12054 18438 12554 18454
rect 12054 18410 12082 18438
rect 12110 18410 12134 18438
rect 12162 18410 12186 18438
rect 12214 18410 12238 18438
rect 12266 18410 12290 18438
rect 12318 18410 12342 18438
rect 12370 18410 12394 18438
rect 12422 18410 12446 18438
rect 12474 18410 12498 18438
rect 12526 18410 12554 18438
rect 12054 17654 12554 18410
rect 12054 17626 12082 17654
rect 12110 17626 12134 17654
rect 12162 17626 12186 17654
rect 12214 17626 12238 17654
rect 12266 17626 12290 17654
rect 12318 17626 12342 17654
rect 12370 17626 12394 17654
rect 12422 17626 12446 17654
rect 12474 17626 12498 17654
rect 12526 17626 12554 17654
rect 12054 16870 12554 17626
rect 12054 16842 12082 16870
rect 12110 16842 12134 16870
rect 12162 16842 12186 16870
rect 12214 16842 12238 16870
rect 12266 16842 12290 16870
rect 12318 16842 12342 16870
rect 12370 16842 12394 16870
rect 12422 16842 12446 16870
rect 12474 16842 12498 16870
rect 12526 16842 12554 16870
rect 9554 15666 9582 15694
rect 9610 15666 9634 15694
rect 9662 15666 9686 15694
rect 9714 15666 9738 15694
rect 9766 15666 9790 15694
rect 9818 15666 9842 15694
rect 9870 15666 9894 15694
rect 9922 15666 9946 15694
rect 9974 15666 9998 15694
rect 10026 15666 10054 15694
rect 9554 14910 10054 15666
rect 10094 16282 10122 16287
rect 10094 15498 10122 16254
rect 10094 15465 10122 15470
rect 12054 16086 12554 16842
rect 12054 16058 12082 16086
rect 12110 16058 12134 16086
rect 12162 16058 12186 16086
rect 12214 16058 12238 16086
rect 12266 16058 12290 16086
rect 12318 16058 12342 16086
rect 12370 16058 12394 16086
rect 12422 16058 12446 16086
rect 12474 16058 12498 16086
rect 12526 16058 12554 16086
rect 9554 14882 9582 14910
rect 9610 14882 9634 14910
rect 9662 14882 9686 14910
rect 9714 14882 9738 14910
rect 9766 14882 9790 14910
rect 9818 14882 9842 14910
rect 9870 14882 9894 14910
rect 9922 14882 9946 14910
rect 9974 14882 9998 14910
rect 10026 14882 10054 14910
rect 9554 14126 10054 14882
rect 9554 14098 9582 14126
rect 9610 14098 9634 14126
rect 9662 14098 9686 14126
rect 9714 14098 9738 14126
rect 9766 14098 9790 14126
rect 9818 14098 9842 14126
rect 9870 14098 9894 14126
rect 9922 14098 9946 14126
rect 9974 14098 9998 14126
rect 10026 14098 10054 14126
rect 9554 13342 10054 14098
rect 9554 13314 9582 13342
rect 9610 13314 9634 13342
rect 9662 13314 9686 13342
rect 9714 13314 9738 13342
rect 9766 13314 9790 13342
rect 9818 13314 9842 13342
rect 9870 13314 9894 13342
rect 9922 13314 9946 13342
rect 9974 13314 9998 13342
rect 10026 13314 10054 13342
rect 9554 12558 10054 13314
rect 9554 12530 9582 12558
rect 9610 12530 9634 12558
rect 9662 12530 9686 12558
rect 9714 12530 9738 12558
rect 9766 12530 9790 12558
rect 9818 12530 9842 12558
rect 9870 12530 9894 12558
rect 9922 12530 9946 12558
rect 9974 12530 9998 12558
rect 10026 12530 10054 12558
rect 9554 11774 10054 12530
rect 9554 11746 9582 11774
rect 9610 11746 9634 11774
rect 9662 11746 9686 11774
rect 9714 11746 9738 11774
rect 9766 11746 9790 11774
rect 9818 11746 9842 11774
rect 9870 11746 9894 11774
rect 9922 11746 9946 11774
rect 9974 11746 9998 11774
rect 10026 11746 10054 11774
rect 9554 10990 10054 11746
rect 9554 10962 9582 10990
rect 9610 10962 9634 10990
rect 9662 10962 9686 10990
rect 9714 10962 9738 10990
rect 9766 10962 9790 10990
rect 9818 10962 9842 10990
rect 9870 10962 9894 10990
rect 9922 10962 9946 10990
rect 9974 10962 9998 10990
rect 10026 10962 10054 10990
rect 9554 10206 10054 10962
rect 9554 10178 9582 10206
rect 9610 10178 9634 10206
rect 9662 10178 9686 10206
rect 9714 10178 9738 10206
rect 9766 10178 9790 10206
rect 9818 10178 9842 10206
rect 9870 10178 9894 10206
rect 9922 10178 9946 10206
rect 9974 10178 9998 10206
rect 10026 10178 10054 10206
rect 9554 9422 10054 10178
rect 9554 9394 9582 9422
rect 9610 9394 9634 9422
rect 9662 9394 9686 9422
rect 9714 9394 9738 9422
rect 9766 9394 9790 9422
rect 9818 9394 9842 9422
rect 9870 9394 9894 9422
rect 9922 9394 9946 9422
rect 9974 9394 9998 9422
rect 10026 9394 10054 9422
rect 9554 8638 10054 9394
rect 9554 8610 9582 8638
rect 9610 8610 9634 8638
rect 9662 8610 9686 8638
rect 9714 8610 9738 8638
rect 9766 8610 9790 8638
rect 9818 8610 9842 8638
rect 9870 8610 9894 8638
rect 9922 8610 9946 8638
rect 9974 8610 9998 8638
rect 10026 8610 10054 8638
rect 9554 7854 10054 8610
rect 9554 7826 9582 7854
rect 9610 7826 9634 7854
rect 9662 7826 9686 7854
rect 9714 7826 9738 7854
rect 9766 7826 9790 7854
rect 9818 7826 9842 7854
rect 9870 7826 9894 7854
rect 9922 7826 9946 7854
rect 9974 7826 9998 7854
rect 10026 7826 10054 7854
rect 9554 7070 10054 7826
rect 9554 7042 9582 7070
rect 9610 7042 9634 7070
rect 9662 7042 9686 7070
rect 9714 7042 9738 7070
rect 9766 7042 9790 7070
rect 9818 7042 9842 7070
rect 9870 7042 9894 7070
rect 9922 7042 9946 7070
rect 9974 7042 9998 7070
rect 10026 7042 10054 7070
rect 9554 6286 10054 7042
rect 9554 6258 9582 6286
rect 9610 6258 9634 6286
rect 9662 6258 9686 6286
rect 9714 6258 9738 6286
rect 9766 6258 9790 6286
rect 9818 6258 9842 6286
rect 9870 6258 9894 6286
rect 9922 6258 9946 6286
rect 9974 6258 9998 6286
rect 10026 6258 10054 6286
rect 9554 5502 10054 6258
rect 9554 5474 9582 5502
rect 9610 5474 9634 5502
rect 9662 5474 9686 5502
rect 9714 5474 9738 5502
rect 9766 5474 9790 5502
rect 9818 5474 9842 5502
rect 9870 5474 9894 5502
rect 9922 5474 9946 5502
rect 9974 5474 9998 5502
rect 10026 5474 10054 5502
rect 9554 4718 10054 5474
rect 9554 4690 9582 4718
rect 9610 4690 9634 4718
rect 9662 4690 9686 4718
rect 9714 4690 9738 4718
rect 9766 4690 9790 4718
rect 9818 4690 9842 4718
rect 9870 4690 9894 4718
rect 9922 4690 9946 4718
rect 9974 4690 9998 4718
rect 10026 4690 10054 4718
rect 9554 3934 10054 4690
rect 9554 3906 9582 3934
rect 9610 3906 9634 3934
rect 9662 3906 9686 3934
rect 9714 3906 9738 3934
rect 9766 3906 9790 3934
rect 9818 3906 9842 3934
rect 9870 3906 9894 3934
rect 9922 3906 9946 3934
rect 9974 3906 9998 3934
rect 10026 3906 10054 3934
rect 9554 3150 10054 3906
rect 9554 3122 9582 3150
rect 9610 3122 9634 3150
rect 9662 3122 9686 3150
rect 9714 3122 9738 3150
rect 9766 3122 9790 3150
rect 9818 3122 9842 3150
rect 9870 3122 9894 3150
rect 9922 3122 9946 3150
rect 9974 3122 9998 3150
rect 10026 3122 10054 3150
rect 9554 2366 10054 3122
rect 9554 2338 9582 2366
rect 9610 2338 9634 2366
rect 9662 2338 9686 2366
rect 9714 2338 9738 2366
rect 9766 2338 9790 2366
rect 9818 2338 9842 2366
rect 9870 2338 9894 2366
rect 9922 2338 9946 2366
rect 9974 2338 9998 2366
rect 10026 2338 10054 2366
rect 9554 1582 10054 2338
rect 9554 1554 9582 1582
rect 9610 1554 9634 1582
rect 9662 1554 9686 1582
rect 9714 1554 9738 1582
rect 9766 1554 9790 1582
rect 9818 1554 9842 1582
rect 9870 1554 9894 1582
rect 9922 1554 9946 1582
rect 9974 1554 9998 1582
rect 10026 1554 10054 1582
rect 9554 1538 10054 1554
rect 12054 15302 12554 16058
rect 12054 15274 12082 15302
rect 12110 15274 12134 15302
rect 12162 15274 12186 15302
rect 12214 15274 12238 15302
rect 12266 15274 12290 15302
rect 12318 15274 12342 15302
rect 12370 15274 12394 15302
rect 12422 15274 12446 15302
rect 12474 15274 12498 15302
rect 12526 15274 12554 15302
rect 12054 14518 12554 15274
rect 12054 14490 12082 14518
rect 12110 14490 12134 14518
rect 12162 14490 12186 14518
rect 12214 14490 12238 14518
rect 12266 14490 12290 14518
rect 12318 14490 12342 14518
rect 12370 14490 12394 14518
rect 12422 14490 12446 14518
rect 12474 14490 12498 14518
rect 12526 14490 12554 14518
rect 12054 13734 12554 14490
rect 12054 13706 12082 13734
rect 12110 13706 12134 13734
rect 12162 13706 12186 13734
rect 12214 13706 12238 13734
rect 12266 13706 12290 13734
rect 12318 13706 12342 13734
rect 12370 13706 12394 13734
rect 12422 13706 12446 13734
rect 12474 13706 12498 13734
rect 12526 13706 12554 13734
rect 12054 12950 12554 13706
rect 12054 12922 12082 12950
rect 12110 12922 12134 12950
rect 12162 12922 12186 12950
rect 12214 12922 12238 12950
rect 12266 12922 12290 12950
rect 12318 12922 12342 12950
rect 12370 12922 12394 12950
rect 12422 12922 12446 12950
rect 12474 12922 12498 12950
rect 12526 12922 12554 12950
rect 12054 12166 12554 12922
rect 12054 12138 12082 12166
rect 12110 12138 12134 12166
rect 12162 12138 12186 12166
rect 12214 12138 12238 12166
rect 12266 12138 12290 12166
rect 12318 12138 12342 12166
rect 12370 12138 12394 12166
rect 12422 12138 12446 12166
rect 12474 12138 12498 12166
rect 12526 12138 12554 12166
rect 12054 11382 12554 12138
rect 12054 11354 12082 11382
rect 12110 11354 12134 11382
rect 12162 11354 12186 11382
rect 12214 11354 12238 11382
rect 12266 11354 12290 11382
rect 12318 11354 12342 11382
rect 12370 11354 12394 11382
rect 12422 11354 12446 11382
rect 12474 11354 12498 11382
rect 12526 11354 12554 11382
rect 12054 10598 12554 11354
rect 12054 10570 12082 10598
rect 12110 10570 12134 10598
rect 12162 10570 12186 10598
rect 12214 10570 12238 10598
rect 12266 10570 12290 10598
rect 12318 10570 12342 10598
rect 12370 10570 12394 10598
rect 12422 10570 12446 10598
rect 12474 10570 12498 10598
rect 12526 10570 12554 10598
rect 12054 9814 12554 10570
rect 12054 9786 12082 9814
rect 12110 9786 12134 9814
rect 12162 9786 12186 9814
rect 12214 9786 12238 9814
rect 12266 9786 12290 9814
rect 12318 9786 12342 9814
rect 12370 9786 12394 9814
rect 12422 9786 12446 9814
rect 12474 9786 12498 9814
rect 12526 9786 12554 9814
rect 12054 9030 12554 9786
rect 12054 9002 12082 9030
rect 12110 9002 12134 9030
rect 12162 9002 12186 9030
rect 12214 9002 12238 9030
rect 12266 9002 12290 9030
rect 12318 9002 12342 9030
rect 12370 9002 12394 9030
rect 12422 9002 12446 9030
rect 12474 9002 12498 9030
rect 12526 9002 12554 9030
rect 12054 8246 12554 9002
rect 12054 8218 12082 8246
rect 12110 8218 12134 8246
rect 12162 8218 12186 8246
rect 12214 8218 12238 8246
rect 12266 8218 12290 8246
rect 12318 8218 12342 8246
rect 12370 8218 12394 8246
rect 12422 8218 12446 8246
rect 12474 8218 12498 8246
rect 12526 8218 12554 8246
rect 12054 7462 12554 8218
rect 12054 7434 12082 7462
rect 12110 7434 12134 7462
rect 12162 7434 12186 7462
rect 12214 7434 12238 7462
rect 12266 7434 12290 7462
rect 12318 7434 12342 7462
rect 12370 7434 12394 7462
rect 12422 7434 12446 7462
rect 12474 7434 12498 7462
rect 12526 7434 12554 7462
rect 12054 6678 12554 7434
rect 12054 6650 12082 6678
rect 12110 6650 12134 6678
rect 12162 6650 12186 6678
rect 12214 6650 12238 6678
rect 12266 6650 12290 6678
rect 12318 6650 12342 6678
rect 12370 6650 12394 6678
rect 12422 6650 12446 6678
rect 12474 6650 12498 6678
rect 12526 6650 12554 6678
rect 12054 5894 12554 6650
rect 12054 5866 12082 5894
rect 12110 5866 12134 5894
rect 12162 5866 12186 5894
rect 12214 5866 12238 5894
rect 12266 5866 12290 5894
rect 12318 5866 12342 5894
rect 12370 5866 12394 5894
rect 12422 5866 12446 5894
rect 12474 5866 12498 5894
rect 12526 5866 12554 5894
rect 12054 5110 12554 5866
rect 12054 5082 12082 5110
rect 12110 5082 12134 5110
rect 12162 5082 12186 5110
rect 12214 5082 12238 5110
rect 12266 5082 12290 5110
rect 12318 5082 12342 5110
rect 12370 5082 12394 5110
rect 12422 5082 12446 5110
rect 12474 5082 12498 5110
rect 12526 5082 12554 5110
rect 12054 4326 12554 5082
rect 12054 4298 12082 4326
rect 12110 4298 12134 4326
rect 12162 4298 12186 4326
rect 12214 4298 12238 4326
rect 12266 4298 12290 4326
rect 12318 4298 12342 4326
rect 12370 4298 12394 4326
rect 12422 4298 12446 4326
rect 12474 4298 12498 4326
rect 12526 4298 12554 4326
rect 12054 3542 12554 4298
rect 12054 3514 12082 3542
rect 12110 3514 12134 3542
rect 12162 3514 12186 3542
rect 12214 3514 12238 3542
rect 12266 3514 12290 3542
rect 12318 3514 12342 3542
rect 12370 3514 12394 3542
rect 12422 3514 12446 3542
rect 12474 3514 12498 3542
rect 12526 3514 12554 3542
rect 12054 2758 12554 3514
rect 12054 2730 12082 2758
rect 12110 2730 12134 2758
rect 12162 2730 12186 2758
rect 12214 2730 12238 2758
rect 12266 2730 12290 2758
rect 12318 2730 12342 2758
rect 12370 2730 12394 2758
rect 12422 2730 12446 2758
rect 12474 2730 12498 2758
rect 12526 2730 12554 2758
rect 12054 1974 12554 2730
rect 12054 1946 12082 1974
rect 12110 1946 12134 1974
rect 12162 1946 12186 1974
rect 12214 1946 12238 1974
rect 12266 1946 12290 1974
rect 12318 1946 12342 1974
rect 12370 1946 12394 1974
rect 12422 1946 12446 1974
rect 12474 1946 12498 1974
rect 12526 1946 12554 1974
rect 12054 1538 12554 1946
rect 14554 18046 15054 18454
rect 14554 18018 14582 18046
rect 14610 18018 14634 18046
rect 14662 18018 14686 18046
rect 14714 18018 14738 18046
rect 14766 18018 14790 18046
rect 14818 18018 14842 18046
rect 14870 18018 14894 18046
rect 14922 18018 14946 18046
rect 14974 18018 14998 18046
rect 15026 18018 15054 18046
rect 14554 17262 15054 18018
rect 14554 17234 14582 17262
rect 14610 17234 14634 17262
rect 14662 17234 14686 17262
rect 14714 17234 14738 17262
rect 14766 17234 14790 17262
rect 14818 17234 14842 17262
rect 14870 17234 14894 17262
rect 14922 17234 14946 17262
rect 14974 17234 14998 17262
rect 15026 17234 15054 17262
rect 14554 16478 15054 17234
rect 14554 16450 14582 16478
rect 14610 16450 14634 16478
rect 14662 16450 14686 16478
rect 14714 16450 14738 16478
rect 14766 16450 14790 16478
rect 14818 16450 14842 16478
rect 14870 16450 14894 16478
rect 14922 16450 14946 16478
rect 14974 16450 14998 16478
rect 15026 16450 15054 16478
rect 14554 15694 15054 16450
rect 14554 15666 14582 15694
rect 14610 15666 14634 15694
rect 14662 15666 14686 15694
rect 14714 15666 14738 15694
rect 14766 15666 14790 15694
rect 14818 15666 14842 15694
rect 14870 15666 14894 15694
rect 14922 15666 14946 15694
rect 14974 15666 14998 15694
rect 15026 15666 15054 15694
rect 14554 14910 15054 15666
rect 14554 14882 14582 14910
rect 14610 14882 14634 14910
rect 14662 14882 14686 14910
rect 14714 14882 14738 14910
rect 14766 14882 14790 14910
rect 14818 14882 14842 14910
rect 14870 14882 14894 14910
rect 14922 14882 14946 14910
rect 14974 14882 14998 14910
rect 15026 14882 15054 14910
rect 14554 14126 15054 14882
rect 14554 14098 14582 14126
rect 14610 14098 14634 14126
rect 14662 14098 14686 14126
rect 14714 14098 14738 14126
rect 14766 14098 14790 14126
rect 14818 14098 14842 14126
rect 14870 14098 14894 14126
rect 14922 14098 14946 14126
rect 14974 14098 14998 14126
rect 15026 14098 15054 14126
rect 14554 13342 15054 14098
rect 14554 13314 14582 13342
rect 14610 13314 14634 13342
rect 14662 13314 14686 13342
rect 14714 13314 14738 13342
rect 14766 13314 14790 13342
rect 14818 13314 14842 13342
rect 14870 13314 14894 13342
rect 14922 13314 14946 13342
rect 14974 13314 14998 13342
rect 15026 13314 15054 13342
rect 14554 12558 15054 13314
rect 14554 12530 14582 12558
rect 14610 12530 14634 12558
rect 14662 12530 14686 12558
rect 14714 12530 14738 12558
rect 14766 12530 14790 12558
rect 14818 12530 14842 12558
rect 14870 12530 14894 12558
rect 14922 12530 14946 12558
rect 14974 12530 14998 12558
rect 15026 12530 15054 12558
rect 14554 11774 15054 12530
rect 14554 11746 14582 11774
rect 14610 11746 14634 11774
rect 14662 11746 14686 11774
rect 14714 11746 14738 11774
rect 14766 11746 14790 11774
rect 14818 11746 14842 11774
rect 14870 11746 14894 11774
rect 14922 11746 14946 11774
rect 14974 11746 14998 11774
rect 15026 11746 15054 11774
rect 14554 10990 15054 11746
rect 14554 10962 14582 10990
rect 14610 10962 14634 10990
rect 14662 10962 14686 10990
rect 14714 10962 14738 10990
rect 14766 10962 14790 10990
rect 14818 10962 14842 10990
rect 14870 10962 14894 10990
rect 14922 10962 14946 10990
rect 14974 10962 14998 10990
rect 15026 10962 15054 10990
rect 14554 10206 15054 10962
rect 14554 10178 14582 10206
rect 14610 10178 14634 10206
rect 14662 10178 14686 10206
rect 14714 10178 14738 10206
rect 14766 10178 14790 10206
rect 14818 10178 14842 10206
rect 14870 10178 14894 10206
rect 14922 10178 14946 10206
rect 14974 10178 14998 10206
rect 15026 10178 15054 10206
rect 14554 9422 15054 10178
rect 14554 9394 14582 9422
rect 14610 9394 14634 9422
rect 14662 9394 14686 9422
rect 14714 9394 14738 9422
rect 14766 9394 14790 9422
rect 14818 9394 14842 9422
rect 14870 9394 14894 9422
rect 14922 9394 14946 9422
rect 14974 9394 14998 9422
rect 15026 9394 15054 9422
rect 14554 8638 15054 9394
rect 14554 8610 14582 8638
rect 14610 8610 14634 8638
rect 14662 8610 14686 8638
rect 14714 8610 14738 8638
rect 14766 8610 14790 8638
rect 14818 8610 14842 8638
rect 14870 8610 14894 8638
rect 14922 8610 14946 8638
rect 14974 8610 14998 8638
rect 15026 8610 15054 8638
rect 14554 7854 15054 8610
rect 14554 7826 14582 7854
rect 14610 7826 14634 7854
rect 14662 7826 14686 7854
rect 14714 7826 14738 7854
rect 14766 7826 14790 7854
rect 14818 7826 14842 7854
rect 14870 7826 14894 7854
rect 14922 7826 14946 7854
rect 14974 7826 14998 7854
rect 15026 7826 15054 7854
rect 14554 7070 15054 7826
rect 14554 7042 14582 7070
rect 14610 7042 14634 7070
rect 14662 7042 14686 7070
rect 14714 7042 14738 7070
rect 14766 7042 14790 7070
rect 14818 7042 14842 7070
rect 14870 7042 14894 7070
rect 14922 7042 14946 7070
rect 14974 7042 14998 7070
rect 15026 7042 15054 7070
rect 14554 6286 15054 7042
rect 14554 6258 14582 6286
rect 14610 6258 14634 6286
rect 14662 6258 14686 6286
rect 14714 6258 14738 6286
rect 14766 6258 14790 6286
rect 14818 6258 14842 6286
rect 14870 6258 14894 6286
rect 14922 6258 14946 6286
rect 14974 6258 14998 6286
rect 15026 6258 15054 6286
rect 14554 5502 15054 6258
rect 14554 5474 14582 5502
rect 14610 5474 14634 5502
rect 14662 5474 14686 5502
rect 14714 5474 14738 5502
rect 14766 5474 14790 5502
rect 14818 5474 14842 5502
rect 14870 5474 14894 5502
rect 14922 5474 14946 5502
rect 14974 5474 14998 5502
rect 15026 5474 15054 5502
rect 14554 4718 15054 5474
rect 14554 4690 14582 4718
rect 14610 4690 14634 4718
rect 14662 4690 14686 4718
rect 14714 4690 14738 4718
rect 14766 4690 14790 4718
rect 14818 4690 14842 4718
rect 14870 4690 14894 4718
rect 14922 4690 14946 4718
rect 14974 4690 14998 4718
rect 15026 4690 15054 4718
rect 14554 3934 15054 4690
rect 14554 3906 14582 3934
rect 14610 3906 14634 3934
rect 14662 3906 14686 3934
rect 14714 3906 14738 3934
rect 14766 3906 14790 3934
rect 14818 3906 14842 3934
rect 14870 3906 14894 3934
rect 14922 3906 14946 3934
rect 14974 3906 14998 3934
rect 15026 3906 15054 3934
rect 14554 3150 15054 3906
rect 14554 3122 14582 3150
rect 14610 3122 14634 3150
rect 14662 3122 14686 3150
rect 14714 3122 14738 3150
rect 14766 3122 14790 3150
rect 14818 3122 14842 3150
rect 14870 3122 14894 3150
rect 14922 3122 14946 3150
rect 14974 3122 14998 3150
rect 15026 3122 15054 3150
rect 14554 2366 15054 3122
rect 14554 2338 14582 2366
rect 14610 2338 14634 2366
rect 14662 2338 14686 2366
rect 14714 2338 14738 2366
rect 14766 2338 14790 2366
rect 14818 2338 14842 2366
rect 14870 2338 14894 2366
rect 14922 2338 14946 2366
rect 14974 2338 14998 2366
rect 15026 2338 15054 2366
rect 14554 1582 15054 2338
rect 14554 1554 14582 1582
rect 14610 1554 14634 1582
rect 14662 1554 14686 1582
rect 14714 1554 14738 1582
rect 14766 1554 14790 1582
rect 14818 1554 14842 1582
rect 14870 1554 14894 1582
rect 14922 1554 14946 1582
rect 14974 1554 14998 1582
rect 15026 1554 15054 1582
rect 14554 1538 15054 1554
rect 17054 18438 17554 18454
rect 17054 18410 17082 18438
rect 17110 18410 17134 18438
rect 17162 18410 17186 18438
rect 17214 18410 17238 18438
rect 17266 18410 17290 18438
rect 17318 18410 17342 18438
rect 17370 18410 17394 18438
rect 17422 18410 17446 18438
rect 17474 18410 17498 18438
rect 17526 18410 17554 18438
rect 17054 17654 17554 18410
rect 17054 17626 17082 17654
rect 17110 17626 17134 17654
rect 17162 17626 17186 17654
rect 17214 17626 17238 17654
rect 17266 17626 17290 17654
rect 17318 17626 17342 17654
rect 17370 17626 17394 17654
rect 17422 17626 17446 17654
rect 17474 17626 17498 17654
rect 17526 17626 17554 17654
rect 17054 16870 17554 17626
rect 17054 16842 17082 16870
rect 17110 16842 17134 16870
rect 17162 16842 17186 16870
rect 17214 16842 17238 16870
rect 17266 16842 17290 16870
rect 17318 16842 17342 16870
rect 17370 16842 17394 16870
rect 17422 16842 17446 16870
rect 17474 16842 17498 16870
rect 17526 16842 17554 16870
rect 17054 16086 17554 16842
rect 17054 16058 17082 16086
rect 17110 16058 17134 16086
rect 17162 16058 17186 16086
rect 17214 16058 17238 16086
rect 17266 16058 17290 16086
rect 17318 16058 17342 16086
rect 17370 16058 17394 16086
rect 17422 16058 17446 16086
rect 17474 16058 17498 16086
rect 17526 16058 17554 16086
rect 17054 15302 17554 16058
rect 17054 15274 17082 15302
rect 17110 15274 17134 15302
rect 17162 15274 17186 15302
rect 17214 15274 17238 15302
rect 17266 15274 17290 15302
rect 17318 15274 17342 15302
rect 17370 15274 17394 15302
rect 17422 15274 17446 15302
rect 17474 15274 17498 15302
rect 17526 15274 17554 15302
rect 17054 14518 17554 15274
rect 17054 14490 17082 14518
rect 17110 14490 17134 14518
rect 17162 14490 17186 14518
rect 17214 14490 17238 14518
rect 17266 14490 17290 14518
rect 17318 14490 17342 14518
rect 17370 14490 17394 14518
rect 17422 14490 17446 14518
rect 17474 14490 17498 14518
rect 17526 14490 17554 14518
rect 17054 13734 17554 14490
rect 17054 13706 17082 13734
rect 17110 13706 17134 13734
rect 17162 13706 17186 13734
rect 17214 13706 17238 13734
rect 17266 13706 17290 13734
rect 17318 13706 17342 13734
rect 17370 13706 17394 13734
rect 17422 13706 17446 13734
rect 17474 13706 17498 13734
rect 17526 13706 17554 13734
rect 17054 12950 17554 13706
rect 17054 12922 17082 12950
rect 17110 12922 17134 12950
rect 17162 12922 17186 12950
rect 17214 12922 17238 12950
rect 17266 12922 17290 12950
rect 17318 12922 17342 12950
rect 17370 12922 17394 12950
rect 17422 12922 17446 12950
rect 17474 12922 17498 12950
rect 17526 12922 17554 12950
rect 17054 12166 17554 12922
rect 17054 12138 17082 12166
rect 17110 12138 17134 12166
rect 17162 12138 17186 12166
rect 17214 12138 17238 12166
rect 17266 12138 17290 12166
rect 17318 12138 17342 12166
rect 17370 12138 17394 12166
rect 17422 12138 17446 12166
rect 17474 12138 17498 12166
rect 17526 12138 17554 12166
rect 17054 11382 17554 12138
rect 17054 11354 17082 11382
rect 17110 11354 17134 11382
rect 17162 11354 17186 11382
rect 17214 11354 17238 11382
rect 17266 11354 17290 11382
rect 17318 11354 17342 11382
rect 17370 11354 17394 11382
rect 17422 11354 17446 11382
rect 17474 11354 17498 11382
rect 17526 11354 17554 11382
rect 17054 10598 17554 11354
rect 17054 10570 17082 10598
rect 17110 10570 17134 10598
rect 17162 10570 17186 10598
rect 17214 10570 17238 10598
rect 17266 10570 17290 10598
rect 17318 10570 17342 10598
rect 17370 10570 17394 10598
rect 17422 10570 17446 10598
rect 17474 10570 17498 10598
rect 17526 10570 17554 10598
rect 17054 9814 17554 10570
rect 17054 9786 17082 9814
rect 17110 9786 17134 9814
rect 17162 9786 17186 9814
rect 17214 9786 17238 9814
rect 17266 9786 17290 9814
rect 17318 9786 17342 9814
rect 17370 9786 17394 9814
rect 17422 9786 17446 9814
rect 17474 9786 17498 9814
rect 17526 9786 17554 9814
rect 17054 9030 17554 9786
rect 17054 9002 17082 9030
rect 17110 9002 17134 9030
rect 17162 9002 17186 9030
rect 17214 9002 17238 9030
rect 17266 9002 17290 9030
rect 17318 9002 17342 9030
rect 17370 9002 17394 9030
rect 17422 9002 17446 9030
rect 17474 9002 17498 9030
rect 17526 9002 17554 9030
rect 17054 8246 17554 9002
rect 17054 8218 17082 8246
rect 17110 8218 17134 8246
rect 17162 8218 17186 8246
rect 17214 8218 17238 8246
rect 17266 8218 17290 8246
rect 17318 8218 17342 8246
rect 17370 8218 17394 8246
rect 17422 8218 17446 8246
rect 17474 8218 17498 8246
rect 17526 8218 17554 8246
rect 17054 7462 17554 8218
rect 17054 7434 17082 7462
rect 17110 7434 17134 7462
rect 17162 7434 17186 7462
rect 17214 7434 17238 7462
rect 17266 7434 17290 7462
rect 17318 7434 17342 7462
rect 17370 7434 17394 7462
rect 17422 7434 17446 7462
rect 17474 7434 17498 7462
rect 17526 7434 17554 7462
rect 17054 6678 17554 7434
rect 17054 6650 17082 6678
rect 17110 6650 17134 6678
rect 17162 6650 17186 6678
rect 17214 6650 17238 6678
rect 17266 6650 17290 6678
rect 17318 6650 17342 6678
rect 17370 6650 17394 6678
rect 17422 6650 17446 6678
rect 17474 6650 17498 6678
rect 17526 6650 17554 6678
rect 17054 5894 17554 6650
rect 17054 5866 17082 5894
rect 17110 5866 17134 5894
rect 17162 5866 17186 5894
rect 17214 5866 17238 5894
rect 17266 5866 17290 5894
rect 17318 5866 17342 5894
rect 17370 5866 17394 5894
rect 17422 5866 17446 5894
rect 17474 5866 17498 5894
rect 17526 5866 17554 5894
rect 17054 5110 17554 5866
rect 17054 5082 17082 5110
rect 17110 5082 17134 5110
rect 17162 5082 17186 5110
rect 17214 5082 17238 5110
rect 17266 5082 17290 5110
rect 17318 5082 17342 5110
rect 17370 5082 17394 5110
rect 17422 5082 17446 5110
rect 17474 5082 17498 5110
rect 17526 5082 17554 5110
rect 17054 4326 17554 5082
rect 17054 4298 17082 4326
rect 17110 4298 17134 4326
rect 17162 4298 17186 4326
rect 17214 4298 17238 4326
rect 17266 4298 17290 4326
rect 17318 4298 17342 4326
rect 17370 4298 17394 4326
rect 17422 4298 17446 4326
rect 17474 4298 17498 4326
rect 17526 4298 17554 4326
rect 17054 3542 17554 4298
rect 17054 3514 17082 3542
rect 17110 3514 17134 3542
rect 17162 3514 17186 3542
rect 17214 3514 17238 3542
rect 17266 3514 17290 3542
rect 17318 3514 17342 3542
rect 17370 3514 17394 3542
rect 17422 3514 17446 3542
rect 17474 3514 17498 3542
rect 17526 3514 17554 3542
rect 17054 2758 17554 3514
rect 17054 2730 17082 2758
rect 17110 2730 17134 2758
rect 17162 2730 17186 2758
rect 17214 2730 17238 2758
rect 17266 2730 17290 2758
rect 17318 2730 17342 2758
rect 17370 2730 17394 2758
rect 17422 2730 17446 2758
rect 17474 2730 17498 2758
rect 17526 2730 17554 2758
rect 17054 1974 17554 2730
rect 17054 1946 17082 1974
rect 17110 1946 17134 1974
rect 17162 1946 17186 1974
rect 17214 1946 17238 1974
rect 17266 1946 17290 1974
rect 17318 1946 17342 1974
rect 17370 1946 17394 1974
rect 17422 1946 17446 1974
rect 17474 1946 17498 1974
rect 17526 1946 17554 1974
rect 17054 1538 17554 1946
rect 19554 18046 20054 18454
rect 19554 18018 19582 18046
rect 19610 18018 19634 18046
rect 19662 18018 19686 18046
rect 19714 18018 19738 18046
rect 19766 18018 19790 18046
rect 19818 18018 19842 18046
rect 19870 18018 19894 18046
rect 19922 18018 19946 18046
rect 19974 18018 19998 18046
rect 20026 18018 20054 18046
rect 19554 17262 20054 18018
rect 19554 17234 19582 17262
rect 19610 17234 19634 17262
rect 19662 17234 19686 17262
rect 19714 17234 19738 17262
rect 19766 17234 19790 17262
rect 19818 17234 19842 17262
rect 19870 17234 19894 17262
rect 19922 17234 19946 17262
rect 19974 17234 19998 17262
rect 20026 17234 20054 17262
rect 19554 16478 20054 17234
rect 19554 16450 19582 16478
rect 19610 16450 19634 16478
rect 19662 16450 19686 16478
rect 19714 16450 19738 16478
rect 19766 16450 19790 16478
rect 19818 16450 19842 16478
rect 19870 16450 19894 16478
rect 19922 16450 19946 16478
rect 19974 16450 19998 16478
rect 20026 16450 20054 16478
rect 19554 15694 20054 16450
rect 19554 15666 19582 15694
rect 19610 15666 19634 15694
rect 19662 15666 19686 15694
rect 19714 15666 19738 15694
rect 19766 15666 19790 15694
rect 19818 15666 19842 15694
rect 19870 15666 19894 15694
rect 19922 15666 19946 15694
rect 19974 15666 19998 15694
rect 20026 15666 20054 15694
rect 19554 14910 20054 15666
rect 19554 14882 19582 14910
rect 19610 14882 19634 14910
rect 19662 14882 19686 14910
rect 19714 14882 19738 14910
rect 19766 14882 19790 14910
rect 19818 14882 19842 14910
rect 19870 14882 19894 14910
rect 19922 14882 19946 14910
rect 19974 14882 19998 14910
rect 20026 14882 20054 14910
rect 19554 14126 20054 14882
rect 19554 14098 19582 14126
rect 19610 14098 19634 14126
rect 19662 14098 19686 14126
rect 19714 14098 19738 14126
rect 19766 14098 19790 14126
rect 19818 14098 19842 14126
rect 19870 14098 19894 14126
rect 19922 14098 19946 14126
rect 19974 14098 19998 14126
rect 20026 14098 20054 14126
rect 19554 13342 20054 14098
rect 19554 13314 19582 13342
rect 19610 13314 19634 13342
rect 19662 13314 19686 13342
rect 19714 13314 19738 13342
rect 19766 13314 19790 13342
rect 19818 13314 19842 13342
rect 19870 13314 19894 13342
rect 19922 13314 19946 13342
rect 19974 13314 19998 13342
rect 20026 13314 20054 13342
rect 19554 12558 20054 13314
rect 19554 12530 19582 12558
rect 19610 12530 19634 12558
rect 19662 12530 19686 12558
rect 19714 12530 19738 12558
rect 19766 12530 19790 12558
rect 19818 12530 19842 12558
rect 19870 12530 19894 12558
rect 19922 12530 19946 12558
rect 19974 12530 19998 12558
rect 20026 12530 20054 12558
rect 19554 11774 20054 12530
rect 19554 11746 19582 11774
rect 19610 11746 19634 11774
rect 19662 11746 19686 11774
rect 19714 11746 19738 11774
rect 19766 11746 19790 11774
rect 19818 11746 19842 11774
rect 19870 11746 19894 11774
rect 19922 11746 19946 11774
rect 19974 11746 19998 11774
rect 20026 11746 20054 11774
rect 19554 10990 20054 11746
rect 19554 10962 19582 10990
rect 19610 10962 19634 10990
rect 19662 10962 19686 10990
rect 19714 10962 19738 10990
rect 19766 10962 19790 10990
rect 19818 10962 19842 10990
rect 19870 10962 19894 10990
rect 19922 10962 19946 10990
rect 19974 10962 19998 10990
rect 20026 10962 20054 10990
rect 19554 10206 20054 10962
rect 19554 10178 19582 10206
rect 19610 10178 19634 10206
rect 19662 10178 19686 10206
rect 19714 10178 19738 10206
rect 19766 10178 19790 10206
rect 19818 10178 19842 10206
rect 19870 10178 19894 10206
rect 19922 10178 19946 10206
rect 19974 10178 19998 10206
rect 20026 10178 20054 10206
rect 19554 9422 20054 10178
rect 19554 9394 19582 9422
rect 19610 9394 19634 9422
rect 19662 9394 19686 9422
rect 19714 9394 19738 9422
rect 19766 9394 19790 9422
rect 19818 9394 19842 9422
rect 19870 9394 19894 9422
rect 19922 9394 19946 9422
rect 19974 9394 19998 9422
rect 20026 9394 20054 9422
rect 19554 8638 20054 9394
rect 19554 8610 19582 8638
rect 19610 8610 19634 8638
rect 19662 8610 19686 8638
rect 19714 8610 19738 8638
rect 19766 8610 19790 8638
rect 19818 8610 19842 8638
rect 19870 8610 19894 8638
rect 19922 8610 19946 8638
rect 19974 8610 19998 8638
rect 20026 8610 20054 8638
rect 19554 7854 20054 8610
rect 19554 7826 19582 7854
rect 19610 7826 19634 7854
rect 19662 7826 19686 7854
rect 19714 7826 19738 7854
rect 19766 7826 19790 7854
rect 19818 7826 19842 7854
rect 19870 7826 19894 7854
rect 19922 7826 19946 7854
rect 19974 7826 19998 7854
rect 20026 7826 20054 7854
rect 19554 7070 20054 7826
rect 19554 7042 19582 7070
rect 19610 7042 19634 7070
rect 19662 7042 19686 7070
rect 19714 7042 19738 7070
rect 19766 7042 19790 7070
rect 19818 7042 19842 7070
rect 19870 7042 19894 7070
rect 19922 7042 19946 7070
rect 19974 7042 19998 7070
rect 20026 7042 20054 7070
rect 19554 6286 20054 7042
rect 19554 6258 19582 6286
rect 19610 6258 19634 6286
rect 19662 6258 19686 6286
rect 19714 6258 19738 6286
rect 19766 6258 19790 6286
rect 19818 6258 19842 6286
rect 19870 6258 19894 6286
rect 19922 6258 19946 6286
rect 19974 6258 19998 6286
rect 20026 6258 20054 6286
rect 19554 5502 20054 6258
rect 19554 5474 19582 5502
rect 19610 5474 19634 5502
rect 19662 5474 19686 5502
rect 19714 5474 19738 5502
rect 19766 5474 19790 5502
rect 19818 5474 19842 5502
rect 19870 5474 19894 5502
rect 19922 5474 19946 5502
rect 19974 5474 19998 5502
rect 20026 5474 20054 5502
rect 19554 4718 20054 5474
rect 19554 4690 19582 4718
rect 19610 4690 19634 4718
rect 19662 4690 19686 4718
rect 19714 4690 19738 4718
rect 19766 4690 19790 4718
rect 19818 4690 19842 4718
rect 19870 4690 19894 4718
rect 19922 4690 19946 4718
rect 19974 4690 19998 4718
rect 20026 4690 20054 4718
rect 19554 3934 20054 4690
rect 19554 3906 19582 3934
rect 19610 3906 19634 3934
rect 19662 3906 19686 3934
rect 19714 3906 19738 3934
rect 19766 3906 19790 3934
rect 19818 3906 19842 3934
rect 19870 3906 19894 3934
rect 19922 3906 19946 3934
rect 19974 3906 19998 3934
rect 20026 3906 20054 3934
rect 19554 3150 20054 3906
rect 19554 3122 19582 3150
rect 19610 3122 19634 3150
rect 19662 3122 19686 3150
rect 19714 3122 19738 3150
rect 19766 3122 19790 3150
rect 19818 3122 19842 3150
rect 19870 3122 19894 3150
rect 19922 3122 19946 3150
rect 19974 3122 19998 3150
rect 20026 3122 20054 3150
rect 19554 2366 20054 3122
rect 19554 2338 19582 2366
rect 19610 2338 19634 2366
rect 19662 2338 19686 2366
rect 19714 2338 19738 2366
rect 19766 2338 19790 2366
rect 19818 2338 19842 2366
rect 19870 2338 19894 2366
rect 19922 2338 19946 2366
rect 19974 2338 19998 2366
rect 20026 2338 20054 2366
rect 19554 1582 20054 2338
rect 19554 1554 19582 1582
rect 19610 1554 19634 1582
rect 19662 1554 19686 1582
rect 19714 1554 19738 1582
rect 19766 1554 19790 1582
rect 19818 1554 19842 1582
rect 19870 1554 19894 1582
rect 19922 1554 19946 1582
rect 19974 1554 19998 1582
rect 20026 1554 20054 1582
rect 19554 1538 20054 1554
rect 22054 18438 22554 18454
rect 22054 18410 22082 18438
rect 22110 18410 22134 18438
rect 22162 18410 22186 18438
rect 22214 18410 22238 18438
rect 22266 18410 22290 18438
rect 22318 18410 22342 18438
rect 22370 18410 22394 18438
rect 22422 18410 22446 18438
rect 22474 18410 22498 18438
rect 22526 18410 22554 18438
rect 22054 17654 22554 18410
rect 22054 17626 22082 17654
rect 22110 17626 22134 17654
rect 22162 17626 22186 17654
rect 22214 17626 22238 17654
rect 22266 17626 22290 17654
rect 22318 17626 22342 17654
rect 22370 17626 22394 17654
rect 22422 17626 22446 17654
rect 22474 17626 22498 17654
rect 22526 17626 22554 17654
rect 22054 16870 22554 17626
rect 22054 16842 22082 16870
rect 22110 16842 22134 16870
rect 22162 16842 22186 16870
rect 22214 16842 22238 16870
rect 22266 16842 22290 16870
rect 22318 16842 22342 16870
rect 22370 16842 22394 16870
rect 22422 16842 22446 16870
rect 22474 16842 22498 16870
rect 22526 16842 22554 16870
rect 22054 16086 22554 16842
rect 22054 16058 22082 16086
rect 22110 16058 22134 16086
rect 22162 16058 22186 16086
rect 22214 16058 22238 16086
rect 22266 16058 22290 16086
rect 22318 16058 22342 16086
rect 22370 16058 22394 16086
rect 22422 16058 22446 16086
rect 22474 16058 22498 16086
rect 22526 16058 22554 16086
rect 22054 15302 22554 16058
rect 22054 15274 22082 15302
rect 22110 15274 22134 15302
rect 22162 15274 22186 15302
rect 22214 15274 22238 15302
rect 22266 15274 22290 15302
rect 22318 15274 22342 15302
rect 22370 15274 22394 15302
rect 22422 15274 22446 15302
rect 22474 15274 22498 15302
rect 22526 15274 22554 15302
rect 22054 14518 22554 15274
rect 22054 14490 22082 14518
rect 22110 14490 22134 14518
rect 22162 14490 22186 14518
rect 22214 14490 22238 14518
rect 22266 14490 22290 14518
rect 22318 14490 22342 14518
rect 22370 14490 22394 14518
rect 22422 14490 22446 14518
rect 22474 14490 22498 14518
rect 22526 14490 22554 14518
rect 22054 13734 22554 14490
rect 22054 13706 22082 13734
rect 22110 13706 22134 13734
rect 22162 13706 22186 13734
rect 22214 13706 22238 13734
rect 22266 13706 22290 13734
rect 22318 13706 22342 13734
rect 22370 13706 22394 13734
rect 22422 13706 22446 13734
rect 22474 13706 22498 13734
rect 22526 13706 22554 13734
rect 22054 12950 22554 13706
rect 22054 12922 22082 12950
rect 22110 12922 22134 12950
rect 22162 12922 22186 12950
rect 22214 12922 22238 12950
rect 22266 12922 22290 12950
rect 22318 12922 22342 12950
rect 22370 12922 22394 12950
rect 22422 12922 22446 12950
rect 22474 12922 22498 12950
rect 22526 12922 22554 12950
rect 22054 12166 22554 12922
rect 22054 12138 22082 12166
rect 22110 12138 22134 12166
rect 22162 12138 22186 12166
rect 22214 12138 22238 12166
rect 22266 12138 22290 12166
rect 22318 12138 22342 12166
rect 22370 12138 22394 12166
rect 22422 12138 22446 12166
rect 22474 12138 22498 12166
rect 22526 12138 22554 12166
rect 22054 11382 22554 12138
rect 22054 11354 22082 11382
rect 22110 11354 22134 11382
rect 22162 11354 22186 11382
rect 22214 11354 22238 11382
rect 22266 11354 22290 11382
rect 22318 11354 22342 11382
rect 22370 11354 22394 11382
rect 22422 11354 22446 11382
rect 22474 11354 22498 11382
rect 22526 11354 22554 11382
rect 22054 10598 22554 11354
rect 22054 10570 22082 10598
rect 22110 10570 22134 10598
rect 22162 10570 22186 10598
rect 22214 10570 22238 10598
rect 22266 10570 22290 10598
rect 22318 10570 22342 10598
rect 22370 10570 22394 10598
rect 22422 10570 22446 10598
rect 22474 10570 22498 10598
rect 22526 10570 22554 10598
rect 22054 9814 22554 10570
rect 22054 9786 22082 9814
rect 22110 9786 22134 9814
rect 22162 9786 22186 9814
rect 22214 9786 22238 9814
rect 22266 9786 22290 9814
rect 22318 9786 22342 9814
rect 22370 9786 22394 9814
rect 22422 9786 22446 9814
rect 22474 9786 22498 9814
rect 22526 9786 22554 9814
rect 22054 9030 22554 9786
rect 22054 9002 22082 9030
rect 22110 9002 22134 9030
rect 22162 9002 22186 9030
rect 22214 9002 22238 9030
rect 22266 9002 22290 9030
rect 22318 9002 22342 9030
rect 22370 9002 22394 9030
rect 22422 9002 22446 9030
rect 22474 9002 22498 9030
rect 22526 9002 22554 9030
rect 22054 8246 22554 9002
rect 22054 8218 22082 8246
rect 22110 8218 22134 8246
rect 22162 8218 22186 8246
rect 22214 8218 22238 8246
rect 22266 8218 22290 8246
rect 22318 8218 22342 8246
rect 22370 8218 22394 8246
rect 22422 8218 22446 8246
rect 22474 8218 22498 8246
rect 22526 8218 22554 8246
rect 22054 7462 22554 8218
rect 22054 7434 22082 7462
rect 22110 7434 22134 7462
rect 22162 7434 22186 7462
rect 22214 7434 22238 7462
rect 22266 7434 22290 7462
rect 22318 7434 22342 7462
rect 22370 7434 22394 7462
rect 22422 7434 22446 7462
rect 22474 7434 22498 7462
rect 22526 7434 22554 7462
rect 22054 6678 22554 7434
rect 22054 6650 22082 6678
rect 22110 6650 22134 6678
rect 22162 6650 22186 6678
rect 22214 6650 22238 6678
rect 22266 6650 22290 6678
rect 22318 6650 22342 6678
rect 22370 6650 22394 6678
rect 22422 6650 22446 6678
rect 22474 6650 22498 6678
rect 22526 6650 22554 6678
rect 22054 5894 22554 6650
rect 22054 5866 22082 5894
rect 22110 5866 22134 5894
rect 22162 5866 22186 5894
rect 22214 5866 22238 5894
rect 22266 5866 22290 5894
rect 22318 5866 22342 5894
rect 22370 5866 22394 5894
rect 22422 5866 22446 5894
rect 22474 5866 22498 5894
rect 22526 5866 22554 5894
rect 22054 5110 22554 5866
rect 22054 5082 22082 5110
rect 22110 5082 22134 5110
rect 22162 5082 22186 5110
rect 22214 5082 22238 5110
rect 22266 5082 22290 5110
rect 22318 5082 22342 5110
rect 22370 5082 22394 5110
rect 22422 5082 22446 5110
rect 22474 5082 22498 5110
rect 22526 5082 22554 5110
rect 22054 4326 22554 5082
rect 22054 4298 22082 4326
rect 22110 4298 22134 4326
rect 22162 4298 22186 4326
rect 22214 4298 22238 4326
rect 22266 4298 22290 4326
rect 22318 4298 22342 4326
rect 22370 4298 22394 4326
rect 22422 4298 22446 4326
rect 22474 4298 22498 4326
rect 22526 4298 22554 4326
rect 22054 3542 22554 4298
rect 22054 3514 22082 3542
rect 22110 3514 22134 3542
rect 22162 3514 22186 3542
rect 22214 3514 22238 3542
rect 22266 3514 22290 3542
rect 22318 3514 22342 3542
rect 22370 3514 22394 3542
rect 22422 3514 22446 3542
rect 22474 3514 22498 3542
rect 22526 3514 22554 3542
rect 22054 2758 22554 3514
rect 22054 2730 22082 2758
rect 22110 2730 22134 2758
rect 22162 2730 22186 2758
rect 22214 2730 22238 2758
rect 22266 2730 22290 2758
rect 22318 2730 22342 2758
rect 22370 2730 22394 2758
rect 22422 2730 22446 2758
rect 22474 2730 22498 2758
rect 22526 2730 22554 2758
rect 22054 1974 22554 2730
rect 22054 1946 22082 1974
rect 22110 1946 22134 1974
rect 22162 1946 22186 1974
rect 22214 1946 22238 1974
rect 22266 1946 22290 1974
rect 22318 1946 22342 1974
rect 22370 1946 22394 1974
rect 22422 1946 22446 1974
rect 22474 1946 22498 1974
rect 22526 1946 22554 1974
rect 22054 1538 22554 1946
rect 24554 18046 25054 18454
rect 24554 18018 24582 18046
rect 24610 18018 24634 18046
rect 24662 18018 24686 18046
rect 24714 18018 24738 18046
rect 24766 18018 24790 18046
rect 24818 18018 24842 18046
rect 24870 18018 24894 18046
rect 24922 18018 24946 18046
rect 24974 18018 24998 18046
rect 25026 18018 25054 18046
rect 24554 17262 25054 18018
rect 24554 17234 24582 17262
rect 24610 17234 24634 17262
rect 24662 17234 24686 17262
rect 24714 17234 24738 17262
rect 24766 17234 24790 17262
rect 24818 17234 24842 17262
rect 24870 17234 24894 17262
rect 24922 17234 24946 17262
rect 24974 17234 24998 17262
rect 25026 17234 25054 17262
rect 24554 16478 25054 17234
rect 24554 16450 24582 16478
rect 24610 16450 24634 16478
rect 24662 16450 24686 16478
rect 24714 16450 24738 16478
rect 24766 16450 24790 16478
rect 24818 16450 24842 16478
rect 24870 16450 24894 16478
rect 24922 16450 24946 16478
rect 24974 16450 24998 16478
rect 25026 16450 25054 16478
rect 24554 15694 25054 16450
rect 24554 15666 24582 15694
rect 24610 15666 24634 15694
rect 24662 15666 24686 15694
rect 24714 15666 24738 15694
rect 24766 15666 24790 15694
rect 24818 15666 24842 15694
rect 24870 15666 24894 15694
rect 24922 15666 24946 15694
rect 24974 15666 24998 15694
rect 25026 15666 25054 15694
rect 24554 14910 25054 15666
rect 24554 14882 24582 14910
rect 24610 14882 24634 14910
rect 24662 14882 24686 14910
rect 24714 14882 24738 14910
rect 24766 14882 24790 14910
rect 24818 14882 24842 14910
rect 24870 14882 24894 14910
rect 24922 14882 24946 14910
rect 24974 14882 24998 14910
rect 25026 14882 25054 14910
rect 24554 14126 25054 14882
rect 24554 14098 24582 14126
rect 24610 14098 24634 14126
rect 24662 14098 24686 14126
rect 24714 14098 24738 14126
rect 24766 14098 24790 14126
rect 24818 14098 24842 14126
rect 24870 14098 24894 14126
rect 24922 14098 24946 14126
rect 24974 14098 24998 14126
rect 25026 14098 25054 14126
rect 24554 13342 25054 14098
rect 24554 13314 24582 13342
rect 24610 13314 24634 13342
rect 24662 13314 24686 13342
rect 24714 13314 24738 13342
rect 24766 13314 24790 13342
rect 24818 13314 24842 13342
rect 24870 13314 24894 13342
rect 24922 13314 24946 13342
rect 24974 13314 24998 13342
rect 25026 13314 25054 13342
rect 24554 12558 25054 13314
rect 24554 12530 24582 12558
rect 24610 12530 24634 12558
rect 24662 12530 24686 12558
rect 24714 12530 24738 12558
rect 24766 12530 24790 12558
rect 24818 12530 24842 12558
rect 24870 12530 24894 12558
rect 24922 12530 24946 12558
rect 24974 12530 24998 12558
rect 25026 12530 25054 12558
rect 24554 11774 25054 12530
rect 24554 11746 24582 11774
rect 24610 11746 24634 11774
rect 24662 11746 24686 11774
rect 24714 11746 24738 11774
rect 24766 11746 24790 11774
rect 24818 11746 24842 11774
rect 24870 11746 24894 11774
rect 24922 11746 24946 11774
rect 24974 11746 24998 11774
rect 25026 11746 25054 11774
rect 24554 10990 25054 11746
rect 24554 10962 24582 10990
rect 24610 10962 24634 10990
rect 24662 10962 24686 10990
rect 24714 10962 24738 10990
rect 24766 10962 24790 10990
rect 24818 10962 24842 10990
rect 24870 10962 24894 10990
rect 24922 10962 24946 10990
rect 24974 10962 24998 10990
rect 25026 10962 25054 10990
rect 24554 10206 25054 10962
rect 24554 10178 24582 10206
rect 24610 10178 24634 10206
rect 24662 10178 24686 10206
rect 24714 10178 24738 10206
rect 24766 10178 24790 10206
rect 24818 10178 24842 10206
rect 24870 10178 24894 10206
rect 24922 10178 24946 10206
rect 24974 10178 24998 10206
rect 25026 10178 25054 10206
rect 24554 9422 25054 10178
rect 24554 9394 24582 9422
rect 24610 9394 24634 9422
rect 24662 9394 24686 9422
rect 24714 9394 24738 9422
rect 24766 9394 24790 9422
rect 24818 9394 24842 9422
rect 24870 9394 24894 9422
rect 24922 9394 24946 9422
rect 24974 9394 24998 9422
rect 25026 9394 25054 9422
rect 24554 8638 25054 9394
rect 24554 8610 24582 8638
rect 24610 8610 24634 8638
rect 24662 8610 24686 8638
rect 24714 8610 24738 8638
rect 24766 8610 24790 8638
rect 24818 8610 24842 8638
rect 24870 8610 24894 8638
rect 24922 8610 24946 8638
rect 24974 8610 24998 8638
rect 25026 8610 25054 8638
rect 24554 7854 25054 8610
rect 24554 7826 24582 7854
rect 24610 7826 24634 7854
rect 24662 7826 24686 7854
rect 24714 7826 24738 7854
rect 24766 7826 24790 7854
rect 24818 7826 24842 7854
rect 24870 7826 24894 7854
rect 24922 7826 24946 7854
rect 24974 7826 24998 7854
rect 25026 7826 25054 7854
rect 24554 7070 25054 7826
rect 24554 7042 24582 7070
rect 24610 7042 24634 7070
rect 24662 7042 24686 7070
rect 24714 7042 24738 7070
rect 24766 7042 24790 7070
rect 24818 7042 24842 7070
rect 24870 7042 24894 7070
rect 24922 7042 24946 7070
rect 24974 7042 24998 7070
rect 25026 7042 25054 7070
rect 24554 6286 25054 7042
rect 24554 6258 24582 6286
rect 24610 6258 24634 6286
rect 24662 6258 24686 6286
rect 24714 6258 24738 6286
rect 24766 6258 24790 6286
rect 24818 6258 24842 6286
rect 24870 6258 24894 6286
rect 24922 6258 24946 6286
rect 24974 6258 24998 6286
rect 25026 6258 25054 6286
rect 24554 5502 25054 6258
rect 24554 5474 24582 5502
rect 24610 5474 24634 5502
rect 24662 5474 24686 5502
rect 24714 5474 24738 5502
rect 24766 5474 24790 5502
rect 24818 5474 24842 5502
rect 24870 5474 24894 5502
rect 24922 5474 24946 5502
rect 24974 5474 24998 5502
rect 25026 5474 25054 5502
rect 24554 4718 25054 5474
rect 24554 4690 24582 4718
rect 24610 4690 24634 4718
rect 24662 4690 24686 4718
rect 24714 4690 24738 4718
rect 24766 4690 24790 4718
rect 24818 4690 24842 4718
rect 24870 4690 24894 4718
rect 24922 4690 24946 4718
rect 24974 4690 24998 4718
rect 25026 4690 25054 4718
rect 24554 3934 25054 4690
rect 24554 3906 24582 3934
rect 24610 3906 24634 3934
rect 24662 3906 24686 3934
rect 24714 3906 24738 3934
rect 24766 3906 24790 3934
rect 24818 3906 24842 3934
rect 24870 3906 24894 3934
rect 24922 3906 24946 3934
rect 24974 3906 24998 3934
rect 25026 3906 25054 3934
rect 24554 3150 25054 3906
rect 24554 3122 24582 3150
rect 24610 3122 24634 3150
rect 24662 3122 24686 3150
rect 24714 3122 24738 3150
rect 24766 3122 24790 3150
rect 24818 3122 24842 3150
rect 24870 3122 24894 3150
rect 24922 3122 24946 3150
rect 24974 3122 24998 3150
rect 25026 3122 25054 3150
rect 24554 2366 25054 3122
rect 24554 2338 24582 2366
rect 24610 2338 24634 2366
rect 24662 2338 24686 2366
rect 24714 2338 24738 2366
rect 24766 2338 24790 2366
rect 24818 2338 24842 2366
rect 24870 2338 24894 2366
rect 24922 2338 24946 2366
rect 24974 2338 24998 2366
rect 25026 2338 25054 2366
rect 24554 1582 25054 2338
rect 24554 1554 24582 1582
rect 24610 1554 24634 1582
rect 24662 1554 24686 1582
rect 24714 1554 24738 1582
rect 24766 1554 24790 1582
rect 24818 1554 24842 1582
rect 24870 1554 24894 1582
rect 24922 1554 24946 1582
rect 24974 1554 24998 1582
rect 25026 1554 25054 1582
rect 24554 1538 25054 1554
rect 27054 18438 27554 18454
rect 27054 18410 27082 18438
rect 27110 18410 27134 18438
rect 27162 18410 27186 18438
rect 27214 18410 27238 18438
rect 27266 18410 27290 18438
rect 27318 18410 27342 18438
rect 27370 18410 27394 18438
rect 27422 18410 27446 18438
rect 27474 18410 27498 18438
rect 27526 18410 27554 18438
rect 27054 17654 27554 18410
rect 27054 17626 27082 17654
rect 27110 17626 27134 17654
rect 27162 17626 27186 17654
rect 27214 17626 27238 17654
rect 27266 17626 27290 17654
rect 27318 17626 27342 17654
rect 27370 17626 27394 17654
rect 27422 17626 27446 17654
rect 27474 17626 27498 17654
rect 27526 17626 27554 17654
rect 27054 16870 27554 17626
rect 27054 16842 27082 16870
rect 27110 16842 27134 16870
rect 27162 16842 27186 16870
rect 27214 16842 27238 16870
rect 27266 16842 27290 16870
rect 27318 16842 27342 16870
rect 27370 16842 27394 16870
rect 27422 16842 27446 16870
rect 27474 16842 27498 16870
rect 27526 16842 27554 16870
rect 27054 16086 27554 16842
rect 27054 16058 27082 16086
rect 27110 16058 27134 16086
rect 27162 16058 27186 16086
rect 27214 16058 27238 16086
rect 27266 16058 27290 16086
rect 27318 16058 27342 16086
rect 27370 16058 27394 16086
rect 27422 16058 27446 16086
rect 27474 16058 27498 16086
rect 27526 16058 27554 16086
rect 27054 15302 27554 16058
rect 27054 15274 27082 15302
rect 27110 15274 27134 15302
rect 27162 15274 27186 15302
rect 27214 15274 27238 15302
rect 27266 15274 27290 15302
rect 27318 15274 27342 15302
rect 27370 15274 27394 15302
rect 27422 15274 27446 15302
rect 27474 15274 27498 15302
rect 27526 15274 27554 15302
rect 27054 14518 27554 15274
rect 27054 14490 27082 14518
rect 27110 14490 27134 14518
rect 27162 14490 27186 14518
rect 27214 14490 27238 14518
rect 27266 14490 27290 14518
rect 27318 14490 27342 14518
rect 27370 14490 27394 14518
rect 27422 14490 27446 14518
rect 27474 14490 27498 14518
rect 27526 14490 27554 14518
rect 27054 13734 27554 14490
rect 27054 13706 27082 13734
rect 27110 13706 27134 13734
rect 27162 13706 27186 13734
rect 27214 13706 27238 13734
rect 27266 13706 27290 13734
rect 27318 13706 27342 13734
rect 27370 13706 27394 13734
rect 27422 13706 27446 13734
rect 27474 13706 27498 13734
rect 27526 13706 27554 13734
rect 27054 12950 27554 13706
rect 27054 12922 27082 12950
rect 27110 12922 27134 12950
rect 27162 12922 27186 12950
rect 27214 12922 27238 12950
rect 27266 12922 27290 12950
rect 27318 12922 27342 12950
rect 27370 12922 27394 12950
rect 27422 12922 27446 12950
rect 27474 12922 27498 12950
rect 27526 12922 27554 12950
rect 27054 12166 27554 12922
rect 27054 12138 27082 12166
rect 27110 12138 27134 12166
rect 27162 12138 27186 12166
rect 27214 12138 27238 12166
rect 27266 12138 27290 12166
rect 27318 12138 27342 12166
rect 27370 12138 27394 12166
rect 27422 12138 27446 12166
rect 27474 12138 27498 12166
rect 27526 12138 27554 12166
rect 27054 11382 27554 12138
rect 27054 11354 27082 11382
rect 27110 11354 27134 11382
rect 27162 11354 27186 11382
rect 27214 11354 27238 11382
rect 27266 11354 27290 11382
rect 27318 11354 27342 11382
rect 27370 11354 27394 11382
rect 27422 11354 27446 11382
rect 27474 11354 27498 11382
rect 27526 11354 27554 11382
rect 27054 10598 27554 11354
rect 27054 10570 27082 10598
rect 27110 10570 27134 10598
rect 27162 10570 27186 10598
rect 27214 10570 27238 10598
rect 27266 10570 27290 10598
rect 27318 10570 27342 10598
rect 27370 10570 27394 10598
rect 27422 10570 27446 10598
rect 27474 10570 27498 10598
rect 27526 10570 27554 10598
rect 27054 9814 27554 10570
rect 27054 9786 27082 9814
rect 27110 9786 27134 9814
rect 27162 9786 27186 9814
rect 27214 9786 27238 9814
rect 27266 9786 27290 9814
rect 27318 9786 27342 9814
rect 27370 9786 27394 9814
rect 27422 9786 27446 9814
rect 27474 9786 27498 9814
rect 27526 9786 27554 9814
rect 27054 9030 27554 9786
rect 27054 9002 27082 9030
rect 27110 9002 27134 9030
rect 27162 9002 27186 9030
rect 27214 9002 27238 9030
rect 27266 9002 27290 9030
rect 27318 9002 27342 9030
rect 27370 9002 27394 9030
rect 27422 9002 27446 9030
rect 27474 9002 27498 9030
rect 27526 9002 27554 9030
rect 27054 8246 27554 9002
rect 27054 8218 27082 8246
rect 27110 8218 27134 8246
rect 27162 8218 27186 8246
rect 27214 8218 27238 8246
rect 27266 8218 27290 8246
rect 27318 8218 27342 8246
rect 27370 8218 27394 8246
rect 27422 8218 27446 8246
rect 27474 8218 27498 8246
rect 27526 8218 27554 8246
rect 27054 7462 27554 8218
rect 27054 7434 27082 7462
rect 27110 7434 27134 7462
rect 27162 7434 27186 7462
rect 27214 7434 27238 7462
rect 27266 7434 27290 7462
rect 27318 7434 27342 7462
rect 27370 7434 27394 7462
rect 27422 7434 27446 7462
rect 27474 7434 27498 7462
rect 27526 7434 27554 7462
rect 27054 6678 27554 7434
rect 27054 6650 27082 6678
rect 27110 6650 27134 6678
rect 27162 6650 27186 6678
rect 27214 6650 27238 6678
rect 27266 6650 27290 6678
rect 27318 6650 27342 6678
rect 27370 6650 27394 6678
rect 27422 6650 27446 6678
rect 27474 6650 27498 6678
rect 27526 6650 27554 6678
rect 27054 5894 27554 6650
rect 27054 5866 27082 5894
rect 27110 5866 27134 5894
rect 27162 5866 27186 5894
rect 27214 5866 27238 5894
rect 27266 5866 27290 5894
rect 27318 5866 27342 5894
rect 27370 5866 27394 5894
rect 27422 5866 27446 5894
rect 27474 5866 27498 5894
rect 27526 5866 27554 5894
rect 27054 5110 27554 5866
rect 27054 5082 27082 5110
rect 27110 5082 27134 5110
rect 27162 5082 27186 5110
rect 27214 5082 27238 5110
rect 27266 5082 27290 5110
rect 27318 5082 27342 5110
rect 27370 5082 27394 5110
rect 27422 5082 27446 5110
rect 27474 5082 27498 5110
rect 27526 5082 27554 5110
rect 27054 4326 27554 5082
rect 27054 4298 27082 4326
rect 27110 4298 27134 4326
rect 27162 4298 27186 4326
rect 27214 4298 27238 4326
rect 27266 4298 27290 4326
rect 27318 4298 27342 4326
rect 27370 4298 27394 4326
rect 27422 4298 27446 4326
rect 27474 4298 27498 4326
rect 27526 4298 27554 4326
rect 27054 3542 27554 4298
rect 27054 3514 27082 3542
rect 27110 3514 27134 3542
rect 27162 3514 27186 3542
rect 27214 3514 27238 3542
rect 27266 3514 27290 3542
rect 27318 3514 27342 3542
rect 27370 3514 27394 3542
rect 27422 3514 27446 3542
rect 27474 3514 27498 3542
rect 27526 3514 27554 3542
rect 27054 2758 27554 3514
rect 27054 2730 27082 2758
rect 27110 2730 27134 2758
rect 27162 2730 27186 2758
rect 27214 2730 27238 2758
rect 27266 2730 27290 2758
rect 27318 2730 27342 2758
rect 27370 2730 27394 2758
rect 27422 2730 27446 2758
rect 27474 2730 27498 2758
rect 27526 2730 27554 2758
rect 27054 1974 27554 2730
rect 27054 1946 27082 1974
rect 27110 1946 27134 1974
rect 27162 1946 27186 1974
rect 27214 1946 27238 1974
rect 27266 1946 27290 1974
rect 27318 1946 27342 1974
rect 27370 1946 27394 1974
rect 27422 1946 27446 1974
rect 27474 1946 27498 1974
rect 27526 1946 27554 1974
rect 27054 1538 27554 1946
rect 29554 18046 30054 18454
rect 29554 18018 29582 18046
rect 29610 18018 29634 18046
rect 29662 18018 29686 18046
rect 29714 18018 29738 18046
rect 29766 18018 29790 18046
rect 29818 18018 29842 18046
rect 29870 18018 29894 18046
rect 29922 18018 29946 18046
rect 29974 18018 29998 18046
rect 30026 18018 30054 18046
rect 29554 17262 30054 18018
rect 29554 17234 29582 17262
rect 29610 17234 29634 17262
rect 29662 17234 29686 17262
rect 29714 17234 29738 17262
rect 29766 17234 29790 17262
rect 29818 17234 29842 17262
rect 29870 17234 29894 17262
rect 29922 17234 29946 17262
rect 29974 17234 29998 17262
rect 30026 17234 30054 17262
rect 29554 16478 30054 17234
rect 29554 16450 29582 16478
rect 29610 16450 29634 16478
rect 29662 16450 29686 16478
rect 29714 16450 29738 16478
rect 29766 16450 29790 16478
rect 29818 16450 29842 16478
rect 29870 16450 29894 16478
rect 29922 16450 29946 16478
rect 29974 16450 29998 16478
rect 30026 16450 30054 16478
rect 29554 15694 30054 16450
rect 29554 15666 29582 15694
rect 29610 15666 29634 15694
rect 29662 15666 29686 15694
rect 29714 15666 29738 15694
rect 29766 15666 29790 15694
rect 29818 15666 29842 15694
rect 29870 15666 29894 15694
rect 29922 15666 29946 15694
rect 29974 15666 29998 15694
rect 30026 15666 30054 15694
rect 29554 14910 30054 15666
rect 29554 14882 29582 14910
rect 29610 14882 29634 14910
rect 29662 14882 29686 14910
rect 29714 14882 29738 14910
rect 29766 14882 29790 14910
rect 29818 14882 29842 14910
rect 29870 14882 29894 14910
rect 29922 14882 29946 14910
rect 29974 14882 29998 14910
rect 30026 14882 30054 14910
rect 29554 14126 30054 14882
rect 29554 14098 29582 14126
rect 29610 14098 29634 14126
rect 29662 14098 29686 14126
rect 29714 14098 29738 14126
rect 29766 14098 29790 14126
rect 29818 14098 29842 14126
rect 29870 14098 29894 14126
rect 29922 14098 29946 14126
rect 29974 14098 29998 14126
rect 30026 14098 30054 14126
rect 29554 13342 30054 14098
rect 29554 13314 29582 13342
rect 29610 13314 29634 13342
rect 29662 13314 29686 13342
rect 29714 13314 29738 13342
rect 29766 13314 29790 13342
rect 29818 13314 29842 13342
rect 29870 13314 29894 13342
rect 29922 13314 29946 13342
rect 29974 13314 29998 13342
rect 30026 13314 30054 13342
rect 29554 12558 30054 13314
rect 29554 12530 29582 12558
rect 29610 12530 29634 12558
rect 29662 12530 29686 12558
rect 29714 12530 29738 12558
rect 29766 12530 29790 12558
rect 29818 12530 29842 12558
rect 29870 12530 29894 12558
rect 29922 12530 29946 12558
rect 29974 12530 29998 12558
rect 30026 12530 30054 12558
rect 29554 11774 30054 12530
rect 29554 11746 29582 11774
rect 29610 11746 29634 11774
rect 29662 11746 29686 11774
rect 29714 11746 29738 11774
rect 29766 11746 29790 11774
rect 29818 11746 29842 11774
rect 29870 11746 29894 11774
rect 29922 11746 29946 11774
rect 29974 11746 29998 11774
rect 30026 11746 30054 11774
rect 29554 10990 30054 11746
rect 29554 10962 29582 10990
rect 29610 10962 29634 10990
rect 29662 10962 29686 10990
rect 29714 10962 29738 10990
rect 29766 10962 29790 10990
rect 29818 10962 29842 10990
rect 29870 10962 29894 10990
rect 29922 10962 29946 10990
rect 29974 10962 29998 10990
rect 30026 10962 30054 10990
rect 29554 10206 30054 10962
rect 29554 10178 29582 10206
rect 29610 10178 29634 10206
rect 29662 10178 29686 10206
rect 29714 10178 29738 10206
rect 29766 10178 29790 10206
rect 29818 10178 29842 10206
rect 29870 10178 29894 10206
rect 29922 10178 29946 10206
rect 29974 10178 29998 10206
rect 30026 10178 30054 10206
rect 29554 9422 30054 10178
rect 29554 9394 29582 9422
rect 29610 9394 29634 9422
rect 29662 9394 29686 9422
rect 29714 9394 29738 9422
rect 29766 9394 29790 9422
rect 29818 9394 29842 9422
rect 29870 9394 29894 9422
rect 29922 9394 29946 9422
rect 29974 9394 29998 9422
rect 30026 9394 30054 9422
rect 29554 8638 30054 9394
rect 29554 8610 29582 8638
rect 29610 8610 29634 8638
rect 29662 8610 29686 8638
rect 29714 8610 29738 8638
rect 29766 8610 29790 8638
rect 29818 8610 29842 8638
rect 29870 8610 29894 8638
rect 29922 8610 29946 8638
rect 29974 8610 29998 8638
rect 30026 8610 30054 8638
rect 29554 7854 30054 8610
rect 32054 18438 32554 18454
rect 32054 18410 32082 18438
rect 32110 18410 32134 18438
rect 32162 18410 32186 18438
rect 32214 18410 32238 18438
rect 32266 18410 32290 18438
rect 32318 18410 32342 18438
rect 32370 18410 32394 18438
rect 32422 18410 32446 18438
rect 32474 18410 32498 18438
rect 32526 18410 32554 18438
rect 32054 17654 32554 18410
rect 32054 17626 32082 17654
rect 32110 17626 32134 17654
rect 32162 17626 32186 17654
rect 32214 17626 32238 17654
rect 32266 17626 32290 17654
rect 32318 17626 32342 17654
rect 32370 17626 32394 17654
rect 32422 17626 32446 17654
rect 32474 17626 32498 17654
rect 32526 17626 32554 17654
rect 32054 16870 32554 17626
rect 32054 16842 32082 16870
rect 32110 16842 32134 16870
rect 32162 16842 32186 16870
rect 32214 16842 32238 16870
rect 32266 16842 32290 16870
rect 32318 16842 32342 16870
rect 32370 16842 32394 16870
rect 32422 16842 32446 16870
rect 32474 16842 32498 16870
rect 32526 16842 32554 16870
rect 32054 16086 32554 16842
rect 32054 16058 32082 16086
rect 32110 16058 32134 16086
rect 32162 16058 32186 16086
rect 32214 16058 32238 16086
rect 32266 16058 32290 16086
rect 32318 16058 32342 16086
rect 32370 16058 32394 16086
rect 32422 16058 32446 16086
rect 32474 16058 32498 16086
rect 32526 16058 32554 16086
rect 32054 15302 32554 16058
rect 32054 15274 32082 15302
rect 32110 15274 32134 15302
rect 32162 15274 32186 15302
rect 32214 15274 32238 15302
rect 32266 15274 32290 15302
rect 32318 15274 32342 15302
rect 32370 15274 32394 15302
rect 32422 15274 32446 15302
rect 32474 15274 32498 15302
rect 32526 15274 32554 15302
rect 32054 14518 32554 15274
rect 32054 14490 32082 14518
rect 32110 14490 32134 14518
rect 32162 14490 32186 14518
rect 32214 14490 32238 14518
rect 32266 14490 32290 14518
rect 32318 14490 32342 14518
rect 32370 14490 32394 14518
rect 32422 14490 32446 14518
rect 32474 14490 32498 14518
rect 32526 14490 32554 14518
rect 32054 13734 32554 14490
rect 32054 13706 32082 13734
rect 32110 13706 32134 13734
rect 32162 13706 32186 13734
rect 32214 13706 32238 13734
rect 32266 13706 32290 13734
rect 32318 13706 32342 13734
rect 32370 13706 32394 13734
rect 32422 13706 32446 13734
rect 32474 13706 32498 13734
rect 32526 13706 32554 13734
rect 32054 12950 32554 13706
rect 32054 12922 32082 12950
rect 32110 12922 32134 12950
rect 32162 12922 32186 12950
rect 32214 12922 32238 12950
rect 32266 12922 32290 12950
rect 32318 12922 32342 12950
rect 32370 12922 32394 12950
rect 32422 12922 32446 12950
rect 32474 12922 32498 12950
rect 32526 12922 32554 12950
rect 32054 12166 32554 12922
rect 32054 12138 32082 12166
rect 32110 12138 32134 12166
rect 32162 12138 32186 12166
rect 32214 12138 32238 12166
rect 32266 12138 32290 12166
rect 32318 12138 32342 12166
rect 32370 12138 32394 12166
rect 32422 12138 32446 12166
rect 32474 12138 32498 12166
rect 32526 12138 32554 12166
rect 32054 11382 32554 12138
rect 32054 11354 32082 11382
rect 32110 11354 32134 11382
rect 32162 11354 32186 11382
rect 32214 11354 32238 11382
rect 32266 11354 32290 11382
rect 32318 11354 32342 11382
rect 32370 11354 32394 11382
rect 32422 11354 32446 11382
rect 32474 11354 32498 11382
rect 32526 11354 32554 11382
rect 32054 10598 32554 11354
rect 32054 10570 32082 10598
rect 32110 10570 32134 10598
rect 32162 10570 32186 10598
rect 32214 10570 32238 10598
rect 32266 10570 32290 10598
rect 32318 10570 32342 10598
rect 32370 10570 32394 10598
rect 32422 10570 32446 10598
rect 32474 10570 32498 10598
rect 32526 10570 32554 10598
rect 32054 9814 32554 10570
rect 32054 9786 32082 9814
rect 32110 9786 32134 9814
rect 32162 9786 32186 9814
rect 32214 9786 32238 9814
rect 32266 9786 32290 9814
rect 32318 9786 32342 9814
rect 32370 9786 32394 9814
rect 32422 9786 32446 9814
rect 32474 9786 32498 9814
rect 32526 9786 32554 9814
rect 32054 9030 32554 9786
rect 32054 9002 32082 9030
rect 32110 9002 32134 9030
rect 32162 9002 32186 9030
rect 32214 9002 32238 9030
rect 32266 9002 32290 9030
rect 32318 9002 32342 9030
rect 32370 9002 32394 9030
rect 32422 9002 32446 9030
rect 32474 9002 32498 9030
rect 32526 9002 32554 9030
rect 29554 7826 29582 7854
rect 29610 7826 29634 7854
rect 29662 7826 29686 7854
rect 29714 7826 29738 7854
rect 29766 7826 29790 7854
rect 29818 7826 29842 7854
rect 29870 7826 29894 7854
rect 29922 7826 29946 7854
rect 29974 7826 29998 7854
rect 30026 7826 30054 7854
rect 29554 7070 30054 7826
rect 29554 7042 29582 7070
rect 29610 7042 29634 7070
rect 29662 7042 29686 7070
rect 29714 7042 29738 7070
rect 29766 7042 29790 7070
rect 29818 7042 29842 7070
rect 29870 7042 29894 7070
rect 29922 7042 29946 7070
rect 29974 7042 29998 7070
rect 30026 7042 30054 7070
rect 29554 6286 30054 7042
rect 29554 6258 29582 6286
rect 29610 6258 29634 6286
rect 29662 6258 29686 6286
rect 29714 6258 29738 6286
rect 29766 6258 29790 6286
rect 29818 6258 29842 6286
rect 29870 6258 29894 6286
rect 29922 6258 29946 6286
rect 29974 6258 29998 6286
rect 30026 6258 30054 6286
rect 29554 5502 30054 6258
rect 31934 8554 31962 8559
rect 31934 6090 31962 8526
rect 32054 8246 32554 9002
rect 32054 8218 32082 8246
rect 32110 8218 32134 8246
rect 32162 8218 32186 8246
rect 32214 8218 32238 8246
rect 32266 8218 32290 8246
rect 32318 8218 32342 8246
rect 32370 8218 32394 8246
rect 32422 8218 32446 8246
rect 32474 8218 32498 8246
rect 32526 8218 32554 8246
rect 31990 7658 32018 7663
rect 31990 6762 32018 7630
rect 31990 6729 32018 6734
rect 32054 7462 32554 8218
rect 32054 7434 32082 7462
rect 32110 7434 32134 7462
rect 32162 7434 32186 7462
rect 32214 7434 32238 7462
rect 32266 7434 32290 7462
rect 32318 7434 32342 7462
rect 32370 7434 32394 7462
rect 32422 7434 32446 7462
rect 32474 7434 32498 7462
rect 32526 7434 32554 7462
rect 32054 6678 32554 7434
rect 32054 6650 32082 6678
rect 32110 6650 32134 6678
rect 32162 6650 32186 6678
rect 32214 6650 32238 6678
rect 32266 6650 32290 6678
rect 32318 6650 32342 6678
rect 32370 6650 32394 6678
rect 32422 6650 32446 6678
rect 32474 6650 32498 6678
rect 32526 6650 32554 6678
rect 31990 6090 32018 6095
rect 31934 6062 31990 6090
rect 29554 5474 29582 5502
rect 29610 5474 29634 5502
rect 29662 5474 29686 5502
rect 29714 5474 29738 5502
rect 29766 5474 29790 5502
rect 29818 5474 29842 5502
rect 29870 5474 29894 5502
rect 29922 5474 29946 5502
rect 29974 5474 29998 5502
rect 30026 5474 30054 5502
rect 29554 4718 30054 5474
rect 31990 5642 32018 6062
rect 31990 5306 32018 5614
rect 31990 5273 32018 5278
rect 32054 5894 32554 6650
rect 32054 5866 32082 5894
rect 32110 5866 32134 5894
rect 32162 5866 32186 5894
rect 32214 5866 32238 5894
rect 32266 5866 32290 5894
rect 32318 5866 32342 5894
rect 32370 5866 32394 5894
rect 32422 5866 32446 5894
rect 32474 5866 32498 5894
rect 32526 5866 32554 5894
rect 32054 5110 32554 5866
rect 32054 5082 32082 5110
rect 32110 5082 32134 5110
rect 32162 5082 32186 5110
rect 32214 5082 32238 5110
rect 32266 5082 32290 5110
rect 32318 5082 32342 5110
rect 32370 5082 32394 5110
rect 32422 5082 32446 5110
rect 32474 5082 32498 5110
rect 32526 5082 32554 5110
rect 29554 4690 29582 4718
rect 29610 4690 29634 4718
rect 29662 4690 29686 4718
rect 29714 4690 29738 4718
rect 29766 4690 29790 4718
rect 29818 4690 29842 4718
rect 29870 4690 29894 4718
rect 29922 4690 29946 4718
rect 29974 4690 29998 4718
rect 30026 4690 30054 4718
rect 29554 3934 30054 4690
rect 29554 3906 29582 3934
rect 29610 3906 29634 3934
rect 29662 3906 29686 3934
rect 29714 3906 29738 3934
rect 29766 3906 29790 3934
rect 29818 3906 29842 3934
rect 29870 3906 29894 3934
rect 29922 3906 29946 3934
rect 29974 3906 29998 3934
rect 30026 3906 30054 3934
rect 29554 3150 30054 3906
rect 31990 4914 32018 4919
rect 31990 4074 32018 4886
rect 31990 3346 32018 4046
rect 31990 3313 32018 3318
rect 32054 4326 32554 5082
rect 32054 4298 32082 4326
rect 32110 4298 32134 4326
rect 32162 4298 32186 4326
rect 32214 4298 32238 4326
rect 32266 4298 32290 4326
rect 32318 4298 32342 4326
rect 32370 4298 32394 4326
rect 32422 4298 32446 4326
rect 32474 4298 32498 4326
rect 32526 4298 32554 4326
rect 32054 3542 32554 4298
rect 32054 3514 32082 3542
rect 32110 3514 32134 3542
rect 32162 3514 32186 3542
rect 32214 3514 32238 3542
rect 32266 3514 32290 3542
rect 32318 3514 32342 3542
rect 32370 3514 32394 3542
rect 32422 3514 32446 3542
rect 32474 3514 32498 3542
rect 32526 3514 32554 3542
rect 29554 3122 29582 3150
rect 29610 3122 29634 3150
rect 29662 3122 29686 3150
rect 29714 3122 29738 3150
rect 29766 3122 29790 3150
rect 29818 3122 29842 3150
rect 29870 3122 29894 3150
rect 29922 3122 29946 3150
rect 29974 3122 29998 3150
rect 30026 3122 30054 3150
rect 29554 2366 30054 3122
rect 29554 2338 29582 2366
rect 29610 2338 29634 2366
rect 29662 2338 29686 2366
rect 29714 2338 29738 2366
rect 29766 2338 29790 2366
rect 29818 2338 29842 2366
rect 29870 2338 29894 2366
rect 29922 2338 29946 2366
rect 29974 2338 29998 2366
rect 30026 2338 30054 2366
rect 29554 1582 30054 2338
rect 29554 1554 29582 1582
rect 29610 1554 29634 1582
rect 29662 1554 29686 1582
rect 29714 1554 29738 1582
rect 29766 1554 29790 1582
rect 29818 1554 29842 1582
rect 29870 1554 29894 1582
rect 29922 1554 29946 1582
rect 29974 1554 29998 1582
rect 30026 1554 30054 1582
rect 29554 1538 30054 1554
rect 32054 2758 32554 3514
rect 32054 2730 32082 2758
rect 32110 2730 32134 2758
rect 32162 2730 32186 2758
rect 32214 2730 32238 2758
rect 32266 2730 32290 2758
rect 32318 2730 32342 2758
rect 32370 2730 32394 2758
rect 32422 2730 32446 2758
rect 32474 2730 32498 2758
rect 32526 2730 32554 2758
rect 32054 1974 32554 2730
rect 32054 1946 32082 1974
rect 32110 1946 32134 1974
rect 32162 1946 32186 1974
rect 32214 1946 32238 1974
rect 32266 1946 32290 1974
rect 32318 1946 32342 1974
rect 32370 1946 32394 1974
rect 32422 1946 32446 1974
rect 32474 1946 32498 1974
rect 32526 1946 32554 1974
rect 32054 1538 32554 1946
rect 34554 18046 35054 18454
rect 34554 18018 34582 18046
rect 34610 18018 34634 18046
rect 34662 18018 34686 18046
rect 34714 18018 34738 18046
rect 34766 18018 34790 18046
rect 34818 18018 34842 18046
rect 34870 18018 34894 18046
rect 34922 18018 34946 18046
rect 34974 18018 34998 18046
rect 35026 18018 35054 18046
rect 34554 17262 35054 18018
rect 34554 17234 34582 17262
rect 34610 17234 34634 17262
rect 34662 17234 34686 17262
rect 34714 17234 34738 17262
rect 34766 17234 34790 17262
rect 34818 17234 34842 17262
rect 34870 17234 34894 17262
rect 34922 17234 34946 17262
rect 34974 17234 34998 17262
rect 35026 17234 35054 17262
rect 34554 16478 35054 17234
rect 34554 16450 34582 16478
rect 34610 16450 34634 16478
rect 34662 16450 34686 16478
rect 34714 16450 34738 16478
rect 34766 16450 34790 16478
rect 34818 16450 34842 16478
rect 34870 16450 34894 16478
rect 34922 16450 34946 16478
rect 34974 16450 34998 16478
rect 35026 16450 35054 16478
rect 34554 15694 35054 16450
rect 34554 15666 34582 15694
rect 34610 15666 34634 15694
rect 34662 15666 34686 15694
rect 34714 15666 34738 15694
rect 34766 15666 34790 15694
rect 34818 15666 34842 15694
rect 34870 15666 34894 15694
rect 34922 15666 34946 15694
rect 34974 15666 34998 15694
rect 35026 15666 35054 15694
rect 34554 14910 35054 15666
rect 34554 14882 34582 14910
rect 34610 14882 34634 14910
rect 34662 14882 34686 14910
rect 34714 14882 34738 14910
rect 34766 14882 34790 14910
rect 34818 14882 34842 14910
rect 34870 14882 34894 14910
rect 34922 14882 34946 14910
rect 34974 14882 34998 14910
rect 35026 14882 35054 14910
rect 34554 14126 35054 14882
rect 34554 14098 34582 14126
rect 34610 14098 34634 14126
rect 34662 14098 34686 14126
rect 34714 14098 34738 14126
rect 34766 14098 34790 14126
rect 34818 14098 34842 14126
rect 34870 14098 34894 14126
rect 34922 14098 34946 14126
rect 34974 14098 34998 14126
rect 35026 14098 35054 14126
rect 34554 13342 35054 14098
rect 34554 13314 34582 13342
rect 34610 13314 34634 13342
rect 34662 13314 34686 13342
rect 34714 13314 34738 13342
rect 34766 13314 34790 13342
rect 34818 13314 34842 13342
rect 34870 13314 34894 13342
rect 34922 13314 34946 13342
rect 34974 13314 34998 13342
rect 35026 13314 35054 13342
rect 34554 12558 35054 13314
rect 34554 12530 34582 12558
rect 34610 12530 34634 12558
rect 34662 12530 34686 12558
rect 34714 12530 34738 12558
rect 34766 12530 34790 12558
rect 34818 12530 34842 12558
rect 34870 12530 34894 12558
rect 34922 12530 34946 12558
rect 34974 12530 34998 12558
rect 35026 12530 35054 12558
rect 34554 11774 35054 12530
rect 34554 11746 34582 11774
rect 34610 11746 34634 11774
rect 34662 11746 34686 11774
rect 34714 11746 34738 11774
rect 34766 11746 34790 11774
rect 34818 11746 34842 11774
rect 34870 11746 34894 11774
rect 34922 11746 34946 11774
rect 34974 11746 34998 11774
rect 35026 11746 35054 11774
rect 34554 10990 35054 11746
rect 34554 10962 34582 10990
rect 34610 10962 34634 10990
rect 34662 10962 34686 10990
rect 34714 10962 34738 10990
rect 34766 10962 34790 10990
rect 34818 10962 34842 10990
rect 34870 10962 34894 10990
rect 34922 10962 34946 10990
rect 34974 10962 34998 10990
rect 35026 10962 35054 10990
rect 34554 10206 35054 10962
rect 34554 10178 34582 10206
rect 34610 10178 34634 10206
rect 34662 10178 34686 10206
rect 34714 10178 34738 10206
rect 34766 10178 34790 10206
rect 34818 10178 34842 10206
rect 34870 10178 34894 10206
rect 34922 10178 34946 10206
rect 34974 10178 34998 10206
rect 35026 10178 35054 10206
rect 34554 9422 35054 10178
rect 34554 9394 34582 9422
rect 34610 9394 34634 9422
rect 34662 9394 34686 9422
rect 34714 9394 34738 9422
rect 34766 9394 34790 9422
rect 34818 9394 34842 9422
rect 34870 9394 34894 9422
rect 34922 9394 34946 9422
rect 34974 9394 34998 9422
rect 35026 9394 35054 9422
rect 34554 8638 35054 9394
rect 34554 8610 34582 8638
rect 34610 8610 34634 8638
rect 34662 8610 34686 8638
rect 34714 8610 34738 8638
rect 34766 8610 34790 8638
rect 34818 8610 34842 8638
rect 34870 8610 34894 8638
rect 34922 8610 34946 8638
rect 34974 8610 34998 8638
rect 35026 8610 35054 8638
rect 34554 7854 35054 8610
rect 34554 7826 34582 7854
rect 34610 7826 34634 7854
rect 34662 7826 34686 7854
rect 34714 7826 34738 7854
rect 34766 7826 34790 7854
rect 34818 7826 34842 7854
rect 34870 7826 34894 7854
rect 34922 7826 34946 7854
rect 34974 7826 34998 7854
rect 35026 7826 35054 7854
rect 34554 7070 35054 7826
rect 34554 7042 34582 7070
rect 34610 7042 34634 7070
rect 34662 7042 34686 7070
rect 34714 7042 34738 7070
rect 34766 7042 34790 7070
rect 34818 7042 34842 7070
rect 34870 7042 34894 7070
rect 34922 7042 34946 7070
rect 34974 7042 34998 7070
rect 35026 7042 35054 7070
rect 34554 6286 35054 7042
rect 34554 6258 34582 6286
rect 34610 6258 34634 6286
rect 34662 6258 34686 6286
rect 34714 6258 34738 6286
rect 34766 6258 34790 6286
rect 34818 6258 34842 6286
rect 34870 6258 34894 6286
rect 34922 6258 34946 6286
rect 34974 6258 34998 6286
rect 35026 6258 35054 6286
rect 34554 5502 35054 6258
rect 34554 5474 34582 5502
rect 34610 5474 34634 5502
rect 34662 5474 34686 5502
rect 34714 5474 34738 5502
rect 34766 5474 34790 5502
rect 34818 5474 34842 5502
rect 34870 5474 34894 5502
rect 34922 5474 34946 5502
rect 34974 5474 34998 5502
rect 35026 5474 35054 5502
rect 34554 4718 35054 5474
rect 34554 4690 34582 4718
rect 34610 4690 34634 4718
rect 34662 4690 34686 4718
rect 34714 4690 34738 4718
rect 34766 4690 34790 4718
rect 34818 4690 34842 4718
rect 34870 4690 34894 4718
rect 34922 4690 34946 4718
rect 34974 4690 34998 4718
rect 35026 4690 35054 4718
rect 34554 3934 35054 4690
rect 34554 3906 34582 3934
rect 34610 3906 34634 3934
rect 34662 3906 34686 3934
rect 34714 3906 34738 3934
rect 34766 3906 34790 3934
rect 34818 3906 34842 3934
rect 34870 3906 34894 3934
rect 34922 3906 34946 3934
rect 34974 3906 34998 3934
rect 35026 3906 35054 3934
rect 34554 3150 35054 3906
rect 34554 3122 34582 3150
rect 34610 3122 34634 3150
rect 34662 3122 34686 3150
rect 34714 3122 34738 3150
rect 34766 3122 34790 3150
rect 34818 3122 34842 3150
rect 34870 3122 34894 3150
rect 34922 3122 34946 3150
rect 34974 3122 34998 3150
rect 35026 3122 35054 3150
rect 34554 2366 35054 3122
rect 34554 2338 34582 2366
rect 34610 2338 34634 2366
rect 34662 2338 34686 2366
rect 34714 2338 34738 2366
rect 34766 2338 34790 2366
rect 34818 2338 34842 2366
rect 34870 2338 34894 2366
rect 34922 2338 34946 2366
rect 34974 2338 34998 2366
rect 35026 2338 35054 2366
rect 34554 1582 35054 2338
rect 34554 1554 34582 1582
rect 34610 1554 34634 1582
rect 34662 1554 34686 1582
rect 34714 1554 34738 1582
rect 34766 1554 34790 1582
rect 34818 1554 34842 1582
rect 34870 1554 34894 1582
rect 34922 1554 34946 1582
rect 34974 1554 34998 1582
rect 35026 1554 35054 1582
rect 34554 1538 35054 1554
rect 37054 18438 37554 18454
rect 37054 18410 37082 18438
rect 37110 18410 37134 18438
rect 37162 18410 37186 18438
rect 37214 18410 37238 18438
rect 37266 18410 37290 18438
rect 37318 18410 37342 18438
rect 37370 18410 37394 18438
rect 37422 18410 37446 18438
rect 37474 18410 37498 18438
rect 37526 18410 37554 18438
rect 37054 17654 37554 18410
rect 37054 17626 37082 17654
rect 37110 17626 37134 17654
rect 37162 17626 37186 17654
rect 37214 17626 37238 17654
rect 37266 17626 37290 17654
rect 37318 17626 37342 17654
rect 37370 17626 37394 17654
rect 37422 17626 37446 17654
rect 37474 17626 37498 17654
rect 37526 17626 37554 17654
rect 37054 16870 37554 17626
rect 37054 16842 37082 16870
rect 37110 16842 37134 16870
rect 37162 16842 37186 16870
rect 37214 16842 37238 16870
rect 37266 16842 37290 16870
rect 37318 16842 37342 16870
rect 37370 16842 37394 16870
rect 37422 16842 37446 16870
rect 37474 16842 37498 16870
rect 37526 16842 37554 16870
rect 37054 16086 37554 16842
rect 37054 16058 37082 16086
rect 37110 16058 37134 16086
rect 37162 16058 37186 16086
rect 37214 16058 37238 16086
rect 37266 16058 37290 16086
rect 37318 16058 37342 16086
rect 37370 16058 37394 16086
rect 37422 16058 37446 16086
rect 37474 16058 37498 16086
rect 37526 16058 37554 16086
rect 37054 15302 37554 16058
rect 37054 15274 37082 15302
rect 37110 15274 37134 15302
rect 37162 15274 37186 15302
rect 37214 15274 37238 15302
rect 37266 15274 37290 15302
rect 37318 15274 37342 15302
rect 37370 15274 37394 15302
rect 37422 15274 37446 15302
rect 37474 15274 37498 15302
rect 37526 15274 37554 15302
rect 37054 14518 37554 15274
rect 37054 14490 37082 14518
rect 37110 14490 37134 14518
rect 37162 14490 37186 14518
rect 37214 14490 37238 14518
rect 37266 14490 37290 14518
rect 37318 14490 37342 14518
rect 37370 14490 37394 14518
rect 37422 14490 37446 14518
rect 37474 14490 37498 14518
rect 37526 14490 37554 14518
rect 37054 13734 37554 14490
rect 37054 13706 37082 13734
rect 37110 13706 37134 13734
rect 37162 13706 37186 13734
rect 37214 13706 37238 13734
rect 37266 13706 37290 13734
rect 37318 13706 37342 13734
rect 37370 13706 37394 13734
rect 37422 13706 37446 13734
rect 37474 13706 37498 13734
rect 37526 13706 37554 13734
rect 37054 12950 37554 13706
rect 37054 12922 37082 12950
rect 37110 12922 37134 12950
rect 37162 12922 37186 12950
rect 37214 12922 37238 12950
rect 37266 12922 37290 12950
rect 37318 12922 37342 12950
rect 37370 12922 37394 12950
rect 37422 12922 37446 12950
rect 37474 12922 37498 12950
rect 37526 12922 37554 12950
rect 37054 12166 37554 12922
rect 37054 12138 37082 12166
rect 37110 12138 37134 12166
rect 37162 12138 37186 12166
rect 37214 12138 37238 12166
rect 37266 12138 37290 12166
rect 37318 12138 37342 12166
rect 37370 12138 37394 12166
rect 37422 12138 37446 12166
rect 37474 12138 37498 12166
rect 37526 12138 37554 12166
rect 37054 11382 37554 12138
rect 37054 11354 37082 11382
rect 37110 11354 37134 11382
rect 37162 11354 37186 11382
rect 37214 11354 37238 11382
rect 37266 11354 37290 11382
rect 37318 11354 37342 11382
rect 37370 11354 37394 11382
rect 37422 11354 37446 11382
rect 37474 11354 37498 11382
rect 37526 11354 37554 11382
rect 37054 10598 37554 11354
rect 37054 10570 37082 10598
rect 37110 10570 37134 10598
rect 37162 10570 37186 10598
rect 37214 10570 37238 10598
rect 37266 10570 37290 10598
rect 37318 10570 37342 10598
rect 37370 10570 37394 10598
rect 37422 10570 37446 10598
rect 37474 10570 37498 10598
rect 37526 10570 37554 10598
rect 37054 9814 37554 10570
rect 37054 9786 37082 9814
rect 37110 9786 37134 9814
rect 37162 9786 37186 9814
rect 37214 9786 37238 9814
rect 37266 9786 37290 9814
rect 37318 9786 37342 9814
rect 37370 9786 37394 9814
rect 37422 9786 37446 9814
rect 37474 9786 37498 9814
rect 37526 9786 37554 9814
rect 37054 9030 37554 9786
rect 37054 9002 37082 9030
rect 37110 9002 37134 9030
rect 37162 9002 37186 9030
rect 37214 9002 37238 9030
rect 37266 9002 37290 9030
rect 37318 9002 37342 9030
rect 37370 9002 37394 9030
rect 37422 9002 37446 9030
rect 37474 9002 37498 9030
rect 37526 9002 37554 9030
rect 37054 8246 37554 9002
rect 37054 8218 37082 8246
rect 37110 8218 37134 8246
rect 37162 8218 37186 8246
rect 37214 8218 37238 8246
rect 37266 8218 37290 8246
rect 37318 8218 37342 8246
rect 37370 8218 37394 8246
rect 37422 8218 37446 8246
rect 37474 8218 37498 8246
rect 37526 8218 37554 8246
rect 37054 7462 37554 8218
rect 37054 7434 37082 7462
rect 37110 7434 37134 7462
rect 37162 7434 37186 7462
rect 37214 7434 37238 7462
rect 37266 7434 37290 7462
rect 37318 7434 37342 7462
rect 37370 7434 37394 7462
rect 37422 7434 37446 7462
rect 37474 7434 37498 7462
rect 37526 7434 37554 7462
rect 37054 6678 37554 7434
rect 37054 6650 37082 6678
rect 37110 6650 37134 6678
rect 37162 6650 37186 6678
rect 37214 6650 37238 6678
rect 37266 6650 37290 6678
rect 37318 6650 37342 6678
rect 37370 6650 37394 6678
rect 37422 6650 37446 6678
rect 37474 6650 37498 6678
rect 37526 6650 37554 6678
rect 37054 5894 37554 6650
rect 37054 5866 37082 5894
rect 37110 5866 37134 5894
rect 37162 5866 37186 5894
rect 37214 5866 37238 5894
rect 37266 5866 37290 5894
rect 37318 5866 37342 5894
rect 37370 5866 37394 5894
rect 37422 5866 37446 5894
rect 37474 5866 37498 5894
rect 37526 5866 37554 5894
rect 37054 5110 37554 5866
rect 37054 5082 37082 5110
rect 37110 5082 37134 5110
rect 37162 5082 37186 5110
rect 37214 5082 37238 5110
rect 37266 5082 37290 5110
rect 37318 5082 37342 5110
rect 37370 5082 37394 5110
rect 37422 5082 37446 5110
rect 37474 5082 37498 5110
rect 37526 5082 37554 5110
rect 37054 4326 37554 5082
rect 37054 4298 37082 4326
rect 37110 4298 37134 4326
rect 37162 4298 37186 4326
rect 37214 4298 37238 4326
rect 37266 4298 37290 4326
rect 37318 4298 37342 4326
rect 37370 4298 37394 4326
rect 37422 4298 37446 4326
rect 37474 4298 37498 4326
rect 37526 4298 37554 4326
rect 37054 3542 37554 4298
rect 37054 3514 37082 3542
rect 37110 3514 37134 3542
rect 37162 3514 37186 3542
rect 37214 3514 37238 3542
rect 37266 3514 37290 3542
rect 37318 3514 37342 3542
rect 37370 3514 37394 3542
rect 37422 3514 37446 3542
rect 37474 3514 37498 3542
rect 37526 3514 37554 3542
rect 37054 2758 37554 3514
rect 37054 2730 37082 2758
rect 37110 2730 37134 2758
rect 37162 2730 37186 2758
rect 37214 2730 37238 2758
rect 37266 2730 37290 2758
rect 37318 2730 37342 2758
rect 37370 2730 37394 2758
rect 37422 2730 37446 2758
rect 37474 2730 37498 2758
rect 37526 2730 37554 2758
rect 37054 1974 37554 2730
rect 37054 1946 37082 1974
rect 37110 1946 37134 1974
rect 37162 1946 37186 1974
rect 37214 1946 37238 1974
rect 37266 1946 37290 1974
rect 37318 1946 37342 1974
rect 37370 1946 37394 1974
rect 37422 1946 37446 1974
rect 37474 1946 37498 1974
rect 37526 1946 37554 1974
rect 37054 1538 37554 1946
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2576 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37
timestamp 1667941163
transform 1 0 2744 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1667941163
transform 1 0 4536 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1667941163
transform 1 0 4704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1667941163
transform 1 0 6496 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1667941163
transform 1 0 6664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1667941163
transform 1 0 8456 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142
timestamp 1667941163
transform 1 0 8624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1667941163
transform 1 0 10416 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_177
timestamp 1667941163
transform 1 0 10584 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1667941163
transform 1 0 12376 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_212
timestamp 1667941163
transform 1 0 12544 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1667941163
transform 1 0 14336 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_247 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 14504 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 14728 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_276
timestamp 1667941163
transform 1 0 16128 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1667941163
transform 1 0 16464 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_307
timestamp 1667941163
transform 1 0 17864 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1667941163
transform 1 0 18424 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_342
timestamp 1667941163
transform 1 0 19824 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_352
timestamp 1667941163
transform 1 0 20384 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1667941163
transform 1 0 22176 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1667941163
transform 1 0 22344 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_412
timestamp 1667941163
transform 1 0 23744 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1667941163
transform 1 0 24304 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_447
timestamp 1667941163
transform 1 0 25704 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1667941163
transform 1 0 26264 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_482
timestamp 1667941163
transform 1 0 27664 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1667941163
transform 1 0 28224 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_517
timestamp 1667941163
transform 1 0 29624 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1667941163
transform 1 0 30184 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_552
timestamp 1667941163
transform 1 0 31584 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1667941163
transform 1 0 32144 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_587
timestamp 1667941163
transform 1 0 33544 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1667941163
transform 1 0 34104 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_622
timestamp 1667941163
transform 1 0 35504 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1667941163
transform 1 0 36064 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_657
timestamp 1667941163
transform 1 0 37464 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1667941163
transform 1 0 38024 0 1 1568
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_676 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 38528 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_686
timestamp 1667941163
transform 1 0 39088 0 1 1568
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 784 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_18
timestamp 1667941163
transform 1 0 1680 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_44
timestamp 1667941163
transform 1 0 3136 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1667941163
transform 1 0 4592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_73
timestamp 1667941163
transform 1 0 4760 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_89
timestamp 1667941163
transform 1 0 5656 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_115
timestamp 1667941163
transform 1 0 7112 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1667941163
transform 1 0 8568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_144
timestamp 1667941163
transform 1 0 8736 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_160
timestamp 1667941163
transform 1 0 9632 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_186
timestamp 1667941163
transform 1 0 11088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1667941163
transform 1 0 12544 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_215
timestamp 1667941163
transform 1 0 12712 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_223
timestamp 1667941163
transform 1 0 13160 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_227
timestamp 1667941163
transform 1 0 13384 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_229
timestamp 1667941163
transform 1 0 13496 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_254
timestamp 1667941163
transform 1 0 14896 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_256
timestamp 1667941163
transform 1 0 15008 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 16408 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1667941163
transform 1 0 16520 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1667941163
transform 1 0 16688 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_311
timestamp 1667941163
transform 1 0 18088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_337
timestamp 1667941163
transform 1 0 19544 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_353
timestamp 1667941163
transform 1 0 20440 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1667941163
transform 1 0 20664 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_382
timestamp 1667941163
transform 1 0 22064 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_408
timestamp 1667941163
transform 1 0 23520 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_416
timestamp 1667941163
transform 1 0 23968 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1667941163
transform 1 0 24472 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1667941163
transform 1 0 24640 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_453
timestamp 1667941163
transform 1 0 26040 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_479
timestamp 1667941163
transform 1 0 27496 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_487
timestamp 1667941163
transform 1 0 27944 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1667941163
transform 1 0 28448 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1667941163
transform 1 0 28616 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_524
timestamp 1667941163
transform 1 0 30016 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_550
timestamp 1667941163
transform 1 0 31472 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_560
timestamp 1667941163
transform 1 0 32032 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1667941163
transform 1 0 32592 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_595
timestamp 1667941163
transform 1 0 33992 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_621
timestamp 1667941163
transform 1 0 35448 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_631
timestamp 1667941163
transform 1 0 36008 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1667941163
transform 1 0 36568 0 -1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_666
timestamp 1667941163
transform 1 0 37968 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_676
timestamp 1667941163
transform 1 0 38528 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_686
timestamp 1667941163
transform 1 0 39088 0 -1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_2
timestamp 1667941163
transform 1 0 784 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1667941163
transform 1 0 2576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_37
timestamp 1667941163
transform 1 0 2744 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_53
timestamp 1667941163
transform 1 0 3640 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_79
timestamp 1667941163
transform 1 0 5096 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1667941163
transform 1 0 6552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_108
timestamp 1667941163
transform 1 0 6720 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_124
timestamp 1667941163
transform 1 0 7616 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_150
timestamp 1667941163
transform 1 0 9072 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1667941163
transform 1 0 10528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_179
timestamp 1667941163
transform 1 0 10696 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_187
timestamp 1667941163
transform 1 0 11144 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_191
timestamp 1667941163
transform 1 0 11368 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_193
timestamp 1667941163
transform 1 0 11480 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_218
timestamp 1667941163
transform 1 0 12880 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_244
timestamp 1667941163
transform 1 0 14336 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_250
timestamp 1667941163
transform 1 0 14672 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_258
timestamp 1667941163
transform 1 0 15120 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_283
timestamp 1667941163
transform 1 0 16520 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_309
timestamp 1667941163
transform 1 0 17976 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_317
timestamp 1667941163
transform 1 0 18424 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_321
timestamp 1667941163
transform 1 0 18648 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_337
timestamp 1667941163
transform 1 0 19544 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_341
timestamp 1667941163
transform 1 0 19768 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_367
timestamp 1667941163
transform 1 0 21224 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_383
timestamp 1667941163
transform 1 0 22120 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_387
timestamp 1667941163
transform 1 0 22344 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1667941163
transform 1 0 22456 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1667941163
transform 1 0 22624 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_417
timestamp 1667941163
transform 1 0 24024 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_443
timestamp 1667941163
transform 1 0 25480 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_451
timestamp 1667941163
transform 1 0 25928 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1667941163
transform 1 0 26432 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1667941163
transform 1 0 26600 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_488
timestamp 1667941163
transform 1 0 28000 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_514
timestamp 1667941163
transform 1 0 29456 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_522
timestamp 1667941163
transform 1 0 29904 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1667941163
transform 1 0 30408 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1667941163
transform 1 0 30576 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_559
timestamp 1667941163
transform 1 0 31976 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_585
timestamp 1667941163
transform 1 0 33432 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_595
timestamp 1667941163
transform 1 0 33992 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1667941163
transform 1 0 34552 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_630
timestamp 1667941163
transform 1 0 35952 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_656
timestamp 1667941163
transform 1 0 37408 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_666
timestamp 1667941163
transform 1 0 37968 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_676
timestamp 1667941163
transform 1 0 38528 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_685
timestamp 1667941163
transform 1 0 39032 0 1 2352
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_687
timestamp 1667941163
transform 1 0 39144 0 1 2352
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_2
timestamp 1667941163
transform 1 0 784 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_18
timestamp 1667941163
transform 1 0 1680 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_44
timestamp 1667941163
transform 1 0 3136 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1667941163
transform 1 0 4592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1667941163
transform 1 0 4760 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_89
timestamp 1667941163
transform 1 0 5656 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_115
timestamp 1667941163
transform 1 0 7112 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1667941163
transform 1 0 8568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_144
timestamp 1667941163
transform 1 0 8736 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_160
timestamp 1667941163
transform 1 0 9632 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_186
timestamp 1667941163
transform 1 0 11088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1667941163
transform 1 0 12544 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_215
timestamp 1667941163
transform 1 0 12712 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_219
timestamp 1667941163
transform 1 0 12936 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_245
timestamp 1667941163
transform 1 0 14392 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_249
timestamp 1667941163
transform 1 0 14616 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_275
timestamp 1667941163
transform 1 0 16072 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1667941163
transform 1 0 16520 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1667941163
transform 1 0 16688 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_311
timestamp 1667941163
transform 1 0 18088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_337
timestamp 1667941163
transform 1 0 19544 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_353
timestamp 1667941163
transform 1 0 20440 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1667941163
transform 1 0 20664 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_382
timestamp 1667941163
transform 1 0 22064 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_408
timestamp 1667941163
transform 1 0 23520 0 -1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_424
timestamp 1667941163
transform 1 0 24416 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1667941163
transform 1 0 24640 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_453
timestamp 1667941163
transform 1 0 26040 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_479
timestamp 1667941163
transform 1 0 27496 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_487
timestamp 1667941163
transform 1 0 27944 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1667941163
transform 1 0 28448 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1667941163
transform 1 0 28616 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_524
timestamp 1667941163
transform 1 0 30016 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_550
timestamp 1667941163
transform 1 0 31472 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_558
timestamp 1667941163
transform 1 0 31920 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1667941163
transform 1 0 32424 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_570
timestamp 1667941163
transform 1 0 32592 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_595
timestamp 1667941163
transform 1 0 33992 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_621
timestamp 1667941163
transform 1 0 35448 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_631
timestamp 1667941163
transform 1 0 36008 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_641
timestamp 1667941163
transform 1 0 36568 0 -1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_666
timestamp 1667941163
transform 1 0 37968 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_676
timestamp 1667941163
transform 1 0 38528 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_686
timestamp 1667941163
transform 1 0 39088 0 -1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_2
timestamp 1667941163
transform 1 0 784 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1667941163
transform 1 0 2576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_37
timestamp 1667941163
transform 1 0 2744 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_53
timestamp 1667941163
transform 1 0 3640 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_79
timestamp 1667941163
transform 1 0 5096 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1667941163
transform 1 0 6552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_108
timestamp 1667941163
transform 1 0 6720 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_124
timestamp 1667941163
transform 1 0 7616 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_150
timestamp 1667941163
transform 1 0 9072 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1667941163
transform 1 0 10528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_179
timestamp 1667941163
transform 1 0 10696 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_195
timestamp 1667941163
transform 1 0 11592 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_221
timestamp 1667941163
transform 1 0 13048 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1667941163
transform 1 0 14504 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_250
timestamp 1667941163
transform 1 0 14672 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_258
timestamp 1667941163
transform 1 0 15120 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_262
timestamp 1667941163
transform 1 0 15344 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_288
timestamp 1667941163
transform 1 0 16800 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 18256 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1667941163
transform 1 0 18480 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1667941163
transform 1 0 18648 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_346
timestamp 1667941163
transform 1 0 20048 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_372
timestamp 1667941163
transform 1 0 21504 0 1 3136
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_388
timestamp 1667941163
transform 1 0 22400 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1667941163
transform 1 0 22624 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_417
timestamp 1667941163
transform 1 0 24024 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_443
timestamp 1667941163
transform 1 0 25480 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_451
timestamp 1667941163
transform 1 0 25928 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1667941163
transform 1 0 26432 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1667941163
transform 1 0 26600 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_488
timestamp 1667941163
transform 1 0 28000 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_514
timestamp 1667941163
transform 1 0 29456 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_522
timestamp 1667941163
transform 1 0 29904 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1667941163
transform 1 0 30408 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_534
timestamp 1667941163
transform 1 0 30576 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_559
timestamp 1667941163
transform 1 0 31976 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_585
timestamp 1667941163
transform 1 0 33432 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_595
timestamp 1667941163
transform 1 0 33992 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_605
timestamp 1667941163
transform 1 0 34552 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_630
timestamp 1667941163
transform 1 0 35952 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_656
timestamp 1667941163
transform 1 0 37408 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_666
timestamp 1667941163
transform 1 0 37968 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_676
timestamp 1667941163
transform 1 0 38528 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_685
timestamp 1667941163
transform 1 0 39032 0 1 3136
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_687
timestamp 1667941163
transform 1 0 39144 0 1 3136
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_2
timestamp 1667941163
transform 1 0 784 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_18
timestamp 1667941163
transform 1 0 1680 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_44
timestamp 1667941163
transform 1 0 3136 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1667941163
transform 1 0 4592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_73
timestamp 1667941163
transform 1 0 4760 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_89
timestamp 1667941163
transform 1 0 5656 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_115
timestamp 1667941163
transform 1 0 7112 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1667941163
transform 1 0 8568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_144
timestamp 1667941163
transform 1 0 8736 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_160
timestamp 1667941163
transform 1 0 9632 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_186
timestamp 1667941163
transform 1 0 11088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1667941163
transform 1 0 12544 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_215
timestamp 1667941163
transform 1 0 12712 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_255
timestamp 1667941163
transform 1 0 14952 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 16408 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1667941163
transform 1 0 16520 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_286
timestamp 1667941163
transform 1 0 16688 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_311
timestamp 1667941163
transform 1 0 18088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_337
timestamp 1667941163
transform 1 0 19544 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_353
timestamp 1667941163
transform 1 0 20440 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1667941163
transform 1 0 20664 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_382
timestamp 1667941163
transform 1 0 22064 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_408
timestamp 1667941163
transform 1 0 23520 0 -1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_424
timestamp 1667941163
transform 1 0 24416 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1667941163
transform 1 0 24640 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_453
timestamp 1667941163
transform 1 0 26040 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_479
timestamp 1667941163
transform 1 0 27496 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_487
timestamp 1667941163
transform 1 0 27944 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1667941163
transform 1 0 28448 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_499
timestamp 1667941163
transform 1 0 28616 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_524
timestamp 1667941163
transform 1 0 30016 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_550
timestamp 1667941163
transform 1 0 31472 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_558
timestamp 1667941163
transform 1 0 31920 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1667941163
transform 1 0 32424 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_570
timestamp 1667941163
transform 1 0 32592 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_595
timestamp 1667941163
transform 1 0 33992 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_621
timestamp 1667941163
transform 1 0 35448 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_631
timestamp 1667941163
transform 1 0 36008 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_641
timestamp 1667941163
transform 1 0 36568 0 -1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_666
timestamp 1667941163
transform 1 0 37968 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_676
timestamp 1667941163
transform 1 0 38528 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_686
timestamp 1667941163
transform 1 0 39088 0 -1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_2
timestamp 1667941163
transform 1 0 784 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1667941163
transform 1 0 2576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1667941163
transform 1 0 2744 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_53
timestamp 1667941163
transform 1 0 3640 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_79
timestamp 1667941163
transform 1 0 5096 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1667941163
transform 1 0 6552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_108
timestamp 1667941163
transform 1 0 6720 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_124
timestamp 1667941163
transform 1 0 7616 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_150
timestamp 1667941163
transform 1 0 9072 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1667941163
transform 1 0 10528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_179
timestamp 1667941163
transform 1 0 10696 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_195
timestamp 1667941163
transform 1 0 11592 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_221
timestamp 1667941163
transform 1 0 13048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1667941163
transform 1 0 14504 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_250
timestamp 1667941163
transform 1 0 14672 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_258
timestamp 1667941163
transform 1 0 15120 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_260
timestamp 1667941163
transform 1 0 15232 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_285
timestamp 1667941163
transform 1 0 16632 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_311
timestamp 1667941163
transform 1 0 18088 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1667941163
transform 1 0 18648 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_346
timestamp 1667941163
transform 1 0 20048 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_372
timestamp 1667941163
transform 1 0 21504 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_388
timestamp 1667941163
transform 1 0 22400 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_392
timestamp 1667941163
transform 1 0 22624 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_417
timestamp 1667941163
transform 1 0 24024 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_443
timestamp 1667941163
transform 1 0 25480 0 1 3920
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_459
timestamp 1667941163
transform 1 0 26376 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1667941163
transform 1 0 26600 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_488
timestamp 1667941163
transform 1 0 28000 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_514
timestamp 1667941163
transform 1 0 29456 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_522
timestamp 1667941163
transform 1 0 29904 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1667941163
transform 1 0 30408 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_534
timestamp 1667941163
transform 1 0 30576 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_559
timestamp 1667941163
transform 1 0 31976 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_585
timestamp 1667941163
transform 1 0 33432 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_595
timestamp 1667941163
transform 1 0 33992 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_605
timestamp 1667941163
transform 1 0 34552 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_630
timestamp 1667941163
transform 1 0 35952 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_656
timestamp 1667941163
transform 1 0 37408 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_666
timestamp 1667941163
transform 1 0 37968 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_676
timestamp 1667941163
transform 1 0 38528 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_685
timestamp 1667941163
transform 1 0 39032 0 1 3920
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_687
timestamp 1667941163
transform 1 0 39144 0 1 3920
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_2
timestamp 1667941163
transform 1 0 784 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_18
timestamp 1667941163
transform 1 0 1680 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_44
timestamp 1667941163
transform 1 0 3136 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 4592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1667941163
transform 1 0 4760 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_89
timestamp 1667941163
transform 1 0 5656 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_115
timestamp 1667941163
transform 1 0 7112 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1667941163
transform 1 0 8568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_144
timestamp 1667941163
transform 1 0 8736 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1667941163
transform 1 0 9632 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_186
timestamp 1667941163
transform 1 0 11088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1667941163
transform 1 0 12544 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_215
timestamp 1667941163
transform 1 0 12712 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_223
timestamp 1667941163
transform 1 0 13160 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_227
timestamp 1667941163
transform 1 0 13384 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_253
timestamp 1667941163
transform 1 0 14840 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1667941163
transform 1 0 16296 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1667941163
transform 1 0 16520 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1667941163
transform 1 0 16688 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_311
timestamp 1667941163
transform 1 0 18088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_337
timestamp 1667941163
transform 1 0 19544 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_353
timestamp 1667941163
transform 1 0 20440 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_357
timestamp 1667941163
transform 1 0 20664 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_382
timestamp 1667941163
transform 1 0 22064 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_408
timestamp 1667941163
transform 1 0 23520 0 -1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_424
timestamp 1667941163
transform 1 0 24416 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1667941163
transform 1 0 24640 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_453
timestamp 1667941163
transform 1 0 26040 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_479
timestamp 1667941163
transform 1 0 27496 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_487
timestamp 1667941163
transform 1 0 27944 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1667941163
transform 1 0 28448 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_499
timestamp 1667941163
transform 1 0 28616 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_524
timestamp 1667941163
transform 1 0 30016 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_550
timestamp 1667941163
transform 1 0 31472 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_558
timestamp 1667941163
transform 1 0 31920 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1667941163
transform 1 0 32424 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_570
timestamp 1667941163
transform 1 0 32592 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_595
timestamp 1667941163
transform 1 0 33992 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_621
timestamp 1667941163
transform 1 0 35448 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_631
timestamp 1667941163
transform 1 0 36008 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_641
timestamp 1667941163
transform 1 0 36568 0 -1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_666
timestamp 1667941163
transform 1 0 37968 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_676
timestamp 1667941163
transform 1 0 38528 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_686
timestamp 1667941163
transform 1 0 39088 0 -1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_2
timestamp 1667941163
transform 1 0 784 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1667941163
transform 1 0 2576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1667941163
transform 1 0 2744 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_53
timestamp 1667941163
transform 1 0 3640 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_79
timestamp 1667941163
transform 1 0 5096 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1667941163
transform 1 0 6552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_108
timestamp 1667941163
transform 1 0 6720 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_124
timestamp 1667941163
transform 1 0 7616 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_150
timestamp 1667941163
transform 1 0 9072 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1667941163
transform 1 0 10528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_179
timestamp 1667941163
transform 1 0 10696 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_195
timestamp 1667941163
transform 1 0 11592 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_221
timestamp 1667941163
transform 1 0 13048 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1667941163
transform 1 0 14504 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_250
timestamp 1667941163
transform 1 0 14672 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_258
timestamp 1667941163
transform 1 0 15120 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_260
timestamp 1667941163
transform 1 0 15232 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_285
timestamp 1667941163
transform 1 0 16632 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_311
timestamp 1667941163
transform 1 0 18088 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1667941163
transform 1 0 18648 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_346
timestamp 1667941163
transform 1 0 20048 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_372
timestamp 1667941163
transform 1 0 21504 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_388
timestamp 1667941163
transform 1 0 22400 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1667941163
transform 1 0 22624 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_417
timestamp 1667941163
transform 1 0 24024 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_443
timestamp 1667941163
transform 1 0 25480 0 1 4704
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_459
timestamp 1667941163
transform 1 0 26376 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_463
timestamp 1667941163
transform 1 0 26600 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_488
timestamp 1667941163
transform 1 0 28000 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_514
timestamp 1667941163
transform 1 0 29456 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_522
timestamp 1667941163
transform 1 0 29904 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1667941163
transform 1 0 30408 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_534
timestamp 1667941163
transform 1 0 30576 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_559
timestamp 1667941163
transform 1 0 31976 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_585
timestamp 1667941163
transform 1 0 33432 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_595
timestamp 1667941163
transform 1 0 33992 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_605
timestamp 1667941163
transform 1 0 34552 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_630
timestamp 1667941163
transform 1 0 35952 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_656
timestamp 1667941163
transform 1 0 37408 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_666
timestamp 1667941163
transform 1 0 37968 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_676
timestamp 1667941163
transform 1 0 38528 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_685
timestamp 1667941163
transform 1 0 39032 0 1 4704
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_687
timestamp 1667941163
transform 1 0 39144 0 1 4704
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_2
timestamp 1667941163
transform 1 0 784 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_18
timestamp 1667941163
transform 1 0 1680 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_44
timestamp 1667941163
transform 1 0 3136 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 4592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_73
timestamp 1667941163
transform 1 0 4760 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_89
timestamp 1667941163
transform 1 0 5656 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_115
timestamp 1667941163
transform 1 0 7112 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1667941163
transform 1 0 8568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_144
timestamp 1667941163
transform 1 0 8736 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_160
timestamp 1667941163
transform 1 0 9632 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_186
timestamp 1667941163
transform 1 0 11088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1667941163
transform 1 0 12544 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_215
timestamp 1667941163
transform 1 0 12712 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_223
timestamp 1667941163
transform 1 0 13160 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_251
timestamp 1667941163
transform 1 0 14728 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_277
timestamp 1667941163
transform 1 0 16184 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 16408 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1667941163
transform 1 0 16520 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_286
timestamp 1667941163
transform 1 0 16688 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_311
timestamp 1667941163
transform 1 0 18088 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_337
timestamp 1667941163
transform 1 0 19544 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_353
timestamp 1667941163
transform 1 0 20440 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1667941163
transform 1 0 20664 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_382
timestamp 1667941163
transform 1 0 22064 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_408
timestamp 1667941163
transform 1 0 23520 0 -1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_424
timestamp 1667941163
transform 1 0 24416 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_428
timestamp 1667941163
transform 1 0 24640 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_453
timestamp 1667941163
transform 1 0 26040 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_479
timestamp 1667941163
transform 1 0 27496 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_487
timestamp 1667941163
transform 1 0 27944 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1667941163
transform 1 0 28448 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_499
timestamp 1667941163
transform 1 0 28616 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_524
timestamp 1667941163
transform 1 0 30016 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_550
timestamp 1667941163
transform 1 0 31472 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_558
timestamp 1667941163
transform 1 0 31920 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1667941163
transform 1 0 32424 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_570
timestamp 1667941163
transform 1 0 32592 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_595
timestamp 1667941163
transform 1 0 33992 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_621
timestamp 1667941163
transform 1 0 35448 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_631
timestamp 1667941163
transform 1 0 36008 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_641
timestamp 1667941163
transform 1 0 36568 0 -1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_666
timestamp 1667941163
transform 1 0 37968 0 -1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_676
timestamp 1667941163
transform 1 0 38528 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_684
timestamp 1667941163
transform 1 0 38976 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1667941163
transform 1 0 784 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1667941163
transform 1 0 2576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1667941163
transform 1 0 2744 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1667941163
transform 1 0 3640 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_79
timestamp 1667941163
transform 1 0 5096 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 6552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_108
timestamp 1667941163
transform 1 0 6720 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_124
timestamp 1667941163
transform 1 0 7616 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_150
timestamp 1667941163
transform 1 0 9072 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1667941163
transform 1 0 10528 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_179
timestamp 1667941163
transform 1 0 10696 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_195
timestamp 1667941163
transform 1 0 11592 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_221
timestamp 1667941163
transform 1 0 13048 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1667941163
transform 1 0 14504 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_250
timestamp 1667941163
transform 1 0 14672 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_254
timestamp 1667941163
transform 1 0 14896 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_280
timestamp 1667941163
transform 1 0 16352 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_306
timestamp 1667941163
transform 1 0 17808 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 18256 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1667941163
transform 1 0 18480 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1667941163
transform 1 0 18648 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_346
timestamp 1667941163
transform 1 0 20048 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_372
timestamp 1667941163
transform 1 0 21504 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_388
timestamp 1667941163
transform 1 0 22400 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_392
timestamp 1667941163
transform 1 0 22624 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_417
timestamp 1667941163
transform 1 0 24024 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_443
timestamp 1667941163
transform 1 0 25480 0 1 5488
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_459
timestamp 1667941163
transform 1 0 26376 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1667941163
transform 1 0 26600 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_488
timestamp 1667941163
transform 1 0 28000 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_514
timestamp 1667941163
transform 1 0 29456 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_522
timestamp 1667941163
transform 1 0 29904 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1667941163
transform 1 0 30408 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_534
timestamp 1667941163
transform 1 0 30576 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_559
timestamp 1667941163
transform 1 0 31976 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_585
timestamp 1667941163
transform 1 0 33432 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_595
timestamp 1667941163
transform 1 0 33992 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_605
timestamp 1667941163
transform 1 0 34552 0 1 5488
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_630
timestamp 1667941163
transform 1 0 35952 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_656
timestamp 1667941163
transform 1 0 37408 0 1 5488
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_666
timestamp 1667941163
transform 1 0 37968 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_676
timestamp 1667941163
transform 1 0 38528 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_684
timestamp 1667941163
transform 1 0 38976 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1667941163
transform 1 0 784 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_18
timestamp 1667941163
transform 1 0 1680 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_44
timestamp 1667941163
transform 1 0 3136 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1667941163
transform 1 0 4592 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_73
timestamp 1667941163
transform 1 0 4760 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_89
timestamp 1667941163
transform 1 0 5656 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_115
timestamp 1667941163
transform 1 0 7112 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1667941163
transform 1 0 8568 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_144
timestamp 1667941163
transform 1 0 8736 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_160
timestamp 1667941163
transform 1 0 9632 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_186
timestamp 1667941163
transform 1 0 11088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1667941163
transform 1 0 12544 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_215
timestamp 1667941163
transform 1 0 12712 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_255
timestamp 1667941163
transform 1 0 14952 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 16408 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1667941163
transform 1 0 16520 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_286
timestamp 1667941163
transform 1 0 16688 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_311
timestamp 1667941163
transform 1 0 18088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_337
timestamp 1667941163
transform 1 0 19544 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_353
timestamp 1667941163
transform 1 0 20440 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1667941163
transform 1 0 20664 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_382
timestamp 1667941163
transform 1 0 22064 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_408
timestamp 1667941163
transform 1 0 23520 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_424
timestamp 1667941163
transform 1 0 24416 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1667941163
transform 1 0 24640 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_453
timestamp 1667941163
transform 1 0 26040 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_479
timestamp 1667941163
transform 1 0 27496 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_495
timestamp 1667941163
transform 1 0 28392 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_499
timestamp 1667941163
transform 1 0 28616 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_524
timestamp 1667941163
transform 1 0 30016 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_550
timestamp 1667941163
transform 1 0 31472 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_558
timestamp 1667941163
transform 1 0 31920 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1667941163
transform 1 0 32424 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_570
timestamp 1667941163
transform 1 0 32592 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_595
timestamp 1667941163
transform 1 0 33992 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_621
timestamp 1667941163
transform 1 0 35448 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_631
timestamp 1667941163
transform 1 0 36008 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_641
timestamp 1667941163
transform 1 0 36568 0 -1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_666
timestamp 1667941163
transform 1 0 37968 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_682
timestamp 1667941163
transform 1 0 38864 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_686
timestamp 1667941163
transform 1 0 39088 0 -1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_2
timestamp 1667941163
transform 1 0 784 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1667941163
transform 1 0 2576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_37
timestamp 1667941163
transform 1 0 2744 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_53
timestamp 1667941163
transform 1 0 3640 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_79
timestamp 1667941163
transform 1 0 5096 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1667941163
transform 1 0 6552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_108
timestamp 1667941163
transform 1 0 6720 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_124
timestamp 1667941163
transform 1 0 7616 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_150
timestamp 1667941163
transform 1 0 9072 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1667941163
transform 1 0 10528 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_179
timestamp 1667941163
transform 1 0 10696 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_195
timestamp 1667941163
transform 1 0 11592 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_221
timestamp 1667941163
transform 1 0 13048 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1667941163
transform 1 0 14504 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_250
timestamp 1667941163
transform 1 0 14672 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_266
timestamp 1667941163
transform 1 0 15568 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_274
timestamp 1667941163
transform 1 0 16016 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_299
timestamp 1667941163
transform 1 0 17416 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_315
timestamp 1667941163
transform 1 0 18312 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1667941163
transform 1 0 18648 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_346
timestamp 1667941163
transform 1 0 20048 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_372
timestamp 1667941163
transform 1 0 21504 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_388
timestamp 1667941163
transform 1 0 22400 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1667941163
transform 1 0 22624 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_417
timestamp 1667941163
transform 1 0 24024 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_443
timestamp 1667941163
transform 1 0 25480 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_459
timestamp 1667941163
transform 1 0 26376 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_463
timestamp 1667941163
transform 1 0 26600 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_488
timestamp 1667941163
transform 1 0 28000 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_514
timestamp 1667941163
transform 1 0 29456 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_522
timestamp 1667941163
transform 1 0 29904 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1667941163
transform 1 0 30408 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_534
timestamp 1667941163
transform 1 0 30576 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_559
timestamp 1667941163
transform 1 0 31976 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_585
timestamp 1667941163
transform 1 0 33432 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_595
timestamp 1667941163
transform 1 0 33992 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_605
timestamp 1667941163
transform 1 0 34552 0 1 6272
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_630
timestamp 1667941163
transform 1 0 35952 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_656
timestamp 1667941163
transform 1 0 37408 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_672
timestamp 1667941163
transform 1 0 38304 0 1 6272
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_676
timestamp 1667941163
transform 1 0 38528 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_684
timestamp 1667941163
transform 1 0 38976 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1667941163
transform 1 0 784 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_18
timestamp 1667941163
transform 1 0 1680 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_44
timestamp 1667941163
transform 1 0 3136 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1667941163
transform 1 0 4592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_73
timestamp 1667941163
transform 1 0 4760 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_89
timestamp 1667941163
transform 1 0 5656 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_115
timestamp 1667941163
transform 1 0 7112 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 8568 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_144
timestamp 1667941163
transform 1 0 8736 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_160
timestamp 1667941163
transform 1 0 9632 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_186
timestamp 1667941163
transform 1 0 11088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 12544 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_215
timestamp 1667941163
transform 1 0 12712 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_231
timestamp 1667941163
transform 1 0 13608 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_256
timestamp 1667941163
transform 1 0 15008 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_258
timestamp 1667941163
transform 1 0 15120 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1667941163
transform 1 0 16520 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1667941163
transform 1 0 16688 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_311
timestamp 1667941163
transform 1 0 18088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_337
timestamp 1667941163
transform 1 0 19544 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_353
timestamp 1667941163
transform 1 0 20440 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_357
timestamp 1667941163
transform 1 0 20664 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_382
timestamp 1667941163
transform 1 0 22064 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_408
timestamp 1667941163
transform 1 0 23520 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_424
timestamp 1667941163
transform 1 0 24416 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1667941163
transform 1 0 24640 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_453
timestamp 1667941163
transform 1 0 26040 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_479
timestamp 1667941163
transform 1 0 27496 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_495
timestamp 1667941163
transform 1 0 28392 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_499
timestamp 1667941163
transform 1 0 28616 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_524
timestamp 1667941163
transform 1 0 30016 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_550
timestamp 1667941163
transform 1 0 31472 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_558
timestamp 1667941163
transform 1 0 31920 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1667941163
transform 1 0 32424 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_570
timestamp 1667941163
transform 1 0 32592 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_595
timestamp 1667941163
transform 1 0 33992 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_621
timestamp 1667941163
transform 1 0 35448 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_631
timestamp 1667941163
transform 1 0 36008 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_641
timestamp 1667941163
transform 1 0 36568 0 -1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_666
timestamp 1667941163
transform 1 0 37968 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_682
timestamp 1667941163
transform 1 0 38864 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_686
timestamp 1667941163
transform 1 0 39088 0 -1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1667941163
transform 1 0 784 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1667941163
transform 1 0 2576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_37
timestamp 1667941163
transform 1 0 2744 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_53
timestamp 1667941163
transform 1 0 3640 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_79
timestamp 1667941163
transform 1 0 5096 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1667941163
transform 1 0 6552 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_108
timestamp 1667941163
transform 1 0 6720 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_124
timestamp 1667941163
transform 1 0 7616 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_150
timestamp 1667941163
transform 1 0 9072 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1667941163
transform 1 0 10528 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_179
timestamp 1667941163
transform 1 0 10696 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_195
timestamp 1667941163
transform 1 0 11592 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_221
timestamp 1667941163
transform 1 0 13048 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1667941163
transform 1 0 14504 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_250
timestamp 1667941163
transform 1 0 14672 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_254
timestamp 1667941163
transform 1 0 14896 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_256
timestamp 1667941163
transform 1 0 15008 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_281
timestamp 1667941163
transform 1 0 16408 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_309
timestamp 1667941163
transform 1 0 17976 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_317
timestamp 1667941163
transform 1 0 18424 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1667941163
transform 1 0 18648 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_346
timestamp 1667941163
transform 1 0 20048 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_372
timestamp 1667941163
transform 1 0 21504 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_388
timestamp 1667941163
transform 1 0 22400 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_392
timestamp 1667941163
transform 1 0 22624 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_417
timestamp 1667941163
transform 1 0 24024 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_443
timestamp 1667941163
transform 1 0 25480 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_459
timestamp 1667941163
transform 1 0 26376 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_463
timestamp 1667941163
transform 1 0 26600 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_488
timestamp 1667941163
transform 1 0 28000 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_514
timestamp 1667941163
transform 1 0 29456 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_530
timestamp 1667941163
transform 1 0 30352 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_534
timestamp 1667941163
transform 1 0 30576 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_559
timestamp 1667941163
transform 1 0 31976 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_585
timestamp 1667941163
transform 1 0 33432 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_595
timestamp 1667941163
transform 1 0 33992 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_605
timestamp 1667941163
transform 1 0 34552 0 1 7056
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_630
timestamp 1667941163
transform 1 0 35952 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_656
timestamp 1667941163
transform 1 0 37408 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_672
timestamp 1667941163
transform 1 0 38304 0 1 7056
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_676
timestamp 1667941163
transform 1 0 38528 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_684
timestamp 1667941163
transform 1 0 38976 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_2
timestamp 1667941163
transform 1 0 784 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_18
timestamp 1667941163
transform 1 0 1680 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_44
timestamp 1667941163
transform 1 0 3136 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1667941163
transform 1 0 4592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_73
timestamp 1667941163
transform 1 0 4760 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_89
timestamp 1667941163
transform 1 0 5656 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_115
timestamp 1667941163
transform 1 0 7112 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1667941163
transform 1 0 8568 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_144
timestamp 1667941163
transform 1 0 8736 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_160
timestamp 1667941163
transform 1 0 9632 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_186
timestamp 1667941163
transform 1 0 11088 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1667941163
transform 1 0 12544 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_215
timestamp 1667941163
transform 1 0 12712 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_231
timestamp 1667941163
transform 1 0 13608 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_257
timestamp 1667941163
transform 1 0 15064 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1667941163
transform 1 0 16520 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1667941163
transform 1 0 16688 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_311
timestamp 1667941163
transform 1 0 18088 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_337
timestamp 1667941163
transform 1 0 19544 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_353
timestamp 1667941163
transform 1 0 20440 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_357
timestamp 1667941163
transform 1 0 20664 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_382
timestamp 1667941163
transform 1 0 22064 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_408
timestamp 1667941163
transform 1 0 23520 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_424
timestamp 1667941163
transform 1 0 24416 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_428
timestamp 1667941163
transform 1 0 24640 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_453
timestamp 1667941163
transform 1 0 26040 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_479
timestamp 1667941163
transform 1 0 27496 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_495
timestamp 1667941163
transform 1 0 28392 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_499
timestamp 1667941163
transform 1 0 28616 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_524
timestamp 1667941163
transform 1 0 30016 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_550
timestamp 1667941163
transform 1 0 31472 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_558
timestamp 1667941163
transform 1 0 31920 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1667941163
transform 1 0 32424 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_570
timestamp 1667941163
transform 1 0 32592 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_595
timestamp 1667941163
transform 1 0 33992 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_621
timestamp 1667941163
transform 1 0 35448 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_637
timestamp 1667941163
transform 1 0 36344 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_641
timestamp 1667941163
transform 1 0 36568 0 -1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_666
timestamp 1667941163
transform 1 0 37968 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_682
timestamp 1667941163
transform 1 0 38864 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_686
timestamp 1667941163
transform 1 0 39088 0 -1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_2
timestamp 1667941163
transform 1 0 784 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1667941163
transform 1 0 2576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_37
timestamp 1667941163
transform 1 0 2744 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_53
timestamp 1667941163
transform 1 0 3640 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_79
timestamp 1667941163
transform 1 0 5096 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1667941163
transform 1 0 6552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_108
timestamp 1667941163
transform 1 0 6720 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_124
timestamp 1667941163
transform 1 0 7616 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_150
timestamp 1667941163
transform 1 0 9072 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1667941163
transform 1 0 10528 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_179
timestamp 1667941163
transform 1 0 10696 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_195
timestamp 1667941163
transform 1 0 11592 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_221
timestamp 1667941163
transform 1 0 13048 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1667941163
transform 1 0 14504 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_250
timestamp 1667941163
transform 1 0 14672 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_258
timestamp 1667941163
transform 1 0 15120 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_284
timestamp 1667941163
transform 1 0 16576 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_310
timestamp 1667941163
transform 1 0 18032 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1667941163
transform 1 0 18480 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_321
timestamp 1667941163
transform 1 0 18648 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_346
timestamp 1667941163
transform 1 0 20048 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_372
timestamp 1667941163
transform 1 0 21504 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_388
timestamp 1667941163
transform 1 0 22400 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_392
timestamp 1667941163
transform 1 0 22624 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_417
timestamp 1667941163
transform 1 0 24024 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_443
timestamp 1667941163
transform 1 0 25480 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_459
timestamp 1667941163
transform 1 0 26376 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_463
timestamp 1667941163
transform 1 0 26600 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_488
timestamp 1667941163
transform 1 0 28000 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_514
timestamp 1667941163
transform 1 0 29456 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_530
timestamp 1667941163
transform 1 0 30352 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_534
timestamp 1667941163
transform 1 0 30576 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_559
timestamp 1667941163
transform 1 0 31976 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_585
timestamp 1667941163
transform 1 0 33432 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_595
timestamp 1667941163
transform 1 0 33992 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_605
timestamp 1667941163
transform 1 0 34552 0 1 7840
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_630
timestamp 1667941163
transform 1 0 35952 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_656
timestamp 1667941163
transform 1 0 37408 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_672
timestamp 1667941163
transform 1 0 38304 0 1 7840
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_676
timestamp 1667941163
transform 1 0 38528 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_684
timestamp 1667941163
transform 1 0 38976 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_2
timestamp 1667941163
transform 1 0 784 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_18
timestamp 1667941163
transform 1 0 1680 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_44
timestamp 1667941163
transform 1 0 3136 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1667941163
transform 1 0 4592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_73
timestamp 1667941163
transform 1 0 4760 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_89
timestamp 1667941163
transform 1 0 5656 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_115
timestamp 1667941163
transform 1 0 7112 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1667941163
transform 1 0 8568 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_144
timestamp 1667941163
transform 1 0 8736 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_160
timestamp 1667941163
transform 1 0 9632 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_186
timestamp 1667941163
transform 1 0 11088 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1667941163
transform 1 0 12544 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_215
timestamp 1667941163
transform 1 0 12712 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_231
timestamp 1667941163
transform 1 0 13608 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_257
timestamp 1667941163
transform 1 0 15064 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1667941163
transform 1 0 16520 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 16688 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_290
timestamp 1667941163
transform 1 0 16912 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_316
timestamp 1667941163
transform 1 0 18368 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_342
timestamp 1667941163
transform 1 0 19824 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1667941163
transform 1 0 20272 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1667941163
transform 1 0 20496 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_357
timestamp 1667941163
transform 1 0 20664 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_382
timestamp 1667941163
transform 1 0 22064 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_408
timestamp 1667941163
transform 1 0 23520 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_424
timestamp 1667941163
transform 1 0 24416 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_428
timestamp 1667941163
transform 1 0 24640 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_453
timestamp 1667941163
transform 1 0 26040 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_479
timestamp 1667941163
transform 1 0 27496 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_495
timestamp 1667941163
transform 1 0 28392 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_499
timestamp 1667941163
transform 1 0 28616 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_524
timestamp 1667941163
transform 1 0 30016 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_550
timestamp 1667941163
transform 1 0 31472 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_558
timestamp 1667941163
transform 1 0 31920 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1667941163
transform 1 0 32424 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_570
timestamp 1667941163
transform 1 0 32592 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_595
timestamp 1667941163
transform 1 0 33992 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_621
timestamp 1667941163
transform 1 0 35448 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_637
timestamp 1667941163
transform 1 0 36344 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_641
timestamp 1667941163
transform 1 0 36568 0 -1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_666
timestamp 1667941163
transform 1 0 37968 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_682
timestamp 1667941163
transform 1 0 38864 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_686
timestamp 1667941163
transform 1 0 39088 0 -1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_2
timestamp 1667941163
transform 1 0 784 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1667941163
transform 1 0 2576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_37
timestamp 1667941163
transform 1 0 2744 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_53
timestamp 1667941163
transform 1 0 3640 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_79
timestamp 1667941163
transform 1 0 5096 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1667941163
transform 1 0 6552 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_108
timestamp 1667941163
transform 1 0 6720 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_124
timestamp 1667941163
transform 1 0 7616 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_150
timestamp 1667941163
transform 1 0 9072 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1667941163
transform 1 0 10528 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_179
timestamp 1667941163
transform 1 0 10696 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_195
timestamp 1667941163
transform 1 0 11592 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_221
timestamp 1667941163
transform 1 0 13048 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1667941163
transform 1 0 14504 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_250
timestamp 1667941163
transform 1 0 14672 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_258
timestamp 1667941163
transform 1 0 15120 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_262
timestamp 1667941163
transform 1 0 15344 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_287
timestamp 1667941163
transform 1 0 16744 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_291
timestamp 1667941163
transform 1 0 16968 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_293
timestamp 1667941163
transform 1 0 17080 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1667941163
transform 1 0 18480 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1667941163
transform 1 0 18648 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_346
timestamp 1667941163
transform 1 0 20048 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_372
timestamp 1667941163
transform 1 0 21504 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_388
timestamp 1667941163
transform 1 0 22400 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_392
timestamp 1667941163
transform 1 0 22624 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_417
timestamp 1667941163
transform 1 0 24024 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_443
timestamp 1667941163
transform 1 0 25480 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_459
timestamp 1667941163
transform 1 0 26376 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_463
timestamp 1667941163
transform 1 0 26600 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_488
timestamp 1667941163
transform 1 0 28000 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_514
timestamp 1667941163
transform 1 0 29456 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_530
timestamp 1667941163
transform 1 0 30352 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_534
timestamp 1667941163
transform 1 0 30576 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_559
timestamp 1667941163
transform 1 0 31976 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_585
timestamp 1667941163
transform 1 0 33432 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_601
timestamp 1667941163
transform 1 0 34328 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_605
timestamp 1667941163
transform 1 0 34552 0 1 8624
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_630
timestamp 1667941163
transform 1 0 35952 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_656
timestamp 1667941163
transform 1 0 37408 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_672
timestamp 1667941163
transform 1 0 38304 0 1 8624
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_676
timestamp 1667941163
transform 1 0 38528 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_684
timestamp 1667941163
transform 1 0 38976 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_2
timestamp 1667941163
transform 1 0 784 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_18
timestamp 1667941163
transform 1 0 1680 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_44
timestamp 1667941163
transform 1 0 3136 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1667941163
transform 1 0 4592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_73
timestamp 1667941163
transform 1 0 4760 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_89
timestamp 1667941163
transform 1 0 5656 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_115
timestamp 1667941163
transform 1 0 7112 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1667941163
transform 1 0 8568 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_144
timestamp 1667941163
transform 1 0 8736 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_160
timestamp 1667941163
transform 1 0 9632 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_186
timestamp 1667941163
transform 1 0 11088 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1667941163
transform 1 0 12544 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_215
timestamp 1667941163
transform 1 0 12712 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_231
timestamp 1667941163
transform 1 0 13608 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_257
timestamp 1667941163
transform 1 0 15064 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1667941163
transform 1 0 16520 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_286
timestamp 1667941163
transform 1 0 16688 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_318
timestamp 1667941163
transform 1 0 18480 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_344
timestamp 1667941163
transform 1 0 19936 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_352
timestamp 1667941163
transform 1 0 20384 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1667941163
transform 1 0 20496 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_357
timestamp 1667941163
transform 1 0 20664 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_382
timestamp 1667941163
transform 1 0 22064 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_408
timestamp 1667941163
transform 1 0 23520 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_424
timestamp 1667941163
transform 1 0 24416 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1667941163
transform 1 0 24640 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_453
timestamp 1667941163
transform 1 0 26040 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_479
timestamp 1667941163
transform 1 0 27496 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_495
timestamp 1667941163
transform 1 0 28392 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_499
timestamp 1667941163
transform 1 0 28616 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_524
timestamp 1667941163
transform 1 0 30016 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_550
timestamp 1667941163
transform 1 0 31472 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_566
timestamp 1667941163
transform 1 0 32368 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_570
timestamp 1667941163
transform 1 0 32592 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_595
timestamp 1667941163
transform 1 0 33992 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_621
timestamp 1667941163
transform 1 0 35448 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_637
timestamp 1667941163
transform 1 0 36344 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_641
timestamp 1667941163
transform 1 0 36568 0 -1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_666
timestamp 1667941163
transform 1 0 37968 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_682
timestamp 1667941163
transform 1 0 38864 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_686
timestamp 1667941163
transform 1 0 39088 0 -1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_2
timestamp 1667941163
transform 1 0 784 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1667941163
transform 1 0 2576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_37
timestamp 1667941163
transform 1 0 2744 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_53
timestamp 1667941163
transform 1 0 3640 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_79
timestamp 1667941163
transform 1 0 5096 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1667941163
transform 1 0 6552 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_108
timestamp 1667941163
transform 1 0 6720 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_124
timestamp 1667941163
transform 1 0 7616 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_150
timestamp 1667941163
transform 1 0 9072 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1667941163
transform 1 0 10528 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_179
timestamp 1667941163
transform 1 0 10696 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_195
timestamp 1667941163
transform 1 0 11592 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_221
timestamp 1667941163
transform 1 0 13048 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1667941163
transform 1 0 14504 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_250
timestamp 1667941163
transform 1 0 14672 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_258
timestamp 1667941163
transform 1 0 15120 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_262
timestamp 1667941163
transform 1 0 15344 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_288
timestamp 1667941163
transform 1 0 16800 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_316
timestamp 1667941163
transform 1 0 18368 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1667941163
transform 1 0 18480 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_321
timestamp 1667941163
transform 1 0 18648 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_346
timestamp 1667941163
transform 1 0 20048 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_372
timestamp 1667941163
transform 1 0 21504 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_388
timestamp 1667941163
transform 1 0 22400 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_392
timestamp 1667941163
transform 1 0 22624 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_417
timestamp 1667941163
transform 1 0 24024 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_443
timestamp 1667941163
transform 1 0 25480 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_459
timestamp 1667941163
transform 1 0 26376 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_463
timestamp 1667941163
transform 1 0 26600 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_488
timestamp 1667941163
transform 1 0 28000 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_514
timestamp 1667941163
transform 1 0 29456 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_530
timestamp 1667941163
transform 1 0 30352 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_534
timestamp 1667941163
transform 1 0 30576 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_559
timestamp 1667941163
transform 1 0 31976 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_585
timestamp 1667941163
transform 1 0 33432 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_601
timestamp 1667941163
transform 1 0 34328 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_605
timestamp 1667941163
transform 1 0 34552 0 1 9408
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_630
timestamp 1667941163
transform 1 0 35952 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_656
timestamp 1667941163
transform 1 0 37408 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_672
timestamp 1667941163
transform 1 0 38304 0 1 9408
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_676
timestamp 1667941163
transform 1 0 38528 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_684
timestamp 1667941163
transform 1 0 38976 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_2
timestamp 1667941163
transform 1 0 784 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_18
timestamp 1667941163
transform 1 0 1680 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_44
timestamp 1667941163
transform 1 0 3136 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1667941163
transform 1 0 4592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_73
timestamp 1667941163
transform 1 0 4760 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_89
timestamp 1667941163
transform 1 0 5656 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_115
timestamp 1667941163
transform 1 0 7112 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1667941163
transform 1 0 8568 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_144
timestamp 1667941163
transform 1 0 8736 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_160
timestamp 1667941163
transform 1 0 9632 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_186
timestamp 1667941163
transform 1 0 11088 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1667941163
transform 1 0 12544 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_215
timestamp 1667941163
transform 1 0 12712 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_231
timestamp 1667941163
transform 1 0 13608 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_257
timestamp 1667941163
transform 1 0 15064 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1667941163
transform 1 0 16520 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1667941163
transform 1 0 16688 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_311
timestamp 1667941163
transform 1 0 18088 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_337
timestamp 1667941163
transform 1 0 19544 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_353
timestamp 1667941163
transform 1 0 20440 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_357
timestamp 1667941163
transform 1 0 20664 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_382
timestamp 1667941163
transform 1 0 22064 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_408
timestamp 1667941163
transform 1 0 23520 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_424
timestamp 1667941163
transform 1 0 24416 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_428
timestamp 1667941163
transform 1 0 24640 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_453
timestamp 1667941163
transform 1 0 26040 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_479
timestamp 1667941163
transform 1 0 27496 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_495
timestamp 1667941163
transform 1 0 28392 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_499
timestamp 1667941163
transform 1 0 28616 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_524
timestamp 1667941163
transform 1 0 30016 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_550
timestamp 1667941163
transform 1 0 31472 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_566
timestamp 1667941163
transform 1 0 32368 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_570
timestamp 1667941163
transform 1 0 32592 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_595
timestamp 1667941163
transform 1 0 33992 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_621
timestamp 1667941163
transform 1 0 35448 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_637
timestamp 1667941163
transform 1 0 36344 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_641
timestamp 1667941163
transform 1 0 36568 0 -1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_666
timestamp 1667941163
transform 1 0 37968 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_682
timestamp 1667941163
transform 1 0 38864 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_686
timestamp 1667941163
transform 1 0 39088 0 -1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_2
timestamp 1667941163
transform 1 0 784 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1667941163
transform 1 0 2576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_37
timestamp 1667941163
transform 1 0 2744 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_53
timestamp 1667941163
transform 1 0 3640 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_79
timestamp 1667941163
transform 1 0 5096 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1667941163
transform 1 0 6552 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_108
timestamp 1667941163
transform 1 0 6720 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_124
timestamp 1667941163
transform 1 0 7616 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_150
timestamp 1667941163
transform 1 0 9072 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1667941163
transform 1 0 10528 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_179
timestamp 1667941163
transform 1 0 10696 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_195
timestamp 1667941163
transform 1 0 11592 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_221
timestamp 1667941163
transform 1 0 13048 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1667941163
transform 1 0 14504 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_250
timestamp 1667941163
transform 1 0 14672 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_266
timestamp 1667941163
transform 1 0 15568 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_291
timestamp 1667941163
transform 1 0 16968 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1667941163
transform 1 0 18424 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1667941163
transform 1 0 18648 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_346
timestamp 1667941163
transform 1 0 20048 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_372
timestamp 1667941163
transform 1 0 21504 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_388
timestamp 1667941163
transform 1 0 22400 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1667941163
transform 1 0 22624 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_417
timestamp 1667941163
transform 1 0 24024 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_443
timestamp 1667941163
transform 1 0 25480 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_459
timestamp 1667941163
transform 1 0 26376 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_463
timestamp 1667941163
transform 1 0 26600 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_488
timestamp 1667941163
transform 1 0 28000 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_514
timestamp 1667941163
transform 1 0 29456 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_530
timestamp 1667941163
transform 1 0 30352 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_534
timestamp 1667941163
transform 1 0 30576 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_559
timestamp 1667941163
transform 1 0 31976 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_585
timestamp 1667941163
transform 1 0 33432 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_601
timestamp 1667941163
transform 1 0 34328 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_605
timestamp 1667941163
transform 1 0 34552 0 1 10192
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_630
timestamp 1667941163
transform 1 0 35952 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_656
timestamp 1667941163
transform 1 0 37408 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_672
timestamp 1667941163
transform 1 0 38304 0 1 10192
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_676
timestamp 1667941163
transform 1 0 38528 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_684
timestamp 1667941163
transform 1 0 38976 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_2
timestamp 1667941163
transform 1 0 784 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_18
timestamp 1667941163
transform 1 0 1680 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_44
timestamp 1667941163
transform 1 0 3136 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1667941163
transform 1 0 4592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_73
timestamp 1667941163
transform 1 0 4760 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_89
timestamp 1667941163
transform 1 0 5656 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_115
timestamp 1667941163
transform 1 0 7112 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1667941163
transform 1 0 8568 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_144
timestamp 1667941163
transform 1 0 8736 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_160
timestamp 1667941163
transform 1 0 9632 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_186
timestamp 1667941163
transform 1 0 11088 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1667941163
transform 1 0 12544 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_215
timestamp 1667941163
transform 1 0 12712 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_231
timestamp 1667941163
transform 1 0 13608 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_257
timestamp 1667941163
transform 1 0 15064 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1667941163
transform 1 0 16520 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1667941163
transform 1 0 16688 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_311
timestamp 1667941163
transform 1 0 18088 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_337
timestamp 1667941163
transform 1 0 19544 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_353
timestamp 1667941163
transform 1 0 20440 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_357
timestamp 1667941163
transform 1 0 20664 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_382
timestamp 1667941163
transform 1 0 22064 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_408
timestamp 1667941163
transform 1 0 23520 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_424
timestamp 1667941163
transform 1 0 24416 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1667941163
transform 1 0 24640 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_453
timestamp 1667941163
transform 1 0 26040 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_479
timestamp 1667941163
transform 1 0 27496 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_495
timestamp 1667941163
transform 1 0 28392 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_499
timestamp 1667941163
transform 1 0 28616 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_524
timestamp 1667941163
transform 1 0 30016 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_550
timestamp 1667941163
transform 1 0 31472 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_566
timestamp 1667941163
transform 1 0 32368 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_570
timestamp 1667941163
transform 1 0 32592 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_595
timestamp 1667941163
transform 1 0 33992 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_621
timestamp 1667941163
transform 1 0 35448 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_637
timestamp 1667941163
transform 1 0 36344 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_641 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 36568 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_673
timestamp 1667941163
transform 1 0 38360 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_681
timestamp 1667941163
transform 1 0 38808 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_685
timestamp 1667941163
transform 1 0 39032 0 -1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_687
timestamp 1667941163
transform 1 0 39144 0 -1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_2
timestamp 1667941163
transform 1 0 784 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1667941163
transform 1 0 2576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_37
timestamp 1667941163
transform 1 0 2744 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_53
timestamp 1667941163
transform 1 0 3640 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_79
timestamp 1667941163
transform 1 0 5096 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1667941163
transform 1 0 6552 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_108
timestamp 1667941163
transform 1 0 6720 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_124
timestamp 1667941163
transform 1 0 7616 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_150
timestamp 1667941163
transform 1 0 9072 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1667941163
transform 1 0 10528 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_179
timestamp 1667941163
transform 1 0 10696 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_195
timestamp 1667941163
transform 1 0 11592 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_221
timestamp 1667941163
transform 1 0 13048 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1667941163
transform 1 0 14504 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_250
timestamp 1667941163
transform 1 0 14672 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_290
timestamp 1667941163
transform 1 0 16912 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_316
timestamp 1667941163
transform 1 0 18368 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1667941163
transform 1 0 18480 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1667941163
transform 1 0 18648 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_346
timestamp 1667941163
transform 1 0 20048 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_372
timestamp 1667941163
transform 1 0 21504 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_388
timestamp 1667941163
transform 1 0 22400 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_392
timestamp 1667941163
transform 1 0 22624 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_417
timestamp 1667941163
transform 1 0 24024 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_443
timestamp 1667941163
transform 1 0 25480 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_459
timestamp 1667941163
transform 1 0 26376 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_463
timestamp 1667941163
transform 1 0 26600 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_488
timestamp 1667941163
transform 1 0 28000 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_514
timestamp 1667941163
transform 1 0 29456 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_530
timestamp 1667941163
transform 1 0 30352 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_534
timestamp 1667941163
transform 1 0 30576 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_559
timestamp 1667941163
transform 1 0 31976 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_585
timestamp 1667941163
transform 1 0 33432 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_601
timestamp 1667941163
transform 1 0 34328 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_605
timestamp 1667941163
transform 1 0 34552 0 1 10976
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_630
timestamp 1667941163
transform 1 0 35952 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_656
timestamp 1667941163
transform 1 0 37408 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_672
timestamp 1667941163
transform 1 0 38304 0 1 10976
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_676
timestamp 1667941163
transform 1 0 38528 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_684
timestamp 1667941163
transform 1 0 38976 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_2
timestamp 1667941163
transform 1 0 784 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_18
timestamp 1667941163
transform 1 0 1680 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_44
timestamp 1667941163
transform 1 0 3136 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1667941163
transform 1 0 4592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_73
timestamp 1667941163
transform 1 0 4760 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_89
timestamp 1667941163
transform 1 0 5656 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_115
timestamp 1667941163
transform 1 0 7112 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1667941163
transform 1 0 8568 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_144
timestamp 1667941163
transform 1 0 8736 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_160
timestamp 1667941163
transform 1 0 9632 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_186
timestamp 1667941163
transform 1 0 11088 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1667941163
transform 1 0 12544 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_215
timestamp 1667941163
transform 1 0 12712 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_231
timestamp 1667941163
transform 1 0 13608 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_257
timestamp 1667941163
transform 1 0 15064 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1667941163
transform 1 0 16520 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1667941163
transform 1 0 16688 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_311
timestamp 1667941163
transform 1 0 18088 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_337
timestamp 1667941163
transform 1 0 19544 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_353
timestamp 1667941163
transform 1 0 20440 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1667941163
transform 1 0 20664 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_382
timestamp 1667941163
transform 1 0 22064 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_408
timestamp 1667941163
transform 1 0 23520 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_424
timestamp 1667941163
transform 1 0 24416 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_428
timestamp 1667941163
transform 1 0 24640 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_453
timestamp 1667941163
transform 1 0 26040 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_479
timestamp 1667941163
transform 1 0 27496 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_495
timestamp 1667941163
transform 1 0 28392 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_499
timestamp 1667941163
transform 1 0 28616 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_524
timestamp 1667941163
transform 1 0 30016 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_550
timestamp 1667941163
transform 1 0 31472 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_566
timestamp 1667941163
transform 1 0 32368 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_570
timestamp 1667941163
transform 1 0 32592 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_595
timestamp 1667941163
transform 1 0 33992 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_627
timestamp 1667941163
transform 1 0 35784 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_635
timestamp 1667941163
transform 1 0 36232 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_641
timestamp 1667941163
transform 1 0 36568 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_673
timestamp 1667941163
transform 1 0 38360 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_681
timestamp 1667941163
transform 1 0 38808 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_685
timestamp 1667941163
transform 1 0 39032 0 -1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_687
timestamp 1667941163
transform 1 0 39144 0 -1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_2
timestamp 1667941163
transform 1 0 784 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1667941163
transform 1 0 2576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_37
timestamp 1667941163
transform 1 0 2744 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_53
timestamp 1667941163
transform 1 0 3640 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_79
timestamp 1667941163
transform 1 0 5096 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1667941163
transform 1 0 6552 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_108
timestamp 1667941163
transform 1 0 6720 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_124
timestamp 1667941163
transform 1 0 7616 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_150
timestamp 1667941163
transform 1 0 9072 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1667941163
transform 1 0 10528 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_179
timestamp 1667941163
transform 1 0 10696 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_195
timestamp 1667941163
transform 1 0 11592 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_221
timestamp 1667941163
transform 1 0 13048 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1667941163
transform 1 0 14504 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_250
timestamp 1667941163
transform 1 0 14672 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_258
timestamp 1667941163
transform 1 0 15120 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_262
timestamp 1667941163
transform 1 0 15344 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_264
timestamp 1667941163
transform 1 0 15456 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_289
timestamp 1667941163
transform 1 0 16856 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_315
timestamp 1667941163
transform 1 0 18312 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1667941163
transform 1 0 18648 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_346
timestamp 1667941163
transform 1 0 20048 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_372
timestamp 1667941163
transform 1 0 21504 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_388
timestamp 1667941163
transform 1 0 22400 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_392
timestamp 1667941163
transform 1 0 22624 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_417
timestamp 1667941163
transform 1 0 24024 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_443
timestamp 1667941163
transform 1 0 25480 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_459
timestamp 1667941163
transform 1 0 26376 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_463
timestamp 1667941163
transform 1 0 26600 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_488
timestamp 1667941163
transform 1 0 28000 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_514
timestamp 1667941163
transform 1 0 29456 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_530
timestamp 1667941163
transform 1 0 30352 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_534
timestamp 1667941163
transform 1 0 30576 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_559
timestamp 1667941163
transform 1 0 31976 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_585
timestamp 1667941163
transform 1 0 33432 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_601
timestamp 1667941163
transform 1 0 34328 0 1 11760
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 34552 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1667941163
transform 1 0 38136 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1667941163
transform 1 0 38360 0 1 11760
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_676
timestamp 1667941163
transform 1 0 38528 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_684
timestamp 1667941163
transform 1 0 38976 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_2
timestamp 1667941163
transform 1 0 784 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_18
timestamp 1667941163
transform 1 0 1680 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_44
timestamp 1667941163
transform 1 0 3136 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1667941163
transform 1 0 4592 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_73
timestamp 1667941163
transform 1 0 4760 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_89
timestamp 1667941163
transform 1 0 5656 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_115
timestamp 1667941163
transform 1 0 7112 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1667941163
transform 1 0 8568 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_144
timestamp 1667941163
transform 1 0 8736 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_160
timestamp 1667941163
transform 1 0 9632 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_186
timestamp 1667941163
transform 1 0 11088 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1667941163
transform 1 0 12544 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_215
timestamp 1667941163
transform 1 0 12712 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_231
timestamp 1667941163
transform 1 0 13608 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_257
timestamp 1667941163
transform 1 0 15064 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1667941163
transform 1 0 16520 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1667941163
transform 1 0 16688 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_311
timestamp 1667941163
transform 1 0 18088 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_337
timestamp 1667941163
transform 1 0 19544 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_353
timestamp 1667941163
transform 1 0 20440 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_357
timestamp 1667941163
transform 1 0 20664 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_382
timestamp 1667941163
transform 1 0 22064 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_408
timestamp 1667941163
transform 1 0 23520 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_424
timestamp 1667941163
transform 1 0 24416 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_428
timestamp 1667941163
transform 1 0 24640 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_453
timestamp 1667941163
transform 1 0 26040 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_479
timestamp 1667941163
transform 1 0 27496 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_495
timestamp 1667941163
transform 1 0 28392 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_499
timestamp 1667941163
transform 1 0 28616 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_524
timestamp 1667941163
transform 1 0 30016 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_550
timestamp 1667941163
transform 1 0 31472 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_566
timestamp 1667941163
transform 1 0 32368 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1667941163
transform 1 0 32592 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1667941163
transform 1 0 36176 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1667941163
transform 1 0 36400 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_641
timestamp 1667941163
transform 1 0 36568 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_673
timestamp 1667941163
transform 1 0 38360 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_681
timestamp 1667941163
transform 1 0 38808 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_685
timestamp 1667941163
transform 1 0 39032 0 -1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1667941163
transform 1 0 39144 0 -1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_2
timestamp 1667941163
transform 1 0 784 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1667941163
transform 1 0 2576 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_37
timestamp 1667941163
transform 1 0 2744 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_53
timestamp 1667941163
transform 1 0 3640 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_79
timestamp 1667941163
transform 1 0 5096 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1667941163
transform 1 0 6552 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_108
timestamp 1667941163
transform 1 0 6720 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_124
timestamp 1667941163
transform 1 0 7616 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_150
timestamp 1667941163
transform 1 0 9072 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1667941163
transform 1 0 10528 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_179
timestamp 1667941163
transform 1 0 10696 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_195
timestamp 1667941163
transform 1 0 11592 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_221
timestamp 1667941163
transform 1 0 13048 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1667941163
transform 1 0 14504 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_250
timestamp 1667941163
transform 1 0 14672 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_258
timestamp 1667941163
transform 1 0 15120 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_262
timestamp 1667941163
transform 1 0 15344 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_287
timestamp 1667941163
transform 1 0 16744 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_313
timestamp 1667941163
transform 1 0 18200 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_317
timestamp 1667941163
transform 1 0 18424 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1667941163
transform 1 0 18648 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_346
timestamp 1667941163
transform 1 0 20048 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_372
timestamp 1667941163
transform 1 0 21504 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_388
timestamp 1667941163
transform 1 0 22400 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1667941163
transform 1 0 22624 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_417
timestamp 1667941163
transform 1 0 24024 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_443
timestamp 1667941163
transform 1 0 25480 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_459
timestamp 1667941163
transform 1 0 26376 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_463
timestamp 1667941163
transform 1 0 26600 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_488
timestamp 1667941163
transform 1 0 28000 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_514
timestamp 1667941163
transform 1 0 29456 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_530
timestamp 1667941163
transform 1 0 30352 0 1 12544
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1667941163
transform 1 0 30576 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1667941163
transform 1 0 34160 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1667941163
transform 1 0 34384 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1667941163
transform 1 0 34552 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1667941163
transform 1 0 38136 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1667941163
transform 1 0 38360 0 1 12544
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_676
timestamp 1667941163
transform 1 0 38528 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_684
timestamp 1667941163
transform 1 0 38976 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_2
timestamp 1667941163
transform 1 0 784 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_18
timestamp 1667941163
transform 1 0 1680 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_44
timestamp 1667941163
transform 1 0 3136 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1667941163
transform 1 0 4592 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_73
timestamp 1667941163
transform 1 0 4760 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_89
timestamp 1667941163
transform 1 0 5656 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_115
timestamp 1667941163
transform 1 0 7112 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1667941163
transform 1 0 8568 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_144
timestamp 1667941163
transform 1 0 8736 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_160
timestamp 1667941163
transform 1 0 9632 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_186
timestamp 1667941163
transform 1 0 11088 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1667941163
transform 1 0 12544 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_215
timestamp 1667941163
transform 1 0 12712 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_223
timestamp 1667941163
transform 1 0 13160 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_225
timestamp 1667941163
transform 1 0 13272 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_250
timestamp 1667941163
transform 1 0 14672 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_276
timestamp 1667941163
transform 1 0 16128 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1667941163
transform 1 0 16688 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_311
timestamp 1667941163
transform 1 0 18088 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_337
timestamp 1667941163
transform 1 0 19544 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_353
timestamp 1667941163
transform 1 0 20440 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1667941163
transform 1 0 20664 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_382
timestamp 1667941163
transform 1 0 22064 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_408
timestamp 1667941163
transform 1 0 23520 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_424
timestamp 1667941163
transform 1 0 24416 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_428
timestamp 1667941163
transform 1 0 24640 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_453
timestamp 1667941163
transform 1 0 26040 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_479
timestamp 1667941163
transform 1 0 27496 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_495
timestamp 1667941163
transform 1 0 28392 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_499
timestamp 1667941163
transform 1 0 28616 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_524
timestamp 1667941163
transform 1 0 30016 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_556
timestamp 1667941163
transform 1 0 31808 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_564
timestamp 1667941163
transform 1 0 32256 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1667941163
transform 1 0 32592 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1667941163
transform 1 0 36176 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1667941163
transform 1 0 36400 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_641
timestamp 1667941163
transform 1 0 36568 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_673
timestamp 1667941163
transform 1 0 38360 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_681
timestamp 1667941163
transform 1 0 38808 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_685
timestamp 1667941163
transform 1 0 39032 0 -1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1667941163
transform 1 0 39144 0 -1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_2
timestamp 1667941163
transform 1 0 784 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1667941163
transform 1 0 2576 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_37
timestamp 1667941163
transform 1 0 2744 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_53
timestamp 1667941163
transform 1 0 3640 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_79
timestamp 1667941163
transform 1 0 5096 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1667941163
transform 1 0 6552 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_108
timestamp 1667941163
transform 1 0 6720 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_124
timestamp 1667941163
transform 1 0 7616 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_150
timestamp 1667941163
transform 1 0 9072 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1667941163
transform 1 0 10528 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_179
timestamp 1667941163
transform 1 0 10696 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_195
timestamp 1667941163
transform 1 0 11592 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_221
timestamp 1667941163
transform 1 0 13048 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1667941163
transform 1 0 14504 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_250
timestamp 1667941163
transform 1 0 14672 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_258
timestamp 1667941163
transform 1 0 15120 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_284
timestamp 1667941163
transform 1 0 16576 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_310
timestamp 1667941163
transform 1 0 18032 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1667941163
transform 1 0 18480 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1667941163
transform 1 0 18648 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_346
timestamp 1667941163
transform 1 0 20048 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_372
timestamp 1667941163
transform 1 0 21504 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_388
timestamp 1667941163
transform 1 0 22400 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_392
timestamp 1667941163
transform 1 0 22624 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_417
timestamp 1667941163
transform 1 0 24024 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_443
timestamp 1667941163
transform 1 0 25480 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_459
timestamp 1667941163
transform 1 0 26376 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_463
timestamp 1667941163
transform 1 0 26600 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_488
timestamp 1667941163
transform 1 0 28000 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_514
timestamp 1667941163
transform 1 0 29456 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_530
timestamp 1667941163
transform 1 0 30352 0 1 13328
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1667941163
transform 1 0 30576 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1667941163
transform 1 0 34160 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1667941163
transform 1 0 34384 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1667941163
transform 1 0 34552 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1667941163
transform 1 0 38136 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1667941163
transform 1 0 38360 0 1 13328
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_676
timestamp 1667941163
transform 1 0 38528 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_684
timestamp 1667941163
transform 1 0 38976 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_2
timestamp 1667941163
transform 1 0 784 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_18
timestamp 1667941163
transform 1 0 1680 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_44
timestamp 1667941163
transform 1 0 3136 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1667941163
transform 1 0 4592 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_73
timestamp 1667941163
transform 1 0 4760 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_89
timestamp 1667941163
transform 1 0 5656 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_115
timestamp 1667941163
transform 1 0 7112 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1667941163
transform 1 0 8568 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_144
timestamp 1667941163
transform 1 0 8736 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_160
timestamp 1667941163
transform 1 0 9632 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_186
timestamp 1667941163
transform 1 0 11088 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1667941163
transform 1 0 12544 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_215
timestamp 1667941163
transform 1 0 12712 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_231
timestamp 1667941163
transform 1 0 13608 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_256
timestamp 1667941163
transform 1 0 15008 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_282
timestamp 1667941163
transform 1 0 16464 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_286
timestamp 1667941163
transform 1 0 16688 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_311
timestamp 1667941163
transform 1 0 18088 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_337
timestamp 1667941163
transform 1 0 19544 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_353
timestamp 1667941163
transform 1 0 20440 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1667941163
transform 1 0 20664 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_382
timestamp 1667941163
transform 1 0 22064 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_408
timestamp 1667941163
transform 1 0 23520 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_424
timestamp 1667941163
transform 1 0 24416 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1667941163
transform 1 0 24640 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_453
timestamp 1667941163
transform 1 0 26040 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_479
timestamp 1667941163
transform 1 0 27496 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_495
timestamp 1667941163
transform 1 0 28392 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1667941163
transform 1 0 28616 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1667941163
transform 1 0 32200 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1667941163
transform 1 0 32424 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1667941163
transform 1 0 32592 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1667941163
transform 1 0 36176 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1667941163
transform 1 0 36400 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_641
timestamp 1667941163
transform 1 0 36568 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_673
timestamp 1667941163
transform 1 0 38360 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_681
timestamp 1667941163
transform 1 0 38808 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_685
timestamp 1667941163
transform 1 0 39032 0 -1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1667941163
transform 1 0 39144 0 -1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_2
timestamp 1667941163
transform 1 0 784 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1667941163
transform 1 0 2576 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_37
timestamp 1667941163
transform 1 0 2744 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_53
timestamp 1667941163
transform 1 0 3640 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_79
timestamp 1667941163
transform 1 0 5096 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1667941163
transform 1 0 6552 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_108
timestamp 1667941163
transform 1 0 6720 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_124
timestamp 1667941163
transform 1 0 7616 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_150
timestamp 1667941163
transform 1 0 9072 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1667941163
transform 1 0 10528 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_179
timestamp 1667941163
transform 1 0 10696 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_195
timestamp 1667941163
transform 1 0 11592 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_221
timestamp 1667941163
transform 1 0 13048 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1667941163
transform 1 0 14504 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1667941163
transform 1 0 14672 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_275
timestamp 1667941163
transform 1 0 16072 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_301
timestamp 1667941163
transform 1 0 17528 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1667941163
transform 1 0 18424 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1667941163
transform 1 0 18648 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_346
timestamp 1667941163
transform 1 0 20048 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_372
timestamp 1667941163
transform 1 0 21504 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_388
timestamp 1667941163
transform 1 0 22400 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1667941163
transform 1 0 22624 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_417
timestamp 1667941163
transform 1 0 24024 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_443
timestamp 1667941163
transform 1 0 25480 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_459
timestamp 1667941163
transform 1 0 26376 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_463
timestamp 1667941163
transform 1 0 26600 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_488
timestamp 1667941163
transform 1 0 28000 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_514
timestamp 1667941163
transform 1 0 29456 0 1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_530
timestamp 1667941163
transform 1 0 30352 0 1 14112
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1667941163
transform 1 0 30576 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1667941163
transform 1 0 34160 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1667941163
transform 1 0 34384 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1667941163
transform 1 0 34552 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1667941163
transform 1 0 38136 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1667941163
transform 1 0 38360 0 1 14112
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_676
timestamp 1667941163
transform 1 0 38528 0 1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_684
timestamp 1667941163
transform 1 0 38976 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_2
timestamp 1667941163
transform 1 0 784 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_18
timestamp 1667941163
transform 1 0 1680 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_44
timestamp 1667941163
transform 1 0 3136 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1667941163
transform 1 0 4592 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_73
timestamp 1667941163
transform 1 0 4760 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_89
timestamp 1667941163
transform 1 0 5656 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_115
timestamp 1667941163
transform 1 0 7112 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1667941163
transform 1 0 8568 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_144
timestamp 1667941163
transform 1 0 8736 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_160
timestamp 1667941163
transform 1 0 9632 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_186
timestamp 1667941163
transform 1 0 11088 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1667941163
transform 1 0 12544 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_215
timestamp 1667941163
transform 1 0 12712 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_231
timestamp 1667941163
transform 1 0 13608 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_256
timestamp 1667941163
transform 1 0 15008 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_282
timestamp 1667941163
transform 1 0 16464 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1667941163
transform 1 0 16688 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_311
timestamp 1667941163
transform 1 0 18088 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_337
timestamp 1667941163
transform 1 0 19544 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_353
timestamp 1667941163
transform 1 0 20440 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1667941163
transform 1 0 20664 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_382
timestamp 1667941163
transform 1 0 22064 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_408
timestamp 1667941163
transform 1 0 23520 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_424
timestamp 1667941163
transform 1 0 24416 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_428
timestamp 1667941163
transform 1 0 24640 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_453
timestamp 1667941163
transform 1 0 26040 0 -1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_485
timestamp 1667941163
transform 1 0 27832 0 -1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_493
timestamp 1667941163
transform 1 0 28280 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1667941163
transform 1 0 28616 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1667941163
transform 1 0 32200 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1667941163
transform 1 0 32424 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1667941163
transform 1 0 32592 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1667941163
transform 1 0 36176 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1667941163
transform 1 0 36400 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_641
timestamp 1667941163
transform 1 0 36568 0 -1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_673
timestamp 1667941163
transform 1 0 38360 0 -1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_681
timestamp 1667941163
transform 1 0 38808 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_685
timestamp 1667941163
transform 1 0 39032 0 -1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_687
timestamp 1667941163
transform 1 0 39144 0 -1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_2
timestamp 1667941163
transform 1 0 784 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1667941163
transform 1 0 2576 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_37
timestamp 1667941163
transform 1 0 2744 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_53
timestamp 1667941163
transform 1 0 3640 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_79
timestamp 1667941163
transform 1 0 5096 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1667941163
transform 1 0 6552 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_108
timestamp 1667941163
transform 1 0 6720 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_124
timestamp 1667941163
transform 1 0 7616 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_150
timestamp 1667941163
transform 1 0 9072 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1667941163
transform 1 0 10528 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_179
timestamp 1667941163
transform 1 0 10696 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_195
timestamp 1667941163
transform 1 0 11592 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_221
timestamp 1667941163
transform 1 0 13048 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1667941163
transform 1 0 14504 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1667941163
transform 1 0 14672 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_275
timestamp 1667941163
transform 1 0 16072 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_301
timestamp 1667941163
transform 1 0 17528 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_317
timestamp 1667941163
transform 1 0 18424 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1667941163
transform 1 0 18648 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_346
timestamp 1667941163
transform 1 0 20048 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_372
timestamp 1667941163
transform 1 0 21504 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_388
timestamp 1667941163
transform 1 0 22400 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_392
timestamp 1667941163
transform 1 0 22624 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_417
timestamp 1667941163
transform 1 0 24024 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_443
timestamp 1667941163
transform 1 0 25480 0 1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_459
timestamp 1667941163
transform 1 0 26376 0 1 14896
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1667941163
transform 1 0 26600 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1667941163
transform 1 0 30184 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1667941163
transform 1 0 30408 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1667941163
transform 1 0 30576 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1667941163
transform 1 0 34160 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1667941163
transform 1 0 34384 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1667941163
transform 1 0 34552 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1667941163
transform 1 0 38136 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1667941163
transform 1 0 38360 0 1 14896
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_676
timestamp 1667941163
transform 1 0 38528 0 1 14896
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_684
timestamp 1667941163
transform 1 0 38976 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_2
timestamp 1667941163
transform 1 0 784 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_18
timestamp 1667941163
transform 1 0 1680 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_44
timestamp 1667941163
transform 1 0 3136 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1667941163
transform 1 0 4592 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_73
timestamp 1667941163
transform 1 0 4760 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_89
timestamp 1667941163
transform 1 0 5656 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_115
timestamp 1667941163
transform 1 0 7112 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1667941163
transform 1 0 8568 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_144
timestamp 1667941163
transform 1 0 8736 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_160
timestamp 1667941163
transform 1 0 9632 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_186
timestamp 1667941163
transform 1 0 11088 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1667941163
transform 1 0 12544 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_215
timestamp 1667941163
transform 1 0 12712 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_231
timestamp 1667941163
transform 1 0 13608 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_256
timestamp 1667941163
transform 1 0 15008 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1667941163
transform 1 0 16464 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_286
timestamp 1667941163
transform 1 0 16688 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_311
timestamp 1667941163
transform 1 0 18088 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_337
timestamp 1667941163
transform 1 0 19544 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_353
timestamp 1667941163
transform 1 0 20440 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1667941163
transform 1 0 20664 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_382
timestamp 1667941163
transform 1 0 22064 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_408
timestamp 1667941163
transform 1 0 23520 0 -1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_424
timestamp 1667941163
transform 1 0 24416 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1667941163
transform 1 0 24640 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1667941163
transform 1 0 28224 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1667941163
transform 1 0 28448 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1667941163
transform 1 0 28616 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1667941163
transform 1 0 32200 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1667941163
transform 1 0 32424 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1667941163
transform 1 0 32592 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1667941163
transform 1 0 36176 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1667941163
transform 1 0 36400 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_641
timestamp 1667941163
transform 1 0 36568 0 -1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_673
timestamp 1667941163
transform 1 0 38360 0 -1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_681
timestamp 1667941163
transform 1 0 38808 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_685
timestamp 1667941163
transform 1 0 39032 0 -1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1667941163
transform 1 0 39144 0 -1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1667941163
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1667941163
transform 1 0 2576 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1667941163
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1667941163
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1667941163
transform 1 0 6552 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_108
timestamp 1667941163
transform 1 0 6720 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_124
timestamp 1667941163
transform 1 0 7616 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_150
timestamp 1667941163
transform 1 0 9072 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1667941163
transform 1 0 10528 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_179
timestamp 1667941163
transform 1 0 10696 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_195
timestamp 1667941163
transform 1 0 11592 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_221
timestamp 1667941163
transform 1 0 13048 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1667941163
transform 1 0 14504 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_250
timestamp 1667941163
transform 1 0 14672 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_275
timestamp 1667941163
transform 1 0 16072 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_301
timestamp 1667941163
transform 1 0 17528 0 1 15680
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_317
timestamp 1667941163
transform 1 0 18424 0 1 15680
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1667941163
transform 1 0 18648 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_346
timestamp 1667941163
transform 1 0 20048 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_378
timestamp 1667941163
transform 1 0 21840 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_386
timestamp 1667941163
transform 1 0 22288 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1667941163
transform 1 0 22624 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1667941163
transform 1 0 26208 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1667941163
transform 1 0 26432 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1667941163
transform 1 0 26600 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1667941163
transform 1 0 30184 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1667941163
transform 1 0 30408 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1667941163
transform 1 0 30576 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1667941163
transform 1 0 34160 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1667941163
transform 1 0 34384 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1667941163
transform 1 0 34552 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1667941163
transform 1 0 38136 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1667941163
transform 1 0 38360 0 1 15680
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_676
timestamp 1667941163
transform 1 0 38528 0 1 15680
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_684
timestamp 1667941163
transform 1 0 38976 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1667941163
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1667941163
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1667941163
transform 1 0 4592 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1667941163
transform 1 0 4760 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1667941163
transform 1 0 8344 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1667941163
transform 1 0 8568 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_144
timestamp 1667941163
transform 1 0 8736 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_160
timestamp 1667941163
transform 1 0 9632 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_186
timestamp 1667941163
transform 1 0 11088 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1667941163
transform 1 0 12544 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_215
timestamp 1667941163
transform 1 0 12712 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_255
timestamp 1667941163
transform 1 0 14952 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 16408 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1667941163
transform 1 0 16520 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1667941163
transform 1 0 16688 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_311
timestamp 1667941163
transform 1 0 18088 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_337
timestamp 1667941163
transform 1 0 19544 0 -1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_353
timestamp 1667941163
transform 1 0 20440 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1667941163
transform 1 0 20664 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1667941163
transform 1 0 24248 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1667941163
transform 1 0 24472 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1667941163
transform 1 0 24640 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1667941163
transform 1 0 28224 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1667941163
transform 1 0 28448 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1667941163
transform 1 0 28616 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1667941163
transform 1 0 32200 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1667941163
transform 1 0 32424 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1667941163
transform 1 0 32592 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1667941163
transform 1 0 36176 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1667941163
transform 1 0 36400 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_641
timestamp 1667941163
transform 1 0 36568 0 -1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_673
timestamp 1667941163
transform 1 0 38360 0 -1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_681
timestamp 1667941163
transform 1 0 38808 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_685
timestamp 1667941163
transform 1 0 39032 0 -1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_687
timestamp 1667941163
transform 1 0 39144 0 -1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1667941163
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1667941163
transform 1 0 2576 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1667941163
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1667941163
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1667941163
transform 1 0 6552 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_108
timestamp 1667941163
transform 1 0 6720 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_124
timestamp 1667941163
transform 1 0 7616 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_150
timestamp 1667941163
transform 1 0 9072 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1667941163
transform 1 0 10528 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_179
timestamp 1667941163
transform 1 0 10696 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_195
timestamp 1667941163
transform 1 0 11592 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_221
timestamp 1667941163
transform 1 0 13048 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1667941163
transform 1 0 14504 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1667941163
transform 1 0 14672 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_275
timestamp 1667941163
transform 1 0 16072 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_301
timestamp 1667941163
transform 1 0 17528 0 1 16464
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_317
timestamp 1667941163
transform 1 0 18424 0 1 16464
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1667941163
transform 1 0 18648 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1667941163
transform 1 0 22232 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1667941163
transform 1 0 22456 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1667941163
transform 1 0 22624 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1667941163
transform 1 0 26208 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1667941163
transform 1 0 26432 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1667941163
transform 1 0 26600 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1667941163
transform 1 0 30184 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1667941163
transform 1 0 30408 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1667941163
transform 1 0 30576 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1667941163
transform 1 0 34160 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1667941163
transform 1 0 34384 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1667941163
transform 1 0 34552 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1667941163
transform 1 0 38136 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1667941163
transform 1 0 38360 0 1 16464
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_676
timestamp 1667941163
transform 1 0 38528 0 1 16464
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_684
timestamp 1667941163
transform 1 0 38976 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1667941163
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1667941163
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1667941163
transform 1 0 4592 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1667941163
transform 1 0 4760 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1667941163
transform 1 0 8344 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1667941163
transform 1 0 8568 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_144
timestamp 1667941163
transform 1 0 8736 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_160
timestamp 1667941163
transform 1 0 9632 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_186
timestamp 1667941163
transform 1 0 11088 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1667941163
transform 1 0 12544 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_215
timestamp 1667941163
transform 1 0 12712 0 -1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_231
timestamp 1667941163
transform 1 0 13608 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_256
timestamp 1667941163
transform 1 0 15008 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_282
timestamp 1667941163
transform 1 0 16464 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1667941163
transform 1 0 16688 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_311
timestamp 1667941163
transform 1 0 18088 0 -1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_343
timestamp 1667941163
transform 1 0 19880 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_351
timestamp 1667941163
transform 1 0 20328 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1667941163
transform 1 0 20664 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1667941163
transform 1 0 24248 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1667941163
transform 1 0 24472 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1667941163
transform 1 0 24640 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1667941163
transform 1 0 28224 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1667941163
transform 1 0 28448 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1667941163
transform 1 0 28616 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1667941163
transform 1 0 32200 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1667941163
transform 1 0 32424 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1667941163
transform 1 0 32592 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1667941163
transform 1 0 36176 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1667941163
transform 1 0 36400 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_641
timestamp 1667941163
transform 1 0 36568 0 -1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_673
timestamp 1667941163
transform 1 0 38360 0 -1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_681
timestamp 1667941163
transform 1 0 38808 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_685
timestamp 1667941163
transform 1 0 39032 0 -1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_687
timestamp 1667941163
transform 1 0 39144 0 -1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1667941163
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1667941163
transform 1 0 2576 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1667941163
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1667941163
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1667941163
transform 1 0 6552 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_108
timestamp 1667941163
transform 1 0 6720 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_140
timestamp 1667941163
transform 1 0 8512 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_148
timestamp 1667941163
transform 1 0 8960 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1667941163
transform 1 0 10528 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_179
timestamp 1667941163
transform 1 0 10696 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_195
timestamp 1667941163
transform 1 0 11592 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_221
timestamp 1667941163
transform 1 0 13048 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1667941163
transform 1 0 14504 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1667941163
transform 1 0 14672 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_275
timestamp 1667941163
transform 1 0 16072 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_301
timestamp 1667941163
transform 1 0 17528 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_317
timestamp 1667941163
transform 1 0 18424 0 1 17248
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1667941163
transform 1 0 18648 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1667941163
transform 1 0 22232 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1667941163
transform 1 0 22456 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1667941163
transform 1 0 22624 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1667941163
transform 1 0 26208 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1667941163
transform 1 0 26432 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1667941163
transform 1 0 26600 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1667941163
transform 1 0 30184 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1667941163
transform 1 0 30408 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1667941163
transform 1 0 30576 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1667941163
transform 1 0 34160 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1667941163
transform 1 0 34384 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1667941163
transform 1 0 34552 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1667941163
transform 1 0 38136 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1667941163
transform 1 0 38360 0 1 17248
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_676
timestamp 1667941163
transform 1 0 38528 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_684
timestamp 1667941163
transform 1 0 38976 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1667941163
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1667941163
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1667941163
transform 1 0 4592 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1667941163
transform 1 0 4760 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1667941163
transform 1 0 8344 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1667941163
transform 1 0 8568 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_144
timestamp 1667941163
transform 1 0 8736 0 -1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_160
timestamp 1667941163
transform 1 0 9632 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_186
timestamp 1667941163
transform 1 0 11088 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1667941163
transform 1 0 12544 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_215
timestamp 1667941163
transform 1 0 12712 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_223
timestamp 1667941163
transform 1 0 13160 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_225
timestamp 1667941163
transform 1 0 13272 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_250
timestamp 1667941163
transform 1 0 14672 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_276
timestamp 1667941163
transform 1 0 16128 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1667941163
transform 1 0 16688 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1667941163
transform 1 0 20272 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1667941163
transform 1 0 20496 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1667941163
transform 1 0 20664 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1667941163
transform 1 0 24248 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1667941163
transform 1 0 24472 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1667941163
transform 1 0 24640 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1667941163
transform 1 0 28224 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1667941163
transform 1 0 28448 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1667941163
transform 1 0 28616 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1667941163
transform 1 0 32200 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1667941163
transform 1 0 32424 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1667941163
transform 1 0 32592 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1667941163
transform 1 0 36176 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1667941163
transform 1 0 36400 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_641
timestamp 1667941163
transform 1 0 36568 0 -1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_673
timestamp 1667941163
transform 1 0 38360 0 -1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_681
timestamp 1667941163
transform 1 0 38808 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_685
timestamp 1667941163
transform 1 0 39032 0 -1 18032
box 0 -30 112 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_687
timestamp 1667941163
transform 1 0 39144 0 -1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1667941163
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1667941163
transform 1 0 2576 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_37
timestamp 1667941163
transform 1 0 2744 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_69
timestamp 1667941163
transform 1 0 4536 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_72
timestamp 1667941163
transform 1 0 4704 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1667941163
transform 1 0 6496 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_107
timestamp 1667941163
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 8456 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_142
timestamp 1667941163
transform 1 0 8624 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1667941163
transform 1 0 10416 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_177
timestamp 1667941163
transform 1 0 10584 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1667941163
transform 1 0 12376 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_212
timestamp 1667941163
transform 1 0 12544 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1667941163
transform 1 0 14336 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1667941163
transform 1 0 14504 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_272
timestamp 1667941163
transform 1 0 15904 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_282
timestamp 1667941163
transform 1 0 16464 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1667941163
transform 1 0 18256 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_317
timestamp 1667941163
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_349
timestamp 1667941163
transform 1 0 20216 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_352
timestamp 1667941163
transform 1 0 20384 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1667941163
transform 1 0 22176 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_387
timestamp 1667941163
transform 1 0 22344 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1667941163
transform 1 0 24136 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_422
timestamp 1667941163
transform 1 0 24304 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1667941163
transform 1 0 26096 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_457
timestamp 1667941163
transform 1 0 26264 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_489
timestamp 1667941163
transform 1 0 28056 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_492
timestamp 1667941163
transform 1 0 28224 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1667941163
transform 1 0 30016 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_527
timestamp 1667941163
transform 1 0 30184 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_559
timestamp 1667941163
transform 1 0 31976 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_562
timestamp 1667941163
transform 1 0 32144 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_594
timestamp 1667941163
transform 1 0 33936 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_597
timestamp 1667941163
transform 1 0 34104 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_629
timestamp 1667941163
transform 1 0 35896 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_632
timestamp 1667941163
transform 1 0 36064 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1667941163
transform 1 0 37856 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_667
timestamp 1667941163
transform 1 0 38024 0 1 18032
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_683
timestamp 1667941163
transform 1 0 38920 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_687
timestamp 1667941163
transform 1 0 39144 0 1 18032
box 0 -30 56 422
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1667941163
transform -1 0 39312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1667941163
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1667941163
transform -1 0 39312 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1667941163
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1667941163
transform -1 0 39312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1667941163
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1667941163
transform -1 0 39312 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1667941163
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1667941163
transform -1 0 39312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1667941163
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1667941163
transform -1 0 39312 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1667941163
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1667941163
transform -1 0 39312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1667941163
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1667941163
transform -1 0 39312 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1667941163
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1667941163
transform -1 0 39312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1667941163
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1667941163
transform -1 0 39312 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1667941163
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1667941163
transform -1 0 39312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1667941163
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1667941163
transform -1 0 39312 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1667941163
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1667941163
transform -1 0 39312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1667941163
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1667941163
transform -1 0 39312 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1667941163
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1667941163
transform -1 0 39312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1667941163
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1667941163
transform -1 0 39312 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1667941163
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1667941163
transform -1 0 39312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1667941163
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1667941163
transform -1 0 39312 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1667941163
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1667941163
transform -1 0 39312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1667941163
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1667941163
transform -1 0 39312 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1667941163
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1667941163
transform -1 0 39312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1667941163
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1667941163
transform -1 0 39312 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1667941163
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1667941163
transform -1 0 39312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1667941163
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1667941163
transform -1 0 39312 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1667941163
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1667941163
transform -1 0 39312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1667941163
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1667941163
transform -1 0 39312 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1667941163
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1667941163
transform -1 0 39312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1667941163
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1667941163
transform -1 0 39312 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1667941163
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1667941163
transform -1 0 39312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1667941163
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1667941163
transform -1 0 39312 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1667941163
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1667941163
transform -1 0 39312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1667941163
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1667941163
transform -1 0 39312 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1667941163
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1667941163
transform -1 0 39312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1667941163
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1667941163
transform -1 0 39312 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1667941163
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1667941163
transform -1 0 39312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1667941163
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1667941163
transform -1 0 39312 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1667941163
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1667941163
transform -1 0 39312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1667941163
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1667941163
transform -1 0 39312 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1667941163
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1667941163
transform -1 0 39312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1667941163
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1667941163
transform -1 0 39312 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1667941163
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1667941163
transform -1 0 39312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1667941163
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1667941163
transform -1 0 39312 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1667941163
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1667941163
transform -1 0 39312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform 1 0 2632 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1667941163
transform 1 0 4592 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1667941163
transform 1 0 6552 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1667941163
transform 1 0 8512 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1667941163
transform 1 0 10472 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1667941163
transform 1 0 12432 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1667941163
transform 1 0 14392 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1667941163
transform 1 0 16352 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1667941163
transform 1 0 18312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1667941163
transform 1 0 20272 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1667941163
transform 1 0 22232 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1667941163
transform 1 0 24192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1667941163
transform 1 0 26152 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1667941163
transform 1 0 28112 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1667941163
transform 1 0 30072 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1667941163
transform 1 0 32032 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1667941163
transform 1 0 33992 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1667941163
transform 1 0 35952 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1667941163
transform 1 0 37912 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1667941163
transform 1 0 4648 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1667941163
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1667941163
transform 1 0 12600 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1667941163
transform 1 0 16576 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1667941163
transform 1 0 20552 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1667941163
transform 1 0 24528 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1667941163
transform 1 0 28504 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1667941163
transform 1 0 32480 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1667941163
transform 1 0 36456 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1667941163
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1667941163
transform 1 0 6608 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1667941163
transform 1 0 10584 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1667941163
transform 1 0 14560 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1667941163
transform 1 0 18536 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1667941163
transform 1 0 22512 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1667941163
transform 1 0 26488 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1667941163
transform 1 0 30464 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1667941163
transform 1 0 34440 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1667941163
transform 1 0 38416 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1667941163
transform 1 0 4648 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1667941163
transform 1 0 8624 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1667941163
transform 1 0 12600 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1667941163
transform 1 0 16576 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1667941163
transform 1 0 20552 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1667941163
transform 1 0 24528 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1667941163
transform 1 0 28504 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1667941163
transform 1 0 32480 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1667941163
transform 1 0 36456 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1667941163
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1667941163
transform 1 0 6608 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1667941163
transform 1 0 10584 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1667941163
transform 1 0 14560 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1667941163
transform 1 0 18536 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1667941163
transform 1 0 22512 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1667941163
transform 1 0 26488 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1667941163
transform 1 0 30464 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1667941163
transform 1 0 34440 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1667941163
transform 1 0 38416 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1667941163
transform 1 0 4648 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1667941163
transform 1 0 8624 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1667941163
transform 1 0 12600 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1667941163
transform 1 0 16576 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1667941163
transform 1 0 20552 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1667941163
transform 1 0 24528 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1667941163
transform 1 0 28504 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1667941163
transform 1 0 32480 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1667941163
transform 1 0 36456 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1667941163
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1667941163
transform 1 0 6608 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1667941163
transform 1 0 10584 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1667941163
transform 1 0 14560 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1667941163
transform 1 0 18536 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1667941163
transform 1 0 22512 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1667941163
transform 1 0 26488 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1667941163
transform 1 0 30464 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1667941163
transform 1 0 34440 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1667941163
transform 1 0 38416 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1667941163
transform 1 0 4648 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1667941163
transform 1 0 8624 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1667941163
transform 1 0 12600 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1667941163
transform 1 0 16576 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1667941163
transform 1 0 20552 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1667941163
transform 1 0 24528 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1667941163
transform 1 0 28504 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1667941163
transform 1 0 32480 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1667941163
transform 1 0 36456 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1667941163
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1667941163
transform 1 0 6608 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1667941163
transform 1 0 10584 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1667941163
transform 1 0 14560 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1667941163
transform 1 0 18536 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1667941163
transform 1 0 22512 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1667941163
transform 1 0 26488 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1667941163
transform 1 0 30464 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1667941163
transform 1 0 34440 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1667941163
transform 1 0 38416 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1667941163
transform 1 0 4648 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1667941163
transform 1 0 8624 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1667941163
transform 1 0 12600 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1667941163
transform 1 0 16576 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1667941163
transform 1 0 20552 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1667941163
transform 1 0 24528 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1667941163
transform 1 0 28504 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1667941163
transform 1 0 32480 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1667941163
transform 1 0 36456 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1667941163
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1667941163
transform 1 0 6608 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1667941163
transform 1 0 10584 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1667941163
transform 1 0 14560 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1667941163
transform 1 0 18536 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1667941163
transform 1 0 22512 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1667941163
transform 1 0 26488 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1667941163
transform 1 0 30464 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1667941163
transform 1 0 34440 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1667941163
transform 1 0 38416 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1667941163
transform 1 0 4648 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1667941163
transform 1 0 8624 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1667941163
transform 1 0 12600 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1667941163
transform 1 0 16576 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1667941163
transform 1 0 20552 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1667941163
transform 1 0 24528 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1667941163
transform 1 0 28504 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1667941163
transform 1 0 32480 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1667941163
transform 1 0 36456 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1667941163
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1667941163
transform 1 0 6608 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1667941163
transform 1 0 10584 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1667941163
transform 1 0 14560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1667941163
transform 1 0 18536 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1667941163
transform 1 0 22512 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1667941163
transform 1 0 26488 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1667941163
transform 1 0 30464 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1667941163
transform 1 0 34440 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1667941163
transform 1 0 38416 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1667941163
transform 1 0 4648 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1667941163
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1667941163
transform 1 0 12600 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1667941163
transform 1 0 16576 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1667941163
transform 1 0 20552 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1667941163
transform 1 0 24528 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1667941163
transform 1 0 28504 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1667941163
transform 1 0 32480 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1667941163
transform 1 0 36456 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1667941163
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1667941163
transform 1 0 6608 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1667941163
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1667941163
transform 1 0 14560 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1667941163
transform 1 0 18536 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1667941163
transform 1 0 22512 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1667941163
transform 1 0 26488 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1667941163
transform 1 0 30464 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1667941163
transform 1 0 34440 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1667941163
transform 1 0 38416 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1667941163
transform 1 0 4648 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1667941163
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1667941163
transform 1 0 12600 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1667941163
transform 1 0 16576 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1667941163
transform 1 0 20552 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1667941163
transform 1 0 24528 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1667941163
transform 1 0 28504 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1667941163
transform 1 0 32480 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1667941163
transform 1 0 36456 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1667941163
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1667941163
transform 1 0 6608 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1667941163
transform 1 0 10584 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1667941163
transform 1 0 14560 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1667941163
transform 1 0 18536 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1667941163
transform 1 0 22512 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1667941163
transform 1 0 26488 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1667941163
transform 1 0 30464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1667941163
transform 1 0 34440 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1667941163
transform 1 0 38416 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1667941163
transform 1 0 4648 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1667941163
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1667941163
transform 1 0 12600 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1667941163
transform 1 0 16576 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1667941163
transform 1 0 20552 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1667941163
transform 1 0 24528 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1667941163
transform 1 0 28504 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1667941163
transform 1 0 32480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1667941163
transform 1 0 36456 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1667941163
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1667941163
transform 1 0 6608 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1667941163
transform 1 0 10584 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1667941163
transform 1 0 14560 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1667941163
transform 1 0 18536 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1667941163
transform 1 0 22512 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1667941163
transform 1 0 26488 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1667941163
transform 1 0 30464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1667941163
transform 1 0 34440 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1667941163
transform 1 0 38416 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1667941163
transform 1 0 4648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1667941163
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1667941163
transform 1 0 12600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1667941163
transform 1 0 16576 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1667941163
transform 1 0 20552 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1667941163
transform 1 0 24528 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1667941163
transform 1 0 28504 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1667941163
transform 1 0 32480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1667941163
transform 1 0 36456 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1667941163
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1667941163
transform 1 0 6608 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1667941163
transform 1 0 10584 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1667941163
transform 1 0 14560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1667941163
transform 1 0 18536 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1667941163
transform 1 0 22512 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1667941163
transform 1 0 26488 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1667941163
transform 1 0 30464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1667941163
transform 1 0 34440 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1667941163
transform 1 0 38416 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1667941163
transform 1 0 4648 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1667941163
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1667941163
transform 1 0 12600 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1667941163
transform 1 0 16576 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1667941163
transform 1 0 20552 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1667941163
transform 1 0 24528 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1667941163
transform 1 0 28504 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1667941163
transform 1 0 32480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1667941163
transform 1 0 36456 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1667941163
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1667941163
transform 1 0 6608 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1667941163
transform 1 0 10584 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1667941163
transform 1 0 14560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1667941163
transform 1 0 18536 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1667941163
transform 1 0 22512 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1667941163
transform 1 0 26488 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1667941163
transform 1 0 30464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1667941163
transform 1 0 34440 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1667941163
transform 1 0 38416 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1667941163
transform 1 0 4648 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1667941163
transform 1 0 8624 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1667941163
transform 1 0 12600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1667941163
transform 1 0 16576 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1667941163
transform 1 0 20552 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1667941163
transform 1 0 24528 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1667941163
transform 1 0 28504 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1667941163
transform 1 0 32480 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1667941163
transform 1 0 36456 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1667941163
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1667941163
transform 1 0 6608 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1667941163
transform 1 0 10584 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1667941163
transform 1 0 14560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1667941163
transform 1 0 18536 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1667941163
transform 1 0 22512 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1667941163
transform 1 0 26488 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1667941163
transform 1 0 30464 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1667941163
transform 1 0 34440 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1667941163
transform 1 0 38416 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1667941163
transform 1 0 4648 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1667941163
transform 1 0 8624 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1667941163
transform 1 0 12600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1667941163
transform 1 0 16576 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1667941163
transform 1 0 20552 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1667941163
transform 1 0 24528 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1667941163
transform 1 0 28504 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1667941163
transform 1 0 32480 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1667941163
transform 1 0 36456 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1667941163
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1667941163
transform 1 0 6608 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1667941163
transform 1 0 10584 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1667941163
transform 1 0 14560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1667941163
transform 1 0 18536 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1667941163
transform 1 0 22512 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1667941163
transform 1 0 26488 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1667941163
transform 1 0 30464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1667941163
transform 1 0 34440 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1667941163
transform 1 0 38416 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1667941163
transform 1 0 4648 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1667941163
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1667941163
transform 1 0 12600 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1667941163
transform 1 0 16576 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1667941163
transform 1 0 20552 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1667941163
transform 1 0 24528 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1667941163
transform 1 0 28504 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1667941163
transform 1 0 32480 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1667941163
transform 1 0 36456 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1667941163
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1667941163
transform 1 0 6608 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1667941163
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1667941163
transform 1 0 14560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1667941163
transform 1 0 18536 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1667941163
transform 1 0 22512 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1667941163
transform 1 0 26488 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1667941163
transform 1 0 30464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1667941163
transform 1 0 34440 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1667941163
transform 1 0 38416 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1667941163
transform 1 0 4648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1667941163
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1667941163
transform 1 0 12600 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1667941163
transform 1 0 16576 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1667941163
transform 1 0 20552 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1667941163
transform 1 0 24528 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1667941163
transform 1 0 28504 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1667941163
transform 1 0 32480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1667941163
transform 1 0 36456 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1667941163
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1667941163
transform 1 0 6608 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1667941163
transform 1 0 10584 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1667941163
transform 1 0 14560 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1667941163
transform 1 0 18536 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1667941163
transform 1 0 22512 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1667941163
transform 1 0 26488 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1667941163
transform 1 0 30464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1667941163
transform 1 0 34440 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1667941163
transform 1 0 38416 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1667941163
transform 1 0 4648 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1667941163
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1667941163
transform 1 0 12600 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1667941163
transform 1 0 16576 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1667941163
transform 1 0 20552 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1667941163
transform 1 0 24528 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1667941163
transform 1 0 28504 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1667941163
transform 1 0 32480 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1667941163
transform 1 0 36456 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1667941163
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1667941163
transform 1 0 6608 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1667941163
transform 1 0 10584 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1667941163
transform 1 0 14560 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1667941163
transform 1 0 18536 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1667941163
transform 1 0 22512 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1667941163
transform 1 0 26488 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1667941163
transform 1 0 30464 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1667941163
transform 1 0 34440 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1667941163
transform 1 0 38416 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1667941163
transform 1 0 4648 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1667941163
transform 1 0 8624 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1667941163
transform 1 0 12600 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1667941163
transform 1 0 16576 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1667941163
transform 1 0 20552 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1667941163
transform 1 0 24528 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1667941163
transform 1 0 28504 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1667941163
transform 1 0 32480 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1667941163
transform 1 0 36456 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1667941163
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1667941163
transform 1 0 6608 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1667941163
transform 1 0 10584 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1667941163
transform 1 0 14560 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1667941163
transform 1 0 18536 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1667941163
transform 1 0 22512 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1667941163
transform 1 0 26488 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1667941163
transform 1 0 30464 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1667941163
transform 1 0 34440 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1667941163
transform 1 0 38416 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1667941163
transform 1 0 4648 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1667941163
transform 1 0 8624 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1667941163
transform 1 0 12600 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1667941163
transform 1 0 16576 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1667941163
transform 1 0 20552 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1667941163
transform 1 0 24528 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1667941163
transform 1 0 28504 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1667941163
transform 1 0 32480 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1667941163
transform 1 0 36456 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1667941163
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1667941163
transform 1 0 6608 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1667941163
transform 1 0 10584 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1667941163
transform 1 0 14560 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1667941163
transform 1 0 18536 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1667941163
transform 1 0 22512 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1667941163
transform 1 0 26488 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1667941163
transform 1 0 30464 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1667941163
transform 1 0 34440 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1667941163
transform 1 0 38416 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1667941163
transform 1 0 4648 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1667941163
transform 1 0 8624 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1667941163
transform 1 0 12600 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1667941163
transform 1 0 16576 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1667941163
transform 1 0 20552 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1667941163
transform 1 0 24528 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1667941163
transform 1 0 28504 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1667941163
transform 1 0 32480 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1667941163
transform 1 0 36456 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1667941163
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1667941163
transform 1 0 6608 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1667941163
transform 1 0 10584 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1667941163
transform 1 0 14560 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1667941163
transform 1 0 18536 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1667941163
transform 1 0 22512 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1667941163
transform 1 0 26488 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1667941163
transform 1 0 30464 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1667941163
transform 1 0 34440 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1667941163
transform 1 0 38416 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1667941163
transform 1 0 4648 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1667941163
transform 1 0 8624 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1667941163
transform 1 0 12600 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1667941163
transform 1 0 16576 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1667941163
transform 1 0 20552 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1667941163
transform 1 0 24528 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1667941163
transform 1 0 28504 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1667941163
transform 1 0 32480 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1667941163
transform 1 0 36456 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1667941163
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1667941163
transform 1 0 6608 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1667941163
transform 1 0 10584 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1667941163
transform 1 0 14560 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1667941163
transform 1 0 18536 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1667941163
transform 1 0 22512 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1667941163
transform 1 0 26488 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1667941163
transform 1 0 30464 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1667941163
transform 1 0 34440 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1667941163
transform 1 0 38416 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1667941163
transform 1 0 4648 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1667941163
transform 1 0 8624 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1667941163
transform 1 0 12600 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1667941163
transform 1 0 16576 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1667941163
transform 1 0 20552 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1667941163
transform 1 0 24528 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1667941163
transform 1 0 28504 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1667941163
transform 1 0 32480 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1667941163
transform 1 0 36456 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1667941163
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1667941163
transform 1 0 4592 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1667941163
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1667941163
transform 1 0 8512 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1667941163
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1667941163
transform 1 0 12432 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1667941163
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1667941163
transform 1 0 16352 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1667941163
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1667941163
transform 1 0 20272 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1667941163
transform 1 0 22232 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1667941163
transform 1 0 24192 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1667941163
transform 1 0 26152 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1667941163
transform 1 0 28112 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1667941163
transform 1 0 30072 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1667941163
transform 1 0 32032 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1667941163
transform 1 0 33992 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1667941163
transform 1 0 35952 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1667941163
transform 1 0 37912 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 5096 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 23744 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[2\].u_series_gyp1
timestamp 1667941163
transform 1 0 1792 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 27496 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[3\].u_series_gyp1
timestamp 1667941163
transform 1 0 1792 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 29624 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 28000 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 27496 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 4536 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[8\].u_series_gyp1
timestamp 1667941163
transform 1 0 1792 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 28000 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 31584 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 31472 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[10\].u_series_gyp1
timestamp 1667941163
transform 1 0 1792 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 4592 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[11\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 28000 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[12\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 30016 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 25704 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[14\].u_series_gyp1
timestamp 1667941163
transform 1 0 1232 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 4592 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[15\].u_series_gyp1
timestamp 1667941163
transform 1 0 1232 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[16\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[16\].u_series_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[17\].u_series_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[17\].u_series_gyp1
timestamp 1667941163
transform -1 0 28000 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[18\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[18\].u_series_gyp1
timestamp 1667941163
transform -1 0 26040 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[19\].u_series_gyn1
timestamp 1667941163
transform -1 0 5096 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[19\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[20\].u_series_gyn1
timestamp 1667941163
transform -1 0 23520 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[20\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[21\].u_series_gyn1
timestamp 1667941163
transform -1 0 27496 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[21\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[22\].u_series_gyn1
timestamp 1667941163
transform -1 0 30016 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[22\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[23\].u_series_gyn1
timestamp 1667941163
transform -1 0 30016 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[23\].u_series_gyp1
timestamp 1667941163
transform 1 0 1232 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[24\].u_series_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[24\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[25\].u_series_gyn1
timestamp 1667941163
transform -1 0 6496 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[25\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[26\].u_series_gyn1
timestamp 1667941163
transform -1 0 27496 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[26\].u_series_gyp1
timestamp 1667941163
transform -1 0 4592 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[27\].u_series_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[27\].u_series_gyp1
timestamp 1667941163
transform -1 0 27496 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[28\].u_series_gyn1
timestamp 1667941163
transform -1 0 28000 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[28\].u_series_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[29\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[29\].u_series_gyp1
timestamp 1667941163
transform 1 0 1232 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[30\].u_series_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[30\].u_series_gyp1
timestamp 1667941163
transform -1 0 25480 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[31\].u_series_gyn1
timestamp 1667941163
transform -1 0 27664 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g1\[31\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 37968 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 37408 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 37968 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 31976 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 31472 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 29456 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyn1
timestamp 1667941163
transform -1 0 33432 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 28000 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g2\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 37408 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 31472 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 37408 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 33992 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 37968 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 35448 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 31976 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g3\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 35952 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 37408 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 37968 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g4\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g5\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 35448 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[0\].u_series_gyn1
timestamp 1667941163
transform -1 0 35448 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[0\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[1\].u_series_gyn1
timestamp 1667941163
transform -1 0 35952 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[1\].u_series_gyp1
timestamp 1667941163
transform -1 0 25480 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[2\].u_series_gyn1
timestamp 1667941163
transform -1 0 35952 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[2\].u_series_gyp1
timestamp 1667941163
transform -1 0 26040 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[3\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[3\].u_series_gyp1
timestamp 1667941163
transform -1 0 29456 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[4\].u_series_gyn1
timestamp 1667941163
transform -1 0 37968 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[4\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[5\].u_series_gyn1
timestamp 1667941163
transform 1 0 1232 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[5\].u_series_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[6\].u_series_gyn1
timestamp 1667941163
transform -1 0 25480 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[6\].u_series_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[7\].u_series_gyn1
timestamp 1667941163
transform -1 0 26040 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[7\].u_series_gyp1
timestamp 1667941163
transform -1 0 37408 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[8\].u_series_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[8\].u_series_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[9\].u_series_gyn1
timestamp 1667941163
transform -1 0 35504 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[9\].u_series_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[10\].u_series_gyn1
timestamp 1667941163
transform -1 0 35448 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[10\].u_series_gyp1
timestamp 1667941163
transform -1 0 27496 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[11\].u_series_gyn1
timestamp 1667941163
transform -1 0 35952 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[11\].u_series_gyp1
timestamp 1667941163
transform -1 0 26040 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[12\].u_series_gyn1
timestamp 1667941163
transform -1 0 24024 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[12\].u_series_gyp1
timestamp 1667941163
transform -1 0 33992 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[13\].u_series_gyn1
timestamp 1667941163
transform -1 0 35448 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[13\].u_series_gyp1
timestamp 1667941163
transform -1 0 35448 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[14\].u_series_gyn1
timestamp 1667941163
transform -1 0 37408 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[14\].u_series_gyp1
timestamp 1667941163
transform -1 0 35952 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[15\].u_series_gyn1
timestamp 1667941163
transform -1 0 37408 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_series_gy_g11\[15\].u_series_gyp1
timestamp 1667941163
transform -1 0 28000 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 16408 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 18368 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 16520 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 12880 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 16296 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 16800 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 19936 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 18480 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 16520 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 18368 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 15064 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 16744 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 19824 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 15064 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 14952 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 14728 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 17808 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 16800 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 17976 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 14392 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 18032 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 18312 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 18424 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[48\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[49\].u_shunt_p
timestamp 1667941163
transform -1 0 15064 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[50\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_n
timestamp 1667941163
transform -1 0 16408 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[51\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[52\].u_shunt_p
timestamp 1667941163
transform -1 0 16408 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[53\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[54\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[55\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[56\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[57\].u_shunt_p
timestamp 1667941163
transform -1 0 15064 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_n
timestamp 1667941163
transform -1 0 14896 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[58\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[59\].u_shunt_p
timestamp 1667941163
transform -1 0 14952 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_n
timestamp 1667941163
transform -1 0 16632 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[60\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[61\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[62\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[63\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[64\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[64\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[65\].u_shunt_n
timestamp 1667941163
transform -1 0 16128 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[65\].u_shunt_p
timestamp 1667941163
transform -1 0 16520 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[66\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[66\].u_shunt_p
timestamp 1667941163
transform -1 0 16520 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[67\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[67\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[68\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[68\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[69\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[69\].u_shunt_p
timestamp 1667941163
transform -1 0 16520 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[70\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[70\].u_shunt_p
timestamp 1667941163
transform -1 0 14336 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[71\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[71\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[72\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[72\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[73\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[73\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[74\].u_shunt_n
timestamp 1667941163
transform -1 0 16520 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[74\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[75\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[75\].u_shunt_p
timestamp 1667941163
transform -1 0 16968 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[76\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[76\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[77\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[77\].u_shunt_p
timestamp 1667941163
transform -1 0 12376 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[78\].u_shunt_n
timestamp 1667941163
transform -1 0 18256 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[78\].u_shunt_p
timestamp 1667941163
transform -1 0 16744 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[79\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[79\].u_shunt_p
timestamp 1667941163
transform -1 0 16184 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[80\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[80\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[81\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[81\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[82\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[82\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[83\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[83\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[84\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[84\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[85\].u_shunt_n
timestamp 1667941163
transform -1 0 12376 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[85\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[86\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[86\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[87\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[87\].u_shunt_p
timestamp 1667941163
transform -1 0 25480 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[88\].u_shunt_n
timestamp 1667941163
transform -1 0 18480 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[88\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[89\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[89\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[90\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[90\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[91\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[91\].u_shunt_p
timestamp 1667941163
transform -1 0 16520 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[92\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[92\].u_shunt_p
timestamp 1667941163
transform -1 0 15064 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[93\].u_shunt_n
timestamp 1667941163
transform -1 0 17976 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[93\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[94\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[94\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[95\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[95\].u_shunt_p
timestamp 1667941163
transform -1 0 18200 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[96\].u_shunt_n
timestamp 1667941163
transform -1 0 14336 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[96\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[97\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[97\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[98\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[98\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[99\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[99\].u_shunt_p
timestamp 1667941163
transform -1 0 16576 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[100\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[100\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[101\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[101\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[102\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[102\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[103\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[103\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[104\].u_shunt_n
timestamp 1667941163
transform -1 0 3136 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[104\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[105\].u_shunt_n
timestamp 1667941163
transform -1 0 17416 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[105\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[106\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[106\].u_shunt_p
timestamp 1667941163
transform -1 0 18368 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[107\].u_shunt_n
timestamp 1667941163
transform -1 0 16520 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[107\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[108\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[108\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[109\].u_shunt_n
timestamp 1667941163
transform -1 0 16632 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[109\].u_shunt_p
timestamp 1667941163
transform -1 0 3136 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[110\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[110\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[111\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[111\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[112\].u_shunt_n
timestamp 1667941163
transform -1 0 2576 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[112\].u_shunt_p
timestamp 1667941163
transform -1 0 16128 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[113\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[113\].u_shunt_p
timestamp 1667941163
transform -1 0 2576 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[114\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[114\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[115\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[115\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[116\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[116\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[117\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[117\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[118\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[118\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[119\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[119\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[120\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[120\].u_shunt_p
timestamp 1667941163
transform -1 0 16856 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[121\].u_shunt_n
timestamp 1667941163
transform -1 0 15064 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[121\].u_shunt_p
timestamp 1667941163
transform -1 0 16352 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[122\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[122\].u_shunt_p
timestamp 1667941163
transform -1 0 16912 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[123\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[123\].u_shunt_p
timestamp 1667941163
transform -1 0 15064 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[124\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[124\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[125\].u_shunt_n
timestamp 1667941163
transform -1 0 16408 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[125\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[126\].u_shunt_n
timestamp 1667941163
transform -1 0 16576 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[126\].u_shunt_p
timestamp 1667941163
transform -1 0 14840 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[127\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g1\[127\].u_shunt_p
timestamp 1667941163
transform -1 0 16520 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 14952 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 18032 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 15008 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[24\].u_shunt_p
timestamp 1667941163
transform -1 0 14504 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 15008 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 9072 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[27\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[32\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[32\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[33\].u_shunt_n
timestamp 1667941163
transform -1 0 14504 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[33\].u_shunt_p
timestamp 1667941163
transform -1 0 14672 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[34\].u_shunt_n
timestamp 1667941163
transform -1 0 16464 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[34\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[35\].u_shunt_n
timestamp 1667941163
transform -1 0 15008 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[35\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[36\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[36\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[37\].u_shunt_n
timestamp 1667941163
transform -1 0 21504 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[37\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[38\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[38\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[39\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[39\].u_shunt_p
timestamp 1667941163
transform -1 0 17528 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[40\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[40\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[41\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[41\].u_shunt_p
timestamp 1667941163
transform -1 0 16128 0 -1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[42\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[42\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[43\].u_shunt_n
timestamp 1667941163
transform -1 0 15008 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[43\].u_shunt_p
timestamp 1667941163
transform -1 0 12544 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[44\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[44\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[45\].u_shunt_n
timestamp 1667941163
transform -1 0 17528 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[45\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[46\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[46\].u_shunt_p
timestamp 1667941163
transform -1 0 16464 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[47\].u_shunt_n
timestamp 1667941163
transform -1 0 16464 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[47\].u_shunt_p
timestamp 1667941163
transform -1 0 10528 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[48\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[48\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[49\].u_shunt_n
timestamp 1667941163
transform -1 0 8568 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[49\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[50\].u_shunt_n
timestamp 1667941163
transform -1 0 11088 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[50\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[51\].u_shunt_n
timestamp 1667941163
transform -1 0 14672 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[51\].u_shunt_p
timestamp 1667941163
transform -1 0 18088 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[52\].u_shunt_n
timestamp 1667941163
transform -1 0 16072 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[52\].u_shunt_p
timestamp 1667941163
transform -1 0 16072 0 1 17248
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[53\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[53\].u_shunt_p
timestamp 1667941163
transform -1 0 16408 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[54\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[54\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[55\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[55\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[56\].u_shunt_n
timestamp 1667941163
transform -1 0 15008 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[56\].u_shunt_p
timestamp 1667941163
transform -1 0 13048 0 1 16464
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[57\].u_shunt_n
timestamp 1667941163
transform -1 0 10528 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[57\].u_shunt_p
timestamp 1667941163
transform -1 0 14336 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[58\].u_shunt_n
timestamp 1667941163
transform -1 0 19544 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[58\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[59\].u_shunt_n
timestamp 1667941163
transform -1 0 18088 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[59\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[60\].u_shunt_n
timestamp 1667941163
transform -1 0 12544 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[60\].u_shunt_p
timestamp 1667941163
transform -1 0 11088 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[61\].u_shunt_n
timestamp 1667941163
transform -1 0 13048 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[61\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[62\].u_shunt_n
timestamp 1667941163
transform -1 0 20048 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[62\].u_shunt_p
timestamp 1667941163
transform -1 0 15904 0 1 18032
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[63\].u_shunt_n
timestamp 1667941163
transform -1 0 16464 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g2\[63\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_n
timestamp 1667941163
transform 1 0 1792 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 26040 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 28000 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 4592 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 19824 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 17864 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_n
timestamp 1667941163
transform 1 0 1792 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 25480 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_n
timestamp 1667941163
transform 1 0 1232 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 25480 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 26040 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 20048 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 10416 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_n
timestamp 1667941163
transform 1 0 1232 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[12\].u_shunt_p
timestamp 1667941163
transform -1 0 25480 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 9072 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 8568 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[15\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[16\].u_shunt_n
timestamp 1667941163
transform -1 0 28000 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[16\].u_shunt_p
timestamp 1667941163
transform -1 0 21504 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[17\].u_shunt_n
timestamp 1667941163
transform -1 0 8456 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[17\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[18\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[18\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[19\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[19\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[20\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[20\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[21\].u_shunt_n
timestamp 1667941163
transform -1 0 5096 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[21\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[22\].u_shunt_n
timestamp 1667941163
transform -1 0 7112 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[22\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[23\].u_shunt_n
timestamp 1667941163
transform -1 0 22064 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[23\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[24\].u_shunt_n
timestamp 1667941163
transform -1 0 6552 0 1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[24\].u_shunt_p
timestamp 1667941163
transform 1 0 1792 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[25\].u_shunt_n
timestamp 1667941163
transform -1 0 28000 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[25\].u_shunt_p
timestamp 1667941163
transform -1 0 26040 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[26\].u_shunt_n
timestamp 1667941163
transform -1 0 29456 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[26\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[27\].u_shunt_n
timestamp 1667941163
transform -1 0 29456 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[27\].u_shunt_p
timestamp 1667941163
transform 1 0 1232 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[28\].u_shunt_n
timestamp 1667941163
transform -1 0 30016 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[28\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[29\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[29\].u_shunt_p
timestamp 1667941163
transform -1 0 19544 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[30\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[30\].u_shunt_p
timestamp 1667941163
transform -1 0 28000 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[31\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g3\[31\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_n
timestamp 1667941163
transform 1 0 1232 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[0\].u_shunt_p
timestamp 1667941163
transform 1 0 1792 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 28000 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 22064 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[3\].u_shunt_p
timestamp 1667941163
transform 1 0 1232 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 23520 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 24024 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_n
timestamp 1667941163
transform 1 0 1232 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[6\].u_shunt_p
timestamp 1667941163
transform 1 0 1792 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 26040 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[8\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[8\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[9\].u_shunt_n
timestamp 1667941163
transform 1 0 1792 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[9\].u_shunt_p
timestamp 1667941163
transform -1 0 6552 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[10\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[10\].u_shunt_p
timestamp 1667941163
transform -1 0 7112 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[11\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[11\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[12\].u_shunt_n
timestamp 1667941163
transform -1 0 27496 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[12\].u_shunt_p
timestamp 1667941163
transform 1 0 1232 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[13\].u_shunt_n
timestamp 1667941163
transform -1 0 25480 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[13\].u_shunt_p
timestamp 1667941163
transform -1 0 5096 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[14\].u_shunt_n
timestamp 1667941163
transform -1 0 23520 0 -1 15680
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[14\].u_shunt_p
timestamp 1667941163
transform -1 0 4592 0 -1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[15\].u_shunt_n
timestamp 1667941163
transform -1 0 24024 0 1 14896
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g4\[15\].u_shunt_p
timestamp 1667941163
transform 1 0 1792 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 35952 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 27496 0 -1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 33992 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 30016 0 -1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 37408 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 29456 0 1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 37968 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 28000 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[4\].u_shunt_n
timestamp 1667941163
transform -1 0 31472 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[4\].u_shunt_p
timestamp 1667941163
transform -1 0 30016 0 -1 12544
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[5\].u_shunt_n
timestamp 1667941163
transform -1 0 31976 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[5\].u_shunt_p
timestamp 1667941163
transform -1 0 31472 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[6\].u_shunt_n
timestamp 1667941163
transform -1 0 29456 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[6\].u_shunt_p
timestamp 1667941163
transform -1 0 29456 0 1 13328
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[7\].u_shunt_n
timestamp 1667941163
transform -1 0 33432 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g5\[7\].u_shunt_p
timestamp 1667941163
transform -1 0 28000 0 1 14112
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 35448 0 -1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 37968 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 35952 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 35448 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[2\].u_shunt_n
timestamp 1667941163
transform -1 0 33432 0 1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[2\].u_shunt_p
timestamp 1667941163
transform -1 0 35952 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[3\].u_shunt_n
timestamp 1667941163
transform -1 0 33992 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g6\[3\].u_shunt_p
timestamp 1667941163
transform -1 0 37408 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 37408 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 35952 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[1\].u_shunt_n
timestamp 1667941163
transform -1 0 37968 0 -1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g7\[1\].u_shunt_p
timestamp 1667941163
transform -1 0 37408 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g8\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 37968 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_g8\[0\].u_shunt_p
timestamp 1667941163
transform -1 0 37408 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn1 pdk_1/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1667941163
transform -1 0 30408 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 33992 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 37968 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 33992 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 32424 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 36008 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 38640 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 36008 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 37968 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 36008 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 36008 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 30408 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[3\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 37968 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 30408 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 38528 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[4\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 38528 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 28000 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 28000 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[5\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 38584 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 32424 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 28000 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[6\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 30408 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 38584 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 33992 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 32424 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g1\[7\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 36008 0 -1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 37968 0 1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 36008 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 37968 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[0\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 38640 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 38584 0 1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 38584 0 1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 38528 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[1\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 28448 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 38640 0 -1 4704
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 25984 0 1 3136
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 33544 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[2\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 32424 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 38528 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 38640 0 -1 3920
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 36008 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g2\[3\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 33992 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 28448 0 -1 5488
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 38528 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 24024 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 38528 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 32424 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyn2
timestamp 1667941163
transform 1 0 38640 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 30408 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g3\[1\].u_shunt_gyp2
timestamp 1667941163
transform 1 0 25984 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_n
timestamp 1667941163
transform -1 0 32032 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  gen_shunt_gy_g4\[0\].u_shunt_p
timestamp 1667941163
transform 1 0 29960 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33992 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 35448 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33992 0 -1 4704
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 30016 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 29456 0 1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 33432 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[3\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 33544 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[4\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 30016 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[5\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 31472 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 26152 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[6\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33992 0 -1 3136
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_shunt_gyn1
timestamp 1667941163
transform 1 0 26656 0 1 9408
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g1\[7\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 31976 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 35448 0 -1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 36624 0 -1 3920
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[1\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 26152 0 -1 11760
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 29456 0 1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[2\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 33432 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 35952 0 1 5488
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g2\[3\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 26656 0 1 10976
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 33992 0 -1 8624
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[0\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 35448 0 -1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 35448 0 -1 7840
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g3\[1\].u_shunt_gyp1
timestamp 1667941163
transform -1 0 35952 0 1 6272
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn1
timestamp 1667941163
transform -1 0 37464 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn2
timestamp 1667941163
transform -1 0 22176 0 1 1568
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyn3
timestamp 1667941163
transform -1 0 30016 0 -1 10192
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp1
timestamp 1667941163
transform 1 0 36624 0 -1 2352
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp2
timestamp 1667941163
transform -1 0 35952 0 1 7056
box -43 -43 1387 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  gen_shunt_gygy_g6\[0\].u_shunt_gyp3
timestamp 1667941163
transform -1 0 21224 0 1 2352
box -43 -43 1387 435
<< labels >>
flabel metal2 s 37408 19600 37464 20000 0 FreeSans 224 90 0 0 cap_series_gygyn
port 0 nsew signal bidirectional
flabel metal2 s 32424 19600 32480 20000 0 FreeSans 224 90 0 0 cap_series_gygyp
port 1 nsew signal bidirectional
flabel metal2 s 27440 19600 27496 20000 0 FreeSans 224 90 0 0 cap_series_gyn
port 2 nsew signal bidirectional
flabel metal2 s 22456 19600 22512 20000 0 FreeSans 224 90 0 0 cap_series_gyp
port 3 nsew signal bidirectional
flabel metal2 s 17472 19600 17528 20000 0 FreeSans 224 90 0 0 cap_shunt_gyn
port 4 nsew signal bidirectional
flabel metal2 s 12488 19600 12544 20000 0 FreeSans 224 90 0 0 cap_shunt_gyp
port 5 nsew signal bidirectional
flabel metal2 s 7504 19600 7560 20000 0 FreeSans 224 90 0 0 cap_shunt_n
port 6 nsew signal bidirectional
flabel metal2 s 2520 19600 2576 20000 0 FreeSans 224 90 0 0 cap_shunt_p
port 7 nsew signal bidirectional
flabel metal2 s 12656 0 12712 400 0 FreeSans 224 90 0 0 tune_series_gy[0]
port 8 nsew signal input
flabel metal2 s 14112 0 14168 400 0 FreeSans 224 90 0 0 tune_series_gy[1]
port 9 nsew signal input
flabel metal2 s 15568 0 15624 400 0 FreeSans 224 90 0 0 tune_series_gy[2]
port 10 nsew signal input
flabel metal2 s 17024 0 17080 400 0 FreeSans 224 90 0 0 tune_series_gy[3]
port 11 nsew signal input
flabel metal2 s 18480 0 18536 400 0 FreeSans 224 90 0 0 tune_series_gy[4]
port 12 nsew signal input
flabel metal2 s 19936 0 19992 400 0 FreeSans 224 90 0 0 tune_series_gy[5]
port 13 nsew signal input
flabel metal2 s 21392 0 21448 400 0 FreeSans 224 90 0 0 tune_series_gygy[0]
port 14 nsew signal input
flabel metal2 s 22848 0 22904 400 0 FreeSans 224 90 0 0 tune_series_gygy[1]
port 15 nsew signal input
flabel metal2 s 24304 0 24360 400 0 FreeSans 224 90 0 0 tune_series_gygy[2]
port 16 nsew signal input
flabel metal2 s 25760 0 25816 400 0 FreeSans 224 90 0 0 tune_series_gygy[3]
port 17 nsew signal input
flabel metal2 s 27216 0 27272 400 0 FreeSans 224 90 0 0 tune_series_gygy[4]
port 18 nsew signal input
flabel metal2 s 28672 0 28728 400 0 FreeSans 224 90 0 0 tune_series_gygy[5]
port 19 nsew signal input
flabel metal2 s 1008 0 1064 400 0 FreeSans 224 90 0 0 tune_shunt[0]
port 20 nsew signal input
flabel metal2 s 2464 0 2520 400 0 FreeSans 224 90 0 0 tune_shunt[1]
port 21 nsew signal input
flabel metal2 s 3920 0 3976 400 0 FreeSans 224 90 0 0 tune_shunt[2]
port 22 nsew signal input
flabel metal2 s 5376 0 5432 400 0 FreeSans 224 90 0 0 tune_shunt[3]
port 23 nsew signal input
flabel metal2 s 6832 0 6888 400 0 FreeSans 224 90 0 0 tune_shunt[4]
port 24 nsew signal input
flabel metal2 s 8288 0 8344 400 0 FreeSans 224 90 0 0 tune_shunt[5]
port 25 nsew signal input
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 tune_shunt[6]
port 26 nsew signal input
flabel metal2 s 11200 0 11256 400 0 FreeSans 224 90 0 0 tune_shunt[7]
port 27 nsew signal input
flabel metal2 s 30128 0 30184 400 0 FreeSans 224 90 0 0 tune_shunt_gy[0]
port 28 nsew signal input
flabel metal2 s 31584 0 31640 400 0 FreeSans 224 90 0 0 tune_shunt_gy[1]
port 29 nsew signal input
flabel metal2 s 33040 0 33096 400 0 FreeSans 224 90 0 0 tune_shunt_gy[2]
port 30 nsew signal input
flabel metal2 s 34496 0 34552 400 0 FreeSans 224 90 0 0 tune_shunt_gy[3]
port 31 nsew signal input
flabel metal2 s 35952 0 36008 400 0 FreeSans 224 90 0 0 tune_shunt_gy[4]
port 32 nsew signal input
flabel metal2 s 37408 0 37464 400 0 FreeSans 224 90 0 0 tune_shunt_gy[5]
port 33 nsew signal input
flabel metal2 s 38864 0 38920 400 0 FreeSans 224 90 0 0 tune_shunt_gy[6]
port 34 nsew signal input
flabel metal4 s 2054 1538 2554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 7054 1538 7554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 12054 1538 12554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 17054 1538 17554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 22054 1538 22554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 27054 1538 27554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 32054 1538 32554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 37054 1538 37554 18454 0 FreeSans 2560 90 0 0 vdd
port 35 nsew power bidirectional
flabel metal4 s 4554 1538 5054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
flabel metal4 s 9554 1538 10054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
flabel metal4 s 14554 1538 15054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
flabel metal4 s 19554 1538 20054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
flabel metal4 s 24554 1538 25054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
flabel metal4 s 29554 1538 30054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
flabel metal4 s 34554 1538 35054 18454 0 FreeSans 2560 90 0 0 vss
port 36 nsew ground bidirectional
rlabel metal1 19992 18424 19992 18424 0 vdd
rlabel metal1 19992 18032 19992 18032 0 vss
rlabel metal3 27356 9604 27356 9604 0 cap_series_gygyn
rlabel metal2 27468 11116 27468 11116 0 cap_series_gygyp
rlabel metal2 1652 2128 1652 2128 0 cap_series_gyn
rlabel metal2 2492 2184 2492 2184 0 cap_series_gyp
rlabel metal2 26124 3332 26124 3332 0 cap_shunt_gyn
rlabel metal2 24220 2184 24220 2184 0 cap_shunt_gyp
rlabel metal2 1652 14252 1652 14252 0 cap_shunt_n
rlabel metal3 2576 14700 2576 14700 0 cap_shunt_p
rlabel metal3 33894 9212 33894 9212 0 tune_series_gy[0]
rlabel metal3 34846 10388 34846 10388 0 tune_series_gy[1]
rlabel metal2 15596 427 15596 427 0 tune_series_gy[2]
rlabel metal2 29064 10780 29064 10780 0 tune_series_gy[3]
rlabel metal2 2520 1764 2520 1764 0 tune_series_gy[4]
rlabel metal2 3500 1792 3500 1792 0 tune_series_gy[5]
rlabel metal2 21420 1715 21420 1715 0 tune_series_gygy[0]
rlabel metal2 22876 1071 22876 1071 0 tune_series_gygy[1]
rlabel metal2 24332 1127 24332 1127 0 tune_series_gygy[2]
rlabel metal2 25788 427 25788 427 0 tune_series_gygy[3]
rlabel metal2 27244 1127 27244 1127 0 tune_series_gygy[4]
rlabel metal2 28700 1519 28700 1519 0 tune_series_gygy[5]
rlabel metal2 1036 4179 1036 4179 0 tune_shunt[0]
rlabel metal2 2492 1015 2492 1015 0 tune_shunt[1]
rlabel metal2 3948 427 3948 427 0 tune_shunt[2]
rlabel metal2 26236 13888 26236 13888 0 tune_shunt[3]
rlabel metal2 2548 13524 2548 13524 0 tune_shunt[4]
rlabel metal3 3864 4116 3864 4116 0 tune_shunt[5]
rlabel metal2 11340 11172 11340 11172 0 tune_shunt[6]
rlabel metal2 1596 10780 1596 10780 0 tune_shunt[7]
rlabel metal2 30296 2492 30296 2492 0 tune_shunt_gy[0]
rlabel metal2 26348 2464 26348 2464 0 tune_shunt_gy[1]
rlabel metal2 24416 2212 24416 2212 0 tune_shunt_gy[2]
rlabel metal2 26348 3920 26348 3920 0 tune_shunt_gy[3]
rlabel metal2 35980 1029 35980 1029 0 tune_shunt_gy[4]
rlabel metal3 29204 3276 29204 3276 0 tune_shunt_gy[5]
rlabel metal3 29232 3780 29232 3780 0 tune_shunt_gy[6]
<< properties >>
string FIXED_BBOX 0 0 40000 20000
<< end >>
