magic
tech gf180mcuC
magscale 1 5
timestamp 1669518838
<< obsm1 >>
rect 672 855 89400 8329
<< metal2 >>
rect 672 9600 728 10000
rect 1456 9600 1512 10000
rect 2240 9600 2296 10000
rect 3024 9600 3080 10000
rect 3808 9600 3864 10000
rect 4592 9600 4648 10000
rect 5376 9600 5432 10000
rect 6160 9600 6216 10000
rect 6944 9600 7000 10000
rect 7728 9600 7784 10000
rect 8512 9600 8568 10000
rect 9296 9600 9352 10000
rect 10080 9600 10136 10000
rect 10864 9600 10920 10000
rect 11648 9600 11704 10000
rect 12432 9600 12488 10000
rect 13216 9600 13272 10000
rect 14000 9600 14056 10000
rect 14784 9600 14840 10000
rect 15568 9600 15624 10000
rect 16352 9600 16408 10000
rect 17136 9600 17192 10000
rect 17920 9600 17976 10000
rect 18704 9600 18760 10000
rect 19488 9600 19544 10000
rect 20272 9600 20328 10000
rect 21056 9600 21112 10000
rect 21840 9600 21896 10000
rect 22624 9600 22680 10000
rect 23408 9600 23464 10000
rect 24192 9600 24248 10000
rect 24976 9600 25032 10000
rect 25760 9600 25816 10000
rect 26544 9600 26600 10000
rect 27328 9600 27384 10000
rect 28112 9600 28168 10000
rect 28896 9600 28952 10000
rect 29680 9600 29736 10000
rect 30464 9600 30520 10000
rect 31248 9600 31304 10000
rect 32032 9600 32088 10000
rect 32816 9600 32872 10000
rect 33600 9600 33656 10000
rect 34384 9600 34440 10000
rect 35168 9600 35224 10000
rect 35952 9600 36008 10000
rect 36736 9600 36792 10000
rect 37520 9600 37576 10000
rect 38304 9600 38360 10000
rect 39088 9600 39144 10000
rect 39872 9600 39928 10000
rect 40656 9600 40712 10000
rect 41440 9600 41496 10000
rect 42224 9600 42280 10000
rect 43008 9600 43064 10000
rect 43792 9600 43848 10000
rect 44576 9600 44632 10000
rect 45360 9600 45416 10000
rect 46144 9600 46200 10000
rect 46928 9600 46984 10000
rect 47712 9600 47768 10000
rect 48496 9600 48552 10000
rect 49280 9600 49336 10000
rect 50064 9600 50120 10000
rect 50848 9600 50904 10000
rect 51632 9600 51688 10000
rect 52416 9600 52472 10000
rect 53200 9600 53256 10000
rect 53984 9600 54040 10000
rect 54768 9600 54824 10000
rect 55552 9600 55608 10000
rect 56336 9600 56392 10000
rect 57120 9600 57176 10000
rect 57904 9600 57960 10000
rect 58688 9600 58744 10000
rect 59472 9600 59528 10000
rect 60256 9600 60312 10000
rect 61040 9600 61096 10000
rect 61824 9600 61880 10000
rect 62608 9600 62664 10000
rect 63392 9600 63448 10000
rect 64176 9600 64232 10000
rect 64960 9600 65016 10000
rect 65744 9600 65800 10000
rect 66528 9600 66584 10000
rect 67312 9600 67368 10000
rect 68096 9600 68152 10000
rect 68880 9600 68936 10000
rect 69664 9600 69720 10000
rect 70448 9600 70504 10000
rect 71232 9600 71288 10000
rect 72016 9600 72072 10000
rect 72800 9600 72856 10000
rect 73584 9600 73640 10000
rect 74368 9600 74424 10000
rect 75152 9600 75208 10000
rect 75936 9600 75992 10000
rect 76720 9600 76776 10000
rect 77504 9600 77560 10000
rect 78288 9600 78344 10000
rect 79072 9600 79128 10000
rect 79856 9600 79912 10000
rect 80640 9600 80696 10000
rect 81424 9600 81480 10000
rect 82208 9600 82264 10000
rect 82992 9600 83048 10000
rect 83776 9600 83832 10000
rect 84560 9600 84616 10000
rect 85344 9600 85400 10000
rect 86128 9600 86184 10000
rect 86912 9600 86968 10000
rect 87696 9600 87752 10000
rect 88480 9600 88536 10000
rect 89264 9600 89320 10000
rect 2968 0 3024 400
rect 3248 0 3304 400
rect 3528 0 3584 400
rect 3808 0 3864 400
rect 4088 0 4144 400
rect 4368 0 4424 400
rect 4648 0 4704 400
rect 4928 0 4984 400
rect 5208 0 5264 400
rect 5488 0 5544 400
rect 5768 0 5824 400
rect 6048 0 6104 400
rect 6328 0 6384 400
rect 6608 0 6664 400
rect 6888 0 6944 400
rect 7168 0 7224 400
rect 7448 0 7504 400
rect 7728 0 7784 400
rect 8008 0 8064 400
rect 8288 0 8344 400
rect 8568 0 8624 400
rect 8848 0 8904 400
rect 9128 0 9184 400
rect 9408 0 9464 400
rect 9688 0 9744 400
rect 9968 0 10024 400
rect 10248 0 10304 400
rect 10528 0 10584 400
rect 10808 0 10864 400
rect 11088 0 11144 400
rect 11368 0 11424 400
rect 11648 0 11704 400
rect 11928 0 11984 400
rect 12208 0 12264 400
rect 12488 0 12544 400
rect 12768 0 12824 400
rect 13048 0 13104 400
rect 13328 0 13384 400
rect 13608 0 13664 400
rect 13888 0 13944 400
rect 14168 0 14224 400
rect 14448 0 14504 400
rect 14728 0 14784 400
rect 15008 0 15064 400
rect 15288 0 15344 400
rect 15568 0 15624 400
rect 15848 0 15904 400
rect 16128 0 16184 400
rect 16408 0 16464 400
rect 16688 0 16744 400
rect 16968 0 17024 400
rect 17248 0 17304 400
rect 17528 0 17584 400
rect 17808 0 17864 400
rect 18088 0 18144 400
rect 18368 0 18424 400
rect 18648 0 18704 400
rect 18928 0 18984 400
rect 19208 0 19264 400
rect 19488 0 19544 400
rect 19768 0 19824 400
rect 20048 0 20104 400
rect 20328 0 20384 400
rect 20608 0 20664 400
rect 20888 0 20944 400
rect 21168 0 21224 400
rect 21448 0 21504 400
rect 21728 0 21784 400
rect 22008 0 22064 400
rect 22288 0 22344 400
rect 22568 0 22624 400
rect 22848 0 22904 400
rect 23128 0 23184 400
rect 23408 0 23464 400
rect 23688 0 23744 400
rect 23968 0 24024 400
rect 24248 0 24304 400
rect 24528 0 24584 400
rect 24808 0 24864 400
rect 25088 0 25144 400
rect 25368 0 25424 400
rect 25648 0 25704 400
rect 25928 0 25984 400
rect 26208 0 26264 400
rect 26488 0 26544 400
rect 26768 0 26824 400
rect 27048 0 27104 400
rect 27328 0 27384 400
rect 27608 0 27664 400
rect 27888 0 27944 400
rect 28168 0 28224 400
rect 28448 0 28504 400
rect 28728 0 28784 400
rect 29008 0 29064 400
rect 29288 0 29344 400
rect 29568 0 29624 400
rect 29848 0 29904 400
rect 30128 0 30184 400
rect 30408 0 30464 400
rect 30688 0 30744 400
rect 30968 0 31024 400
rect 31248 0 31304 400
rect 31528 0 31584 400
rect 31808 0 31864 400
rect 32088 0 32144 400
rect 32368 0 32424 400
rect 32648 0 32704 400
rect 32928 0 32984 400
rect 33208 0 33264 400
rect 33488 0 33544 400
rect 33768 0 33824 400
rect 34048 0 34104 400
rect 34328 0 34384 400
rect 34608 0 34664 400
rect 34888 0 34944 400
rect 35168 0 35224 400
rect 35448 0 35504 400
rect 35728 0 35784 400
rect 36008 0 36064 400
rect 36288 0 36344 400
rect 36568 0 36624 400
rect 36848 0 36904 400
rect 37128 0 37184 400
rect 37408 0 37464 400
rect 37688 0 37744 400
rect 37968 0 38024 400
rect 38248 0 38304 400
rect 38528 0 38584 400
rect 38808 0 38864 400
rect 39088 0 39144 400
rect 39368 0 39424 400
rect 39648 0 39704 400
rect 39928 0 39984 400
rect 40208 0 40264 400
rect 40488 0 40544 400
rect 40768 0 40824 400
rect 41048 0 41104 400
rect 41328 0 41384 400
rect 41608 0 41664 400
rect 41888 0 41944 400
rect 42168 0 42224 400
rect 42448 0 42504 400
rect 42728 0 42784 400
rect 43008 0 43064 400
rect 43288 0 43344 400
rect 43568 0 43624 400
rect 43848 0 43904 400
rect 44128 0 44184 400
rect 44408 0 44464 400
rect 44688 0 44744 400
rect 44968 0 45024 400
rect 45248 0 45304 400
rect 45528 0 45584 400
rect 45808 0 45864 400
rect 46088 0 46144 400
rect 46368 0 46424 400
rect 46648 0 46704 400
rect 46928 0 46984 400
rect 47208 0 47264 400
rect 47488 0 47544 400
rect 47768 0 47824 400
rect 48048 0 48104 400
rect 48328 0 48384 400
rect 48608 0 48664 400
rect 48888 0 48944 400
rect 49168 0 49224 400
rect 49448 0 49504 400
rect 49728 0 49784 400
rect 50008 0 50064 400
rect 50288 0 50344 400
rect 50568 0 50624 400
rect 50848 0 50904 400
rect 51128 0 51184 400
rect 51408 0 51464 400
rect 51688 0 51744 400
rect 51968 0 52024 400
rect 52248 0 52304 400
rect 52528 0 52584 400
rect 52808 0 52864 400
rect 53088 0 53144 400
rect 53368 0 53424 400
rect 53648 0 53704 400
rect 53928 0 53984 400
rect 54208 0 54264 400
rect 54488 0 54544 400
rect 54768 0 54824 400
rect 55048 0 55104 400
rect 55328 0 55384 400
rect 55608 0 55664 400
rect 55888 0 55944 400
rect 56168 0 56224 400
rect 56448 0 56504 400
rect 56728 0 56784 400
rect 57008 0 57064 400
rect 57288 0 57344 400
rect 57568 0 57624 400
rect 57848 0 57904 400
rect 58128 0 58184 400
rect 58408 0 58464 400
rect 58688 0 58744 400
rect 58968 0 59024 400
rect 59248 0 59304 400
rect 59528 0 59584 400
rect 59808 0 59864 400
rect 60088 0 60144 400
rect 60368 0 60424 400
rect 60648 0 60704 400
rect 60928 0 60984 400
rect 61208 0 61264 400
rect 61488 0 61544 400
rect 61768 0 61824 400
rect 62048 0 62104 400
rect 62328 0 62384 400
rect 62608 0 62664 400
rect 62888 0 62944 400
rect 63168 0 63224 400
rect 63448 0 63504 400
rect 63728 0 63784 400
rect 64008 0 64064 400
rect 64288 0 64344 400
rect 64568 0 64624 400
rect 64848 0 64904 400
rect 65128 0 65184 400
rect 65408 0 65464 400
rect 65688 0 65744 400
rect 65968 0 66024 400
rect 66248 0 66304 400
rect 66528 0 66584 400
rect 66808 0 66864 400
rect 67088 0 67144 400
rect 67368 0 67424 400
rect 67648 0 67704 400
rect 67928 0 67984 400
rect 68208 0 68264 400
rect 68488 0 68544 400
rect 68768 0 68824 400
rect 69048 0 69104 400
rect 69328 0 69384 400
rect 69608 0 69664 400
rect 69888 0 69944 400
rect 70168 0 70224 400
rect 70448 0 70504 400
rect 70728 0 70784 400
rect 71008 0 71064 400
rect 71288 0 71344 400
rect 71568 0 71624 400
rect 71848 0 71904 400
rect 72128 0 72184 400
rect 72408 0 72464 400
rect 72688 0 72744 400
rect 72968 0 73024 400
rect 73248 0 73304 400
rect 73528 0 73584 400
rect 73808 0 73864 400
rect 74088 0 74144 400
rect 74368 0 74424 400
rect 74648 0 74704 400
rect 74928 0 74984 400
rect 75208 0 75264 400
rect 75488 0 75544 400
rect 75768 0 75824 400
rect 76048 0 76104 400
rect 76328 0 76384 400
rect 76608 0 76664 400
rect 76888 0 76944 400
rect 77168 0 77224 400
rect 77448 0 77504 400
rect 77728 0 77784 400
rect 78008 0 78064 400
rect 78288 0 78344 400
rect 78568 0 78624 400
rect 78848 0 78904 400
rect 79128 0 79184 400
rect 79408 0 79464 400
rect 79688 0 79744 400
rect 79968 0 80024 400
rect 80248 0 80304 400
rect 80528 0 80584 400
rect 80808 0 80864 400
rect 81088 0 81144 400
rect 81368 0 81424 400
rect 81648 0 81704 400
rect 81928 0 81984 400
rect 82208 0 82264 400
rect 82488 0 82544 400
rect 82768 0 82824 400
rect 83048 0 83104 400
rect 83328 0 83384 400
rect 83608 0 83664 400
rect 83888 0 83944 400
rect 84168 0 84224 400
rect 84448 0 84504 400
rect 84728 0 84784 400
rect 85008 0 85064 400
rect 85288 0 85344 400
rect 85568 0 85624 400
rect 85848 0 85904 400
rect 86128 0 86184 400
rect 86408 0 86464 400
rect 86688 0 86744 400
rect 86968 0 87024 400
<< obsm2 >>
rect 758 9570 1426 9600
rect 1542 9570 2210 9600
rect 2326 9570 2994 9600
rect 3110 9570 3778 9600
rect 3894 9570 4562 9600
rect 4678 9570 5346 9600
rect 5462 9570 6130 9600
rect 6246 9570 6914 9600
rect 7030 9570 7698 9600
rect 7814 9570 8482 9600
rect 8598 9570 9266 9600
rect 9382 9570 10050 9600
rect 10166 9570 10834 9600
rect 10950 9570 11618 9600
rect 11734 9570 12402 9600
rect 12518 9570 13186 9600
rect 13302 9570 13970 9600
rect 14086 9570 14754 9600
rect 14870 9570 15538 9600
rect 15654 9570 16322 9600
rect 16438 9570 17106 9600
rect 17222 9570 17890 9600
rect 18006 9570 18674 9600
rect 18790 9570 19458 9600
rect 19574 9570 20242 9600
rect 20358 9570 21026 9600
rect 21142 9570 21810 9600
rect 21926 9570 22594 9600
rect 22710 9570 23378 9600
rect 23494 9570 24162 9600
rect 24278 9570 24946 9600
rect 25062 9570 25730 9600
rect 25846 9570 26514 9600
rect 26630 9570 27298 9600
rect 27414 9570 28082 9600
rect 28198 9570 28866 9600
rect 28982 9570 29650 9600
rect 29766 9570 30434 9600
rect 30550 9570 31218 9600
rect 31334 9570 32002 9600
rect 32118 9570 32786 9600
rect 32902 9570 33570 9600
rect 33686 9570 34354 9600
rect 34470 9570 35138 9600
rect 35254 9570 35922 9600
rect 36038 9570 36706 9600
rect 36822 9570 37490 9600
rect 37606 9570 38274 9600
rect 38390 9570 39058 9600
rect 39174 9570 39842 9600
rect 39958 9570 40626 9600
rect 40742 9570 41410 9600
rect 41526 9570 42194 9600
rect 42310 9570 42978 9600
rect 43094 9570 43762 9600
rect 43878 9570 44546 9600
rect 44662 9570 45330 9600
rect 45446 9570 46114 9600
rect 46230 9570 46898 9600
rect 47014 9570 47682 9600
rect 47798 9570 48466 9600
rect 48582 9570 49250 9600
rect 49366 9570 50034 9600
rect 50150 9570 50818 9600
rect 50934 9570 51602 9600
rect 51718 9570 52386 9600
rect 52502 9570 53170 9600
rect 53286 9570 53954 9600
rect 54070 9570 54738 9600
rect 54854 9570 55522 9600
rect 55638 9570 56306 9600
rect 56422 9570 57090 9600
rect 57206 9570 57874 9600
rect 57990 9570 58658 9600
rect 58774 9570 59442 9600
rect 59558 9570 60226 9600
rect 60342 9570 61010 9600
rect 61126 9570 61794 9600
rect 61910 9570 62578 9600
rect 62694 9570 63362 9600
rect 63478 9570 64146 9600
rect 64262 9570 64930 9600
rect 65046 9570 65714 9600
rect 65830 9570 66498 9600
rect 66614 9570 67282 9600
rect 67398 9570 68066 9600
rect 68182 9570 68850 9600
rect 68966 9570 69634 9600
rect 69750 9570 70418 9600
rect 70534 9570 71202 9600
rect 71318 9570 71986 9600
rect 72102 9570 72770 9600
rect 72886 9570 73554 9600
rect 73670 9570 74338 9600
rect 74454 9570 75122 9600
rect 75238 9570 75906 9600
rect 76022 9570 76690 9600
rect 76806 9570 77474 9600
rect 77590 9570 78258 9600
rect 78374 9570 79042 9600
rect 79158 9570 79826 9600
rect 79942 9570 80610 9600
rect 80726 9570 81394 9600
rect 81510 9570 82178 9600
rect 82294 9570 82962 9600
rect 83078 9570 83746 9600
rect 83862 9570 84530 9600
rect 84646 9570 85314 9600
rect 85430 9570 86098 9600
rect 86214 9570 86882 9600
rect 86998 9570 87666 9600
rect 87782 9570 88450 9600
rect 88566 9570 89234 9600
rect 89350 9570 89386 9600
rect 686 430 89386 9570
rect 686 400 2938 430
rect 3054 400 3218 430
rect 3334 400 3498 430
rect 3614 400 3778 430
rect 3894 400 4058 430
rect 4174 400 4338 430
rect 4454 400 4618 430
rect 4734 400 4898 430
rect 5014 400 5178 430
rect 5294 400 5458 430
rect 5574 400 5738 430
rect 5854 400 6018 430
rect 6134 400 6298 430
rect 6414 400 6578 430
rect 6694 400 6858 430
rect 6974 400 7138 430
rect 7254 400 7418 430
rect 7534 400 7698 430
rect 7814 400 7978 430
rect 8094 400 8258 430
rect 8374 400 8538 430
rect 8654 400 8818 430
rect 8934 400 9098 430
rect 9214 400 9378 430
rect 9494 400 9658 430
rect 9774 400 9938 430
rect 10054 400 10218 430
rect 10334 400 10498 430
rect 10614 400 10778 430
rect 10894 400 11058 430
rect 11174 400 11338 430
rect 11454 400 11618 430
rect 11734 400 11898 430
rect 12014 400 12178 430
rect 12294 400 12458 430
rect 12574 400 12738 430
rect 12854 400 13018 430
rect 13134 400 13298 430
rect 13414 400 13578 430
rect 13694 400 13858 430
rect 13974 400 14138 430
rect 14254 400 14418 430
rect 14534 400 14698 430
rect 14814 400 14978 430
rect 15094 400 15258 430
rect 15374 400 15538 430
rect 15654 400 15818 430
rect 15934 400 16098 430
rect 16214 400 16378 430
rect 16494 400 16658 430
rect 16774 400 16938 430
rect 17054 400 17218 430
rect 17334 400 17498 430
rect 17614 400 17778 430
rect 17894 400 18058 430
rect 18174 400 18338 430
rect 18454 400 18618 430
rect 18734 400 18898 430
rect 19014 400 19178 430
rect 19294 400 19458 430
rect 19574 400 19738 430
rect 19854 400 20018 430
rect 20134 400 20298 430
rect 20414 400 20578 430
rect 20694 400 20858 430
rect 20974 400 21138 430
rect 21254 400 21418 430
rect 21534 400 21698 430
rect 21814 400 21978 430
rect 22094 400 22258 430
rect 22374 400 22538 430
rect 22654 400 22818 430
rect 22934 400 23098 430
rect 23214 400 23378 430
rect 23494 400 23658 430
rect 23774 400 23938 430
rect 24054 400 24218 430
rect 24334 400 24498 430
rect 24614 400 24778 430
rect 24894 400 25058 430
rect 25174 400 25338 430
rect 25454 400 25618 430
rect 25734 400 25898 430
rect 26014 400 26178 430
rect 26294 400 26458 430
rect 26574 400 26738 430
rect 26854 400 27018 430
rect 27134 400 27298 430
rect 27414 400 27578 430
rect 27694 400 27858 430
rect 27974 400 28138 430
rect 28254 400 28418 430
rect 28534 400 28698 430
rect 28814 400 28978 430
rect 29094 400 29258 430
rect 29374 400 29538 430
rect 29654 400 29818 430
rect 29934 400 30098 430
rect 30214 400 30378 430
rect 30494 400 30658 430
rect 30774 400 30938 430
rect 31054 400 31218 430
rect 31334 400 31498 430
rect 31614 400 31778 430
rect 31894 400 32058 430
rect 32174 400 32338 430
rect 32454 400 32618 430
rect 32734 400 32898 430
rect 33014 400 33178 430
rect 33294 400 33458 430
rect 33574 400 33738 430
rect 33854 400 34018 430
rect 34134 400 34298 430
rect 34414 400 34578 430
rect 34694 400 34858 430
rect 34974 400 35138 430
rect 35254 400 35418 430
rect 35534 400 35698 430
rect 35814 400 35978 430
rect 36094 400 36258 430
rect 36374 400 36538 430
rect 36654 400 36818 430
rect 36934 400 37098 430
rect 37214 400 37378 430
rect 37494 400 37658 430
rect 37774 400 37938 430
rect 38054 400 38218 430
rect 38334 400 38498 430
rect 38614 400 38778 430
rect 38894 400 39058 430
rect 39174 400 39338 430
rect 39454 400 39618 430
rect 39734 400 39898 430
rect 40014 400 40178 430
rect 40294 400 40458 430
rect 40574 400 40738 430
rect 40854 400 41018 430
rect 41134 400 41298 430
rect 41414 400 41578 430
rect 41694 400 41858 430
rect 41974 400 42138 430
rect 42254 400 42418 430
rect 42534 400 42698 430
rect 42814 400 42978 430
rect 43094 400 43258 430
rect 43374 400 43538 430
rect 43654 400 43818 430
rect 43934 400 44098 430
rect 44214 400 44378 430
rect 44494 400 44658 430
rect 44774 400 44938 430
rect 45054 400 45218 430
rect 45334 400 45498 430
rect 45614 400 45778 430
rect 45894 400 46058 430
rect 46174 400 46338 430
rect 46454 400 46618 430
rect 46734 400 46898 430
rect 47014 400 47178 430
rect 47294 400 47458 430
rect 47574 400 47738 430
rect 47854 400 48018 430
rect 48134 400 48298 430
rect 48414 400 48578 430
rect 48694 400 48858 430
rect 48974 400 49138 430
rect 49254 400 49418 430
rect 49534 400 49698 430
rect 49814 400 49978 430
rect 50094 400 50258 430
rect 50374 400 50538 430
rect 50654 400 50818 430
rect 50934 400 51098 430
rect 51214 400 51378 430
rect 51494 400 51658 430
rect 51774 400 51938 430
rect 52054 400 52218 430
rect 52334 400 52498 430
rect 52614 400 52778 430
rect 52894 400 53058 430
rect 53174 400 53338 430
rect 53454 400 53618 430
rect 53734 400 53898 430
rect 54014 400 54178 430
rect 54294 400 54458 430
rect 54574 400 54738 430
rect 54854 400 55018 430
rect 55134 400 55298 430
rect 55414 400 55578 430
rect 55694 400 55858 430
rect 55974 400 56138 430
rect 56254 400 56418 430
rect 56534 400 56698 430
rect 56814 400 56978 430
rect 57094 400 57258 430
rect 57374 400 57538 430
rect 57654 400 57818 430
rect 57934 400 58098 430
rect 58214 400 58378 430
rect 58494 400 58658 430
rect 58774 400 58938 430
rect 59054 400 59218 430
rect 59334 400 59498 430
rect 59614 400 59778 430
rect 59894 400 60058 430
rect 60174 400 60338 430
rect 60454 400 60618 430
rect 60734 400 60898 430
rect 61014 400 61178 430
rect 61294 400 61458 430
rect 61574 400 61738 430
rect 61854 400 62018 430
rect 62134 400 62298 430
rect 62414 400 62578 430
rect 62694 400 62858 430
rect 62974 400 63138 430
rect 63254 400 63418 430
rect 63534 400 63698 430
rect 63814 400 63978 430
rect 64094 400 64258 430
rect 64374 400 64538 430
rect 64654 400 64818 430
rect 64934 400 65098 430
rect 65214 400 65378 430
rect 65494 400 65658 430
rect 65774 400 65938 430
rect 66054 400 66218 430
rect 66334 400 66498 430
rect 66614 400 66778 430
rect 66894 400 67058 430
rect 67174 400 67338 430
rect 67454 400 67618 430
rect 67734 400 67898 430
rect 68014 400 68178 430
rect 68294 400 68458 430
rect 68574 400 68738 430
rect 68854 400 69018 430
rect 69134 400 69298 430
rect 69414 400 69578 430
rect 69694 400 69858 430
rect 69974 400 70138 430
rect 70254 400 70418 430
rect 70534 400 70698 430
rect 70814 400 70978 430
rect 71094 400 71258 430
rect 71374 400 71538 430
rect 71654 400 71818 430
rect 71934 400 72098 430
rect 72214 400 72378 430
rect 72494 400 72658 430
rect 72774 400 72938 430
rect 73054 400 73218 430
rect 73334 400 73498 430
rect 73614 400 73778 430
rect 73894 400 74058 430
rect 74174 400 74338 430
rect 74454 400 74618 430
rect 74734 400 74898 430
rect 75014 400 75178 430
rect 75294 400 75458 430
rect 75574 400 75738 430
rect 75854 400 76018 430
rect 76134 400 76298 430
rect 76414 400 76578 430
rect 76694 400 76858 430
rect 76974 400 77138 430
rect 77254 400 77418 430
rect 77534 400 77698 430
rect 77814 400 77978 430
rect 78094 400 78258 430
rect 78374 400 78538 430
rect 78654 400 78818 430
rect 78934 400 79098 430
rect 79214 400 79378 430
rect 79494 400 79658 430
rect 79774 400 79938 430
rect 80054 400 80218 430
rect 80334 400 80498 430
rect 80614 400 80778 430
rect 80894 400 81058 430
rect 81174 400 81338 430
rect 81454 400 81618 430
rect 81734 400 81898 430
rect 82014 400 82178 430
rect 82294 400 82458 430
rect 82574 400 82738 430
rect 82854 400 83018 430
rect 83134 400 83298 430
rect 83414 400 83578 430
rect 83694 400 83858 430
rect 83974 400 84138 430
rect 84254 400 84418 430
rect 84534 400 84698 430
rect 84814 400 84978 430
rect 85094 400 85258 430
rect 85374 400 85538 430
rect 85654 400 85818 430
rect 85934 400 86098 430
rect 86214 400 86378 430
rect 86494 400 86658 430
rect 86774 400 86938 430
rect 87054 400 89386 430
<< obsm3 >>
rect 1073 1554 89391 8246
<< metal4 >>
rect 11673 1538 11833 8262
rect 22754 1538 22914 8262
rect 33835 1538 33995 8262
rect 44916 1538 45076 8262
rect 55997 1538 56157 8262
rect 67078 1538 67238 8262
rect 78159 1538 78319 8262
rect 89240 1538 89400 8262
<< labels >>
rlabel metal2 s 672 9600 728 10000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24192 9600 24248 10000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 26544 9600 26600 10000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 28896 9600 28952 10000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 31248 9600 31304 10000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 33600 9600 33656 10000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 35952 9600 36008 10000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38304 9600 38360 10000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40656 9600 40712 10000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43008 9600 43064 10000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45360 9600 45416 10000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3024 9600 3080 10000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47712 9600 47768 10000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50064 9600 50120 10000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 52416 9600 52472 10000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 54768 9600 54824 10000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57120 9600 57176 10000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 59472 9600 59528 10000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 61824 9600 61880 10000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 64176 9600 64232 10000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 66528 9600 66584 10000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 68880 9600 68936 10000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5376 9600 5432 10000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 71232 9600 71288 10000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 73584 9600 73640 10000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 75936 9600 75992 10000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 78288 9600 78344 10000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 80640 9600 80696 10000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 82992 9600 83048 10000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 85344 9600 85400 10000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 87696 9600 87752 10000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7728 9600 7784 10000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10080 9600 10136 10000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12432 9600 12488 10000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14784 9600 14840 10000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17136 9600 17192 10000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19488 9600 19544 10000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 21840 9600 21896 10000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1456 9600 1512 10000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 24976 9600 25032 10000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27328 9600 27384 10000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29680 9600 29736 10000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32032 9600 32088 10000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34384 9600 34440 10000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36736 9600 36792 10000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39088 9600 39144 10000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41440 9600 41496 10000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 43792 9600 43848 10000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46144 9600 46200 10000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3808 9600 3864 10000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48496 9600 48552 10000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 50848 9600 50904 10000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 53200 9600 53256 10000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 55552 9600 55608 10000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 57904 9600 57960 10000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 60256 9600 60312 10000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 62608 9600 62664 10000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 64960 9600 65016 10000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 67312 9600 67368 10000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 69664 9600 69720 10000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6160 9600 6216 10000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 72016 9600 72072 10000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 74368 9600 74424 10000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 76720 9600 76776 10000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 79072 9600 79128 10000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 81424 9600 81480 10000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 83776 9600 83832 10000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 86128 9600 86184 10000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 88480 9600 88536 10000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8512 9600 8568 10000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10864 9600 10920 10000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13216 9600 13272 10000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15568 9600 15624 10000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17920 9600 17976 10000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20272 9600 20328 10000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 22624 9600 22680 10000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2240 9600 2296 10000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 25760 9600 25816 10000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28112 9600 28168 10000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 30464 9600 30520 10000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 32816 9600 32872 10000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35168 9600 35224 10000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37520 9600 37576 10000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 39872 9600 39928 10000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42224 9600 42280 10000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44576 9600 44632 10000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 46928 9600 46984 10000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4592 9600 4648 10000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 49280 9600 49336 10000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 51632 9600 51688 10000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 53984 9600 54040 10000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 56336 9600 56392 10000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 58688 9600 58744 10000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 61040 9600 61096 10000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 63392 9600 63448 10000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 65744 9600 65800 10000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 68096 9600 68152 10000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 70448 9600 70504 10000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6944 9600 7000 10000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 72800 9600 72856 10000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 75152 9600 75208 10000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 77504 9600 77560 10000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 79856 9600 79912 10000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 82208 9600 82264 10000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 84560 9600 84616 10000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 86912 9600 86968 10000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 89264 9600 89320 10000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9296 9600 9352 10000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11648 9600 11704 10000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14000 9600 14056 10000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16352 9600 16408 10000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18704 9600 18760 10000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 21056 9600 21112 10000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23408 9600 23464 10000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 86408 0 86464 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 86688 0 86744 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 86968 0 87024 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 32648 0 32704 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 41048 0 41104 400 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 42728 0 42784 400 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 44408 0 44464 400 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 46088 0 46144 400 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 47768 0 47824 400 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 49448 0 49504 400 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 51128 0 51184 400 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 51968 0 52024 400 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 52808 0 52864 400 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 54488 0 54544 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 56168 0 56224 400 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 34328 0 34384 400 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 57848 0 57904 400 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 58688 0 58744 400 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 59528 0 59584 400 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 61208 0 61264 400 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 62888 0 62944 400 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 63728 0 63784 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 64568 0 64624 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 65408 0 65464 400 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 66248 0 66304 400 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 67088 0 67144 400 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 67928 0 67984 400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 68768 0 68824 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 69608 0 69664 400 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 70448 0 70504 400 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 71288 0 71344 400 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 72968 0 73024 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 73808 0 73864 400 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 36008 0 36064 400 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 74648 0 74704 400 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 76328 0 76384 400 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 78008 0 78064 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 78848 0 78904 400 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 79688 0 79744 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 80528 0 80584 400 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 81368 0 81424 400 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 82208 0 82264 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 83048 0 83104 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 84728 0 84784 400 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 85568 0 85624 400 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 37688 0 37744 400 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 39368 0 39424 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 42168 0 42224 400 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 43008 0 43064 400 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 43848 0 43904 400 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 44688 0 44744 400 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 45528 0 45584 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 46368 0 46424 400 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 47208 0 47264 400 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 48888 0 48944 400 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 33768 0 33824 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 49728 0 49784 400 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 50568 0 50624 400 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 51408 0 51464 400 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 52248 0 52304 400 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 53928 0 53984 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 55608 0 55664 400 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 56448 0 56504 400 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 57288 0 57344 400 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 58968 0 59024 400 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 59808 0 59864 400 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 60648 0 60704 400 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 62328 0 62384 400 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 64008 0 64064 400 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 65688 0 65744 400 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 35448 0 35504 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 66528 0 66584 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 67368 0 67424 400 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 69048 0 69104 400 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 69888 0 69944 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 70728 0 70784 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 71568 0 71624 400 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 72408 0 72464 400 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 73248 0 73304 400 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 74088 0 74144 400 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 74928 0 74984 400 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 75768 0 75824 400 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 76608 0 76664 400 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 77448 0 77504 400 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 78288 0 78344 400 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 79128 0 79184 400 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 79968 0 80024 400 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 80808 0 80864 400 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 81648 0 81704 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 82488 0 82544 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 37128 0 37184 400 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 83328 0 83384 400 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 84168 0 84224 400 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 85008 0 85064 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 85848 0 85904 400 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 38808 0 38864 400 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 39648 0 39704 400 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 40488 0 40544 400 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 33208 0 33264 400 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 41608 0 41664 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 43288 0 43344 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 44968 0 45024 400 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 46648 0 46704 400 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 48328 0 48384 400 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 50008 0 50064 400 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 51688 0 51744 400 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 53368 0 53424 400 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 54208 0 54264 400 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 55048 0 55104 400 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 56728 0 56784 400 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 34888 0 34944 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 58408 0 58464 400 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 60088 0 60144 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 61768 0 61824 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 62608 0 62664 400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 63448 0 63504 400 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 65128 0 65184 400 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 66808 0 66864 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 67648 0 67704 400 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 68488 0 68544 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 70168 0 70224 400 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 71848 0 71904 400 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 73528 0 73584 400 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 36568 0 36624 400 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 75208 0 75264 400 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 76048 0 76104 400 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 76888 0 76944 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 78568 0 78624 400 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 80248 0 80304 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 81088 0 81144 400 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 81928 0 81984 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 82768 0 82824 400 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 83608 0 83664 400 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 85288 0 85344 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 38248 0 38304 400 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 39928 0 39984 400 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 11673 1538 11833 8262 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 33835 1538 33995 8262 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 55997 1538 56157 8262 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 78159 1538 78319 8262 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 22754 1538 22914 8262 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 44916 1538 45076 8262 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 67078 1538 67238 8262 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 89240 1538 89400 8262 6 vss
port 311 nsew ground bidirectional
rlabel metal2 s 2968 0 3024 400 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 3248 0 3304 400 6 wb_rst_i
port 313 nsew signal input
rlabel metal2 s 3528 0 3584 400 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 4648 0 4704 400 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 14168 0 14224 400 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 15848 0 15904 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal2 s 17528 0 17584 400 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal2 s 18368 0 18424 400 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 19208 0 19264 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal2 s 20888 0 20944 400 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal2 s 5768 0 5824 400 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal2 s 22568 0 22624 400 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 24248 0 24304 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 25928 0 25984 400 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 27608 0 27664 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal2 s 29288 0 29344 400 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal2 s 6888 0 6944 400 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal2 s 30968 0 31024 400 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 9128 0 9184 400 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal2 s 10808 0 10864 400 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal2 s 12488 0 12544 400 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal2 s 4928 0 4984 400 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal2 s 15288 0 15344 400 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 16968 0 17024 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal2 s 18648 0 18704 400 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 20328 0 20384 400 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 22008 0 22064 400 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 23688 0 23744 400 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal2 s 25368 0 25424 400 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 27048 0 27104 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 28728 0 28784 400 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal2 s 30408 0 30464 400 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal2 s 32088 0 32144 400 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 10248 0 10304 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 11928 0 11984 400 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal2 s 13608 0 13664 400 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal2 s 5208 0 5264 400 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal2 s 14728 0 14784 400 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal2 s 16408 0 16464 400 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 17248 0 17304 400 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal2 s 18088 0 18144 400 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal2 s 19768 0 19824 400 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal2 s 20608 0 20664 400 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 21448 0 21504 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 6328 0 6384 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal2 s 23128 0 23184 400 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal2 s 23968 0 24024 400 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 24808 0 24864 400 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 26488 0 26544 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 27328 0 27384 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 28168 0 28224 400 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 29008 0 29064 400 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 29848 0 29904 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal2 s 7448 0 7504 400 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal2 s 31528 0 31584 400 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 8568 0 8624 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 9688 0 9744 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal2 s 11368 0 11424 400 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 12208 0 12264 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 13048 0 13104 400 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 13888 0 13944 400 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal2 s 5488 0 5544 400 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal2 s 4088 0 4144 400 6 wbs_stb_i
port 416 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 642518
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/user_proj_example/runs/22_11_26_22_13/results/signoff/user_proj_example.magic.gds
string GDS_START 94304
<< end >>

