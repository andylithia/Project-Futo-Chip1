magic
tech gf180mcuC
magscale 1 5
timestamp 1669922098
<< obsm1 >>
rect 672 1538 19320 28254
<< metal2 >>
rect 1344 29600 1400 30000
rect 3808 29600 3864 30000
rect 6272 29600 6328 30000
rect 8736 29600 8792 30000
rect 11200 29600 11256 30000
rect 13664 29600 13720 30000
rect 16128 29600 16184 30000
rect 18592 29600 18648 30000
rect 1680 0 1736 400
rect 4984 0 5040 400
rect 8288 0 8344 400
rect 11592 0 11648 400
rect 14896 0 14952 400
rect 18200 0 18256 400
<< obsm2 >>
rect 910 29570 1314 29600
rect 1430 29570 3778 29600
rect 3894 29570 6242 29600
rect 6358 29570 8706 29600
rect 8822 29570 11170 29600
rect 11286 29570 13634 29600
rect 13750 29570 16098 29600
rect 16214 29570 18562 29600
rect 18678 29570 19082 29600
rect 910 430 19082 29570
rect 910 350 1650 430
rect 1766 350 4954 430
rect 5070 350 8258 430
rect 8374 350 11562 430
rect 11678 350 14866 430
rect 14982 350 18170 430
rect 18286 350 19082 430
<< metal3 >>
rect 19600 28728 20000 28784
rect 0 27888 400 27944
rect 19600 26432 20000 26488
rect 0 24192 400 24248
rect 19600 24136 20000 24192
rect 19600 21840 20000 21896
rect 0 20496 400 20552
rect 19600 19544 20000 19600
rect 19600 17248 20000 17304
rect 0 16800 400 16856
rect 19600 14952 20000 15008
rect 0 13104 400 13160
rect 19600 12656 20000 12712
rect 19600 10360 20000 10416
rect 0 9408 400 9464
rect 19600 8064 20000 8120
rect 0 5712 400 5768
rect 19600 5768 20000 5824
rect 19600 3472 20000 3528
rect 0 2016 400 2072
rect 19600 1176 20000 1232
<< obsm3 >>
rect 400 28698 19570 28770
rect 400 27974 19600 28698
rect 430 27858 19600 27974
rect 400 26518 19600 27858
rect 400 26402 19570 26518
rect 400 24278 19600 26402
rect 430 24222 19600 24278
rect 430 24162 19570 24222
rect 400 24106 19570 24162
rect 400 21926 19600 24106
rect 400 21810 19570 21926
rect 400 20582 19600 21810
rect 430 20466 19600 20582
rect 400 19630 19600 20466
rect 400 19514 19570 19630
rect 400 17334 19600 19514
rect 400 17218 19570 17334
rect 400 16886 19600 17218
rect 430 16770 19600 16886
rect 400 15038 19600 16770
rect 400 14922 19570 15038
rect 400 13190 19600 14922
rect 430 13074 19600 13190
rect 400 12742 19600 13074
rect 400 12626 19570 12742
rect 400 10446 19600 12626
rect 400 10330 19570 10446
rect 400 9494 19600 10330
rect 430 9378 19600 9494
rect 400 8150 19600 9378
rect 400 8034 19570 8150
rect 400 5854 19600 8034
rect 400 5798 19570 5854
rect 430 5738 19570 5798
rect 430 5682 19600 5738
rect 400 3558 19600 5682
rect 400 3442 19570 3558
rect 400 2102 19600 3442
rect 430 1986 19600 2102
rect 400 1262 19600 1986
rect 400 1190 19570 1262
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
<< obsm4 >>
rect 17822 3313 17850 5815
<< labels >>
rlabel metal2 s 18592 29600 18648 30000 6 cap_series_gygyn
port 1 nsew signal bidirectional
rlabel metal2 s 16128 29600 16184 30000 6 cap_series_gygyp
port 2 nsew signal bidirectional
rlabel metal2 s 13664 29600 13720 30000 6 cap_series_gyn
port 3 nsew signal bidirectional
rlabel metal2 s 11200 29600 11256 30000 6 cap_series_gyp
port 4 nsew signal bidirectional
rlabel metal2 s 8736 29600 8792 30000 6 cap_shunt_gyn
port 5 nsew signal bidirectional
rlabel metal2 s 6272 29600 6328 30000 6 cap_shunt_gyp
port 6 nsew signal bidirectional
rlabel metal2 s 3808 29600 3864 30000 6 cap_shunt_n
port 7 nsew signal bidirectional
rlabel metal2 s 1344 29600 1400 30000 6 cap_shunt_p
port 8 nsew signal bidirectional
rlabel metal2 s 1680 0 1736 400 6 tune_series_gy[0]
port 9 nsew signal input
rlabel metal2 s 4984 0 5040 400 6 tune_series_gy[1]
port 10 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 tune_series_gy[2]
port 11 nsew signal input
rlabel metal2 s 11592 0 11648 400 6 tune_series_gy[3]
port 12 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 tune_series_gy[4]
port 13 nsew signal input
rlabel metal2 s 18200 0 18256 400 6 tune_series_gy[5]
port 14 nsew signal input
rlabel metal3 s 19600 1176 20000 1232 6 tune_series_gygy[0]
port 15 nsew signal input
rlabel metal3 s 19600 3472 20000 3528 6 tune_series_gygy[1]
port 16 nsew signal input
rlabel metal3 s 19600 5768 20000 5824 6 tune_series_gygy[2]
port 17 nsew signal input
rlabel metal3 s 19600 8064 20000 8120 6 tune_series_gygy[3]
port 18 nsew signal input
rlabel metal3 s 19600 10360 20000 10416 6 tune_series_gygy[4]
port 19 nsew signal input
rlabel metal3 s 19600 12656 20000 12712 6 tune_series_gygy[5]
port 20 nsew signal input
rlabel metal3 s 0 2016 400 2072 6 tune_shunt[0]
port 21 nsew signal input
rlabel metal3 s 0 5712 400 5768 6 tune_shunt[1]
port 22 nsew signal input
rlabel metal3 s 0 9408 400 9464 6 tune_shunt[2]
port 23 nsew signal input
rlabel metal3 s 0 13104 400 13160 6 tune_shunt[3]
port 24 nsew signal input
rlabel metal3 s 0 16800 400 16856 6 tune_shunt[4]
port 25 nsew signal input
rlabel metal3 s 0 20496 400 20552 6 tune_shunt[5]
port 26 nsew signal input
rlabel metal3 s 0 24192 400 24248 6 tune_shunt[6]
port 27 nsew signal input
rlabel metal3 s 0 27888 400 27944 6 tune_shunt[7]
port 28 nsew signal input
rlabel metal3 s 19600 14952 20000 15008 6 tune_shunt_gy[0]
port 29 nsew signal input
rlabel metal3 s 19600 17248 20000 17304 6 tune_shunt_gy[1]
port 30 nsew signal input
rlabel metal3 s 19600 19544 20000 19600 6 tune_shunt_gy[2]
port 31 nsew signal input
rlabel metal3 s 19600 21840 20000 21896 6 tune_shunt_gy[3]
port 32 nsew signal input
rlabel metal3 s 19600 24136 20000 24192 6 tune_shunt_gy[4]
port 33 nsew signal input
rlabel metal3 s 19600 26432 20000 26488 6 tune_shunt_gy[5]
port 34 nsew signal input
rlabel metal3 s 19600 28728 20000 28784 6 tune_shunt_gy[6]
port 35 nsew signal input
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 36 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 36 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 37 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 768870
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/caparray_s1/runs/22_12_01_14_14/results/signoff/caparray_s1.magic.gds
string GDS_START 54730
<< end >>

