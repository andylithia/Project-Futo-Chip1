magic
tech gf180mcuC
magscale 1 10
timestamp 1669525571
<< error_p >>
rect -258 -244 -224 196
rect -48 109 -37 155
rect -138 -124 -104 76
rect 104 -124 138 76
rect 224 -244 258 196
<< nwell >>
rect -224 -254 224 254
<< mvpmos >>
rect -50 -124 50 76
<< mvpdiff >>
rect -138 63 -50 76
rect -138 -111 -125 63
rect -79 -111 -50 63
rect -138 -124 -50 -111
rect 50 63 138 76
rect 50 -111 79 63
rect 125 -111 138 63
rect 50 -124 138 -111
<< mvpdiffc >>
rect -125 -111 -79 63
rect 79 -111 125 63
<< polysilicon >>
rect -50 155 50 168
rect -50 109 -37 155
rect 37 109 50 155
rect -50 76 50 109
rect -50 -168 50 -124
<< polycontact >>
rect -37 109 37 155
<< metal1 >>
rect -48 109 -37 155
rect 37 109 48 155
rect -125 63 -79 74
rect -125 -122 -79 -111
rect 79 63 125 74
rect 79 -122 125 -111
<< properties >>
string gencell pmos_6p0
string library gf180mcu
string parameters w 1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
