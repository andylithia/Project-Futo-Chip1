magic
tech gf180mcuC
magscale 1 5
timestamp 1669692784
<< obsm1 >>
rect 672 1538 19400 18454
<< metal2 >>
rect 1344 0 1400 400
rect 3808 0 3864 400
rect 6272 0 6328 400
rect 8736 0 8792 400
rect 11200 0 11256 400
rect 13664 0 13720 400
rect 16128 0 16184 400
rect 18592 0 18648 400
<< obsm2 >>
rect 1358 430 19386 18443
rect 1430 350 3778 430
rect 3894 350 6242 430
rect 6358 350 8706 430
rect 8822 350 11170 430
rect 11286 350 13634 430
rect 13750 350 16098 430
rect 16214 350 18562 430
rect 18678 350 19386 430
<< obsm3 >>
rect 1353 1554 19391 18438
<< metal4 >>
rect 2923 1538 3083 18454
rect 5254 1538 5414 18454
rect 7585 1538 7745 18454
rect 9916 1538 10076 18454
rect 12247 1538 12407 18454
rect 14578 1538 14738 18454
rect 16909 1538 17069 18454
rect 19240 1538 19400 18454
<< labels >>
rlabel metal2 s 1344 0 1400 400 6 clk
port 1 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 clko
port 2 nsew signal output
rlabel metal2 s 8736 0 8792 400 6 latch
port 3 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 on
port 4 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 op
port 5 nsew signal output
rlabel metal2 s 3808 0 3864 400 6 rst
port 6 nsew signal input
rlabel metal2 s 6272 0 6328 400 6 sdi
port 7 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 sig
port 8 nsew signal input
rlabel metal4 s 2923 1538 3083 18454 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 7585 1538 7745 18454 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 12247 1538 12407 18454 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 16909 1538 17069 18454 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 5254 1538 5414 18454 6 vss
port 10 nsew ground bidirectional
rlabel metal4 s 9916 1538 10076 18454 6 vss
port 10 nsew ground bidirectional
rlabel metal4 s 14578 1538 14738 18454 6 vss
port 10 nsew ground bidirectional
rlabel metal4 s 19240 1538 19400 18454 6 vss
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 365658
string GDS_FILE /home/andylithia/openmpw/Project-Futo-Chip1/openlane/dlc/runs/22_11_28_22_32/results/signoff/dlc.magic.gds
string GDS_START 51750
<< end >>

