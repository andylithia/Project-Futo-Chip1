magic
tech gf180mcuC
magscale 1 10
timestamp 1669860689
<< nwell >>
rect 1258 8192 10726 8710
rect 1258 6624 10726 7488
rect 1258 5056 10726 5920
rect 1258 3488 10726 4352
<< pwell >>
rect 1258 7488 10726 8192
rect 1258 5920 10726 6624
rect 1258 4352 10726 5056
rect 1258 3050 10726 3488
<< mvnmos >>
rect 1692 7908 1892 8072
rect 2140 7908 2260 8072
rect 2812 7908 2932 8072
rect 3484 7908 3604 8072
rect 4156 7908 4276 8072
rect 4828 7908 4948 8072
rect 5612 7908 5812 8072
rect 6060 7908 6260 8072
rect 6508 7908 6708 8072
rect 6956 7908 7156 8072
rect 7404 7908 7604 8072
rect 7852 7908 8052 8072
rect 8300 7908 8500 8072
rect 8748 7908 8948 8072
rect 9532 7908 9732 8072
rect 9980 7908 10180 8072
rect 1692 7608 1892 7772
rect 2140 7608 2260 7772
rect 2812 7608 2932 7772
rect 3484 7608 3604 7772
rect 4156 7608 4276 7772
rect 4828 7608 4948 7772
rect 5580 7608 5700 7772
rect 6252 7608 6372 7772
rect 6620 7608 6820 7772
rect 7068 7608 7268 7772
rect 7516 7608 7716 7772
rect 7964 7608 8164 7772
rect 8412 7608 8612 7772
rect 8860 7608 9060 7772
rect 10060 7608 10180 7772
rect 1916 6340 2036 6504
rect 2588 6340 2708 6504
rect 3260 6340 3380 6504
rect 3932 6340 4052 6504
rect 4604 6340 4724 6504
rect 5724 6340 5844 6504
rect 6396 6340 6516 6504
rect 7068 6340 7188 6504
rect 7516 6340 7716 6504
rect 7964 6340 8164 6504
rect 8412 6340 8532 6504
rect 9084 6365 9204 6437
rect 9308 6365 9428 6437
rect 9568 6340 9688 6504
rect 9792 6340 9912 6504
rect 9976 6340 10096 6504
rect 1804 6040 1924 6204
rect 2476 6040 2596 6204
rect 3148 6040 3268 6204
rect 3820 6040 3940 6204
rect 4492 6040 4612 6204
rect 5164 6040 5284 6204
rect 5836 6040 5956 6204
rect 6508 6040 6628 6204
rect 6956 6040 7156 6204
rect 7740 6040 7860 6204
rect 8412 6040 8532 6204
rect 8860 6040 9060 6204
rect 10060 6040 10180 6204
rect 1692 4772 1892 4936
rect 2140 4772 2260 4936
rect 2812 4772 2932 4936
rect 3484 4772 3604 4936
rect 4156 4772 4276 4936
rect 4828 4772 4948 4936
rect 5724 4772 5844 4936
rect 6172 4772 6372 4936
rect 6956 4772 7076 4936
rect 7628 4772 7748 4936
rect 8300 4772 8420 4936
rect 8748 4772 8948 4936
rect 9308 4772 9428 4936
rect 10060 4772 10180 4936
rect 1916 4472 2036 4636
rect 2588 4472 2708 4636
rect 3260 4472 3380 4636
rect 3932 4472 4052 4636
rect 4604 4472 4724 4636
rect 5052 4472 5252 4636
rect 5724 4472 5844 4636
rect 6396 4472 6516 4636
rect 7068 4472 7188 4636
rect 7740 4472 7860 4636
rect 8412 4472 8532 4636
rect 8860 4472 9060 4636
rect 9980 4472 10100 4636
rect 1996 3204 2116 3368
rect 2588 3204 2708 3368
rect 3260 3204 3380 3368
rect 3932 3204 4052 3368
rect 4604 3204 4724 3368
rect 5724 3204 5844 3368
rect 6172 3204 6372 3368
rect 6620 3204 6740 3368
rect 7292 3204 7412 3368
rect 8044 3204 8164 3368
rect 8636 3204 8756 3368
rect 9532 3204 9732 3368
rect 9980 3204 10100 3368
<< mvpmos >>
rect 1692 8312 1892 8556
rect 2160 8312 2260 8556
rect 2832 8312 2932 8556
rect 3504 8312 3604 8556
rect 4176 8312 4276 8556
rect 4848 8312 4948 8556
rect 5612 8312 5812 8556
rect 6060 8312 6260 8556
rect 6508 8312 6708 8556
rect 6956 8312 7156 8556
rect 7404 8312 7604 8556
rect 7852 8312 8052 8556
rect 8300 8312 8500 8556
rect 8748 8312 8948 8556
rect 9532 8312 9732 8556
rect 9980 8312 10180 8556
rect 1692 7124 1892 7368
rect 2160 7124 2260 7368
rect 2832 7124 2932 7368
rect 3504 7124 3604 7368
rect 4176 7124 4276 7368
rect 4848 7124 4948 7368
rect 5580 7124 5680 7368
rect 6252 7124 6352 7368
rect 6620 7124 6820 7368
rect 7068 7124 7268 7368
rect 7516 7124 7716 7368
rect 7964 7124 8164 7368
rect 8412 7124 8612 7368
rect 8860 7124 9060 7368
rect 10060 7124 10160 7368
rect 1936 6744 2036 6988
rect 2608 6744 2708 6988
rect 3280 6744 3380 6988
rect 3952 6744 4052 6988
rect 4624 6744 4724 6988
rect 5744 6744 5844 6988
rect 6416 6744 6516 6988
rect 7088 6744 7188 6988
rect 7516 6744 7716 6988
rect 7964 6744 8164 6988
rect 8432 6744 8532 6988
rect 9104 6876 9204 6988
rect 9308 6876 9408 6988
rect 9588 6744 9688 6988
rect 9792 6744 9892 6988
rect 9996 6744 10096 6988
rect 1824 5556 1924 5800
rect 2496 5556 2596 5800
rect 3168 5556 3268 5800
rect 3840 5556 3940 5800
rect 4512 5556 4612 5800
rect 5184 5556 5284 5800
rect 5856 5556 5956 5800
rect 6528 5556 6628 5800
rect 6956 5556 7156 5800
rect 7760 5556 7860 5800
rect 8432 5556 8532 5800
rect 8860 5556 9060 5800
rect 10060 5556 10160 5800
rect 1692 5176 1892 5420
rect 2160 5176 2260 5420
rect 2832 5176 2932 5420
rect 3504 5176 3604 5420
rect 4176 5176 4276 5420
rect 4848 5176 4948 5420
rect 5744 5176 5844 5420
rect 6172 5176 6372 5420
rect 6976 5176 7076 5420
rect 7648 5176 7748 5420
rect 8320 5176 8420 5420
rect 8748 5176 8948 5420
rect 9328 5176 9428 5420
rect 10060 5176 10160 5420
rect 1936 3988 2036 4232
rect 2608 3988 2708 4232
rect 3280 3988 3380 4232
rect 3952 3988 4052 4232
rect 4624 3988 4724 4232
rect 5052 3988 5252 4232
rect 5744 3988 5844 4232
rect 6416 3988 6516 4232
rect 7088 3988 7188 4232
rect 7760 3988 7860 4232
rect 8432 3988 8532 4232
rect 8860 3988 9060 4232
rect 10000 3988 10100 4232
rect 1996 3608 2096 3852
rect 2608 3608 2708 3852
rect 3280 3608 3380 3852
rect 3952 3608 4052 3852
rect 4624 3608 4724 3852
rect 5744 3608 5844 3852
rect 6172 3608 6372 3852
rect 6640 3608 6740 3852
rect 7312 3608 7412 3852
rect 8044 3608 8144 3852
rect 8656 3608 8756 3852
rect 9532 3608 9732 3852
rect 10000 3608 10100 3852
<< mvndiff >>
rect 1604 8032 1692 8072
rect 1604 7986 1617 8032
rect 1663 7986 1692 8032
rect 1604 7908 1692 7986
rect 1892 8032 1980 8072
rect 1892 7986 1921 8032
rect 1967 7986 1980 8032
rect 1892 7908 1980 7986
rect 2052 8032 2140 8072
rect 2052 7986 2065 8032
rect 2111 7986 2140 8032
rect 2052 7908 2140 7986
rect 2260 8032 2348 8072
rect 2260 7986 2289 8032
rect 2335 7986 2348 8032
rect 2260 7908 2348 7986
rect 2724 8032 2812 8072
rect 2724 7986 2737 8032
rect 2783 7986 2812 8032
rect 2724 7908 2812 7986
rect 2932 8032 3020 8072
rect 2932 7986 2961 8032
rect 3007 7986 3020 8032
rect 2932 7908 3020 7986
rect 3396 8032 3484 8072
rect 3396 7986 3409 8032
rect 3455 7986 3484 8032
rect 3396 7908 3484 7986
rect 3604 8032 3692 8072
rect 3604 7986 3633 8032
rect 3679 7986 3692 8032
rect 3604 7908 3692 7986
rect 4068 8032 4156 8072
rect 4068 7986 4081 8032
rect 4127 7986 4156 8032
rect 4068 7908 4156 7986
rect 4276 8032 4364 8072
rect 4276 7986 4305 8032
rect 4351 7986 4364 8032
rect 4276 7908 4364 7986
rect 4740 8032 4828 8072
rect 4740 7986 4753 8032
rect 4799 7986 4828 8032
rect 4740 7908 4828 7986
rect 4948 8032 5036 8072
rect 4948 7986 4977 8032
rect 5023 7986 5036 8032
rect 4948 7908 5036 7986
rect 5524 8032 5612 8072
rect 5524 7986 5537 8032
rect 5583 7986 5612 8032
rect 5524 7908 5612 7986
rect 5812 8032 5900 8072
rect 5812 7986 5841 8032
rect 5887 7986 5900 8032
rect 5812 7908 5900 7986
rect 5972 8032 6060 8072
rect 5972 7986 5985 8032
rect 6031 7986 6060 8032
rect 5972 7908 6060 7986
rect 6260 8032 6348 8072
rect 6260 7986 6289 8032
rect 6335 7986 6348 8032
rect 6260 7908 6348 7986
rect 6420 8032 6508 8072
rect 6420 7986 6433 8032
rect 6479 7986 6508 8032
rect 6420 7908 6508 7986
rect 6708 8032 6796 8072
rect 6708 7986 6737 8032
rect 6783 7986 6796 8032
rect 6708 7908 6796 7986
rect 6868 8032 6956 8072
rect 6868 7986 6881 8032
rect 6927 7986 6956 8032
rect 6868 7908 6956 7986
rect 7156 8032 7244 8072
rect 7156 7986 7185 8032
rect 7231 7986 7244 8032
rect 7156 7908 7244 7986
rect 7316 8032 7404 8072
rect 7316 7986 7329 8032
rect 7375 7986 7404 8032
rect 7316 7908 7404 7986
rect 7604 8032 7692 8072
rect 7604 7986 7633 8032
rect 7679 7986 7692 8032
rect 7604 7908 7692 7986
rect 7764 8032 7852 8072
rect 7764 7986 7777 8032
rect 7823 7986 7852 8032
rect 7764 7908 7852 7986
rect 8052 8032 8140 8072
rect 8052 7986 8081 8032
rect 8127 7986 8140 8032
rect 8052 7908 8140 7986
rect 8212 8032 8300 8072
rect 8212 7986 8225 8032
rect 8271 7986 8300 8032
rect 8212 7908 8300 7986
rect 8500 8032 8588 8072
rect 8500 7986 8529 8032
rect 8575 7986 8588 8032
rect 8500 7908 8588 7986
rect 8660 8032 8748 8072
rect 8660 7986 8673 8032
rect 8719 7986 8748 8032
rect 8660 7908 8748 7986
rect 8948 8032 9036 8072
rect 8948 7986 8977 8032
rect 9023 7986 9036 8032
rect 8948 7908 9036 7986
rect 9444 8032 9532 8072
rect 9444 7986 9457 8032
rect 9503 7986 9532 8032
rect 9444 7908 9532 7986
rect 9732 8032 9820 8072
rect 9732 7986 9761 8032
rect 9807 7986 9820 8032
rect 9732 7908 9820 7986
rect 9892 8032 9980 8072
rect 9892 7986 9905 8032
rect 9951 7986 9980 8032
rect 9892 7908 9980 7986
rect 10180 8032 10268 8072
rect 10180 7986 10209 8032
rect 10255 7986 10268 8032
rect 10180 7908 10268 7986
rect 1604 7694 1692 7772
rect 1604 7648 1617 7694
rect 1663 7648 1692 7694
rect 1604 7608 1692 7648
rect 1892 7694 1980 7772
rect 1892 7648 1921 7694
rect 1967 7648 1980 7694
rect 1892 7608 1980 7648
rect 2052 7694 2140 7772
rect 2052 7648 2065 7694
rect 2111 7648 2140 7694
rect 2052 7608 2140 7648
rect 2260 7694 2348 7772
rect 2260 7648 2289 7694
rect 2335 7648 2348 7694
rect 2260 7608 2348 7648
rect 2724 7694 2812 7772
rect 2724 7648 2737 7694
rect 2783 7648 2812 7694
rect 2724 7608 2812 7648
rect 2932 7694 3020 7772
rect 2932 7648 2961 7694
rect 3007 7648 3020 7694
rect 2932 7608 3020 7648
rect 3396 7694 3484 7772
rect 3396 7648 3409 7694
rect 3455 7648 3484 7694
rect 3396 7608 3484 7648
rect 3604 7694 3692 7772
rect 3604 7648 3633 7694
rect 3679 7648 3692 7694
rect 3604 7608 3692 7648
rect 4068 7694 4156 7772
rect 4068 7648 4081 7694
rect 4127 7648 4156 7694
rect 4068 7608 4156 7648
rect 4276 7694 4364 7772
rect 4276 7648 4305 7694
rect 4351 7648 4364 7694
rect 4276 7608 4364 7648
rect 4740 7694 4828 7772
rect 4740 7648 4753 7694
rect 4799 7648 4828 7694
rect 4740 7608 4828 7648
rect 4948 7694 5036 7772
rect 4948 7648 4977 7694
rect 5023 7648 5036 7694
rect 4948 7608 5036 7648
rect 5492 7694 5580 7772
rect 5492 7648 5505 7694
rect 5551 7648 5580 7694
rect 5492 7608 5580 7648
rect 5700 7694 5788 7772
rect 5700 7648 5729 7694
rect 5775 7648 5788 7694
rect 5700 7608 5788 7648
rect 6164 7694 6252 7772
rect 6164 7648 6177 7694
rect 6223 7648 6252 7694
rect 6164 7608 6252 7648
rect 6372 7694 6460 7772
rect 6372 7648 6401 7694
rect 6447 7648 6460 7694
rect 6372 7608 6460 7648
rect 6532 7694 6620 7772
rect 6532 7648 6545 7694
rect 6591 7648 6620 7694
rect 6532 7608 6620 7648
rect 6820 7694 6908 7772
rect 6820 7648 6849 7694
rect 6895 7648 6908 7694
rect 6820 7608 6908 7648
rect 6980 7694 7068 7772
rect 6980 7648 6993 7694
rect 7039 7648 7068 7694
rect 6980 7608 7068 7648
rect 7268 7694 7356 7772
rect 7268 7648 7297 7694
rect 7343 7648 7356 7694
rect 7268 7608 7356 7648
rect 7428 7694 7516 7772
rect 7428 7648 7441 7694
rect 7487 7648 7516 7694
rect 7428 7608 7516 7648
rect 7716 7694 7804 7772
rect 7716 7648 7745 7694
rect 7791 7648 7804 7694
rect 7716 7608 7804 7648
rect 7876 7694 7964 7772
rect 7876 7648 7889 7694
rect 7935 7648 7964 7694
rect 7876 7608 7964 7648
rect 8164 7694 8252 7772
rect 8164 7648 8193 7694
rect 8239 7648 8252 7694
rect 8164 7608 8252 7648
rect 8324 7694 8412 7772
rect 8324 7648 8337 7694
rect 8383 7648 8412 7694
rect 8324 7608 8412 7648
rect 8612 7694 8700 7772
rect 8612 7648 8641 7694
rect 8687 7648 8700 7694
rect 8612 7608 8700 7648
rect 8772 7694 8860 7772
rect 8772 7648 8785 7694
rect 8831 7648 8860 7694
rect 8772 7608 8860 7648
rect 9060 7694 9148 7772
rect 9060 7648 9089 7694
rect 9135 7648 9148 7694
rect 9060 7608 9148 7648
rect 9972 7694 10060 7772
rect 9972 7648 9985 7694
rect 10031 7648 10060 7694
rect 9972 7608 10060 7648
rect 10180 7694 10268 7772
rect 10180 7648 10209 7694
rect 10255 7648 10268 7694
rect 10180 7608 10268 7648
rect 1828 6464 1916 6504
rect 1828 6418 1841 6464
rect 1887 6418 1916 6464
rect 1828 6340 1916 6418
rect 2036 6464 2124 6504
rect 2036 6418 2065 6464
rect 2111 6418 2124 6464
rect 2036 6340 2124 6418
rect 2500 6464 2588 6504
rect 2500 6418 2513 6464
rect 2559 6418 2588 6464
rect 2500 6340 2588 6418
rect 2708 6464 2796 6504
rect 2708 6418 2737 6464
rect 2783 6418 2796 6464
rect 2708 6340 2796 6418
rect 3172 6464 3260 6504
rect 3172 6418 3185 6464
rect 3231 6418 3260 6464
rect 3172 6340 3260 6418
rect 3380 6464 3468 6504
rect 3380 6418 3409 6464
rect 3455 6418 3468 6464
rect 3380 6340 3468 6418
rect 3844 6464 3932 6504
rect 3844 6418 3857 6464
rect 3903 6418 3932 6464
rect 3844 6340 3932 6418
rect 4052 6464 4140 6504
rect 4052 6418 4081 6464
rect 4127 6418 4140 6464
rect 4052 6340 4140 6418
rect 4516 6464 4604 6504
rect 4516 6418 4529 6464
rect 4575 6418 4604 6464
rect 4516 6340 4604 6418
rect 4724 6464 4812 6504
rect 4724 6418 4753 6464
rect 4799 6418 4812 6464
rect 4724 6340 4812 6418
rect 5636 6464 5724 6504
rect 5636 6418 5649 6464
rect 5695 6418 5724 6464
rect 5636 6340 5724 6418
rect 5844 6464 5932 6504
rect 5844 6418 5873 6464
rect 5919 6418 5932 6464
rect 5844 6340 5932 6418
rect 6308 6464 6396 6504
rect 6308 6418 6321 6464
rect 6367 6418 6396 6464
rect 6308 6340 6396 6418
rect 6516 6464 6604 6504
rect 6516 6418 6545 6464
rect 6591 6418 6604 6464
rect 6516 6340 6604 6418
rect 6980 6464 7068 6504
rect 6980 6418 6993 6464
rect 7039 6418 7068 6464
rect 6980 6340 7068 6418
rect 7188 6464 7276 6504
rect 7188 6418 7217 6464
rect 7263 6418 7276 6464
rect 7188 6340 7276 6418
rect 7428 6464 7516 6504
rect 7428 6418 7441 6464
rect 7487 6418 7516 6464
rect 7428 6340 7516 6418
rect 7716 6464 7804 6504
rect 7716 6418 7745 6464
rect 7791 6418 7804 6464
rect 7716 6340 7804 6418
rect 7876 6464 7964 6504
rect 7876 6418 7889 6464
rect 7935 6418 7964 6464
rect 7876 6340 7964 6418
rect 8164 6464 8252 6504
rect 8164 6418 8193 6464
rect 8239 6418 8252 6464
rect 8164 6340 8252 6418
rect 8324 6464 8412 6504
rect 8324 6418 8337 6464
rect 8383 6418 8412 6464
rect 8324 6340 8412 6418
rect 8532 6464 8620 6504
rect 8532 6418 8561 6464
rect 8607 6418 8620 6464
rect 9488 6437 9568 6504
rect 8532 6340 8620 6418
rect 8996 6424 9084 6437
rect 8996 6378 9009 6424
rect 9055 6378 9084 6424
rect 8996 6365 9084 6378
rect 9204 6424 9308 6437
rect 9204 6378 9233 6424
rect 9279 6378 9308 6424
rect 9204 6365 9308 6378
rect 9428 6424 9568 6437
rect 9428 6378 9493 6424
rect 9539 6378 9568 6424
rect 9428 6365 9568 6378
rect 9488 6340 9568 6365
rect 9688 6441 9792 6504
rect 9688 6395 9717 6441
rect 9763 6395 9792 6441
rect 9688 6340 9792 6395
rect 9912 6340 9976 6504
rect 10096 6399 10184 6504
rect 10096 6353 10125 6399
rect 10171 6353 10184 6399
rect 10096 6340 10184 6353
rect 1716 6126 1804 6204
rect 1716 6080 1729 6126
rect 1775 6080 1804 6126
rect 1716 6040 1804 6080
rect 1924 6126 2012 6204
rect 1924 6080 1953 6126
rect 1999 6080 2012 6126
rect 1924 6040 2012 6080
rect 2388 6126 2476 6204
rect 2388 6080 2401 6126
rect 2447 6080 2476 6126
rect 2388 6040 2476 6080
rect 2596 6126 2684 6204
rect 2596 6080 2625 6126
rect 2671 6080 2684 6126
rect 2596 6040 2684 6080
rect 3060 6126 3148 6204
rect 3060 6080 3073 6126
rect 3119 6080 3148 6126
rect 3060 6040 3148 6080
rect 3268 6126 3356 6204
rect 3268 6080 3297 6126
rect 3343 6080 3356 6126
rect 3268 6040 3356 6080
rect 3732 6126 3820 6204
rect 3732 6080 3745 6126
rect 3791 6080 3820 6126
rect 3732 6040 3820 6080
rect 3940 6126 4028 6204
rect 3940 6080 3969 6126
rect 4015 6080 4028 6126
rect 3940 6040 4028 6080
rect 4404 6126 4492 6204
rect 4404 6080 4417 6126
rect 4463 6080 4492 6126
rect 4404 6040 4492 6080
rect 4612 6126 4700 6204
rect 4612 6080 4641 6126
rect 4687 6080 4700 6126
rect 4612 6040 4700 6080
rect 5076 6126 5164 6204
rect 5076 6080 5089 6126
rect 5135 6080 5164 6126
rect 5076 6040 5164 6080
rect 5284 6126 5372 6204
rect 5284 6080 5313 6126
rect 5359 6080 5372 6126
rect 5284 6040 5372 6080
rect 5748 6126 5836 6204
rect 5748 6080 5761 6126
rect 5807 6080 5836 6126
rect 5748 6040 5836 6080
rect 5956 6126 6044 6204
rect 5956 6080 5985 6126
rect 6031 6080 6044 6126
rect 5956 6040 6044 6080
rect 6420 6126 6508 6204
rect 6420 6080 6433 6126
rect 6479 6080 6508 6126
rect 6420 6040 6508 6080
rect 6628 6126 6716 6204
rect 6628 6080 6657 6126
rect 6703 6080 6716 6126
rect 6628 6040 6716 6080
rect 6868 6126 6956 6204
rect 6868 6080 6881 6126
rect 6927 6080 6956 6126
rect 6868 6040 6956 6080
rect 7156 6126 7244 6204
rect 7156 6080 7185 6126
rect 7231 6080 7244 6126
rect 7156 6040 7244 6080
rect 7652 6126 7740 6204
rect 7652 6080 7665 6126
rect 7711 6080 7740 6126
rect 7652 6040 7740 6080
rect 7860 6126 7948 6204
rect 7860 6080 7889 6126
rect 7935 6080 7948 6126
rect 7860 6040 7948 6080
rect 8324 6126 8412 6204
rect 8324 6080 8337 6126
rect 8383 6080 8412 6126
rect 8324 6040 8412 6080
rect 8532 6126 8620 6204
rect 8532 6080 8561 6126
rect 8607 6080 8620 6126
rect 8532 6040 8620 6080
rect 8772 6126 8860 6204
rect 8772 6080 8785 6126
rect 8831 6080 8860 6126
rect 8772 6040 8860 6080
rect 9060 6126 9148 6204
rect 9060 6080 9089 6126
rect 9135 6080 9148 6126
rect 9060 6040 9148 6080
rect 9972 6126 10060 6204
rect 9972 6080 9985 6126
rect 10031 6080 10060 6126
rect 9972 6040 10060 6080
rect 10180 6126 10268 6204
rect 10180 6080 10209 6126
rect 10255 6080 10268 6126
rect 10180 6040 10268 6080
rect 1604 4896 1692 4936
rect 1604 4850 1617 4896
rect 1663 4850 1692 4896
rect 1604 4772 1692 4850
rect 1892 4896 1980 4936
rect 1892 4850 1921 4896
rect 1967 4850 1980 4896
rect 1892 4772 1980 4850
rect 2052 4896 2140 4936
rect 2052 4850 2065 4896
rect 2111 4850 2140 4896
rect 2052 4772 2140 4850
rect 2260 4896 2348 4936
rect 2260 4850 2289 4896
rect 2335 4850 2348 4896
rect 2260 4772 2348 4850
rect 2724 4896 2812 4936
rect 2724 4850 2737 4896
rect 2783 4850 2812 4896
rect 2724 4772 2812 4850
rect 2932 4896 3020 4936
rect 2932 4850 2961 4896
rect 3007 4850 3020 4896
rect 2932 4772 3020 4850
rect 3396 4896 3484 4936
rect 3396 4850 3409 4896
rect 3455 4850 3484 4896
rect 3396 4772 3484 4850
rect 3604 4896 3692 4936
rect 3604 4850 3633 4896
rect 3679 4850 3692 4896
rect 3604 4772 3692 4850
rect 4068 4896 4156 4936
rect 4068 4850 4081 4896
rect 4127 4850 4156 4896
rect 4068 4772 4156 4850
rect 4276 4896 4364 4936
rect 4276 4850 4305 4896
rect 4351 4850 4364 4896
rect 4276 4772 4364 4850
rect 4740 4896 4828 4936
rect 4740 4850 4753 4896
rect 4799 4850 4828 4896
rect 4740 4772 4828 4850
rect 4948 4896 5036 4936
rect 4948 4850 4977 4896
rect 5023 4850 5036 4896
rect 4948 4772 5036 4850
rect 5636 4896 5724 4936
rect 5636 4850 5649 4896
rect 5695 4850 5724 4896
rect 5636 4772 5724 4850
rect 5844 4896 5932 4936
rect 5844 4850 5873 4896
rect 5919 4850 5932 4896
rect 5844 4772 5932 4850
rect 6084 4896 6172 4936
rect 6084 4850 6097 4896
rect 6143 4850 6172 4896
rect 6084 4772 6172 4850
rect 6372 4896 6460 4936
rect 6372 4850 6401 4896
rect 6447 4850 6460 4896
rect 6372 4772 6460 4850
rect 6868 4896 6956 4936
rect 6868 4850 6881 4896
rect 6927 4850 6956 4896
rect 6868 4772 6956 4850
rect 7076 4896 7164 4936
rect 7076 4850 7105 4896
rect 7151 4850 7164 4896
rect 7076 4772 7164 4850
rect 7540 4896 7628 4936
rect 7540 4850 7553 4896
rect 7599 4850 7628 4896
rect 7540 4772 7628 4850
rect 7748 4896 7836 4936
rect 7748 4850 7777 4896
rect 7823 4850 7836 4896
rect 7748 4772 7836 4850
rect 8212 4896 8300 4936
rect 8212 4850 8225 4896
rect 8271 4850 8300 4896
rect 8212 4772 8300 4850
rect 8420 4896 8508 4936
rect 8420 4850 8449 4896
rect 8495 4850 8508 4896
rect 8420 4772 8508 4850
rect 8660 4896 8748 4936
rect 8660 4850 8673 4896
rect 8719 4850 8748 4896
rect 8660 4772 8748 4850
rect 8948 4896 9036 4936
rect 8948 4850 8977 4896
rect 9023 4850 9036 4896
rect 8948 4772 9036 4850
rect 9220 4896 9308 4936
rect 9220 4850 9233 4896
rect 9279 4850 9308 4896
rect 9220 4772 9308 4850
rect 9428 4896 9516 4936
rect 9428 4850 9457 4896
rect 9503 4850 9516 4896
rect 9428 4772 9516 4850
rect 9972 4896 10060 4936
rect 9972 4850 9985 4896
rect 10031 4850 10060 4896
rect 9972 4772 10060 4850
rect 10180 4896 10268 4936
rect 10180 4850 10209 4896
rect 10255 4850 10268 4896
rect 10180 4772 10268 4850
rect 1828 4558 1916 4636
rect 1828 4512 1841 4558
rect 1887 4512 1916 4558
rect 1828 4472 1916 4512
rect 2036 4558 2124 4636
rect 2036 4512 2065 4558
rect 2111 4512 2124 4558
rect 2036 4472 2124 4512
rect 2500 4558 2588 4636
rect 2500 4512 2513 4558
rect 2559 4512 2588 4558
rect 2500 4472 2588 4512
rect 2708 4558 2796 4636
rect 2708 4512 2737 4558
rect 2783 4512 2796 4558
rect 2708 4472 2796 4512
rect 3172 4558 3260 4636
rect 3172 4512 3185 4558
rect 3231 4512 3260 4558
rect 3172 4472 3260 4512
rect 3380 4558 3468 4636
rect 3380 4512 3409 4558
rect 3455 4512 3468 4558
rect 3380 4472 3468 4512
rect 3844 4558 3932 4636
rect 3844 4512 3857 4558
rect 3903 4512 3932 4558
rect 3844 4472 3932 4512
rect 4052 4558 4140 4636
rect 4052 4512 4081 4558
rect 4127 4512 4140 4558
rect 4052 4472 4140 4512
rect 4516 4558 4604 4636
rect 4516 4512 4529 4558
rect 4575 4512 4604 4558
rect 4516 4472 4604 4512
rect 4724 4558 4812 4636
rect 4724 4512 4753 4558
rect 4799 4512 4812 4558
rect 4724 4472 4812 4512
rect 4964 4558 5052 4636
rect 4964 4512 4977 4558
rect 5023 4512 5052 4558
rect 4964 4472 5052 4512
rect 5252 4558 5340 4636
rect 5252 4512 5281 4558
rect 5327 4512 5340 4558
rect 5252 4472 5340 4512
rect 5636 4558 5724 4636
rect 5636 4512 5649 4558
rect 5695 4512 5724 4558
rect 5636 4472 5724 4512
rect 5844 4558 5932 4636
rect 5844 4512 5873 4558
rect 5919 4512 5932 4558
rect 5844 4472 5932 4512
rect 6308 4558 6396 4636
rect 6308 4512 6321 4558
rect 6367 4512 6396 4558
rect 6308 4472 6396 4512
rect 6516 4558 6604 4636
rect 6516 4512 6545 4558
rect 6591 4512 6604 4558
rect 6516 4472 6604 4512
rect 6980 4558 7068 4636
rect 6980 4512 6993 4558
rect 7039 4512 7068 4558
rect 6980 4472 7068 4512
rect 7188 4558 7276 4636
rect 7188 4512 7217 4558
rect 7263 4512 7276 4558
rect 7188 4472 7276 4512
rect 7652 4558 7740 4636
rect 7652 4512 7665 4558
rect 7711 4512 7740 4558
rect 7652 4472 7740 4512
rect 7860 4558 7948 4636
rect 7860 4512 7889 4558
rect 7935 4512 7948 4558
rect 7860 4472 7948 4512
rect 8324 4558 8412 4636
rect 8324 4512 8337 4558
rect 8383 4512 8412 4558
rect 8324 4472 8412 4512
rect 8532 4558 8620 4636
rect 8532 4512 8561 4558
rect 8607 4512 8620 4558
rect 8532 4472 8620 4512
rect 8772 4558 8860 4636
rect 8772 4512 8785 4558
rect 8831 4512 8860 4558
rect 8772 4472 8860 4512
rect 9060 4558 9148 4636
rect 9060 4512 9089 4558
rect 9135 4512 9148 4558
rect 9060 4472 9148 4512
rect 9892 4558 9980 4636
rect 9892 4512 9905 4558
rect 9951 4512 9980 4558
rect 9892 4472 9980 4512
rect 10100 4558 10188 4636
rect 10100 4512 10129 4558
rect 10175 4512 10188 4558
rect 10100 4472 10188 4512
rect 1908 3328 1996 3368
rect 1908 3282 1921 3328
rect 1967 3282 1996 3328
rect 1908 3204 1996 3282
rect 2116 3328 2204 3368
rect 2116 3282 2145 3328
rect 2191 3282 2204 3328
rect 2116 3204 2204 3282
rect 2500 3328 2588 3368
rect 2500 3282 2513 3328
rect 2559 3282 2588 3328
rect 2500 3204 2588 3282
rect 2708 3328 2796 3368
rect 2708 3282 2737 3328
rect 2783 3282 2796 3328
rect 2708 3204 2796 3282
rect 3172 3328 3260 3368
rect 3172 3282 3185 3328
rect 3231 3282 3260 3328
rect 3172 3204 3260 3282
rect 3380 3328 3468 3368
rect 3380 3282 3409 3328
rect 3455 3282 3468 3328
rect 3380 3204 3468 3282
rect 3844 3328 3932 3368
rect 3844 3282 3857 3328
rect 3903 3282 3932 3328
rect 3844 3204 3932 3282
rect 4052 3328 4140 3368
rect 4052 3282 4081 3328
rect 4127 3282 4140 3328
rect 4052 3204 4140 3282
rect 4516 3328 4604 3368
rect 4516 3282 4529 3328
rect 4575 3282 4604 3328
rect 4516 3204 4604 3282
rect 4724 3328 4812 3368
rect 4724 3282 4753 3328
rect 4799 3282 4812 3328
rect 4724 3204 4812 3282
rect 5636 3328 5724 3368
rect 5636 3282 5649 3328
rect 5695 3282 5724 3328
rect 5636 3204 5724 3282
rect 5844 3328 5932 3368
rect 5844 3282 5873 3328
rect 5919 3282 5932 3328
rect 5844 3204 5932 3282
rect 6084 3328 6172 3368
rect 6084 3282 6097 3328
rect 6143 3282 6172 3328
rect 6084 3204 6172 3282
rect 6372 3328 6460 3368
rect 6372 3282 6401 3328
rect 6447 3282 6460 3328
rect 6372 3204 6460 3282
rect 6532 3328 6620 3368
rect 6532 3282 6545 3328
rect 6591 3282 6620 3328
rect 6532 3204 6620 3282
rect 6740 3328 6828 3368
rect 6740 3282 6769 3328
rect 6815 3282 6828 3328
rect 6740 3204 6828 3282
rect 7204 3328 7292 3368
rect 7204 3282 7217 3328
rect 7263 3282 7292 3328
rect 7204 3204 7292 3282
rect 7412 3328 7500 3368
rect 7412 3282 7441 3328
rect 7487 3282 7500 3328
rect 7412 3204 7500 3282
rect 7956 3328 8044 3368
rect 7956 3282 7969 3328
rect 8015 3282 8044 3328
rect 7956 3204 8044 3282
rect 8164 3328 8252 3368
rect 8164 3282 8193 3328
rect 8239 3282 8252 3328
rect 8164 3204 8252 3282
rect 8548 3328 8636 3368
rect 8548 3282 8561 3328
rect 8607 3282 8636 3328
rect 8548 3204 8636 3282
rect 8756 3328 8844 3368
rect 8756 3282 8785 3328
rect 8831 3282 8844 3328
rect 8756 3204 8844 3282
rect 9444 3328 9532 3368
rect 9444 3282 9457 3328
rect 9503 3282 9532 3328
rect 9444 3204 9532 3282
rect 9732 3328 9820 3368
rect 9732 3282 9761 3328
rect 9807 3282 9820 3328
rect 9732 3204 9820 3282
rect 9892 3328 9980 3368
rect 9892 3282 9905 3328
rect 9951 3282 9980 3328
rect 9892 3204 9980 3282
rect 10100 3328 10188 3368
rect 10100 3282 10129 3328
rect 10175 3282 10188 3328
rect 10100 3204 10188 3282
<< mvpdiff >>
rect 1604 8497 1692 8556
rect 1604 8357 1617 8497
rect 1663 8357 1692 8497
rect 1604 8312 1692 8357
rect 1892 8497 1980 8556
rect 1892 8357 1921 8497
rect 1967 8357 1980 8497
rect 1892 8312 1980 8357
rect 2072 8505 2160 8556
rect 2072 8365 2085 8505
rect 2131 8365 2160 8505
rect 2072 8312 2160 8365
rect 2260 8505 2348 8556
rect 2260 8365 2289 8505
rect 2335 8365 2348 8505
rect 2260 8312 2348 8365
rect 2744 8505 2832 8556
rect 2744 8365 2757 8505
rect 2803 8365 2832 8505
rect 2744 8312 2832 8365
rect 2932 8505 3020 8556
rect 2932 8365 2961 8505
rect 3007 8365 3020 8505
rect 2932 8312 3020 8365
rect 3416 8505 3504 8556
rect 3416 8365 3429 8505
rect 3475 8365 3504 8505
rect 3416 8312 3504 8365
rect 3604 8505 3692 8556
rect 3604 8365 3633 8505
rect 3679 8365 3692 8505
rect 3604 8312 3692 8365
rect 4088 8505 4176 8556
rect 4088 8365 4101 8505
rect 4147 8365 4176 8505
rect 4088 8312 4176 8365
rect 4276 8505 4364 8556
rect 4276 8365 4305 8505
rect 4351 8365 4364 8505
rect 4276 8312 4364 8365
rect 4760 8505 4848 8556
rect 4760 8365 4773 8505
rect 4819 8365 4848 8505
rect 4760 8312 4848 8365
rect 4948 8505 5036 8556
rect 4948 8365 4977 8505
rect 5023 8365 5036 8505
rect 4948 8312 5036 8365
rect 5524 8497 5612 8556
rect 5524 8357 5537 8497
rect 5583 8357 5612 8497
rect 5524 8312 5612 8357
rect 5812 8497 5900 8556
rect 5812 8357 5841 8497
rect 5887 8357 5900 8497
rect 5812 8312 5900 8357
rect 5972 8497 6060 8556
rect 5972 8357 5985 8497
rect 6031 8357 6060 8497
rect 5972 8312 6060 8357
rect 6260 8497 6348 8556
rect 6260 8357 6289 8497
rect 6335 8357 6348 8497
rect 6260 8312 6348 8357
rect 6420 8497 6508 8556
rect 6420 8357 6433 8497
rect 6479 8357 6508 8497
rect 6420 8312 6508 8357
rect 6708 8497 6796 8556
rect 6708 8357 6737 8497
rect 6783 8357 6796 8497
rect 6708 8312 6796 8357
rect 6868 8497 6956 8556
rect 6868 8357 6881 8497
rect 6927 8357 6956 8497
rect 6868 8312 6956 8357
rect 7156 8497 7244 8556
rect 7156 8357 7185 8497
rect 7231 8357 7244 8497
rect 7156 8312 7244 8357
rect 7316 8497 7404 8556
rect 7316 8357 7329 8497
rect 7375 8357 7404 8497
rect 7316 8312 7404 8357
rect 7604 8497 7692 8556
rect 7604 8357 7633 8497
rect 7679 8357 7692 8497
rect 7604 8312 7692 8357
rect 7764 8497 7852 8556
rect 7764 8357 7777 8497
rect 7823 8357 7852 8497
rect 7764 8312 7852 8357
rect 8052 8497 8140 8556
rect 8052 8357 8081 8497
rect 8127 8357 8140 8497
rect 8052 8312 8140 8357
rect 8212 8497 8300 8556
rect 8212 8357 8225 8497
rect 8271 8357 8300 8497
rect 8212 8312 8300 8357
rect 8500 8497 8588 8556
rect 8500 8357 8529 8497
rect 8575 8357 8588 8497
rect 8500 8312 8588 8357
rect 8660 8497 8748 8556
rect 8660 8357 8673 8497
rect 8719 8357 8748 8497
rect 8660 8312 8748 8357
rect 8948 8497 9036 8556
rect 8948 8357 8977 8497
rect 9023 8357 9036 8497
rect 8948 8312 9036 8357
rect 9444 8497 9532 8556
rect 9444 8357 9457 8497
rect 9503 8357 9532 8497
rect 9444 8312 9532 8357
rect 9732 8497 9820 8556
rect 9732 8357 9761 8497
rect 9807 8357 9820 8497
rect 9732 8312 9820 8357
rect 9892 8497 9980 8556
rect 9892 8357 9905 8497
rect 9951 8357 9980 8497
rect 9892 8312 9980 8357
rect 10180 8497 10268 8556
rect 10180 8357 10209 8497
rect 10255 8357 10268 8497
rect 10180 8312 10268 8357
rect 1604 7323 1692 7368
rect 1604 7183 1617 7323
rect 1663 7183 1692 7323
rect 1604 7124 1692 7183
rect 1892 7323 1980 7368
rect 1892 7183 1921 7323
rect 1967 7183 1980 7323
rect 1892 7124 1980 7183
rect 2072 7315 2160 7368
rect 2072 7175 2085 7315
rect 2131 7175 2160 7315
rect 2072 7124 2160 7175
rect 2260 7315 2348 7368
rect 2260 7175 2289 7315
rect 2335 7175 2348 7315
rect 2260 7124 2348 7175
rect 2744 7315 2832 7368
rect 2744 7175 2757 7315
rect 2803 7175 2832 7315
rect 2744 7124 2832 7175
rect 2932 7315 3020 7368
rect 2932 7175 2961 7315
rect 3007 7175 3020 7315
rect 2932 7124 3020 7175
rect 3416 7315 3504 7368
rect 3416 7175 3429 7315
rect 3475 7175 3504 7315
rect 3416 7124 3504 7175
rect 3604 7315 3692 7368
rect 3604 7175 3633 7315
rect 3679 7175 3692 7315
rect 3604 7124 3692 7175
rect 4088 7315 4176 7368
rect 4088 7175 4101 7315
rect 4147 7175 4176 7315
rect 4088 7124 4176 7175
rect 4276 7315 4364 7368
rect 4276 7175 4305 7315
rect 4351 7175 4364 7315
rect 4276 7124 4364 7175
rect 4760 7315 4848 7368
rect 4760 7175 4773 7315
rect 4819 7175 4848 7315
rect 4760 7124 4848 7175
rect 4948 7315 5036 7368
rect 4948 7175 4977 7315
rect 5023 7175 5036 7315
rect 4948 7124 5036 7175
rect 5492 7315 5580 7368
rect 5492 7175 5505 7315
rect 5551 7175 5580 7315
rect 5492 7124 5580 7175
rect 5680 7315 5768 7368
rect 5680 7175 5709 7315
rect 5755 7175 5768 7315
rect 5680 7124 5768 7175
rect 6164 7315 6252 7368
rect 6164 7175 6177 7315
rect 6223 7175 6252 7315
rect 6164 7124 6252 7175
rect 6352 7315 6440 7368
rect 6352 7175 6381 7315
rect 6427 7175 6440 7315
rect 6352 7124 6440 7175
rect 6532 7323 6620 7368
rect 6532 7183 6545 7323
rect 6591 7183 6620 7323
rect 6532 7124 6620 7183
rect 6820 7323 6908 7368
rect 6820 7183 6849 7323
rect 6895 7183 6908 7323
rect 6820 7124 6908 7183
rect 6980 7323 7068 7368
rect 6980 7183 6993 7323
rect 7039 7183 7068 7323
rect 6980 7124 7068 7183
rect 7268 7323 7356 7368
rect 7268 7183 7297 7323
rect 7343 7183 7356 7323
rect 7268 7124 7356 7183
rect 7428 7323 7516 7368
rect 7428 7183 7441 7323
rect 7487 7183 7516 7323
rect 7428 7124 7516 7183
rect 7716 7323 7804 7368
rect 7716 7183 7745 7323
rect 7791 7183 7804 7323
rect 7716 7124 7804 7183
rect 7876 7323 7964 7368
rect 7876 7183 7889 7323
rect 7935 7183 7964 7323
rect 7876 7124 7964 7183
rect 8164 7323 8252 7368
rect 8164 7183 8193 7323
rect 8239 7183 8252 7323
rect 8164 7124 8252 7183
rect 8324 7323 8412 7368
rect 8324 7183 8337 7323
rect 8383 7183 8412 7323
rect 8324 7124 8412 7183
rect 8612 7323 8700 7368
rect 8612 7183 8641 7323
rect 8687 7183 8700 7323
rect 8612 7124 8700 7183
rect 8772 7323 8860 7368
rect 8772 7183 8785 7323
rect 8831 7183 8860 7323
rect 8772 7124 8860 7183
rect 9060 7323 9148 7368
rect 9060 7183 9089 7323
rect 9135 7183 9148 7323
rect 9060 7124 9148 7183
rect 9972 7315 10060 7368
rect 9972 7175 9985 7315
rect 10031 7175 10060 7315
rect 9972 7124 10060 7175
rect 10160 7315 10248 7368
rect 10160 7175 10189 7315
rect 10235 7175 10248 7315
rect 10160 7124 10248 7175
rect 1848 6937 1936 6988
rect 1848 6797 1861 6937
rect 1907 6797 1936 6937
rect 1848 6744 1936 6797
rect 2036 6937 2124 6988
rect 2036 6797 2065 6937
rect 2111 6797 2124 6937
rect 2036 6744 2124 6797
rect 2520 6937 2608 6988
rect 2520 6797 2533 6937
rect 2579 6797 2608 6937
rect 2520 6744 2608 6797
rect 2708 6937 2796 6988
rect 2708 6797 2737 6937
rect 2783 6797 2796 6937
rect 2708 6744 2796 6797
rect 3192 6937 3280 6988
rect 3192 6797 3205 6937
rect 3251 6797 3280 6937
rect 3192 6744 3280 6797
rect 3380 6937 3468 6988
rect 3380 6797 3409 6937
rect 3455 6797 3468 6937
rect 3380 6744 3468 6797
rect 3864 6937 3952 6988
rect 3864 6797 3877 6937
rect 3923 6797 3952 6937
rect 3864 6744 3952 6797
rect 4052 6937 4140 6988
rect 4052 6797 4081 6937
rect 4127 6797 4140 6937
rect 4052 6744 4140 6797
rect 4536 6937 4624 6988
rect 4536 6797 4549 6937
rect 4595 6797 4624 6937
rect 4536 6744 4624 6797
rect 4724 6937 4812 6988
rect 4724 6797 4753 6937
rect 4799 6797 4812 6937
rect 4724 6744 4812 6797
rect 5656 6937 5744 6988
rect 5656 6797 5669 6937
rect 5715 6797 5744 6937
rect 5656 6744 5744 6797
rect 5844 6937 5932 6988
rect 5844 6797 5873 6937
rect 5919 6797 5932 6937
rect 5844 6744 5932 6797
rect 6328 6937 6416 6988
rect 6328 6797 6341 6937
rect 6387 6797 6416 6937
rect 6328 6744 6416 6797
rect 6516 6937 6604 6988
rect 6516 6797 6545 6937
rect 6591 6797 6604 6937
rect 6516 6744 6604 6797
rect 7000 6937 7088 6988
rect 7000 6797 7013 6937
rect 7059 6797 7088 6937
rect 7000 6744 7088 6797
rect 7188 6937 7276 6988
rect 7188 6797 7217 6937
rect 7263 6797 7276 6937
rect 7188 6744 7276 6797
rect 7428 6929 7516 6988
rect 7428 6789 7441 6929
rect 7487 6789 7516 6929
rect 7428 6744 7516 6789
rect 7716 6929 7804 6988
rect 7716 6789 7745 6929
rect 7791 6789 7804 6929
rect 7716 6744 7804 6789
rect 7876 6929 7964 6988
rect 7876 6789 7889 6929
rect 7935 6789 7964 6929
rect 7876 6744 7964 6789
rect 8164 6929 8252 6988
rect 8164 6789 8193 6929
rect 8239 6789 8252 6929
rect 8164 6744 8252 6789
rect 8344 6937 8432 6988
rect 8344 6797 8357 6937
rect 8403 6797 8432 6937
rect 8344 6744 8432 6797
rect 8532 6937 8620 6988
rect 8532 6797 8561 6937
rect 8607 6797 8620 6937
rect 9016 6941 9104 6988
rect 9016 6895 9029 6941
rect 9075 6895 9104 6941
rect 9016 6876 9104 6895
rect 9204 6876 9308 6988
rect 9408 6975 9588 6988
rect 9408 6876 9513 6975
rect 8532 6744 8620 6797
rect 9498 6835 9513 6876
rect 9559 6835 9588 6975
rect 9498 6744 9588 6835
rect 9688 6950 9792 6988
rect 9688 6904 9717 6950
rect 9763 6904 9792 6950
rect 9688 6744 9792 6904
rect 9892 6857 9996 6988
rect 9892 6811 9921 6857
rect 9967 6811 9996 6857
rect 9892 6744 9996 6811
rect 10096 6950 10184 6988
rect 10096 6904 10125 6950
rect 10171 6904 10184 6950
rect 10096 6744 10184 6904
rect 1736 5747 1824 5800
rect 1736 5607 1749 5747
rect 1795 5607 1824 5747
rect 1736 5556 1824 5607
rect 1924 5747 2012 5800
rect 1924 5607 1953 5747
rect 1999 5607 2012 5747
rect 1924 5556 2012 5607
rect 2408 5747 2496 5800
rect 2408 5607 2421 5747
rect 2467 5607 2496 5747
rect 2408 5556 2496 5607
rect 2596 5747 2684 5800
rect 2596 5607 2625 5747
rect 2671 5607 2684 5747
rect 2596 5556 2684 5607
rect 3080 5747 3168 5800
rect 3080 5607 3093 5747
rect 3139 5607 3168 5747
rect 3080 5556 3168 5607
rect 3268 5747 3356 5800
rect 3268 5607 3297 5747
rect 3343 5607 3356 5747
rect 3268 5556 3356 5607
rect 3752 5747 3840 5800
rect 3752 5607 3765 5747
rect 3811 5607 3840 5747
rect 3752 5556 3840 5607
rect 3940 5747 4028 5800
rect 3940 5607 3969 5747
rect 4015 5607 4028 5747
rect 3940 5556 4028 5607
rect 4424 5747 4512 5800
rect 4424 5607 4437 5747
rect 4483 5607 4512 5747
rect 4424 5556 4512 5607
rect 4612 5747 4700 5800
rect 4612 5607 4641 5747
rect 4687 5607 4700 5747
rect 4612 5556 4700 5607
rect 5096 5747 5184 5800
rect 5096 5607 5109 5747
rect 5155 5607 5184 5747
rect 5096 5556 5184 5607
rect 5284 5747 5372 5800
rect 5284 5607 5313 5747
rect 5359 5607 5372 5747
rect 5284 5556 5372 5607
rect 5768 5747 5856 5800
rect 5768 5607 5781 5747
rect 5827 5607 5856 5747
rect 5768 5556 5856 5607
rect 5956 5747 6044 5800
rect 5956 5607 5985 5747
rect 6031 5607 6044 5747
rect 5956 5556 6044 5607
rect 6440 5747 6528 5800
rect 6440 5607 6453 5747
rect 6499 5607 6528 5747
rect 6440 5556 6528 5607
rect 6628 5747 6716 5800
rect 6628 5607 6657 5747
rect 6703 5607 6716 5747
rect 6628 5556 6716 5607
rect 6868 5755 6956 5800
rect 6868 5615 6881 5755
rect 6927 5615 6956 5755
rect 6868 5556 6956 5615
rect 7156 5755 7244 5800
rect 7156 5615 7185 5755
rect 7231 5615 7244 5755
rect 7156 5556 7244 5615
rect 7672 5747 7760 5800
rect 7672 5607 7685 5747
rect 7731 5607 7760 5747
rect 7672 5556 7760 5607
rect 7860 5747 7948 5800
rect 7860 5607 7889 5747
rect 7935 5607 7948 5747
rect 7860 5556 7948 5607
rect 8344 5747 8432 5800
rect 8344 5607 8357 5747
rect 8403 5607 8432 5747
rect 8344 5556 8432 5607
rect 8532 5747 8620 5800
rect 8532 5607 8561 5747
rect 8607 5607 8620 5747
rect 8532 5556 8620 5607
rect 8772 5755 8860 5800
rect 8772 5615 8785 5755
rect 8831 5615 8860 5755
rect 8772 5556 8860 5615
rect 9060 5755 9148 5800
rect 9060 5615 9089 5755
rect 9135 5615 9148 5755
rect 9060 5556 9148 5615
rect 9972 5747 10060 5800
rect 9972 5607 9985 5747
rect 10031 5607 10060 5747
rect 9972 5556 10060 5607
rect 10160 5747 10248 5800
rect 10160 5607 10189 5747
rect 10235 5607 10248 5747
rect 10160 5556 10248 5607
rect 1604 5361 1692 5420
rect 1604 5221 1617 5361
rect 1663 5221 1692 5361
rect 1604 5176 1692 5221
rect 1892 5361 1980 5420
rect 1892 5221 1921 5361
rect 1967 5221 1980 5361
rect 1892 5176 1980 5221
rect 2072 5369 2160 5420
rect 2072 5229 2085 5369
rect 2131 5229 2160 5369
rect 2072 5176 2160 5229
rect 2260 5369 2348 5420
rect 2260 5229 2289 5369
rect 2335 5229 2348 5369
rect 2260 5176 2348 5229
rect 2744 5369 2832 5420
rect 2744 5229 2757 5369
rect 2803 5229 2832 5369
rect 2744 5176 2832 5229
rect 2932 5369 3020 5420
rect 2932 5229 2961 5369
rect 3007 5229 3020 5369
rect 2932 5176 3020 5229
rect 3416 5369 3504 5420
rect 3416 5229 3429 5369
rect 3475 5229 3504 5369
rect 3416 5176 3504 5229
rect 3604 5369 3692 5420
rect 3604 5229 3633 5369
rect 3679 5229 3692 5369
rect 3604 5176 3692 5229
rect 4088 5369 4176 5420
rect 4088 5229 4101 5369
rect 4147 5229 4176 5369
rect 4088 5176 4176 5229
rect 4276 5369 4364 5420
rect 4276 5229 4305 5369
rect 4351 5229 4364 5369
rect 4276 5176 4364 5229
rect 4760 5369 4848 5420
rect 4760 5229 4773 5369
rect 4819 5229 4848 5369
rect 4760 5176 4848 5229
rect 4948 5369 5036 5420
rect 4948 5229 4977 5369
rect 5023 5229 5036 5369
rect 4948 5176 5036 5229
rect 5656 5369 5744 5420
rect 5656 5229 5669 5369
rect 5715 5229 5744 5369
rect 5656 5176 5744 5229
rect 5844 5369 5932 5420
rect 5844 5229 5873 5369
rect 5919 5229 5932 5369
rect 5844 5176 5932 5229
rect 6084 5361 6172 5420
rect 6084 5221 6097 5361
rect 6143 5221 6172 5361
rect 6084 5176 6172 5221
rect 6372 5361 6460 5420
rect 6372 5221 6401 5361
rect 6447 5221 6460 5361
rect 6372 5176 6460 5221
rect 6888 5369 6976 5420
rect 6888 5229 6901 5369
rect 6947 5229 6976 5369
rect 6888 5176 6976 5229
rect 7076 5369 7164 5420
rect 7076 5229 7105 5369
rect 7151 5229 7164 5369
rect 7076 5176 7164 5229
rect 7560 5369 7648 5420
rect 7560 5229 7573 5369
rect 7619 5229 7648 5369
rect 7560 5176 7648 5229
rect 7748 5369 7836 5420
rect 7748 5229 7777 5369
rect 7823 5229 7836 5369
rect 7748 5176 7836 5229
rect 8232 5369 8320 5420
rect 8232 5229 8245 5369
rect 8291 5229 8320 5369
rect 8232 5176 8320 5229
rect 8420 5369 8508 5420
rect 8420 5229 8449 5369
rect 8495 5229 8508 5369
rect 8420 5176 8508 5229
rect 8660 5361 8748 5420
rect 8660 5221 8673 5361
rect 8719 5221 8748 5361
rect 8660 5176 8748 5221
rect 8948 5361 9036 5420
rect 8948 5221 8977 5361
rect 9023 5221 9036 5361
rect 8948 5176 9036 5221
rect 9240 5369 9328 5420
rect 9240 5229 9253 5369
rect 9299 5229 9328 5369
rect 9240 5176 9328 5229
rect 9428 5369 9516 5420
rect 9428 5229 9457 5369
rect 9503 5229 9516 5369
rect 9428 5176 9516 5229
rect 9972 5369 10060 5420
rect 9972 5229 9985 5369
rect 10031 5229 10060 5369
rect 9972 5176 10060 5229
rect 10160 5369 10248 5420
rect 10160 5229 10189 5369
rect 10235 5229 10248 5369
rect 10160 5176 10248 5229
rect 1848 4179 1936 4232
rect 1848 4039 1861 4179
rect 1907 4039 1936 4179
rect 1848 3988 1936 4039
rect 2036 4179 2124 4232
rect 2036 4039 2065 4179
rect 2111 4039 2124 4179
rect 2036 3988 2124 4039
rect 2520 4179 2608 4232
rect 2520 4039 2533 4179
rect 2579 4039 2608 4179
rect 2520 3988 2608 4039
rect 2708 4179 2796 4232
rect 2708 4039 2737 4179
rect 2783 4039 2796 4179
rect 2708 3988 2796 4039
rect 3192 4179 3280 4232
rect 3192 4039 3205 4179
rect 3251 4039 3280 4179
rect 3192 3988 3280 4039
rect 3380 4179 3468 4232
rect 3380 4039 3409 4179
rect 3455 4039 3468 4179
rect 3380 3988 3468 4039
rect 3864 4179 3952 4232
rect 3864 4039 3877 4179
rect 3923 4039 3952 4179
rect 3864 3988 3952 4039
rect 4052 4179 4140 4232
rect 4052 4039 4081 4179
rect 4127 4039 4140 4179
rect 4052 3988 4140 4039
rect 4536 4179 4624 4232
rect 4536 4039 4549 4179
rect 4595 4039 4624 4179
rect 4536 3988 4624 4039
rect 4724 4179 4812 4232
rect 4724 4039 4753 4179
rect 4799 4039 4812 4179
rect 4724 3988 4812 4039
rect 4964 4187 5052 4232
rect 4964 4047 4977 4187
rect 5023 4047 5052 4187
rect 4964 3988 5052 4047
rect 5252 4187 5340 4232
rect 5252 4047 5281 4187
rect 5327 4047 5340 4187
rect 5252 3988 5340 4047
rect 5656 4179 5744 4232
rect 5656 4039 5669 4179
rect 5715 4039 5744 4179
rect 5656 3988 5744 4039
rect 5844 4179 5932 4232
rect 5844 4039 5873 4179
rect 5919 4039 5932 4179
rect 5844 3988 5932 4039
rect 6328 4179 6416 4232
rect 6328 4039 6341 4179
rect 6387 4039 6416 4179
rect 6328 3988 6416 4039
rect 6516 4179 6604 4232
rect 6516 4039 6545 4179
rect 6591 4039 6604 4179
rect 6516 3988 6604 4039
rect 7000 4179 7088 4232
rect 7000 4039 7013 4179
rect 7059 4039 7088 4179
rect 7000 3988 7088 4039
rect 7188 4179 7276 4232
rect 7188 4039 7217 4179
rect 7263 4039 7276 4179
rect 7188 3988 7276 4039
rect 7672 4179 7760 4232
rect 7672 4039 7685 4179
rect 7731 4039 7760 4179
rect 7672 3988 7760 4039
rect 7860 4179 7948 4232
rect 7860 4039 7889 4179
rect 7935 4039 7948 4179
rect 7860 3988 7948 4039
rect 8344 4179 8432 4232
rect 8344 4039 8357 4179
rect 8403 4039 8432 4179
rect 8344 3988 8432 4039
rect 8532 4179 8620 4232
rect 8532 4039 8561 4179
rect 8607 4039 8620 4179
rect 8532 3988 8620 4039
rect 8772 4187 8860 4232
rect 8772 4047 8785 4187
rect 8831 4047 8860 4187
rect 8772 3988 8860 4047
rect 9060 4187 9148 4232
rect 9060 4047 9089 4187
rect 9135 4047 9148 4187
rect 9060 3988 9148 4047
rect 9912 4179 10000 4232
rect 9912 4039 9925 4179
rect 9971 4039 10000 4179
rect 9912 3988 10000 4039
rect 10100 4179 10188 4232
rect 10100 4039 10129 4179
rect 10175 4039 10188 4179
rect 10100 3988 10188 4039
rect 1908 3801 1996 3852
rect 1908 3661 1921 3801
rect 1967 3661 1996 3801
rect 1908 3608 1996 3661
rect 2096 3801 2184 3852
rect 2096 3661 2125 3801
rect 2171 3661 2184 3801
rect 2096 3608 2184 3661
rect 2520 3801 2608 3852
rect 2520 3661 2533 3801
rect 2579 3661 2608 3801
rect 2520 3608 2608 3661
rect 2708 3801 2796 3852
rect 2708 3661 2737 3801
rect 2783 3661 2796 3801
rect 2708 3608 2796 3661
rect 3192 3801 3280 3852
rect 3192 3661 3205 3801
rect 3251 3661 3280 3801
rect 3192 3608 3280 3661
rect 3380 3801 3468 3852
rect 3380 3661 3409 3801
rect 3455 3661 3468 3801
rect 3380 3608 3468 3661
rect 3864 3801 3952 3852
rect 3864 3661 3877 3801
rect 3923 3661 3952 3801
rect 3864 3608 3952 3661
rect 4052 3801 4140 3852
rect 4052 3661 4081 3801
rect 4127 3661 4140 3801
rect 4052 3608 4140 3661
rect 4536 3801 4624 3852
rect 4536 3661 4549 3801
rect 4595 3661 4624 3801
rect 4536 3608 4624 3661
rect 4724 3801 4812 3852
rect 4724 3661 4753 3801
rect 4799 3661 4812 3801
rect 4724 3608 4812 3661
rect 5656 3801 5744 3852
rect 5656 3661 5669 3801
rect 5715 3661 5744 3801
rect 5656 3608 5744 3661
rect 5844 3801 5932 3852
rect 5844 3661 5873 3801
rect 5919 3661 5932 3801
rect 5844 3608 5932 3661
rect 6084 3793 6172 3852
rect 6084 3653 6097 3793
rect 6143 3653 6172 3793
rect 6084 3608 6172 3653
rect 6372 3793 6460 3852
rect 6372 3653 6401 3793
rect 6447 3653 6460 3793
rect 6372 3608 6460 3653
rect 6552 3801 6640 3852
rect 6552 3661 6565 3801
rect 6611 3661 6640 3801
rect 6552 3608 6640 3661
rect 6740 3801 6828 3852
rect 6740 3661 6769 3801
rect 6815 3661 6828 3801
rect 6740 3608 6828 3661
rect 7224 3801 7312 3852
rect 7224 3661 7237 3801
rect 7283 3661 7312 3801
rect 7224 3608 7312 3661
rect 7412 3801 7500 3852
rect 7412 3661 7441 3801
rect 7487 3661 7500 3801
rect 7412 3608 7500 3661
rect 7956 3801 8044 3852
rect 7956 3661 7969 3801
rect 8015 3661 8044 3801
rect 7956 3608 8044 3661
rect 8144 3801 8232 3852
rect 8144 3661 8173 3801
rect 8219 3661 8232 3801
rect 8144 3608 8232 3661
rect 8568 3801 8656 3852
rect 8568 3661 8581 3801
rect 8627 3661 8656 3801
rect 8568 3608 8656 3661
rect 8756 3801 8844 3852
rect 8756 3661 8785 3801
rect 8831 3661 8844 3801
rect 8756 3608 8844 3661
rect 9444 3793 9532 3852
rect 9444 3653 9457 3793
rect 9503 3653 9532 3793
rect 9444 3608 9532 3653
rect 9732 3793 9820 3852
rect 9732 3653 9761 3793
rect 9807 3653 9820 3793
rect 9732 3608 9820 3653
rect 9912 3801 10000 3852
rect 9912 3661 9925 3801
rect 9971 3661 10000 3801
rect 9912 3608 10000 3661
rect 10100 3801 10188 3852
rect 10100 3661 10129 3801
rect 10175 3661 10188 3801
rect 10100 3608 10188 3661
<< mvndiffc >>
rect 1617 7986 1663 8032
rect 1921 7986 1967 8032
rect 2065 7986 2111 8032
rect 2289 7986 2335 8032
rect 2737 7986 2783 8032
rect 2961 7986 3007 8032
rect 3409 7986 3455 8032
rect 3633 7986 3679 8032
rect 4081 7986 4127 8032
rect 4305 7986 4351 8032
rect 4753 7986 4799 8032
rect 4977 7986 5023 8032
rect 5537 7986 5583 8032
rect 5841 7986 5887 8032
rect 5985 7986 6031 8032
rect 6289 7986 6335 8032
rect 6433 7986 6479 8032
rect 6737 7986 6783 8032
rect 6881 7986 6927 8032
rect 7185 7986 7231 8032
rect 7329 7986 7375 8032
rect 7633 7986 7679 8032
rect 7777 7986 7823 8032
rect 8081 7986 8127 8032
rect 8225 7986 8271 8032
rect 8529 7986 8575 8032
rect 8673 7986 8719 8032
rect 8977 7986 9023 8032
rect 9457 7986 9503 8032
rect 9761 7986 9807 8032
rect 9905 7986 9951 8032
rect 10209 7986 10255 8032
rect 1617 7648 1663 7694
rect 1921 7648 1967 7694
rect 2065 7648 2111 7694
rect 2289 7648 2335 7694
rect 2737 7648 2783 7694
rect 2961 7648 3007 7694
rect 3409 7648 3455 7694
rect 3633 7648 3679 7694
rect 4081 7648 4127 7694
rect 4305 7648 4351 7694
rect 4753 7648 4799 7694
rect 4977 7648 5023 7694
rect 5505 7648 5551 7694
rect 5729 7648 5775 7694
rect 6177 7648 6223 7694
rect 6401 7648 6447 7694
rect 6545 7648 6591 7694
rect 6849 7648 6895 7694
rect 6993 7648 7039 7694
rect 7297 7648 7343 7694
rect 7441 7648 7487 7694
rect 7745 7648 7791 7694
rect 7889 7648 7935 7694
rect 8193 7648 8239 7694
rect 8337 7648 8383 7694
rect 8641 7648 8687 7694
rect 8785 7648 8831 7694
rect 9089 7648 9135 7694
rect 9985 7648 10031 7694
rect 10209 7648 10255 7694
rect 1841 6418 1887 6464
rect 2065 6418 2111 6464
rect 2513 6418 2559 6464
rect 2737 6418 2783 6464
rect 3185 6418 3231 6464
rect 3409 6418 3455 6464
rect 3857 6418 3903 6464
rect 4081 6418 4127 6464
rect 4529 6418 4575 6464
rect 4753 6418 4799 6464
rect 5649 6418 5695 6464
rect 5873 6418 5919 6464
rect 6321 6418 6367 6464
rect 6545 6418 6591 6464
rect 6993 6418 7039 6464
rect 7217 6418 7263 6464
rect 7441 6418 7487 6464
rect 7745 6418 7791 6464
rect 7889 6418 7935 6464
rect 8193 6418 8239 6464
rect 8337 6418 8383 6464
rect 8561 6418 8607 6464
rect 9009 6378 9055 6424
rect 9233 6378 9279 6424
rect 9493 6378 9539 6424
rect 9717 6395 9763 6441
rect 10125 6353 10171 6399
rect 1729 6080 1775 6126
rect 1953 6080 1999 6126
rect 2401 6080 2447 6126
rect 2625 6080 2671 6126
rect 3073 6080 3119 6126
rect 3297 6080 3343 6126
rect 3745 6080 3791 6126
rect 3969 6080 4015 6126
rect 4417 6080 4463 6126
rect 4641 6080 4687 6126
rect 5089 6080 5135 6126
rect 5313 6080 5359 6126
rect 5761 6080 5807 6126
rect 5985 6080 6031 6126
rect 6433 6080 6479 6126
rect 6657 6080 6703 6126
rect 6881 6080 6927 6126
rect 7185 6080 7231 6126
rect 7665 6080 7711 6126
rect 7889 6080 7935 6126
rect 8337 6080 8383 6126
rect 8561 6080 8607 6126
rect 8785 6080 8831 6126
rect 9089 6080 9135 6126
rect 9985 6080 10031 6126
rect 10209 6080 10255 6126
rect 1617 4850 1663 4896
rect 1921 4850 1967 4896
rect 2065 4850 2111 4896
rect 2289 4850 2335 4896
rect 2737 4850 2783 4896
rect 2961 4850 3007 4896
rect 3409 4850 3455 4896
rect 3633 4850 3679 4896
rect 4081 4850 4127 4896
rect 4305 4850 4351 4896
rect 4753 4850 4799 4896
rect 4977 4850 5023 4896
rect 5649 4850 5695 4896
rect 5873 4850 5919 4896
rect 6097 4850 6143 4896
rect 6401 4850 6447 4896
rect 6881 4850 6927 4896
rect 7105 4850 7151 4896
rect 7553 4850 7599 4896
rect 7777 4850 7823 4896
rect 8225 4850 8271 4896
rect 8449 4850 8495 4896
rect 8673 4850 8719 4896
rect 8977 4850 9023 4896
rect 9233 4850 9279 4896
rect 9457 4850 9503 4896
rect 9985 4850 10031 4896
rect 10209 4850 10255 4896
rect 1841 4512 1887 4558
rect 2065 4512 2111 4558
rect 2513 4512 2559 4558
rect 2737 4512 2783 4558
rect 3185 4512 3231 4558
rect 3409 4512 3455 4558
rect 3857 4512 3903 4558
rect 4081 4512 4127 4558
rect 4529 4512 4575 4558
rect 4753 4512 4799 4558
rect 4977 4512 5023 4558
rect 5281 4512 5327 4558
rect 5649 4512 5695 4558
rect 5873 4512 5919 4558
rect 6321 4512 6367 4558
rect 6545 4512 6591 4558
rect 6993 4512 7039 4558
rect 7217 4512 7263 4558
rect 7665 4512 7711 4558
rect 7889 4512 7935 4558
rect 8337 4512 8383 4558
rect 8561 4512 8607 4558
rect 8785 4512 8831 4558
rect 9089 4512 9135 4558
rect 9905 4512 9951 4558
rect 10129 4512 10175 4558
rect 1921 3282 1967 3328
rect 2145 3282 2191 3328
rect 2513 3282 2559 3328
rect 2737 3282 2783 3328
rect 3185 3282 3231 3328
rect 3409 3282 3455 3328
rect 3857 3282 3903 3328
rect 4081 3282 4127 3328
rect 4529 3282 4575 3328
rect 4753 3282 4799 3328
rect 5649 3282 5695 3328
rect 5873 3282 5919 3328
rect 6097 3282 6143 3328
rect 6401 3282 6447 3328
rect 6545 3282 6591 3328
rect 6769 3282 6815 3328
rect 7217 3282 7263 3328
rect 7441 3282 7487 3328
rect 7969 3282 8015 3328
rect 8193 3282 8239 3328
rect 8561 3282 8607 3328
rect 8785 3282 8831 3328
rect 9457 3282 9503 3328
rect 9761 3282 9807 3328
rect 9905 3282 9951 3328
rect 10129 3282 10175 3328
<< mvpdiffc >>
rect 1617 8357 1663 8497
rect 1921 8357 1967 8497
rect 2085 8365 2131 8505
rect 2289 8365 2335 8505
rect 2757 8365 2803 8505
rect 2961 8365 3007 8505
rect 3429 8365 3475 8505
rect 3633 8365 3679 8505
rect 4101 8365 4147 8505
rect 4305 8365 4351 8505
rect 4773 8365 4819 8505
rect 4977 8365 5023 8505
rect 5537 8357 5583 8497
rect 5841 8357 5887 8497
rect 5985 8357 6031 8497
rect 6289 8357 6335 8497
rect 6433 8357 6479 8497
rect 6737 8357 6783 8497
rect 6881 8357 6927 8497
rect 7185 8357 7231 8497
rect 7329 8357 7375 8497
rect 7633 8357 7679 8497
rect 7777 8357 7823 8497
rect 8081 8357 8127 8497
rect 8225 8357 8271 8497
rect 8529 8357 8575 8497
rect 8673 8357 8719 8497
rect 8977 8357 9023 8497
rect 9457 8357 9503 8497
rect 9761 8357 9807 8497
rect 9905 8357 9951 8497
rect 10209 8357 10255 8497
rect 1617 7183 1663 7323
rect 1921 7183 1967 7323
rect 2085 7175 2131 7315
rect 2289 7175 2335 7315
rect 2757 7175 2803 7315
rect 2961 7175 3007 7315
rect 3429 7175 3475 7315
rect 3633 7175 3679 7315
rect 4101 7175 4147 7315
rect 4305 7175 4351 7315
rect 4773 7175 4819 7315
rect 4977 7175 5023 7315
rect 5505 7175 5551 7315
rect 5709 7175 5755 7315
rect 6177 7175 6223 7315
rect 6381 7175 6427 7315
rect 6545 7183 6591 7323
rect 6849 7183 6895 7323
rect 6993 7183 7039 7323
rect 7297 7183 7343 7323
rect 7441 7183 7487 7323
rect 7745 7183 7791 7323
rect 7889 7183 7935 7323
rect 8193 7183 8239 7323
rect 8337 7183 8383 7323
rect 8641 7183 8687 7323
rect 8785 7183 8831 7323
rect 9089 7183 9135 7323
rect 9985 7175 10031 7315
rect 10189 7175 10235 7315
rect 1861 6797 1907 6937
rect 2065 6797 2111 6937
rect 2533 6797 2579 6937
rect 2737 6797 2783 6937
rect 3205 6797 3251 6937
rect 3409 6797 3455 6937
rect 3877 6797 3923 6937
rect 4081 6797 4127 6937
rect 4549 6797 4595 6937
rect 4753 6797 4799 6937
rect 5669 6797 5715 6937
rect 5873 6797 5919 6937
rect 6341 6797 6387 6937
rect 6545 6797 6591 6937
rect 7013 6797 7059 6937
rect 7217 6797 7263 6937
rect 7441 6789 7487 6929
rect 7745 6789 7791 6929
rect 7889 6789 7935 6929
rect 8193 6789 8239 6929
rect 8357 6797 8403 6937
rect 8561 6797 8607 6937
rect 9029 6895 9075 6941
rect 9513 6835 9559 6975
rect 9717 6904 9763 6950
rect 9921 6811 9967 6857
rect 10125 6904 10171 6950
rect 1749 5607 1795 5747
rect 1953 5607 1999 5747
rect 2421 5607 2467 5747
rect 2625 5607 2671 5747
rect 3093 5607 3139 5747
rect 3297 5607 3343 5747
rect 3765 5607 3811 5747
rect 3969 5607 4015 5747
rect 4437 5607 4483 5747
rect 4641 5607 4687 5747
rect 5109 5607 5155 5747
rect 5313 5607 5359 5747
rect 5781 5607 5827 5747
rect 5985 5607 6031 5747
rect 6453 5607 6499 5747
rect 6657 5607 6703 5747
rect 6881 5615 6927 5755
rect 7185 5615 7231 5755
rect 7685 5607 7731 5747
rect 7889 5607 7935 5747
rect 8357 5607 8403 5747
rect 8561 5607 8607 5747
rect 8785 5615 8831 5755
rect 9089 5615 9135 5755
rect 9985 5607 10031 5747
rect 10189 5607 10235 5747
rect 1617 5221 1663 5361
rect 1921 5221 1967 5361
rect 2085 5229 2131 5369
rect 2289 5229 2335 5369
rect 2757 5229 2803 5369
rect 2961 5229 3007 5369
rect 3429 5229 3475 5369
rect 3633 5229 3679 5369
rect 4101 5229 4147 5369
rect 4305 5229 4351 5369
rect 4773 5229 4819 5369
rect 4977 5229 5023 5369
rect 5669 5229 5715 5369
rect 5873 5229 5919 5369
rect 6097 5221 6143 5361
rect 6401 5221 6447 5361
rect 6901 5229 6947 5369
rect 7105 5229 7151 5369
rect 7573 5229 7619 5369
rect 7777 5229 7823 5369
rect 8245 5229 8291 5369
rect 8449 5229 8495 5369
rect 8673 5221 8719 5361
rect 8977 5221 9023 5361
rect 9253 5229 9299 5369
rect 9457 5229 9503 5369
rect 9985 5229 10031 5369
rect 10189 5229 10235 5369
rect 1861 4039 1907 4179
rect 2065 4039 2111 4179
rect 2533 4039 2579 4179
rect 2737 4039 2783 4179
rect 3205 4039 3251 4179
rect 3409 4039 3455 4179
rect 3877 4039 3923 4179
rect 4081 4039 4127 4179
rect 4549 4039 4595 4179
rect 4753 4039 4799 4179
rect 4977 4047 5023 4187
rect 5281 4047 5327 4187
rect 5669 4039 5715 4179
rect 5873 4039 5919 4179
rect 6341 4039 6387 4179
rect 6545 4039 6591 4179
rect 7013 4039 7059 4179
rect 7217 4039 7263 4179
rect 7685 4039 7731 4179
rect 7889 4039 7935 4179
rect 8357 4039 8403 4179
rect 8561 4039 8607 4179
rect 8785 4047 8831 4187
rect 9089 4047 9135 4187
rect 9925 4039 9971 4179
rect 10129 4039 10175 4179
rect 1921 3661 1967 3801
rect 2125 3661 2171 3801
rect 2533 3661 2579 3801
rect 2737 3661 2783 3801
rect 3205 3661 3251 3801
rect 3409 3661 3455 3801
rect 3877 3661 3923 3801
rect 4081 3661 4127 3801
rect 4549 3661 4595 3801
rect 4753 3661 4799 3801
rect 5669 3661 5715 3801
rect 5873 3661 5919 3801
rect 6097 3653 6143 3793
rect 6401 3653 6447 3793
rect 6565 3661 6611 3801
rect 6769 3661 6815 3801
rect 7237 3661 7283 3801
rect 7441 3661 7487 3801
rect 7969 3661 8015 3801
rect 8173 3661 8219 3801
rect 8581 3661 8627 3801
rect 8785 3661 8831 3801
rect 9457 3653 9503 3793
rect 9761 3653 9807 3793
rect 9925 3661 9971 3801
rect 10129 3661 10175 3801
<< mvpsubdiff >>
rect 1400 8066 1504 8096
rect 1400 7919 1429 8066
rect 1475 7919 1504 8066
rect 1400 7896 1504 7919
rect 5320 8066 5432 8096
rect 5320 7919 5353 8066
rect 5399 7919 5432 8066
rect 5320 7896 5432 7919
rect 9240 8066 9352 8096
rect 9240 7919 9273 8066
rect 9319 7919 9352 8066
rect 9240 7896 9352 7919
rect 10480 8066 10584 8096
rect 10480 7919 10509 8066
rect 10555 7919 10584 8066
rect 10480 7896 10584 7919
rect 1400 7761 1504 7784
rect 1400 7614 1429 7761
rect 1475 7614 1504 7761
rect 1400 7584 1504 7614
rect 9352 7761 9464 7784
rect 9352 7614 9385 7761
rect 9431 7614 9464 7761
rect 9352 7584 9464 7614
rect 10480 7761 10584 7784
rect 10480 7614 10509 7761
rect 10555 7614 10584 7761
rect 10480 7584 10584 7614
rect 1400 6498 1504 6528
rect 1400 6351 1429 6498
rect 1475 6351 1504 6498
rect 1400 6328 1504 6351
rect 5320 6498 5432 6528
rect 5320 6351 5353 6498
rect 5399 6351 5432 6498
rect 5320 6328 5432 6351
rect 10480 6498 10584 6528
rect 10480 6351 10509 6498
rect 10555 6351 10584 6498
rect 10480 6328 10584 6351
rect 1400 6193 1504 6216
rect 1400 6046 1429 6193
rect 1475 6046 1504 6193
rect 1400 6016 1504 6046
rect 9352 6193 9464 6216
rect 9352 6046 9385 6193
rect 9431 6046 9464 6193
rect 9352 6016 9464 6046
rect 10480 6193 10584 6216
rect 10480 6046 10509 6193
rect 10555 6046 10584 6193
rect 10480 6016 10584 6046
rect 1400 4930 1504 4960
rect 1400 4783 1429 4930
rect 1475 4783 1504 4930
rect 1400 4760 1504 4783
rect 5320 4930 5432 4960
rect 5320 4783 5353 4930
rect 5399 4783 5432 4930
rect 5320 4760 5432 4783
rect 10480 4930 10584 4960
rect 10480 4783 10509 4930
rect 10555 4783 10584 4930
rect 10480 4760 10584 4783
rect 1400 4625 1504 4648
rect 1400 4478 1429 4625
rect 1475 4478 1504 4625
rect 1400 4448 1504 4478
rect 9352 4625 9464 4648
rect 9352 4478 9385 4625
rect 9431 4478 9464 4625
rect 9352 4448 9464 4478
rect 10480 4625 10584 4648
rect 10480 4478 10509 4625
rect 10555 4478 10584 4625
rect 10480 4448 10584 4478
rect 1400 3362 1504 3392
rect 1400 3215 1429 3362
rect 1475 3215 1504 3362
rect 1400 3192 1504 3215
rect 5320 3362 5432 3392
rect 5320 3215 5353 3362
rect 5399 3215 5432 3362
rect 5320 3192 5432 3215
rect 9240 3362 9352 3392
rect 9240 3215 9273 3362
rect 9319 3215 9352 3362
rect 9240 3192 9352 3215
rect 10480 3362 10584 3392
rect 10480 3215 10509 3362
rect 10555 3215 10584 3362
rect 10480 3192 10584 3215
<< mvnsubdiff >>
rect 1416 8539 1488 8552
rect 1416 8493 1429 8539
rect 1475 8493 1488 8539
rect 1416 8411 1488 8493
rect 1416 8365 1429 8411
rect 1475 8365 1488 8411
rect 1416 8283 1488 8365
rect 5336 8539 5416 8552
rect 5336 8493 5353 8539
rect 5399 8493 5416 8539
rect 5336 8411 5416 8493
rect 5336 8365 5353 8411
rect 5399 8365 5416 8411
rect 1416 8237 1429 8283
rect 1475 8237 1488 8283
rect 1416 8224 1488 8237
rect 5336 8283 5416 8365
rect 9256 8539 9336 8552
rect 9256 8493 9273 8539
rect 9319 8493 9336 8539
rect 9256 8411 9336 8493
rect 9256 8365 9273 8411
rect 9319 8365 9336 8411
rect 5336 8237 5353 8283
rect 5399 8237 5416 8283
rect 5336 8224 5416 8237
rect 9256 8283 9336 8365
rect 10496 8539 10568 8552
rect 10496 8493 10509 8539
rect 10555 8493 10568 8539
rect 10496 8411 10568 8493
rect 10496 8365 10509 8411
rect 10555 8365 10568 8411
rect 9256 8237 9273 8283
rect 9319 8237 9336 8283
rect 9256 8224 9336 8237
rect 10496 8283 10568 8365
rect 10496 8237 10509 8283
rect 10555 8237 10568 8283
rect 10496 8224 10568 8237
rect 1416 7443 1488 7456
rect 1416 7397 1429 7443
rect 1475 7397 1488 7443
rect 1416 7315 1488 7397
rect 9368 7443 9448 7456
rect 9368 7397 9385 7443
rect 9431 7397 9448 7443
rect 1416 7269 1429 7315
rect 1475 7269 1488 7315
rect 1416 7187 1488 7269
rect 1416 7141 1429 7187
rect 1475 7141 1488 7187
rect 1416 7128 1488 7141
rect 9368 7315 9448 7397
rect 10496 7443 10568 7456
rect 10496 7397 10509 7443
rect 10555 7397 10568 7443
rect 9368 7269 9385 7315
rect 9431 7269 9448 7315
rect 9368 7187 9448 7269
rect 9368 7141 9385 7187
rect 9431 7141 9448 7187
rect 9368 7128 9448 7141
rect 10496 7315 10568 7397
rect 10496 7269 10509 7315
rect 10555 7269 10568 7315
rect 10496 7187 10568 7269
rect 10496 7141 10509 7187
rect 10555 7141 10568 7187
rect 10496 7128 10568 7141
rect 1416 6971 1488 6984
rect 1416 6925 1429 6971
rect 1475 6925 1488 6971
rect 1416 6843 1488 6925
rect 1416 6797 1429 6843
rect 1475 6797 1488 6843
rect 1416 6715 1488 6797
rect 5336 6971 5416 6984
rect 5336 6925 5353 6971
rect 5399 6925 5416 6971
rect 5336 6843 5416 6925
rect 5336 6797 5353 6843
rect 5399 6797 5416 6843
rect 1416 6669 1429 6715
rect 1475 6669 1488 6715
rect 1416 6656 1488 6669
rect 5336 6715 5416 6797
rect 5336 6669 5353 6715
rect 5399 6669 5416 6715
rect 5336 6656 5416 6669
rect 10496 6971 10568 6984
rect 10496 6925 10509 6971
rect 10555 6925 10568 6971
rect 10496 6843 10568 6925
rect 10496 6797 10509 6843
rect 10555 6797 10568 6843
rect 10496 6715 10568 6797
rect 10496 6669 10509 6715
rect 10555 6669 10568 6715
rect 10496 6656 10568 6669
rect 1416 5875 1488 5888
rect 1416 5829 1429 5875
rect 1475 5829 1488 5875
rect 1416 5747 1488 5829
rect 9368 5875 9448 5888
rect 9368 5829 9385 5875
rect 9431 5829 9448 5875
rect 1416 5701 1429 5747
rect 1475 5701 1488 5747
rect 1416 5619 1488 5701
rect 1416 5573 1429 5619
rect 1475 5573 1488 5619
rect 1416 5560 1488 5573
rect 9368 5747 9448 5829
rect 10496 5875 10568 5888
rect 10496 5829 10509 5875
rect 10555 5829 10568 5875
rect 9368 5701 9385 5747
rect 9431 5701 9448 5747
rect 9368 5619 9448 5701
rect 9368 5573 9385 5619
rect 9431 5573 9448 5619
rect 9368 5560 9448 5573
rect 10496 5747 10568 5829
rect 10496 5701 10509 5747
rect 10555 5701 10568 5747
rect 10496 5619 10568 5701
rect 10496 5573 10509 5619
rect 10555 5573 10568 5619
rect 10496 5560 10568 5573
rect 1416 5403 1488 5416
rect 1416 5357 1429 5403
rect 1475 5357 1488 5403
rect 1416 5275 1488 5357
rect 1416 5229 1429 5275
rect 1475 5229 1488 5275
rect 1416 5147 1488 5229
rect 5336 5403 5416 5416
rect 5336 5357 5353 5403
rect 5399 5357 5416 5403
rect 5336 5275 5416 5357
rect 5336 5229 5353 5275
rect 5399 5229 5416 5275
rect 1416 5101 1429 5147
rect 1475 5101 1488 5147
rect 1416 5088 1488 5101
rect 5336 5147 5416 5229
rect 10496 5403 10568 5416
rect 10496 5357 10509 5403
rect 10555 5357 10568 5403
rect 10496 5275 10568 5357
rect 10496 5229 10509 5275
rect 10555 5229 10568 5275
rect 5336 5101 5353 5147
rect 5399 5101 5416 5147
rect 5336 5088 5416 5101
rect 10496 5147 10568 5229
rect 10496 5101 10509 5147
rect 10555 5101 10568 5147
rect 10496 5088 10568 5101
rect 1416 4307 1488 4320
rect 1416 4261 1429 4307
rect 1475 4261 1488 4307
rect 1416 4179 1488 4261
rect 9368 4307 9448 4320
rect 9368 4261 9385 4307
rect 9431 4261 9448 4307
rect 1416 4133 1429 4179
rect 1475 4133 1488 4179
rect 1416 4051 1488 4133
rect 1416 4005 1429 4051
rect 1475 4005 1488 4051
rect 1416 3992 1488 4005
rect 9368 4179 9448 4261
rect 10496 4307 10568 4320
rect 10496 4261 10509 4307
rect 10555 4261 10568 4307
rect 9368 4133 9385 4179
rect 9431 4133 9448 4179
rect 9368 4051 9448 4133
rect 9368 4005 9385 4051
rect 9431 4005 9448 4051
rect 9368 3992 9448 4005
rect 10496 4179 10568 4261
rect 10496 4133 10509 4179
rect 10555 4133 10568 4179
rect 10496 4051 10568 4133
rect 10496 4005 10509 4051
rect 10555 4005 10568 4051
rect 10496 3992 10568 4005
rect 1416 3835 1488 3848
rect 1416 3789 1429 3835
rect 1475 3789 1488 3835
rect 1416 3707 1488 3789
rect 1416 3661 1429 3707
rect 1475 3661 1488 3707
rect 1416 3579 1488 3661
rect 5336 3835 5416 3848
rect 5336 3789 5353 3835
rect 5399 3789 5416 3835
rect 5336 3707 5416 3789
rect 5336 3661 5353 3707
rect 5399 3661 5416 3707
rect 1416 3533 1429 3579
rect 1475 3533 1488 3579
rect 1416 3520 1488 3533
rect 5336 3579 5416 3661
rect 9256 3835 9336 3848
rect 9256 3789 9273 3835
rect 9319 3789 9336 3835
rect 9256 3707 9336 3789
rect 9256 3661 9273 3707
rect 9319 3661 9336 3707
rect 5336 3533 5353 3579
rect 5399 3533 5416 3579
rect 5336 3520 5416 3533
rect 9256 3579 9336 3661
rect 10496 3835 10568 3848
rect 10496 3789 10509 3835
rect 10555 3789 10568 3835
rect 10496 3707 10568 3789
rect 10496 3661 10509 3707
rect 10555 3661 10568 3707
rect 9256 3533 9273 3579
rect 9319 3533 9336 3579
rect 9256 3520 9336 3533
rect 10496 3579 10568 3661
rect 10496 3533 10509 3579
rect 10555 3533 10568 3579
rect 10496 3520 10568 3533
<< mvpsubdiffcont >>
rect 1429 7919 1475 8066
rect 5353 7919 5399 8066
rect 9273 7919 9319 8066
rect 10509 7919 10555 8066
rect 1429 7614 1475 7761
rect 9385 7614 9431 7761
rect 10509 7614 10555 7761
rect 1429 6351 1475 6498
rect 5353 6351 5399 6498
rect 10509 6351 10555 6498
rect 1429 6046 1475 6193
rect 9385 6046 9431 6193
rect 10509 6046 10555 6193
rect 1429 4783 1475 4930
rect 5353 4783 5399 4930
rect 10509 4783 10555 4930
rect 1429 4478 1475 4625
rect 9385 4478 9431 4625
rect 10509 4478 10555 4625
rect 1429 3215 1475 3362
rect 5353 3215 5399 3362
rect 9273 3215 9319 3362
rect 10509 3215 10555 3362
<< mvnsubdiffcont >>
rect 1429 8493 1475 8539
rect 1429 8365 1475 8411
rect 5353 8493 5399 8539
rect 5353 8365 5399 8411
rect 1429 8237 1475 8283
rect 9273 8493 9319 8539
rect 9273 8365 9319 8411
rect 5353 8237 5399 8283
rect 10509 8493 10555 8539
rect 10509 8365 10555 8411
rect 9273 8237 9319 8283
rect 10509 8237 10555 8283
rect 1429 7397 1475 7443
rect 9385 7397 9431 7443
rect 1429 7269 1475 7315
rect 1429 7141 1475 7187
rect 10509 7397 10555 7443
rect 9385 7269 9431 7315
rect 9385 7141 9431 7187
rect 10509 7269 10555 7315
rect 10509 7141 10555 7187
rect 1429 6925 1475 6971
rect 1429 6797 1475 6843
rect 5353 6925 5399 6971
rect 5353 6797 5399 6843
rect 1429 6669 1475 6715
rect 5353 6669 5399 6715
rect 10509 6925 10555 6971
rect 10509 6797 10555 6843
rect 10509 6669 10555 6715
rect 1429 5829 1475 5875
rect 9385 5829 9431 5875
rect 1429 5701 1475 5747
rect 1429 5573 1475 5619
rect 10509 5829 10555 5875
rect 9385 5701 9431 5747
rect 9385 5573 9431 5619
rect 10509 5701 10555 5747
rect 10509 5573 10555 5619
rect 1429 5357 1475 5403
rect 1429 5229 1475 5275
rect 5353 5357 5399 5403
rect 5353 5229 5399 5275
rect 1429 5101 1475 5147
rect 10509 5357 10555 5403
rect 10509 5229 10555 5275
rect 5353 5101 5399 5147
rect 10509 5101 10555 5147
rect 1429 4261 1475 4307
rect 9385 4261 9431 4307
rect 1429 4133 1475 4179
rect 1429 4005 1475 4051
rect 10509 4261 10555 4307
rect 9385 4133 9431 4179
rect 9385 4005 9431 4051
rect 10509 4133 10555 4179
rect 10509 4005 10555 4051
rect 1429 3789 1475 3835
rect 1429 3661 1475 3707
rect 5353 3789 5399 3835
rect 5353 3661 5399 3707
rect 1429 3533 1475 3579
rect 9273 3789 9319 3835
rect 9273 3661 9319 3707
rect 5353 3533 5399 3579
rect 10509 3789 10555 3835
rect 10509 3661 10555 3707
rect 9273 3533 9319 3579
rect 10509 3533 10555 3579
<< polysilicon >>
rect 1692 8556 1892 8600
rect 2160 8556 2260 8600
rect 2832 8556 2932 8600
rect 3504 8556 3604 8600
rect 4176 8556 4276 8600
rect 4848 8556 4948 8600
rect 5612 8556 5812 8600
rect 6060 8556 6260 8600
rect 6508 8556 6708 8600
rect 6956 8556 7156 8600
rect 7404 8556 7604 8600
rect 7852 8556 8052 8600
rect 8300 8556 8500 8600
rect 8748 8556 8948 8600
rect 9532 8556 9732 8600
rect 9980 8556 10180 8600
rect 1692 8278 1892 8312
rect 1692 8232 1728 8278
rect 1868 8232 1892 8278
rect 1692 8215 1892 8232
rect 2160 8263 2260 8312
rect 2160 8226 2173 8263
rect 1692 8151 1892 8164
rect 1692 8105 1720 8151
rect 1860 8105 1892 8151
rect 1692 8072 1892 8105
rect 2140 8123 2173 8226
rect 2219 8123 2260 8263
rect 2832 8263 2932 8312
rect 2832 8226 2845 8263
rect 2140 8072 2260 8123
rect 2812 8123 2845 8226
rect 2891 8123 2932 8263
rect 3504 8263 3604 8312
rect 3504 8226 3517 8263
rect 2812 8072 2932 8123
rect 3484 8123 3517 8226
rect 3563 8123 3604 8263
rect 4176 8263 4276 8312
rect 4176 8226 4189 8263
rect 3484 8072 3604 8123
rect 4156 8123 4189 8226
rect 4235 8123 4276 8263
rect 4848 8263 4948 8312
rect 4848 8226 4861 8263
rect 4156 8072 4276 8123
rect 4828 8123 4861 8226
rect 4907 8123 4948 8263
rect 5612 8278 5812 8312
rect 5612 8232 5648 8278
rect 5788 8232 5812 8278
rect 5612 8215 5812 8232
rect 6060 8278 6260 8312
rect 6060 8232 6096 8278
rect 6236 8232 6260 8278
rect 6060 8215 6260 8232
rect 6508 8278 6708 8312
rect 6508 8232 6544 8278
rect 6684 8232 6708 8278
rect 6508 8215 6708 8232
rect 6956 8278 7156 8312
rect 6956 8232 6992 8278
rect 7132 8232 7156 8278
rect 6956 8215 7156 8232
rect 7404 8278 7604 8312
rect 7404 8232 7440 8278
rect 7580 8232 7604 8278
rect 7404 8215 7604 8232
rect 7852 8278 8052 8312
rect 7852 8232 7888 8278
rect 8028 8232 8052 8278
rect 7852 8215 8052 8232
rect 8300 8278 8500 8312
rect 8300 8232 8336 8278
rect 8476 8232 8500 8278
rect 8300 8215 8500 8232
rect 8748 8278 8948 8312
rect 8748 8232 8784 8278
rect 8924 8232 8948 8278
rect 8748 8215 8948 8232
rect 9532 8278 9732 8312
rect 9532 8232 9568 8278
rect 9708 8232 9732 8278
rect 9532 8215 9732 8232
rect 9980 8278 10180 8312
rect 9980 8232 10016 8278
rect 10156 8232 10180 8278
rect 9980 8215 10180 8232
rect 4828 8072 4948 8123
rect 5612 8151 5812 8164
rect 5612 8105 5640 8151
rect 5780 8105 5812 8151
rect 5612 8072 5812 8105
rect 6060 8151 6260 8164
rect 6060 8105 6088 8151
rect 6228 8105 6260 8151
rect 6060 8072 6260 8105
rect 6508 8151 6708 8164
rect 6508 8105 6536 8151
rect 6676 8105 6708 8151
rect 6508 8072 6708 8105
rect 6956 8151 7156 8164
rect 6956 8105 6984 8151
rect 7124 8105 7156 8151
rect 6956 8072 7156 8105
rect 7404 8151 7604 8164
rect 7404 8105 7432 8151
rect 7572 8105 7604 8151
rect 7404 8072 7604 8105
rect 7852 8151 8052 8164
rect 7852 8105 7880 8151
rect 8020 8105 8052 8151
rect 7852 8072 8052 8105
rect 8300 8151 8500 8164
rect 8300 8105 8328 8151
rect 8468 8105 8500 8151
rect 8300 8072 8500 8105
rect 8748 8151 8948 8164
rect 8748 8105 8776 8151
rect 8916 8105 8948 8151
rect 8748 8072 8948 8105
rect 9532 8151 9732 8164
rect 9532 8105 9560 8151
rect 9700 8105 9732 8151
rect 1692 7864 1892 7908
rect 2140 7864 2260 7908
rect 2812 7864 2932 7908
rect 3484 7864 3604 7908
rect 4156 7864 4276 7908
rect 4828 7864 4948 7908
rect 9532 8072 9732 8105
rect 9980 8151 10180 8164
rect 9980 8105 10008 8151
rect 10148 8105 10180 8151
rect 9980 8072 10180 8105
rect 5612 7864 5812 7908
rect 6060 7864 6260 7908
rect 6508 7864 6708 7908
rect 6956 7864 7156 7908
rect 7404 7864 7604 7908
rect 7852 7864 8052 7908
rect 8300 7864 8500 7908
rect 8748 7864 8948 7908
rect 9532 7864 9732 7908
rect 9980 7864 10180 7908
rect 1692 7772 1892 7816
rect 2140 7772 2260 7816
rect 2812 7772 2932 7816
rect 3484 7772 3604 7816
rect 4156 7772 4276 7816
rect 4828 7772 4948 7816
rect 5580 7772 5700 7816
rect 6252 7772 6372 7816
rect 6620 7772 6820 7816
rect 7068 7772 7268 7816
rect 7516 7772 7716 7816
rect 7964 7772 8164 7816
rect 8412 7772 8612 7816
rect 8860 7772 9060 7816
rect 10060 7772 10180 7816
rect 1692 7575 1892 7608
rect 1692 7529 1720 7575
rect 1860 7529 1892 7575
rect 1692 7516 1892 7529
rect 2140 7557 2260 7608
rect 1692 7448 1892 7465
rect 2140 7454 2173 7557
rect 1692 7402 1728 7448
rect 1868 7402 1892 7448
rect 1692 7368 1892 7402
rect 2160 7417 2173 7454
rect 2219 7417 2260 7557
rect 2812 7557 2932 7608
rect 2812 7454 2845 7557
rect 2160 7368 2260 7417
rect 2832 7417 2845 7454
rect 2891 7417 2932 7557
rect 3484 7557 3604 7608
rect 3484 7454 3517 7557
rect 2832 7368 2932 7417
rect 3504 7417 3517 7454
rect 3563 7417 3604 7557
rect 4156 7557 4276 7608
rect 4156 7454 4189 7557
rect 3504 7368 3604 7417
rect 4176 7417 4189 7454
rect 4235 7417 4276 7557
rect 4828 7557 4948 7608
rect 4828 7454 4861 7557
rect 4176 7368 4276 7417
rect 4848 7417 4861 7454
rect 4907 7417 4948 7557
rect 4848 7368 4948 7417
rect 5580 7557 5700 7608
rect 5580 7417 5621 7557
rect 5667 7454 5700 7557
rect 6252 7557 6372 7608
rect 5667 7417 5680 7454
rect 5580 7368 5680 7417
rect 6252 7417 6293 7557
rect 6339 7454 6372 7557
rect 6620 7575 6820 7608
rect 6620 7529 6648 7575
rect 6788 7529 6820 7575
rect 6620 7516 6820 7529
rect 7068 7575 7268 7608
rect 7068 7529 7096 7575
rect 7236 7529 7268 7575
rect 7068 7516 7268 7529
rect 7516 7575 7716 7608
rect 7516 7529 7544 7575
rect 7684 7529 7716 7575
rect 7516 7516 7716 7529
rect 7964 7575 8164 7608
rect 7964 7529 7992 7575
rect 8132 7529 8164 7575
rect 7964 7516 8164 7529
rect 8412 7575 8612 7608
rect 8412 7529 8440 7575
rect 8580 7529 8612 7575
rect 8412 7516 8612 7529
rect 8860 7575 9060 7608
rect 8860 7529 8888 7575
rect 9028 7529 9060 7575
rect 8860 7516 9060 7529
rect 10060 7557 10180 7608
rect 6339 7417 6352 7454
rect 6252 7368 6352 7417
rect 6620 7448 6820 7465
rect 6620 7402 6656 7448
rect 6796 7402 6820 7448
rect 6620 7368 6820 7402
rect 7068 7448 7268 7465
rect 7068 7402 7104 7448
rect 7244 7402 7268 7448
rect 7068 7368 7268 7402
rect 7516 7448 7716 7465
rect 7516 7402 7552 7448
rect 7692 7402 7716 7448
rect 7516 7368 7716 7402
rect 7964 7448 8164 7465
rect 7964 7402 8000 7448
rect 8140 7402 8164 7448
rect 7964 7368 8164 7402
rect 8412 7448 8612 7465
rect 8412 7402 8448 7448
rect 8588 7402 8612 7448
rect 8412 7368 8612 7402
rect 8860 7448 9060 7465
rect 8860 7402 8896 7448
rect 9036 7402 9060 7448
rect 8860 7368 9060 7402
rect 10060 7417 10101 7557
rect 10147 7454 10180 7557
rect 10147 7417 10160 7454
rect 10060 7368 10160 7417
rect 1692 7080 1892 7124
rect 2160 7080 2260 7124
rect 2832 7080 2932 7124
rect 3504 7080 3604 7124
rect 4176 7080 4276 7124
rect 4848 7080 4948 7124
rect 5580 7080 5680 7124
rect 6252 7080 6352 7124
rect 6620 7080 6820 7124
rect 7068 7080 7268 7124
rect 7516 7080 7716 7124
rect 7964 7080 8164 7124
rect 8412 7080 8612 7124
rect 8860 7080 9060 7124
rect 10060 7080 10160 7124
rect 1936 6988 2036 7032
rect 2608 6988 2708 7032
rect 3280 6988 3380 7032
rect 3952 6988 4052 7032
rect 4624 6988 4724 7032
rect 5744 6988 5844 7032
rect 6416 6988 6516 7032
rect 7088 6988 7188 7032
rect 7516 6988 7716 7032
rect 7964 6988 8164 7032
rect 8432 6988 8532 7032
rect 9104 6988 9204 7032
rect 9308 6988 9408 7032
rect 9588 6988 9688 7032
rect 9792 6988 9892 7032
rect 9996 6988 10096 7032
rect 1936 6695 2036 6744
rect 1936 6658 1949 6695
rect 1916 6555 1949 6658
rect 1995 6555 2036 6695
rect 2608 6695 2708 6744
rect 2608 6658 2621 6695
rect 1916 6504 2036 6555
rect 2588 6555 2621 6658
rect 2667 6555 2708 6695
rect 3280 6695 3380 6744
rect 3280 6658 3293 6695
rect 2588 6504 2708 6555
rect 3260 6555 3293 6658
rect 3339 6555 3380 6695
rect 3952 6695 4052 6744
rect 3952 6658 3965 6695
rect 3260 6504 3380 6555
rect 3932 6555 3965 6658
rect 4011 6555 4052 6695
rect 4624 6695 4724 6744
rect 4624 6658 4637 6695
rect 3932 6504 4052 6555
rect 4604 6555 4637 6658
rect 4683 6555 4724 6695
rect 5744 6695 5844 6744
rect 5744 6658 5757 6695
rect 4604 6504 4724 6555
rect 5724 6555 5757 6658
rect 5803 6555 5844 6695
rect 6416 6695 6516 6744
rect 6416 6658 6429 6695
rect 5724 6504 5844 6555
rect 6396 6555 6429 6658
rect 6475 6555 6516 6695
rect 7088 6695 7188 6744
rect 7088 6658 7101 6695
rect 6396 6504 6516 6555
rect 7068 6555 7101 6658
rect 7147 6555 7188 6695
rect 7516 6710 7716 6744
rect 7516 6664 7552 6710
rect 7692 6664 7716 6710
rect 7516 6647 7716 6664
rect 7964 6710 8164 6744
rect 7964 6664 8000 6710
rect 8140 6664 8164 6710
rect 7964 6647 8164 6664
rect 8432 6695 8532 6744
rect 8432 6658 8445 6695
rect 7068 6504 7188 6555
rect 7516 6583 7716 6596
rect 7516 6537 7544 6583
rect 7684 6537 7716 6583
rect 7516 6504 7716 6537
rect 7964 6583 8164 6596
rect 7964 6537 7992 6583
rect 8132 6537 8164 6583
rect 7964 6504 8164 6537
rect 8412 6555 8445 6658
rect 8491 6555 8532 6695
rect 8412 6504 8532 6555
rect 9104 6687 9204 6876
rect 9104 6641 9139 6687
rect 9185 6641 9204 6687
rect 1916 6296 2036 6340
rect 2588 6296 2708 6340
rect 3260 6296 3380 6340
rect 3932 6296 4052 6340
rect 4604 6296 4724 6340
rect 9104 6481 9204 6641
rect 9084 6437 9204 6481
rect 9308 6687 9408 6876
rect 9308 6641 9346 6687
rect 9392 6641 9408 6687
rect 9308 6481 9408 6641
rect 9588 6583 9688 6744
rect 9588 6548 9605 6583
rect 9568 6537 9605 6548
rect 9651 6537 9688 6583
rect 9568 6504 9688 6537
rect 9792 6586 9892 6744
rect 9792 6540 9805 6586
rect 9851 6548 9892 6586
rect 9996 6692 10096 6744
rect 9996 6646 10009 6692
rect 10055 6646 10096 6692
rect 9996 6548 10096 6646
rect 9851 6540 9912 6548
rect 9792 6504 9912 6540
rect 9976 6504 10096 6548
rect 9308 6437 9428 6481
rect 5724 6296 5844 6340
rect 6396 6296 6516 6340
rect 7068 6296 7188 6340
rect 7516 6296 7716 6340
rect 7964 6296 8164 6340
rect 8412 6296 8532 6340
rect 9084 6321 9204 6365
rect 9308 6321 9428 6365
rect 9568 6296 9688 6340
rect 9792 6296 9912 6340
rect 9976 6296 10096 6340
rect 1804 6204 1924 6248
rect 2476 6204 2596 6248
rect 3148 6204 3268 6248
rect 3820 6204 3940 6248
rect 4492 6204 4612 6248
rect 5164 6204 5284 6248
rect 5836 6204 5956 6248
rect 6508 6204 6628 6248
rect 6956 6204 7156 6248
rect 7740 6204 7860 6248
rect 8412 6204 8532 6248
rect 8860 6204 9060 6248
rect 10060 6204 10180 6248
rect 1804 5989 1924 6040
rect 1804 5886 1837 5989
rect 1824 5849 1837 5886
rect 1883 5849 1924 5989
rect 2476 5989 2596 6040
rect 2476 5886 2509 5989
rect 1824 5800 1924 5849
rect 2496 5849 2509 5886
rect 2555 5849 2596 5989
rect 3148 5989 3268 6040
rect 3148 5886 3181 5989
rect 2496 5800 2596 5849
rect 3168 5849 3181 5886
rect 3227 5849 3268 5989
rect 3820 5989 3940 6040
rect 3820 5886 3853 5989
rect 3168 5800 3268 5849
rect 3840 5849 3853 5886
rect 3899 5849 3940 5989
rect 4492 5989 4612 6040
rect 4492 5886 4525 5989
rect 3840 5800 3940 5849
rect 4512 5849 4525 5886
rect 4571 5849 4612 5989
rect 5164 5989 5284 6040
rect 5164 5886 5197 5989
rect 4512 5800 4612 5849
rect 5184 5849 5197 5886
rect 5243 5849 5284 5989
rect 5836 5989 5956 6040
rect 5836 5886 5869 5989
rect 5184 5800 5284 5849
rect 5856 5849 5869 5886
rect 5915 5849 5956 5989
rect 6508 5989 6628 6040
rect 6508 5886 6541 5989
rect 5856 5800 5956 5849
rect 6528 5849 6541 5886
rect 6587 5849 6628 5989
rect 6956 6007 7156 6040
rect 6956 5961 6984 6007
rect 7124 5961 7156 6007
rect 6956 5948 7156 5961
rect 7740 5989 7860 6040
rect 6528 5800 6628 5849
rect 6956 5880 7156 5897
rect 7740 5886 7773 5989
rect 6956 5834 6992 5880
rect 7132 5834 7156 5880
rect 6956 5800 7156 5834
rect 7760 5849 7773 5886
rect 7819 5849 7860 5989
rect 8412 5989 8532 6040
rect 8412 5886 8445 5989
rect 7760 5800 7860 5849
rect 8432 5849 8445 5886
rect 8491 5849 8532 5989
rect 8860 6007 9060 6040
rect 8860 5961 8888 6007
rect 9028 5961 9060 6007
rect 8860 5948 9060 5961
rect 10060 5989 10180 6040
rect 8432 5800 8532 5849
rect 8860 5880 9060 5897
rect 8860 5834 8896 5880
rect 9036 5834 9060 5880
rect 8860 5800 9060 5834
rect 10060 5849 10101 5989
rect 10147 5886 10180 5989
rect 10147 5849 10160 5886
rect 10060 5800 10160 5849
rect 1824 5512 1924 5556
rect 2496 5512 2596 5556
rect 3168 5512 3268 5556
rect 3840 5512 3940 5556
rect 4512 5512 4612 5556
rect 5184 5512 5284 5556
rect 5856 5512 5956 5556
rect 6528 5512 6628 5556
rect 6956 5512 7156 5556
rect 7760 5512 7860 5556
rect 8432 5512 8532 5556
rect 8860 5512 9060 5556
rect 10060 5512 10160 5556
rect 1692 5420 1892 5464
rect 2160 5420 2260 5464
rect 2832 5420 2932 5464
rect 3504 5420 3604 5464
rect 4176 5420 4276 5464
rect 4848 5420 4948 5464
rect 5744 5420 5844 5464
rect 6172 5420 6372 5464
rect 6976 5420 7076 5464
rect 7648 5420 7748 5464
rect 8320 5420 8420 5464
rect 8748 5420 8948 5464
rect 9328 5420 9428 5464
rect 10060 5420 10160 5464
rect 1692 5142 1892 5176
rect 1692 5096 1728 5142
rect 1868 5096 1892 5142
rect 1692 5079 1892 5096
rect 2160 5127 2260 5176
rect 2160 5090 2173 5127
rect 1692 5015 1892 5028
rect 1692 4969 1720 5015
rect 1860 4969 1892 5015
rect 1692 4936 1892 4969
rect 2140 4987 2173 5090
rect 2219 4987 2260 5127
rect 2832 5127 2932 5176
rect 2832 5090 2845 5127
rect 2140 4936 2260 4987
rect 2812 4987 2845 5090
rect 2891 4987 2932 5127
rect 3504 5127 3604 5176
rect 3504 5090 3517 5127
rect 2812 4936 2932 4987
rect 3484 4987 3517 5090
rect 3563 4987 3604 5127
rect 4176 5127 4276 5176
rect 4176 5090 4189 5127
rect 3484 4936 3604 4987
rect 4156 4987 4189 5090
rect 4235 4987 4276 5127
rect 4848 5127 4948 5176
rect 4848 5090 4861 5127
rect 4156 4936 4276 4987
rect 4828 4987 4861 5090
rect 4907 4987 4948 5127
rect 5744 5127 5844 5176
rect 5744 5090 5757 5127
rect 4828 4936 4948 4987
rect 5724 4987 5757 5090
rect 5803 4987 5844 5127
rect 6172 5142 6372 5176
rect 6172 5096 6208 5142
rect 6348 5096 6372 5142
rect 6172 5079 6372 5096
rect 6976 5127 7076 5176
rect 6976 5090 6989 5127
rect 5724 4936 5844 4987
rect 6172 5015 6372 5028
rect 6172 4969 6200 5015
rect 6340 4969 6372 5015
rect 6172 4936 6372 4969
rect 6956 4987 6989 5090
rect 7035 4987 7076 5127
rect 7648 5127 7748 5176
rect 7648 5090 7661 5127
rect 6956 4936 7076 4987
rect 7628 4987 7661 5090
rect 7707 4987 7748 5127
rect 8320 5127 8420 5176
rect 8320 5090 8333 5127
rect 7628 4936 7748 4987
rect 8300 4987 8333 5090
rect 8379 4987 8420 5127
rect 8748 5142 8948 5176
rect 8748 5096 8784 5142
rect 8924 5096 8948 5142
rect 8748 5079 8948 5096
rect 9328 5127 9428 5176
rect 9328 5090 9341 5127
rect 8300 4936 8420 4987
rect 8748 5015 8948 5028
rect 8748 4969 8776 5015
rect 8916 4969 8948 5015
rect 8748 4936 8948 4969
rect 9308 4987 9341 5090
rect 9387 4987 9428 5127
rect 9308 4936 9428 4987
rect 10060 5127 10160 5176
rect 10060 4987 10101 5127
rect 10147 5090 10160 5127
rect 10147 4987 10180 5090
rect 10060 4936 10180 4987
rect 1692 4728 1892 4772
rect 2140 4728 2260 4772
rect 2812 4728 2932 4772
rect 3484 4728 3604 4772
rect 4156 4728 4276 4772
rect 4828 4728 4948 4772
rect 5724 4728 5844 4772
rect 6172 4728 6372 4772
rect 6956 4728 7076 4772
rect 7628 4728 7748 4772
rect 8300 4728 8420 4772
rect 8748 4728 8948 4772
rect 9308 4728 9428 4772
rect 10060 4728 10180 4772
rect 1916 4636 2036 4680
rect 2588 4636 2708 4680
rect 3260 4636 3380 4680
rect 3932 4636 4052 4680
rect 4604 4636 4724 4680
rect 5052 4636 5252 4680
rect 5724 4636 5844 4680
rect 6396 4636 6516 4680
rect 7068 4636 7188 4680
rect 7740 4636 7860 4680
rect 8412 4636 8532 4680
rect 8860 4636 9060 4680
rect 9980 4636 10100 4680
rect 1916 4421 2036 4472
rect 1916 4318 1949 4421
rect 1936 4281 1949 4318
rect 1995 4281 2036 4421
rect 2588 4421 2708 4472
rect 2588 4318 2621 4421
rect 1936 4232 2036 4281
rect 2608 4281 2621 4318
rect 2667 4281 2708 4421
rect 3260 4421 3380 4472
rect 3260 4318 3293 4421
rect 2608 4232 2708 4281
rect 3280 4281 3293 4318
rect 3339 4281 3380 4421
rect 3932 4421 4052 4472
rect 3932 4318 3965 4421
rect 3280 4232 3380 4281
rect 3952 4281 3965 4318
rect 4011 4281 4052 4421
rect 4604 4421 4724 4472
rect 4604 4318 4637 4421
rect 3952 4232 4052 4281
rect 4624 4281 4637 4318
rect 4683 4281 4724 4421
rect 5052 4439 5252 4472
rect 5052 4393 5080 4439
rect 5220 4393 5252 4439
rect 5052 4380 5252 4393
rect 5724 4421 5844 4472
rect 4624 4232 4724 4281
rect 5052 4312 5252 4329
rect 5724 4318 5757 4421
rect 5052 4266 5088 4312
rect 5228 4266 5252 4312
rect 5052 4232 5252 4266
rect 5744 4281 5757 4318
rect 5803 4281 5844 4421
rect 6396 4421 6516 4472
rect 6396 4318 6429 4421
rect 5744 4232 5844 4281
rect 6416 4281 6429 4318
rect 6475 4281 6516 4421
rect 7068 4421 7188 4472
rect 7068 4318 7101 4421
rect 6416 4232 6516 4281
rect 7088 4281 7101 4318
rect 7147 4281 7188 4421
rect 7740 4421 7860 4472
rect 7740 4318 7773 4421
rect 7088 4232 7188 4281
rect 7760 4281 7773 4318
rect 7819 4281 7860 4421
rect 8412 4421 8532 4472
rect 8412 4318 8445 4421
rect 7760 4232 7860 4281
rect 8432 4281 8445 4318
rect 8491 4281 8532 4421
rect 8860 4439 9060 4472
rect 8860 4393 8888 4439
rect 9028 4393 9060 4439
rect 8860 4380 9060 4393
rect 9980 4421 10100 4472
rect 8432 4232 8532 4281
rect 8860 4312 9060 4329
rect 8860 4266 8896 4312
rect 9036 4266 9060 4312
rect 8860 4232 9060 4266
rect 9980 4318 10013 4421
rect 10000 4281 10013 4318
rect 10059 4281 10100 4421
rect 10000 4232 10100 4281
rect 1936 3944 2036 3988
rect 2608 3944 2708 3988
rect 3280 3944 3380 3988
rect 3952 3944 4052 3988
rect 4624 3944 4724 3988
rect 5052 3944 5252 3988
rect 5744 3944 5844 3988
rect 6416 3944 6516 3988
rect 7088 3944 7188 3988
rect 7760 3944 7860 3988
rect 8432 3944 8532 3988
rect 8860 3944 9060 3988
rect 10000 3944 10100 3988
rect 1996 3852 2096 3896
rect 2608 3852 2708 3896
rect 3280 3852 3380 3896
rect 3952 3852 4052 3896
rect 4624 3852 4724 3896
rect 5744 3852 5844 3896
rect 6172 3852 6372 3896
rect 6640 3852 6740 3896
rect 7312 3852 7412 3896
rect 8044 3852 8144 3896
rect 8656 3852 8756 3896
rect 9532 3852 9732 3896
rect 10000 3852 10100 3896
rect 1996 3559 2096 3608
rect 1996 3419 2037 3559
rect 2083 3522 2096 3559
rect 2608 3559 2708 3608
rect 2608 3522 2621 3559
rect 2083 3419 2116 3522
rect 1996 3368 2116 3419
rect 2588 3419 2621 3522
rect 2667 3419 2708 3559
rect 3280 3559 3380 3608
rect 3280 3522 3293 3559
rect 2588 3368 2708 3419
rect 3260 3419 3293 3522
rect 3339 3419 3380 3559
rect 3952 3559 4052 3608
rect 3952 3522 3965 3559
rect 3260 3368 3380 3419
rect 3932 3419 3965 3522
rect 4011 3419 4052 3559
rect 4624 3559 4724 3608
rect 4624 3522 4637 3559
rect 3932 3368 4052 3419
rect 4604 3419 4637 3522
rect 4683 3419 4724 3559
rect 5744 3559 5844 3608
rect 5744 3522 5757 3559
rect 4604 3368 4724 3419
rect 5724 3419 5757 3522
rect 5803 3419 5844 3559
rect 6172 3574 6372 3608
rect 6172 3528 6208 3574
rect 6348 3528 6372 3574
rect 6172 3511 6372 3528
rect 6640 3559 6740 3608
rect 6640 3522 6653 3559
rect 5724 3368 5844 3419
rect 6172 3447 6372 3460
rect 6172 3401 6200 3447
rect 6340 3401 6372 3447
rect 6172 3368 6372 3401
rect 6620 3419 6653 3522
rect 6699 3419 6740 3559
rect 7312 3559 7412 3608
rect 7312 3522 7325 3559
rect 6620 3368 6740 3419
rect 7292 3419 7325 3522
rect 7371 3419 7412 3559
rect 7292 3368 7412 3419
rect 8044 3559 8144 3608
rect 8044 3419 8085 3559
rect 8131 3522 8144 3559
rect 8656 3559 8756 3608
rect 8656 3522 8669 3559
rect 8131 3419 8164 3522
rect 8044 3368 8164 3419
rect 8636 3419 8669 3522
rect 8715 3419 8756 3559
rect 9532 3574 9732 3608
rect 9532 3528 9568 3574
rect 9708 3528 9732 3574
rect 9532 3511 9732 3528
rect 10000 3559 10100 3608
rect 10000 3522 10013 3559
rect 8636 3368 8756 3419
rect 9532 3447 9732 3460
rect 9532 3401 9560 3447
rect 9700 3401 9732 3447
rect 1996 3160 2116 3204
rect 2588 3160 2708 3204
rect 3260 3160 3380 3204
rect 3932 3160 4052 3204
rect 4604 3160 4724 3204
rect 9532 3368 9732 3401
rect 9980 3419 10013 3522
rect 10059 3419 10100 3559
rect 9980 3368 10100 3419
rect 5724 3160 5844 3204
rect 6172 3160 6372 3204
rect 6620 3160 6740 3204
rect 7292 3160 7412 3204
rect 8044 3160 8164 3204
rect 8636 3160 8756 3204
rect 9532 3160 9732 3204
rect 9980 3160 10100 3204
<< polycontact >>
rect 1728 8232 1868 8278
rect 1720 8105 1860 8151
rect 2173 8123 2219 8263
rect 2845 8123 2891 8263
rect 3517 8123 3563 8263
rect 4189 8123 4235 8263
rect 4861 8123 4907 8263
rect 5648 8232 5788 8278
rect 6096 8232 6236 8278
rect 6544 8232 6684 8278
rect 6992 8232 7132 8278
rect 7440 8232 7580 8278
rect 7888 8232 8028 8278
rect 8336 8232 8476 8278
rect 8784 8232 8924 8278
rect 9568 8232 9708 8278
rect 10016 8232 10156 8278
rect 5640 8105 5780 8151
rect 6088 8105 6228 8151
rect 6536 8105 6676 8151
rect 6984 8105 7124 8151
rect 7432 8105 7572 8151
rect 7880 8105 8020 8151
rect 8328 8105 8468 8151
rect 8776 8105 8916 8151
rect 9560 8105 9700 8151
rect 10008 8105 10148 8151
rect 1720 7529 1860 7575
rect 1728 7402 1868 7448
rect 2173 7417 2219 7557
rect 2845 7417 2891 7557
rect 3517 7417 3563 7557
rect 4189 7417 4235 7557
rect 4861 7417 4907 7557
rect 5621 7417 5667 7557
rect 6293 7417 6339 7557
rect 6648 7529 6788 7575
rect 7096 7529 7236 7575
rect 7544 7529 7684 7575
rect 7992 7529 8132 7575
rect 8440 7529 8580 7575
rect 8888 7529 9028 7575
rect 6656 7402 6796 7448
rect 7104 7402 7244 7448
rect 7552 7402 7692 7448
rect 8000 7402 8140 7448
rect 8448 7402 8588 7448
rect 8896 7402 9036 7448
rect 10101 7417 10147 7557
rect 1949 6555 1995 6695
rect 2621 6555 2667 6695
rect 3293 6555 3339 6695
rect 3965 6555 4011 6695
rect 4637 6555 4683 6695
rect 5757 6555 5803 6695
rect 6429 6555 6475 6695
rect 7101 6555 7147 6695
rect 7552 6664 7692 6710
rect 8000 6664 8140 6710
rect 7544 6537 7684 6583
rect 7992 6537 8132 6583
rect 8445 6555 8491 6695
rect 9139 6641 9185 6687
rect 9346 6641 9392 6687
rect 9605 6537 9651 6583
rect 9805 6540 9851 6586
rect 10009 6646 10055 6692
rect 1837 5849 1883 5989
rect 2509 5849 2555 5989
rect 3181 5849 3227 5989
rect 3853 5849 3899 5989
rect 4525 5849 4571 5989
rect 5197 5849 5243 5989
rect 5869 5849 5915 5989
rect 6541 5849 6587 5989
rect 6984 5961 7124 6007
rect 6992 5834 7132 5880
rect 7773 5849 7819 5989
rect 8445 5849 8491 5989
rect 8888 5961 9028 6007
rect 8896 5834 9036 5880
rect 10101 5849 10147 5989
rect 1728 5096 1868 5142
rect 1720 4969 1860 5015
rect 2173 4987 2219 5127
rect 2845 4987 2891 5127
rect 3517 4987 3563 5127
rect 4189 4987 4235 5127
rect 4861 4987 4907 5127
rect 5757 4987 5803 5127
rect 6208 5096 6348 5142
rect 6200 4969 6340 5015
rect 6989 4987 7035 5127
rect 7661 4987 7707 5127
rect 8333 4987 8379 5127
rect 8784 5096 8924 5142
rect 8776 4969 8916 5015
rect 9341 4987 9387 5127
rect 10101 4987 10147 5127
rect 1949 4281 1995 4421
rect 2621 4281 2667 4421
rect 3293 4281 3339 4421
rect 3965 4281 4011 4421
rect 4637 4281 4683 4421
rect 5080 4393 5220 4439
rect 5088 4266 5228 4312
rect 5757 4281 5803 4421
rect 6429 4281 6475 4421
rect 7101 4281 7147 4421
rect 7773 4281 7819 4421
rect 8445 4281 8491 4421
rect 8888 4393 9028 4439
rect 8896 4266 9036 4312
rect 10013 4281 10059 4421
rect 2037 3419 2083 3559
rect 2621 3419 2667 3559
rect 3293 3419 3339 3559
rect 3965 3419 4011 3559
rect 4637 3419 4683 3559
rect 5757 3419 5803 3559
rect 6208 3528 6348 3574
rect 6200 3401 6340 3447
rect 6653 3419 6699 3559
rect 7325 3419 7371 3559
rect 8085 3419 8131 3559
rect 8669 3419 8715 3559
rect 9568 3528 9708 3574
rect 9560 3401 9700 3447
rect 10013 3419 10059 3559
<< metal1 >>
rect 1344 8650 10640 8684
rect 1344 8598 2376 8650
rect 2636 8598 4700 8650
rect 4960 8598 7024 8650
rect 7284 8598 9348 8650
rect 9608 8598 10640 8650
rect 1344 8564 10640 8598
rect 1418 8539 1486 8564
rect 1418 8493 1429 8539
rect 1475 8493 1486 8539
rect 1418 8411 1486 8493
rect 1418 8365 1429 8411
rect 1475 8365 1486 8411
rect 1418 8283 1486 8365
rect 1418 8237 1429 8283
rect 1475 8237 1486 8283
rect 1418 8224 1486 8237
rect 1617 8497 1663 8518
rect 1617 8151 1663 8357
rect 1921 8497 1967 8564
rect 1921 8338 1967 8357
rect 2085 8505 2131 8564
rect 2085 8346 2131 8365
rect 2269 8505 2335 8518
rect 2269 8365 2289 8505
rect 1714 8232 1728 8278
rect 1868 8232 1967 8278
rect 1617 8105 1720 8151
rect 1860 8105 1872 8151
rect 1418 8066 1486 8078
rect 1418 7919 1429 8066
rect 1475 7919 1486 8066
rect 1418 7900 1486 7919
rect 1617 8032 1663 8059
rect 1617 7900 1663 7986
rect 1921 8032 1967 8232
rect 2158 8263 2223 8280
rect 2158 8146 2173 8263
rect 2219 8123 2223 8263
rect 2210 8094 2223 8123
rect 2158 8080 2223 8094
rect 1921 7946 1967 7986
rect 2065 8032 2111 8072
rect 2065 7900 2111 7986
rect 2269 8034 2335 8365
rect 2757 8505 2803 8564
rect 2757 8346 2803 8365
rect 2941 8505 3007 8518
rect 2941 8365 2961 8505
rect 2830 8263 2895 8280
rect 2830 8146 2845 8263
rect 2891 8123 2895 8263
rect 2882 8094 2895 8123
rect 2830 8080 2895 8094
rect 2269 7982 2270 8034
rect 2322 8032 2335 8034
rect 2322 7982 2335 7986
rect 2269 7946 2335 7982
rect 2737 8032 2783 8072
rect 2737 7900 2783 7986
rect 2941 8034 3007 8365
rect 3429 8505 3475 8564
rect 3429 8346 3475 8365
rect 3613 8505 3679 8518
rect 3613 8365 3633 8505
rect 3502 8263 3567 8280
rect 3502 8146 3517 8263
rect 3563 8123 3567 8263
rect 3554 8094 3567 8123
rect 3502 8080 3567 8094
rect 3613 8146 3679 8365
rect 4101 8505 4147 8564
rect 4101 8346 4147 8365
rect 4285 8505 4351 8518
rect 4285 8365 4305 8505
rect 3613 8094 3614 8146
rect 3666 8094 3679 8146
rect 2941 7982 2942 8034
rect 2994 8032 3007 8034
rect 2994 7982 3007 7986
rect 2941 7946 3007 7982
rect 3409 8032 3455 8072
rect 3409 7900 3455 7986
rect 3613 8032 3679 8094
rect 4174 8263 4239 8280
rect 4174 8146 4189 8263
rect 4235 8123 4239 8263
rect 4226 8094 4239 8123
rect 4174 8080 4239 8094
rect 3613 7986 3633 8032
rect 3613 7946 3679 7986
rect 4081 8032 4127 8072
rect 4081 7900 4127 7986
rect 4285 8034 4351 8365
rect 4773 8505 4819 8564
rect 5342 8539 5410 8564
rect 4773 8346 4819 8365
rect 4957 8505 5023 8518
rect 4957 8365 4977 8505
rect 4846 8263 4911 8280
rect 4846 8146 4861 8263
rect 4907 8123 4911 8263
rect 4898 8094 4911 8123
rect 4846 8080 4911 8094
rect 4285 7982 4286 8034
rect 4338 8032 4351 8034
rect 4338 7982 4351 7986
rect 4285 7946 4351 7982
rect 4753 8032 4799 8072
rect 4753 7900 4799 7986
rect 4957 8034 5023 8365
rect 5342 8493 5353 8539
rect 5399 8493 5410 8539
rect 5342 8411 5410 8493
rect 5342 8365 5353 8411
rect 5399 8365 5410 8411
rect 5342 8283 5410 8365
rect 5342 8237 5353 8283
rect 5399 8237 5410 8283
rect 5342 8226 5410 8237
rect 5537 8497 5583 8518
rect 5537 8151 5583 8357
rect 5841 8497 5887 8564
rect 5841 8338 5887 8357
rect 5985 8497 6031 8518
rect 5634 8232 5648 8278
rect 5788 8232 5887 8278
rect 5537 8105 5640 8151
rect 5780 8105 5792 8151
rect 4957 7982 4958 8034
rect 5010 8032 5023 8034
rect 5010 7982 5023 7986
rect 4957 7946 5023 7982
rect 5342 8066 5410 8077
rect 5342 7919 5353 8066
rect 5399 7919 5410 8066
rect 5342 7900 5410 7919
rect 5537 8032 5583 8049
rect 5537 7900 5583 7986
rect 5841 8032 5887 8232
rect 5985 8151 6031 8357
rect 6289 8497 6335 8564
rect 6289 8338 6335 8357
rect 6433 8497 6479 8518
rect 6082 8232 6096 8278
rect 6236 8232 6335 8278
rect 5985 8105 6088 8151
rect 6228 8105 6240 8151
rect 5841 7946 5887 7986
rect 5985 8032 6031 8049
rect 5985 7900 6031 7986
rect 6289 8032 6335 8232
rect 6433 8151 6479 8357
rect 6737 8497 6783 8564
rect 6737 8338 6783 8357
rect 6881 8497 6927 8518
rect 6530 8232 6544 8278
rect 6684 8232 6783 8278
rect 6433 8105 6536 8151
rect 6676 8105 6688 8151
rect 6289 7946 6335 7986
rect 6433 8032 6479 8049
rect 6433 7900 6479 7986
rect 6737 8032 6783 8232
rect 6881 8151 6927 8357
rect 7185 8497 7231 8564
rect 7185 8338 7231 8357
rect 7329 8497 7375 8518
rect 6978 8232 6992 8278
rect 7132 8232 7231 8278
rect 6881 8105 6984 8151
rect 7124 8105 7136 8151
rect 6737 7946 6783 7986
rect 6881 8032 6927 8049
rect 6881 7900 6927 7986
rect 7185 8032 7231 8232
rect 7329 8151 7375 8357
rect 7633 8497 7679 8564
rect 7633 8338 7679 8357
rect 7777 8497 7823 8518
rect 7426 8232 7440 8278
rect 7580 8232 7679 8278
rect 7329 8105 7432 8151
rect 7572 8105 7584 8151
rect 7185 7946 7231 7986
rect 7329 8032 7375 8049
rect 7329 7900 7375 7986
rect 7633 8032 7679 8232
rect 7777 8151 7823 8357
rect 8081 8497 8127 8564
rect 8081 8338 8127 8357
rect 8225 8497 8271 8518
rect 7874 8232 7888 8278
rect 8028 8232 8127 8278
rect 7777 8105 7880 8151
rect 8020 8105 8032 8151
rect 7633 7946 7679 7986
rect 7777 8032 7823 8049
rect 7777 7900 7823 7986
rect 8081 8032 8127 8232
rect 8225 8151 8271 8357
rect 8529 8497 8575 8564
rect 8529 8338 8575 8357
rect 8673 8497 8719 8518
rect 8322 8232 8336 8278
rect 8476 8232 8575 8278
rect 8225 8105 8328 8151
rect 8468 8105 8480 8151
rect 8081 7946 8127 7986
rect 8225 8032 8271 8049
rect 8225 7900 8271 7986
rect 8529 8032 8575 8232
rect 8673 8151 8719 8357
rect 8977 8497 9023 8564
rect 8977 8338 9023 8357
rect 9262 8539 9330 8564
rect 9262 8493 9273 8539
rect 9319 8493 9330 8539
rect 9262 8411 9330 8493
rect 9262 8365 9273 8411
rect 9319 8365 9330 8411
rect 9262 8283 9330 8365
rect 8770 8232 8784 8278
rect 8924 8232 9023 8278
rect 8673 8105 8776 8151
rect 8916 8105 8928 8151
rect 8529 7946 8575 7986
rect 8673 8032 8719 8049
rect 8673 7900 8719 7986
rect 8977 8032 9023 8232
rect 9262 8237 9273 8283
rect 9319 8237 9330 8283
rect 9262 8226 9330 8237
rect 9457 8497 9503 8518
rect 9457 8151 9503 8357
rect 9761 8497 9807 8564
rect 9761 8338 9807 8357
rect 9905 8497 9951 8518
rect 9554 8232 9568 8278
rect 9708 8232 9807 8278
rect 9457 8105 9560 8151
rect 9700 8105 9712 8151
rect 8977 7946 9023 7986
rect 9262 8066 9330 8077
rect 9262 7919 9273 8066
rect 9319 7919 9330 8066
rect 9262 7900 9330 7919
rect 9457 8032 9503 8057
rect 9457 7900 9503 7986
rect 9761 8032 9807 8232
rect 9905 8151 9951 8357
rect 10209 8497 10255 8564
rect 10209 8338 10255 8357
rect 10498 8539 10566 8564
rect 10498 8493 10509 8539
rect 10555 8493 10566 8539
rect 10498 8411 10566 8493
rect 10498 8365 10509 8411
rect 10555 8365 10566 8411
rect 10498 8283 10566 8365
rect 10002 8232 10016 8278
rect 10156 8232 10255 8278
rect 9905 8105 10008 8151
rect 10148 8105 10160 8151
rect 9761 7946 9807 7986
rect 9905 8032 9951 8057
rect 9905 7900 9951 7986
rect 10209 8032 10255 8232
rect 10498 8237 10509 8283
rect 10555 8237 10566 8283
rect 10498 8224 10566 8237
rect 10209 7946 10255 7986
rect 10498 8066 10566 8078
rect 10498 7919 10509 8066
rect 10555 7919 10566 8066
rect 10498 7900 10566 7919
rect 1344 7866 10800 7900
rect 1344 7814 3538 7866
rect 3798 7814 5862 7866
rect 6122 7814 8186 7866
rect 8446 7814 10510 7866
rect 10770 7814 10800 7866
rect 1344 7780 10800 7814
rect 1418 7761 1486 7780
rect 1418 7614 1429 7761
rect 1475 7614 1486 7761
rect 1617 7694 1663 7780
rect 1617 7621 1663 7648
rect 1921 7694 1967 7734
rect 1418 7602 1486 7614
rect 1617 7529 1720 7575
rect 1860 7529 1872 7575
rect 1418 7443 1486 7456
rect 1418 7397 1429 7443
rect 1475 7397 1486 7443
rect 1418 7315 1486 7397
rect 1418 7269 1429 7315
rect 1475 7269 1486 7315
rect 1418 7187 1486 7269
rect 1418 7141 1429 7187
rect 1475 7141 1486 7187
rect 1617 7323 1663 7529
rect 1921 7448 1967 7648
rect 2065 7694 2111 7780
rect 2065 7608 2111 7648
rect 2269 7694 2335 7734
rect 2269 7648 2289 7694
rect 1714 7402 1728 7448
rect 1868 7402 1967 7448
rect 2158 7557 2223 7600
rect 2158 7474 2173 7557
rect 2158 7417 2173 7422
rect 2219 7417 2223 7557
rect 2158 7400 2223 7417
rect 1617 7162 1663 7183
rect 1921 7323 1967 7342
rect 1418 7116 1486 7141
rect 1921 7116 1967 7183
rect 2085 7315 2131 7334
rect 2085 7116 2131 7175
rect 2269 7315 2335 7648
rect 2737 7694 2783 7780
rect 2737 7608 2783 7648
rect 2941 7694 3007 7734
rect 2941 7648 2961 7694
rect 2830 7557 2895 7600
rect 2830 7474 2845 7557
rect 2830 7417 2845 7422
rect 2891 7417 2895 7557
rect 2830 7400 2895 7417
rect 2941 7474 3007 7648
rect 3409 7694 3455 7780
rect 3409 7608 3455 7648
rect 3613 7694 3679 7734
rect 3613 7648 3633 7694
rect 2941 7422 2942 7474
rect 2994 7422 3007 7474
rect 2269 7250 2289 7315
rect 2269 7198 2270 7250
rect 2269 7175 2289 7198
rect 2269 7162 2335 7175
rect 2757 7315 2803 7334
rect 2757 7116 2803 7175
rect 2941 7315 3007 7422
rect 3502 7557 3567 7600
rect 3502 7474 3517 7557
rect 3502 7417 3517 7422
rect 3563 7417 3567 7557
rect 3502 7400 3567 7417
rect 2941 7175 2961 7315
rect 2941 7162 3007 7175
rect 3429 7315 3475 7334
rect 3429 7116 3475 7175
rect 3613 7315 3679 7648
rect 4081 7694 4127 7780
rect 4081 7608 4127 7648
rect 4285 7694 4351 7734
rect 4285 7648 4305 7694
rect 4174 7557 4239 7600
rect 4174 7474 4189 7557
rect 4174 7417 4189 7422
rect 4235 7417 4239 7557
rect 4174 7400 4239 7417
rect 4285 7474 4351 7648
rect 4753 7694 4799 7780
rect 4753 7608 4799 7648
rect 4957 7694 5023 7734
rect 4957 7648 4977 7694
rect 4285 7422 4286 7474
rect 4338 7422 4351 7474
rect 3613 7250 3633 7315
rect 3613 7198 3614 7250
rect 3613 7175 3633 7198
rect 3613 7162 3679 7175
rect 4101 7315 4147 7334
rect 4101 7116 4147 7175
rect 4285 7315 4351 7422
rect 4846 7557 4911 7600
rect 4846 7474 4861 7557
rect 4846 7417 4861 7422
rect 4907 7417 4911 7557
rect 4846 7400 4911 7417
rect 4957 7474 5023 7648
rect 4957 7422 4958 7474
rect 5010 7422 5023 7474
rect 4285 7175 4305 7315
rect 4285 7162 4351 7175
rect 4773 7315 4819 7334
rect 4773 7116 4819 7175
rect 4957 7315 5023 7422
rect 4957 7175 4977 7315
rect 4957 7162 5023 7175
rect 5505 7694 5571 7734
rect 5551 7648 5571 7694
rect 5505 7315 5571 7648
rect 5729 7694 5775 7780
rect 5729 7608 5775 7648
rect 6177 7694 6243 7734
rect 6223 7648 6243 7694
rect 5617 7557 5682 7600
rect 5617 7417 5621 7557
rect 5667 7474 5682 7557
rect 5667 7417 5682 7422
rect 5617 7400 5682 7417
rect 5551 7250 5571 7315
rect 5570 7198 5571 7250
rect 5551 7175 5571 7198
rect 5505 7162 5571 7175
rect 5709 7315 5755 7334
rect 5709 7116 5755 7175
rect 6177 7315 6243 7648
rect 6401 7694 6447 7780
rect 6401 7608 6447 7648
rect 6545 7694 6591 7780
rect 6545 7626 6591 7648
rect 6849 7694 6895 7734
rect 6289 7557 6354 7600
rect 6289 7417 6293 7557
rect 6339 7474 6354 7557
rect 6339 7417 6354 7422
rect 6289 7400 6354 7417
rect 6545 7529 6648 7575
rect 6788 7529 6800 7575
rect 6223 7250 6243 7315
rect 6242 7198 6243 7250
rect 6223 7175 6243 7198
rect 6177 7162 6243 7175
rect 6381 7315 6427 7334
rect 6381 7116 6427 7175
rect 6545 7323 6591 7529
rect 6849 7448 6895 7648
rect 6993 7694 7039 7780
rect 6993 7626 7039 7648
rect 7297 7694 7343 7734
rect 6642 7402 6656 7448
rect 6796 7402 6895 7448
rect 6993 7529 7096 7575
rect 7236 7529 7248 7575
rect 6545 7162 6591 7183
rect 6849 7323 6895 7342
rect 6849 7116 6895 7183
rect 6993 7323 7039 7529
rect 7297 7448 7343 7648
rect 7441 7694 7487 7780
rect 7441 7626 7487 7648
rect 7745 7694 7791 7734
rect 7090 7402 7104 7448
rect 7244 7402 7343 7448
rect 7441 7529 7544 7575
rect 7684 7529 7696 7575
rect 6993 7162 7039 7183
rect 7297 7323 7343 7342
rect 7297 7116 7343 7183
rect 7441 7323 7487 7529
rect 7745 7448 7791 7648
rect 7889 7694 7935 7780
rect 7889 7626 7935 7648
rect 8193 7694 8239 7734
rect 7538 7402 7552 7448
rect 7692 7402 7791 7448
rect 7889 7529 7992 7575
rect 8132 7529 8144 7575
rect 7441 7162 7487 7183
rect 7745 7323 7791 7342
rect 7745 7116 7791 7183
rect 7889 7323 7935 7529
rect 8193 7448 8239 7648
rect 8337 7694 8383 7780
rect 8337 7623 8383 7648
rect 8641 7694 8687 7734
rect 7986 7402 8000 7448
rect 8140 7402 8239 7448
rect 8337 7529 8440 7575
rect 8580 7529 8592 7575
rect 7889 7162 7935 7183
rect 8193 7323 8239 7342
rect 8193 7116 8239 7183
rect 8337 7323 8383 7529
rect 8641 7448 8687 7648
rect 8785 7694 8831 7780
rect 9374 7761 9442 7780
rect 8785 7623 8831 7648
rect 9089 7694 9135 7734
rect 8434 7402 8448 7448
rect 8588 7402 8687 7448
rect 8785 7529 8888 7575
rect 9028 7529 9040 7575
rect 8337 7162 8383 7183
rect 8641 7323 8687 7342
rect 8641 7116 8687 7183
rect 8785 7323 8831 7529
rect 9089 7448 9135 7648
rect 9374 7614 9385 7761
rect 9431 7614 9442 7761
rect 9374 7603 9442 7614
rect 9985 7694 10051 7734
rect 10031 7648 10051 7694
rect 8882 7402 8896 7448
rect 9036 7402 9135 7448
rect 9374 7443 9442 7454
rect 9374 7397 9385 7443
rect 9431 7397 9442 7443
rect 8785 7162 8831 7183
rect 9089 7323 9135 7342
rect 9089 7116 9135 7183
rect 9374 7315 9442 7397
rect 9374 7269 9385 7315
rect 9431 7269 9442 7315
rect 9374 7187 9442 7269
rect 9374 7141 9385 7187
rect 9431 7141 9442 7187
rect 9985 7315 10051 7648
rect 10209 7694 10255 7780
rect 10209 7608 10255 7648
rect 10498 7761 10566 7780
rect 10498 7614 10509 7761
rect 10555 7614 10566 7761
rect 10498 7602 10566 7614
rect 10097 7557 10162 7600
rect 10097 7417 10101 7557
rect 10147 7474 10162 7557
rect 10147 7417 10162 7422
rect 10097 7400 10162 7417
rect 10498 7443 10566 7456
rect 10498 7397 10509 7443
rect 10555 7397 10566 7443
rect 10031 7250 10051 7315
rect 10050 7198 10051 7250
rect 10031 7175 10051 7198
rect 9985 7162 10051 7175
rect 10189 7315 10235 7334
rect 9374 7116 9442 7141
rect 10189 7116 10235 7175
rect 10498 7315 10566 7397
rect 10498 7269 10509 7315
rect 10555 7269 10566 7315
rect 10498 7187 10566 7269
rect 10498 7141 10509 7187
rect 10555 7141 10566 7187
rect 10498 7116 10566 7141
rect 1344 7082 10640 7116
rect 1344 7030 2376 7082
rect 2636 7030 4700 7082
rect 4960 7030 7024 7082
rect 7284 7030 9348 7082
rect 9608 7030 10640 7082
rect 1344 6996 10640 7030
rect 1418 6971 1486 6996
rect 1418 6925 1429 6971
rect 1475 6925 1486 6971
rect 1418 6843 1486 6925
rect 1418 6797 1429 6843
rect 1475 6797 1486 6843
rect 1418 6715 1486 6797
rect 1861 6937 1907 6996
rect 1861 6778 1907 6797
rect 2045 6937 2111 6950
rect 2045 6797 2065 6937
rect 1418 6669 1429 6715
rect 1475 6669 1486 6715
rect 1418 6656 1486 6669
rect 1934 6695 1999 6712
rect 1934 6578 1949 6695
rect 1995 6555 1999 6695
rect 1986 6526 1999 6555
rect 1934 6512 1999 6526
rect 1418 6498 1486 6510
rect 1418 6351 1429 6498
rect 1475 6351 1486 6498
rect 1418 6332 1486 6351
rect 1841 6464 1887 6504
rect 1841 6332 1887 6418
rect 2045 6466 2111 6797
rect 2533 6937 2579 6996
rect 2533 6778 2579 6797
rect 2717 6937 2783 6950
rect 2717 6797 2737 6937
rect 2606 6695 2671 6712
rect 2606 6578 2621 6695
rect 2667 6555 2671 6695
rect 2658 6526 2671 6555
rect 2606 6512 2671 6526
rect 2045 6414 2046 6466
rect 2098 6464 2111 6466
rect 2098 6414 2111 6418
rect 2045 6378 2111 6414
rect 2513 6464 2559 6504
rect 2513 6332 2559 6418
rect 2717 6466 2783 6797
rect 3205 6937 3251 6996
rect 3205 6778 3251 6797
rect 3389 6937 3455 6950
rect 3389 6797 3409 6937
rect 3278 6695 3343 6712
rect 3278 6578 3293 6695
rect 3339 6555 3343 6695
rect 3330 6526 3343 6555
rect 3278 6512 3343 6526
rect 3389 6578 3455 6797
rect 3877 6937 3923 6996
rect 3877 6778 3923 6797
rect 4061 6937 4127 6950
rect 4061 6797 4081 6937
rect 3389 6526 3390 6578
rect 3442 6526 3455 6578
rect 2717 6414 2718 6466
rect 2770 6464 2783 6466
rect 2770 6414 2783 6418
rect 2717 6378 2783 6414
rect 3185 6464 3231 6504
rect 3185 6332 3231 6418
rect 3389 6464 3455 6526
rect 3950 6695 4015 6712
rect 3950 6578 3965 6695
rect 4011 6555 4015 6695
rect 4002 6526 4015 6555
rect 3950 6512 4015 6526
rect 3389 6418 3409 6464
rect 3389 6378 3455 6418
rect 3857 6464 3903 6504
rect 3857 6332 3903 6418
rect 4061 6466 4127 6797
rect 4549 6937 4595 6996
rect 5342 6971 5410 6996
rect 4549 6778 4595 6797
rect 4733 6937 4799 6950
rect 4733 6797 4753 6937
rect 4622 6695 4687 6712
rect 4622 6578 4637 6695
rect 4683 6555 4687 6695
rect 4674 6526 4687 6555
rect 4622 6512 4687 6526
rect 4061 6414 4062 6466
rect 4114 6464 4127 6466
rect 4114 6414 4127 6418
rect 4061 6378 4127 6414
rect 4529 6464 4575 6504
rect 4529 6332 4575 6418
rect 4733 6466 4799 6797
rect 5342 6925 5353 6971
rect 5399 6925 5410 6971
rect 5342 6843 5410 6925
rect 5342 6797 5353 6843
rect 5399 6797 5410 6843
rect 5342 6715 5410 6797
rect 5669 6937 5715 6996
rect 5669 6778 5715 6797
rect 5853 6937 5919 6950
rect 5853 6797 5873 6937
rect 5342 6669 5353 6715
rect 5399 6669 5410 6715
rect 5342 6658 5410 6669
rect 5742 6695 5807 6712
rect 5742 6578 5757 6695
rect 5803 6555 5807 6695
rect 5794 6526 5807 6555
rect 5742 6512 5807 6526
rect 4733 6414 4734 6466
rect 4786 6464 4799 6466
rect 4786 6414 4799 6418
rect 4733 6378 4799 6414
rect 5342 6498 5410 6509
rect 5342 6351 5353 6498
rect 5399 6351 5410 6498
rect 5342 6332 5410 6351
rect 5649 6464 5695 6504
rect 5649 6332 5695 6418
rect 5853 6466 5919 6797
rect 6341 6937 6387 6996
rect 6341 6778 6387 6797
rect 6525 6937 6591 6950
rect 6525 6797 6545 6937
rect 6414 6695 6479 6712
rect 6414 6578 6429 6695
rect 6475 6555 6479 6695
rect 6466 6526 6479 6555
rect 6414 6512 6479 6526
rect 5853 6414 5854 6466
rect 5906 6464 5919 6466
rect 5906 6414 5919 6418
rect 5853 6378 5919 6414
rect 6321 6464 6367 6504
rect 6321 6332 6367 6418
rect 6525 6466 6591 6797
rect 7013 6937 7059 6996
rect 7013 6778 7059 6797
rect 7197 6937 7263 6950
rect 7197 6797 7217 6937
rect 7086 6695 7151 6712
rect 7086 6578 7101 6695
rect 7147 6555 7151 6695
rect 7138 6526 7151 6555
rect 7086 6512 7151 6526
rect 7197 6578 7263 6797
rect 7197 6526 7198 6578
rect 7250 6526 7263 6578
rect 7441 6929 7487 6950
rect 7441 6583 7487 6789
rect 7745 6929 7791 6996
rect 7745 6770 7791 6789
rect 7889 6929 7935 6950
rect 7538 6664 7552 6710
rect 7692 6664 7791 6710
rect 7441 6537 7544 6583
rect 7684 6537 7696 6583
rect 6525 6414 6526 6466
rect 6578 6464 6591 6466
rect 6578 6414 6591 6418
rect 6525 6378 6591 6414
rect 6993 6464 7039 6504
rect 6993 6332 7039 6418
rect 7197 6464 7263 6526
rect 7197 6418 7217 6464
rect 7197 6378 7263 6418
rect 7441 6464 7487 6489
rect 7441 6332 7487 6418
rect 7745 6464 7791 6664
rect 7889 6583 7935 6789
rect 8193 6929 8239 6996
rect 8193 6770 8239 6789
rect 8357 6937 8403 6996
rect 9502 6975 9570 6996
rect 8357 6778 8403 6797
rect 8541 6937 8607 6950
rect 8541 6797 8561 6937
rect 7986 6664 8000 6710
rect 8140 6664 8239 6710
rect 7889 6537 7992 6583
rect 8132 6537 8144 6583
rect 7745 6378 7791 6418
rect 7889 6464 7935 6489
rect 7889 6332 7935 6418
rect 8193 6464 8239 6664
rect 8430 6695 8495 6712
rect 8430 6578 8445 6695
rect 8491 6555 8495 6695
rect 8482 6526 8495 6555
rect 8430 6512 8495 6526
rect 8193 6378 8239 6418
rect 8337 6464 8383 6504
rect 8337 6332 8383 6418
rect 8541 6466 8607 6797
rect 9018 6941 9086 6942
rect 9018 6895 9029 6941
rect 9075 6895 9086 6941
rect 9018 6530 9086 6895
rect 9502 6835 9513 6975
rect 9559 6835 9570 6975
rect 10498 6971 10566 6996
rect 9678 6904 9717 6950
rect 9763 6904 10125 6950
rect 10171 6904 10184 6950
rect 9678 6903 10184 6904
rect 10498 6925 10509 6971
rect 10555 6925 10566 6971
rect 9502 6830 9570 6835
rect 9136 6784 9425 6818
rect 9910 6811 9921 6857
rect 9967 6811 10168 6857
rect 10104 6802 10168 6811
rect 9762 6784 9774 6802
rect 9136 6750 9774 6784
rect 9826 6784 9838 6802
rect 9826 6750 9859 6784
rect 9136 6738 9859 6750
rect 9136 6687 9272 6738
rect 9811 6703 9859 6738
rect 10104 6750 10110 6802
rect 10162 6750 10168 6802
rect 9811 6692 10058 6703
rect 9136 6641 9139 6687
rect 9185 6641 9272 6687
rect 9136 6610 9272 6641
rect 9335 6690 9763 6692
rect 9335 6687 9662 6690
rect 9335 6641 9346 6687
rect 9392 6641 9662 6687
rect 9335 6638 9662 6641
rect 9714 6638 9763 6690
rect 9335 6636 9763 6638
rect 9717 6586 9763 6636
rect 9811 6646 10009 6692
rect 10055 6646 10058 6692
rect 9811 6632 10058 6646
rect 9594 6537 9605 6583
rect 9651 6537 9662 6583
rect 9717 6540 9805 6586
rect 9851 6540 9865 6586
rect 9594 6530 9662 6537
rect 9018 6470 9662 6530
rect 10104 6494 10168 6750
rect 10498 6843 10566 6925
rect 10498 6797 10509 6843
rect 10555 6797 10566 6843
rect 10498 6715 10566 6797
rect 10498 6669 10509 6715
rect 10555 6669 10566 6715
rect 10498 6656 10566 6669
rect 8541 6414 8542 6466
rect 8594 6464 8607 6466
rect 9222 6424 9290 6470
rect 9717 6447 10168 6494
rect 10498 6498 10566 6510
rect 9717 6441 9763 6447
rect 8594 6414 8607 6418
rect 8541 6378 8607 6414
rect 8998 6378 9009 6424
rect 9055 6378 9066 6424
rect 9222 6378 9233 6424
rect 9279 6378 9290 6424
rect 9482 6378 9493 6424
rect 9539 6378 9550 6424
rect 9717 6378 9763 6395
rect 8998 6332 9066 6378
rect 9482 6332 9550 6378
rect 10114 6353 10125 6399
rect 10171 6353 10182 6399
rect 10114 6332 10182 6353
rect 10498 6351 10509 6498
rect 10555 6351 10566 6498
rect 10498 6332 10566 6351
rect 1344 6298 10800 6332
rect 1344 6246 3538 6298
rect 3798 6246 5862 6298
rect 6122 6246 8186 6298
rect 8446 6246 10510 6298
rect 10770 6246 10800 6298
rect 1344 6212 10800 6246
rect 1418 6193 1486 6212
rect 1418 6046 1429 6193
rect 1475 6046 1486 6193
rect 1418 6034 1486 6046
rect 1729 6126 1775 6212
rect 1729 6040 1775 6080
rect 1933 6126 1999 6166
rect 1933 6080 1953 6126
rect 1822 6018 1887 6032
rect 1874 5989 1887 6018
rect 1418 5875 1486 5888
rect 1418 5829 1429 5875
rect 1475 5829 1486 5875
rect 1822 5849 1837 5966
rect 1883 5849 1887 5989
rect 1822 5832 1887 5849
rect 1933 6018 1999 6080
rect 2401 6126 2447 6212
rect 2401 6040 2447 6080
rect 2605 6126 2671 6166
rect 2605 6080 2625 6126
rect 1933 5966 1934 6018
rect 1986 5966 1999 6018
rect 1418 5747 1486 5829
rect 1418 5701 1429 5747
rect 1475 5701 1486 5747
rect 1418 5619 1486 5701
rect 1418 5573 1429 5619
rect 1475 5573 1486 5619
rect 1418 5548 1486 5573
rect 1749 5747 1795 5766
rect 1749 5548 1795 5607
rect 1933 5747 1999 5966
rect 2494 6018 2559 6032
rect 2546 5989 2559 6018
rect 2494 5849 2509 5966
rect 2555 5849 2559 5989
rect 2494 5832 2559 5849
rect 2605 6018 2671 6080
rect 3073 6126 3119 6212
rect 3073 6040 3119 6080
rect 3277 6126 3343 6166
rect 3277 6080 3297 6126
rect 2605 5966 2606 6018
rect 2658 5966 2671 6018
rect 1933 5607 1953 5747
rect 1933 5594 1999 5607
rect 2421 5747 2467 5766
rect 2421 5548 2467 5607
rect 2605 5747 2671 5966
rect 3166 6018 3231 6032
rect 3218 5989 3231 6018
rect 3166 5849 3181 5966
rect 3227 5849 3231 5989
rect 3166 5832 3231 5849
rect 2605 5607 2625 5747
rect 2605 5594 2671 5607
rect 3093 5747 3139 5766
rect 3093 5548 3139 5607
rect 3277 5747 3343 6080
rect 3745 6126 3791 6212
rect 3745 6040 3791 6080
rect 3949 6126 4015 6166
rect 3949 6080 3969 6126
rect 3838 6018 3903 6032
rect 3890 5989 3903 6018
rect 3838 5849 3853 5966
rect 3899 5849 3903 5989
rect 3838 5832 3903 5849
rect 3277 5682 3297 5747
rect 3277 5630 3278 5682
rect 3277 5607 3297 5630
rect 3277 5594 3343 5607
rect 3765 5747 3811 5766
rect 3765 5548 3811 5607
rect 3949 5747 4015 6080
rect 4417 6126 4463 6212
rect 4417 6040 4463 6080
rect 4621 6126 4687 6166
rect 4621 6080 4641 6126
rect 4510 5989 4575 6032
rect 4510 5906 4525 5989
rect 4510 5849 4525 5854
rect 4571 5849 4575 5989
rect 4510 5832 4575 5849
rect 3949 5682 3969 5747
rect 3949 5630 3950 5682
rect 3949 5607 3969 5630
rect 3949 5594 4015 5607
rect 4437 5747 4483 5766
rect 4437 5548 4483 5607
rect 4621 5747 4687 6080
rect 5089 6126 5135 6212
rect 5089 6040 5135 6080
rect 5293 6126 5359 6166
rect 5293 6080 5313 6126
rect 5182 5989 5247 6032
rect 5182 5906 5197 5989
rect 5182 5849 5197 5854
rect 5243 5849 5247 5989
rect 5182 5832 5247 5849
rect 4621 5682 4641 5747
rect 4621 5630 4622 5682
rect 4621 5607 4641 5630
rect 4621 5594 4687 5607
rect 5109 5747 5155 5766
rect 5109 5548 5155 5607
rect 5293 5747 5359 6080
rect 5761 6126 5807 6212
rect 5761 6040 5807 6080
rect 5965 6126 6031 6166
rect 5965 6080 5985 6126
rect 5854 6018 5919 6032
rect 5906 5989 5919 6018
rect 5854 5849 5869 5966
rect 5915 5849 5919 5989
rect 5854 5832 5919 5849
rect 5293 5682 5313 5747
rect 5293 5630 5294 5682
rect 5293 5607 5313 5630
rect 5293 5594 5359 5607
rect 5781 5747 5827 5766
rect 5781 5548 5827 5607
rect 5965 5747 6031 6080
rect 6433 6126 6479 6212
rect 6433 6040 6479 6080
rect 6637 6126 6703 6166
rect 6637 6080 6657 6126
rect 6526 6018 6591 6032
rect 6578 5989 6591 6018
rect 6526 5849 6541 5966
rect 6587 5849 6591 5989
rect 6526 5832 6591 5849
rect 6637 6018 6703 6080
rect 6881 6126 6927 6212
rect 6881 6053 6927 6080
rect 7185 6126 7231 6166
rect 6637 5966 6638 6018
rect 6690 5966 6703 6018
rect 5965 5682 5985 5747
rect 5965 5630 5966 5682
rect 5965 5607 5985 5630
rect 5965 5594 6031 5607
rect 6453 5747 6499 5766
rect 6453 5548 6499 5607
rect 6637 5747 6703 5966
rect 6637 5607 6657 5747
rect 6637 5594 6703 5607
rect 6881 5961 6984 6007
rect 7124 5961 7136 6007
rect 6881 5755 6927 5961
rect 7185 5880 7231 6080
rect 7665 6126 7711 6212
rect 7665 6040 7711 6080
rect 7869 6126 7935 6166
rect 7869 6080 7889 6126
rect 6978 5834 6992 5880
rect 7132 5834 7231 5880
rect 7758 6018 7823 6032
rect 7810 5989 7823 6018
rect 7758 5849 7773 5966
rect 7819 5849 7823 5989
rect 7758 5832 7823 5849
rect 6881 5594 6927 5615
rect 7185 5755 7231 5774
rect 7185 5548 7231 5615
rect 7685 5747 7731 5766
rect 7685 5548 7731 5607
rect 7869 5747 7935 6080
rect 8337 6126 8383 6212
rect 8337 6040 8383 6080
rect 8541 6126 8607 6166
rect 8541 6080 8561 6126
rect 8430 6018 8495 6032
rect 8482 5989 8495 6018
rect 8430 5849 8445 5966
rect 8491 5849 8495 5989
rect 8430 5832 8495 5849
rect 7869 5682 7889 5747
rect 7869 5630 7870 5682
rect 7869 5607 7889 5630
rect 7869 5594 7935 5607
rect 8357 5747 8403 5766
rect 8357 5548 8403 5607
rect 8541 5747 8607 6080
rect 8785 6126 8831 6212
rect 9374 6193 9442 6212
rect 8785 6053 8831 6080
rect 9089 6126 9135 6166
rect 8541 5682 8561 5747
rect 8541 5630 8542 5682
rect 8541 5607 8561 5630
rect 8541 5594 8607 5607
rect 8785 5961 8888 6007
rect 9028 5961 9040 6007
rect 8785 5755 8831 5961
rect 9089 5880 9135 6080
rect 9374 6046 9385 6193
rect 9431 6046 9442 6193
rect 9374 6035 9442 6046
rect 9985 6130 10051 6166
rect 9985 6126 9998 6130
rect 9985 6078 9998 6080
rect 10050 6078 10051 6130
rect 8882 5834 8896 5880
rect 9036 5834 9135 5880
rect 9374 5875 9442 5886
rect 9374 5829 9385 5875
rect 9431 5829 9442 5875
rect 8785 5594 8831 5615
rect 9089 5755 9135 5774
rect 9089 5548 9135 5615
rect 9374 5747 9442 5829
rect 9374 5701 9385 5747
rect 9431 5701 9442 5747
rect 9374 5619 9442 5701
rect 9374 5573 9385 5619
rect 9431 5573 9442 5619
rect 9985 5747 10051 6078
rect 10209 6126 10255 6212
rect 10209 6040 10255 6080
rect 10498 6193 10566 6212
rect 10498 6046 10509 6193
rect 10555 6046 10566 6193
rect 10498 6034 10566 6046
rect 10097 5989 10162 6032
rect 10097 5849 10101 5989
rect 10147 5906 10162 5989
rect 10147 5849 10162 5854
rect 10097 5832 10162 5849
rect 10498 5875 10566 5888
rect 10498 5829 10509 5875
rect 10555 5829 10566 5875
rect 10031 5607 10051 5747
rect 9985 5594 10051 5607
rect 10189 5747 10235 5766
rect 9374 5548 9442 5573
rect 10189 5548 10235 5607
rect 10498 5747 10566 5829
rect 10498 5701 10509 5747
rect 10555 5701 10566 5747
rect 10498 5619 10566 5701
rect 10498 5573 10509 5619
rect 10555 5573 10566 5619
rect 10498 5548 10566 5573
rect 1344 5514 10640 5548
rect 1344 5462 2376 5514
rect 2636 5462 4700 5514
rect 4960 5462 7024 5514
rect 7284 5462 9348 5514
rect 9608 5462 10640 5514
rect 1344 5428 10640 5462
rect 1418 5403 1486 5428
rect 1418 5357 1429 5403
rect 1475 5357 1486 5403
rect 1418 5275 1486 5357
rect 1418 5229 1429 5275
rect 1475 5229 1486 5275
rect 1418 5147 1486 5229
rect 1418 5101 1429 5147
rect 1475 5101 1486 5147
rect 1418 5088 1486 5101
rect 1617 5361 1663 5382
rect 1617 5015 1663 5221
rect 1921 5361 1967 5428
rect 1921 5202 1967 5221
rect 2085 5369 2131 5428
rect 2085 5210 2131 5229
rect 2269 5369 2335 5382
rect 2269 5346 2289 5369
rect 2269 5294 2270 5346
rect 2269 5229 2289 5294
rect 1714 5096 1728 5142
rect 1868 5096 1967 5142
rect 1617 4969 1720 5015
rect 1860 4969 1872 5015
rect 1418 4930 1486 4942
rect 1418 4783 1429 4930
rect 1475 4783 1486 4930
rect 1418 4764 1486 4783
rect 1617 4896 1663 4923
rect 1617 4764 1663 4850
rect 1921 4896 1967 5096
rect 2158 5127 2223 5144
rect 2158 5122 2173 5127
rect 2158 4987 2173 5070
rect 2219 4987 2223 5127
rect 2158 4944 2223 4987
rect 1921 4810 1967 4850
rect 2065 4896 2111 4936
rect 2065 4764 2111 4850
rect 2269 4896 2335 5229
rect 2757 5369 2803 5428
rect 2757 5210 2803 5229
rect 2941 5369 3007 5382
rect 2941 5346 2961 5369
rect 2941 5294 2942 5346
rect 2941 5229 2961 5294
rect 2830 5127 2895 5144
rect 2830 5122 2845 5127
rect 2830 4987 2845 5070
rect 2891 4987 2895 5127
rect 2830 4944 2895 4987
rect 2269 4850 2289 4896
rect 2269 4810 2335 4850
rect 2737 4896 2783 4936
rect 2737 4764 2783 4850
rect 2941 4896 3007 5229
rect 3429 5369 3475 5428
rect 3429 5210 3475 5229
rect 3613 5369 3679 5382
rect 3613 5229 3633 5369
rect 3502 5127 3567 5144
rect 3502 5122 3517 5127
rect 3502 4987 3517 5070
rect 3563 4987 3567 5127
rect 3502 4944 3567 4987
rect 3613 5122 3679 5229
rect 4101 5369 4147 5428
rect 4101 5210 4147 5229
rect 4285 5369 4351 5382
rect 4285 5346 4305 5369
rect 4285 5294 4286 5346
rect 4285 5229 4305 5294
rect 3613 5070 3614 5122
rect 3666 5070 3679 5122
rect 2941 4850 2961 4896
rect 2941 4810 3007 4850
rect 3409 4896 3455 4936
rect 3409 4764 3455 4850
rect 3613 4896 3679 5070
rect 4174 5127 4239 5144
rect 4174 5010 4189 5127
rect 4235 4987 4239 5127
rect 4226 4958 4239 4987
rect 4174 4944 4239 4958
rect 3613 4850 3633 4896
rect 3613 4810 3679 4850
rect 4081 4896 4127 4936
rect 4081 4764 4127 4850
rect 4285 4896 4351 5229
rect 4773 5369 4819 5428
rect 5342 5403 5410 5428
rect 4773 5210 4819 5229
rect 4957 5369 5023 5382
rect 4957 5229 4977 5369
rect 4846 5127 4911 5144
rect 4846 5010 4861 5127
rect 4907 4987 4911 5127
rect 4898 4958 4911 4987
rect 4846 4944 4911 4958
rect 4957 5010 5023 5229
rect 5342 5357 5353 5403
rect 5399 5357 5410 5403
rect 5342 5275 5410 5357
rect 5342 5229 5353 5275
rect 5399 5229 5410 5275
rect 5342 5147 5410 5229
rect 5669 5369 5715 5428
rect 5669 5210 5715 5229
rect 5853 5369 5919 5382
rect 5853 5229 5873 5369
rect 5342 5101 5353 5147
rect 5399 5101 5410 5147
rect 5342 5090 5410 5101
rect 5742 5127 5807 5144
rect 4957 4958 4958 5010
rect 5010 4958 5023 5010
rect 4285 4850 4305 4896
rect 4285 4810 4351 4850
rect 4753 4896 4799 4936
rect 4753 4764 4799 4850
rect 4957 4896 5023 4958
rect 5742 5010 5757 5127
rect 5803 4987 5807 5127
rect 5794 4958 5807 4987
rect 5742 4944 5807 4958
rect 5853 5010 5919 5229
rect 5853 4958 5854 5010
rect 5906 4958 5919 5010
rect 6097 5361 6143 5382
rect 6097 5015 6143 5221
rect 6401 5361 6447 5428
rect 6401 5202 6447 5221
rect 6901 5369 6947 5428
rect 6901 5210 6947 5229
rect 7085 5369 7151 5382
rect 7085 5346 7105 5369
rect 7085 5294 7086 5346
rect 7085 5229 7105 5294
rect 6194 5096 6208 5142
rect 6348 5096 6447 5142
rect 6097 4969 6200 5015
rect 6340 4969 6352 5015
rect 4957 4850 4977 4896
rect 4957 4810 5023 4850
rect 5342 4930 5410 4941
rect 5342 4783 5353 4930
rect 5399 4783 5410 4930
rect 5342 4764 5410 4783
rect 5649 4896 5695 4936
rect 5649 4764 5695 4850
rect 5853 4896 5919 4958
rect 5853 4850 5873 4896
rect 5853 4810 5919 4850
rect 6097 4896 6143 4923
rect 6097 4764 6143 4850
rect 6401 4896 6447 5096
rect 6974 5127 7039 5144
rect 6974 5122 6989 5127
rect 6974 4987 6989 5070
rect 7035 4987 7039 5127
rect 6974 4944 7039 4987
rect 6401 4810 6447 4850
rect 6881 4896 6927 4936
rect 6881 4764 6927 4850
rect 7085 4896 7151 5229
rect 7573 5369 7619 5428
rect 7573 5210 7619 5229
rect 7757 5369 7823 5382
rect 7757 5346 7777 5369
rect 7757 5294 7758 5346
rect 7757 5229 7777 5294
rect 7646 5127 7711 5144
rect 7646 5010 7661 5127
rect 7707 4987 7711 5127
rect 7698 4958 7711 4987
rect 7646 4944 7711 4958
rect 7085 4850 7105 4896
rect 7085 4810 7151 4850
rect 7553 4896 7599 4936
rect 7553 4764 7599 4850
rect 7757 4896 7823 5229
rect 8245 5369 8291 5428
rect 8245 5210 8291 5229
rect 8429 5369 8495 5382
rect 8429 5229 8449 5369
rect 8318 5127 8383 5144
rect 8318 5122 8333 5127
rect 8318 4987 8333 5070
rect 8379 4987 8383 5127
rect 8318 4944 8383 4987
rect 8429 5122 8495 5229
rect 8429 5070 8430 5122
rect 8482 5070 8495 5122
rect 7757 4850 7777 4896
rect 7757 4810 7823 4850
rect 8225 4896 8271 4936
rect 8225 4764 8271 4850
rect 8429 4896 8495 5070
rect 8673 5361 8719 5382
rect 8673 5015 8719 5221
rect 8977 5361 9023 5428
rect 8977 5202 9023 5221
rect 9253 5369 9299 5428
rect 9253 5210 9299 5229
rect 9437 5369 9503 5382
rect 9437 5229 9457 5369
rect 8770 5096 8784 5142
rect 8924 5096 9023 5142
rect 8673 4969 8776 5015
rect 8916 4969 8928 5015
rect 8429 4850 8449 4896
rect 8429 4810 8495 4850
rect 8673 4896 8719 4923
rect 8673 4764 8719 4850
rect 8977 4896 9023 5096
rect 9326 5127 9391 5144
rect 9326 5010 9341 5127
rect 9387 4987 9391 5127
rect 9378 4958 9391 4987
rect 9326 4944 9391 4958
rect 8977 4810 9023 4850
rect 9233 4896 9279 4936
rect 9233 4764 9279 4850
rect 9437 4898 9503 5229
rect 9437 4846 9438 4898
rect 9490 4896 9503 4898
rect 9490 4846 9503 4850
rect 9437 4810 9503 4846
rect 9985 5369 10051 5382
rect 10031 5346 10051 5369
rect 10050 5294 10051 5346
rect 10031 5229 10051 5294
rect 9985 4896 10051 5229
rect 10189 5369 10235 5428
rect 10189 5210 10235 5229
rect 10498 5403 10566 5428
rect 10498 5357 10509 5403
rect 10555 5357 10566 5403
rect 10498 5275 10566 5357
rect 10498 5229 10509 5275
rect 10555 5229 10566 5275
rect 10498 5147 10566 5229
rect 10097 5127 10162 5144
rect 10097 4987 10101 5127
rect 10147 5122 10162 5127
rect 10498 5101 10509 5147
rect 10555 5101 10566 5147
rect 10498 5088 10566 5101
rect 10147 4987 10162 5070
rect 10097 4944 10162 4987
rect 10031 4850 10051 4896
rect 9985 4810 10051 4850
rect 10209 4896 10255 4936
rect 10209 4764 10255 4850
rect 10498 4930 10566 4942
rect 10498 4783 10509 4930
rect 10555 4783 10566 4930
rect 10498 4764 10566 4783
rect 1344 4730 10800 4764
rect 1344 4678 3538 4730
rect 3798 4678 5862 4730
rect 6122 4678 8186 4730
rect 8446 4678 10510 4730
rect 10770 4678 10800 4730
rect 1344 4644 10800 4678
rect 1418 4625 1486 4644
rect 1418 4478 1429 4625
rect 1475 4478 1486 4625
rect 1418 4466 1486 4478
rect 1841 4558 1887 4644
rect 1841 4472 1887 4512
rect 2045 4562 2111 4598
rect 2045 4510 2046 4562
rect 2098 4558 2111 4562
rect 2098 4510 2111 4512
rect 1934 4450 1999 4464
rect 1986 4421 1999 4450
rect 1418 4307 1486 4320
rect 1418 4261 1429 4307
rect 1475 4261 1486 4307
rect 1934 4281 1949 4398
rect 1995 4281 1999 4421
rect 1934 4264 1999 4281
rect 1418 4179 1486 4261
rect 1418 4133 1429 4179
rect 1475 4133 1486 4179
rect 1418 4051 1486 4133
rect 1418 4005 1429 4051
rect 1475 4005 1486 4051
rect 1418 3980 1486 4005
rect 1861 4179 1907 4198
rect 1861 3980 1907 4039
rect 2045 4179 2111 4510
rect 2513 4558 2559 4644
rect 2513 4472 2559 4512
rect 2717 4558 2783 4598
rect 2717 4512 2737 4558
rect 2606 4450 2671 4464
rect 2658 4421 2671 4450
rect 2606 4281 2621 4398
rect 2667 4281 2671 4421
rect 2606 4264 2671 4281
rect 2045 4039 2065 4179
rect 2045 4026 2111 4039
rect 2533 4179 2579 4198
rect 2533 3980 2579 4039
rect 2717 4179 2783 4512
rect 3185 4558 3231 4644
rect 3185 4472 3231 4512
rect 3389 4562 3455 4598
rect 3389 4510 3390 4562
rect 3442 4558 3455 4562
rect 3442 4510 3455 4512
rect 3278 4421 3343 4464
rect 3278 4338 3293 4421
rect 3278 4281 3293 4286
rect 3339 4281 3343 4421
rect 3278 4264 3343 4281
rect 2717 4114 2737 4179
rect 2717 4062 2718 4114
rect 2717 4039 2737 4062
rect 2717 4026 2783 4039
rect 3205 4179 3251 4198
rect 3205 3980 3251 4039
rect 3389 4179 3455 4510
rect 3857 4558 3903 4644
rect 3857 4472 3903 4512
rect 4061 4558 4127 4598
rect 4061 4512 4081 4558
rect 3950 4450 4015 4464
rect 4002 4421 4015 4450
rect 3950 4281 3965 4398
rect 4011 4281 4015 4421
rect 3950 4264 4015 4281
rect 3389 4039 3409 4179
rect 3389 4026 3455 4039
rect 3877 4179 3923 4198
rect 3877 3980 3923 4039
rect 4061 4179 4127 4512
rect 4529 4558 4575 4644
rect 4529 4472 4575 4512
rect 4733 4558 4799 4598
rect 4733 4512 4753 4558
rect 4622 4421 4687 4464
rect 4622 4338 4637 4421
rect 4622 4281 4637 4286
rect 4683 4281 4687 4421
rect 4622 4264 4687 4281
rect 4061 4114 4081 4179
rect 4061 4062 4062 4114
rect 4061 4039 4081 4062
rect 4061 4026 4127 4039
rect 4549 4179 4595 4198
rect 4549 3980 4595 4039
rect 4733 4179 4799 4512
rect 4977 4558 5023 4644
rect 4977 4485 5023 4512
rect 5281 4558 5327 4598
rect 4733 4114 4753 4179
rect 4733 4062 4734 4114
rect 4733 4039 4753 4062
rect 4733 4026 4799 4039
rect 4977 4393 5080 4439
rect 5220 4393 5232 4439
rect 4977 4187 5023 4393
rect 5281 4312 5327 4512
rect 5649 4558 5695 4644
rect 5649 4472 5695 4512
rect 5853 4558 5919 4598
rect 5853 4512 5873 4558
rect 5074 4266 5088 4312
rect 5228 4266 5327 4312
rect 5742 4421 5807 4464
rect 5742 4338 5757 4421
rect 5742 4281 5757 4286
rect 5803 4281 5807 4421
rect 5742 4264 5807 4281
rect 4977 4026 5023 4047
rect 5281 4187 5327 4206
rect 5281 3980 5327 4047
rect 5669 4179 5715 4198
rect 5669 3980 5715 4039
rect 5853 4179 5919 4512
rect 6321 4558 6367 4644
rect 6321 4472 6367 4512
rect 6525 4562 6591 4598
rect 6525 4510 6526 4562
rect 6578 4558 6591 4562
rect 6578 4510 6591 4512
rect 6414 4450 6479 4464
rect 6466 4421 6479 4450
rect 6414 4281 6429 4398
rect 6475 4281 6479 4421
rect 6414 4264 6479 4281
rect 5853 4114 5873 4179
rect 5853 4062 5854 4114
rect 5853 4039 5873 4062
rect 5853 4026 5919 4039
rect 6341 4179 6387 4198
rect 6341 3980 6387 4039
rect 6525 4179 6591 4510
rect 6993 4558 7039 4644
rect 6993 4472 7039 4512
rect 7197 4562 7263 4598
rect 7197 4510 7198 4562
rect 7250 4558 7263 4562
rect 7250 4510 7263 4512
rect 7086 4450 7151 4464
rect 7138 4421 7151 4450
rect 7086 4281 7101 4398
rect 7147 4281 7151 4421
rect 7086 4264 7151 4281
rect 6525 4039 6545 4179
rect 6525 4026 6591 4039
rect 7013 4179 7059 4198
rect 7013 3980 7059 4039
rect 7197 4179 7263 4510
rect 7665 4558 7711 4644
rect 7665 4472 7711 4512
rect 7869 4558 7935 4598
rect 7869 4512 7889 4558
rect 7758 4450 7823 4464
rect 7810 4421 7823 4450
rect 7758 4281 7773 4398
rect 7819 4281 7823 4421
rect 7758 4264 7823 4281
rect 7197 4039 7217 4179
rect 7197 4026 7263 4039
rect 7685 4179 7731 4198
rect 7685 3980 7731 4039
rect 7869 4179 7935 4512
rect 8337 4558 8383 4644
rect 8337 4472 8383 4512
rect 8541 4558 8607 4598
rect 8541 4512 8561 4558
rect 8430 4421 8495 4464
rect 8430 4338 8445 4421
rect 8430 4281 8445 4286
rect 8491 4281 8495 4421
rect 8430 4264 8495 4281
rect 7869 4114 7889 4179
rect 7869 4062 7870 4114
rect 7869 4039 7889 4062
rect 7869 4026 7935 4039
rect 8357 4179 8403 4198
rect 8357 3980 8403 4039
rect 8541 4179 8607 4512
rect 8785 4558 8831 4644
rect 9374 4625 9442 4644
rect 8785 4485 8831 4512
rect 9089 4558 9135 4598
rect 8541 4114 8561 4179
rect 8541 4062 8542 4114
rect 8541 4039 8561 4062
rect 8541 4026 8607 4039
rect 8785 4393 8888 4439
rect 9028 4393 9040 4439
rect 8785 4187 8831 4393
rect 9089 4312 9135 4512
rect 9374 4478 9385 4625
rect 9431 4478 9442 4625
rect 9374 4467 9442 4478
rect 9905 4558 9951 4644
rect 10498 4625 10566 4644
rect 9905 4472 9951 4512
rect 10109 4558 10175 4598
rect 10109 4512 10129 4558
rect 9998 4421 10063 4464
rect 9998 4338 10013 4421
rect 8882 4266 8896 4312
rect 9036 4266 9135 4312
rect 9374 4307 9442 4318
rect 9374 4261 9385 4307
rect 9431 4261 9442 4307
rect 9998 4281 10013 4286
rect 10059 4281 10063 4421
rect 9998 4264 10063 4281
rect 8785 4026 8831 4047
rect 9089 4187 9135 4206
rect 9089 3980 9135 4047
rect 9374 4179 9442 4261
rect 9374 4133 9385 4179
rect 9431 4133 9442 4179
rect 9374 4051 9442 4133
rect 9374 4005 9385 4051
rect 9431 4005 9442 4051
rect 9374 3980 9442 4005
rect 9925 4179 9971 4198
rect 9925 3980 9971 4039
rect 10109 4179 10175 4512
rect 10498 4478 10509 4625
rect 10555 4478 10566 4625
rect 10498 4466 10566 4478
rect 10109 4114 10129 4179
rect 10109 4062 10110 4114
rect 10109 4039 10129 4062
rect 10109 4026 10175 4039
rect 10498 4307 10566 4320
rect 10498 4261 10509 4307
rect 10555 4261 10566 4307
rect 10498 4179 10566 4261
rect 10498 4133 10509 4179
rect 10555 4133 10566 4179
rect 10498 4051 10566 4133
rect 10498 4005 10509 4051
rect 10555 4005 10566 4051
rect 10498 3980 10566 4005
rect 1344 3946 10640 3980
rect 1344 3894 2376 3946
rect 2636 3894 4700 3946
rect 4960 3894 7024 3946
rect 7284 3894 9348 3946
rect 9608 3894 10640 3946
rect 1344 3860 10640 3894
rect 1418 3835 1486 3860
rect 1418 3789 1429 3835
rect 1475 3789 1486 3835
rect 1418 3707 1486 3789
rect 1418 3661 1429 3707
rect 1475 3661 1486 3707
rect 1418 3579 1486 3661
rect 1418 3533 1429 3579
rect 1475 3533 1486 3579
rect 1418 3520 1486 3533
rect 1921 3801 1987 3814
rect 1967 3661 1987 3801
rect 1921 3442 1987 3661
rect 2125 3801 2171 3860
rect 2125 3642 2171 3661
rect 2533 3801 2579 3860
rect 2533 3642 2579 3661
rect 2717 3801 2783 3814
rect 2717 3661 2737 3801
rect 1921 3390 1934 3442
rect 1986 3390 1987 3442
rect 1418 3362 1486 3374
rect 1418 3215 1429 3362
rect 1475 3215 1486 3362
rect 1921 3328 1987 3390
rect 2033 3559 2098 3576
rect 2033 3419 2037 3559
rect 2083 3554 2098 3559
rect 2083 3419 2098 3502
rect 2033 3376 2098 3419
rect 2606 3559 2671 3576
rect 2606 3442 2621 3559
rect 2667 3419 2671 3559
rect 2658 3390 2671 3419
rect 2606 3376 2671 3390
rect 2717 3554 2783 3661
rect 3205 3801 3251 3860
rect 3205 3642 3251 3661
rect 3389 3801 3455 3814
rect 3389 3661 3409 3801
rect 2717 3502 2718 3554
rect 2770 3502 2783 3554
rect 1967 3282 1987 3328
rect 1921 3242 1987 3282
rect 2145 3328 2191 3368
rect 1418 3196 1486 3215
rect 2145 3196 2191 3282
rect 2513 3328 2559 3368
rect 2513 3196 2559 3282
rect 2717 3328 2783 3502
rect 3278 3559 3343 3576
rect 3278 3442 3293 3559
rect 3339 3419 3343 3559
rect 3330 3390 3343 3419
rect 3278 3376 3343 3390
rect 3389 3442 3455 3661
rect 3877 3801 3923 3860
rect 3877 3642 3923 3661
rect 4061 3801 4127 3814
rect 4061 3661 4081 3801
rect 3389 3390 3390 3442
rect 3442 3390 3455 3442
rect 2717 3282 2737 3328
rect 2717 3242 2783 3282
rect 3185 3328 3231 3368
rect 3185 3196 3231 3282
rect 3389 3328 3455 3390
rect 3950 3559 4015 3576
rect 3950 3442 3965 3559
rect 4011 3419 4015 3559
rect 4002 3390 4015 3419
rect 3950 3376 4015 3390
rect 4061 3442 4127 3661
rect 4549 3801 4595 3860
rect 5342 3835 5410 3860
rect 4549 3642 4595 3661
rect 4733 3801 4799 3814
rect 4733 3661 4753 3801
rect 4061 3390 4062 3442
rect 4114 3390 4127 3442
rect 3389 3282 3409 3328
rect 3389 3242 3455 3282
rect 3857 3328 3903 3368
rect 3857 3196 3903 3282
rect 4061 3328 4127 3390
rect 4622 3559 4687 3576
rect 4622 3442 4637 3559
rect 4683 3419 4687 3559
rect 4674 3390 4687 3419
rect 4622 3376 4687 3390
rect 4733 3442 4799 3661
rect 5342 3789 5353 3835
rect 5399 3789 5410 3835
rect 5342 3707 5410 3789
rect 5342 3661 5353 3707
rect 5399 3661 5410 3707
rect 5342 3579 5410 3661
rect 5669 3801 5715 3860
rect 5669 3642 5715 3661
rect 5853 3801 5919 3814
rect 5853 3778 5873 3801
rect 5853 3726 5854 3778
rect 5853 3661 5873 3726
rect 5342 3533 5353 3579
rect 5399 3533 5410 3579
rect 5342 3522 5410 3533
rect 5742 3559 5807 3576
rect 4733 3390 4734 3442
rect 4786 3390 4799 3442
rect 4061 3282 4081 3328
rect 4061 3242 4127 3282
rect 4529 3328 4575 3368
rect 4529 3196 4575 3282
rect 4733 3328 4799 3390
rect 5742 3442 5757 3559
rect 5803 3419 5807 3559
rect 5794 3390 5807 3419
rect 5742 3376 5807 3390
rect 4733 3282 4753 3328
rect 4733 3242 4799 3282
rect 5342 3362 5410 3373
rect 5342 3215 5353 3362
rect 5399 3215 5410 3362
rect 5342 3196 5410 3215
rect 5649 3328 5695 3368
rect 5649 3196 5695 3282
rect 5853 3328 5919 3661
rect 6097 3793 6143 3814
rect 6097 3447 6143 3653
rect 6401 3793 6447 3860
rect 6401 3634 6447 3653
rect 6565 3801 6611 3860
rect 6565 3642 6611 3661
rect 6749 3801 6815 3814
rect 6749 3778 6769 3801
rect 6749 3726 6750 3778
rect 6749 3661 6769 3726
rect 6194 3528 6208 3574
rect 6348 3528 6447 3574
rect 6097 3401 6200 3447
rect 6340 3401 6352 3447
rect 5853 3282 5873 3328
rect 5853 3242 5919 3282
rect 6097 3328 6143 3355
rect 6097 3196 6143 3282
rect 6401 3328 6447 3528
rect 6638 3559 6703 3576
rect 6638 3554 6653 3559
rect 6638 3419 6653 3502
rect 6699 3419 6703 3559
rect 6638 3376 6703 3419
rect 6401 3242 6447 3282
rect 6545 3328 6591 3368
rect 6545 3196 6591 3282
rect 6749 3328 6815 3661
rect 7237 3801 7283 3860
rect 7237 3642 7283 3661
rect 7421 3801 7487 3814
rect 7421 3778 7441 3801
rect 7421 3726 7422 3778
rect 7421 3661 7441 3726
rect 7310 3559 7375 3576
rect 7310 3554 7325 3559
rect 7310 3419 7325 3502
rect 7371 3419 7375 3559
rect 7310 3376 7375 3419
rect 6749 3282 6769 3328
rect 6749 3242 6815 3282
rect 7217 3328 7263 3368
rect 7217 3196 7263 3282
rect 7421 3328 7487 3661
rect 7421 3282 7441 3328
rect 7421 3242 7487 3282
rect 7969 3801 8035 3814
rect 8015 3778 8035 3801
rect 8034 3726 8035 3778
rect 8015 3661 8035 3726
rect 7969 3328 8035 3661
rect 8173 3801 8219 3860
rect 8173 3642 8219 3661
rect 8581 3801 8627 3860
rect 9262 3835 9330 3860
rect 8581 3642 8627 3661
rect 8765 3801 8831 3814
rect 8765 3666 8785 3801
rect 8765 3614 8766 3666
rect 8818 3614 8831 3661
rect 8081 3559 8146 3576
rect 8081 3419 8085 3559
rect 8131 3554 8146 3559
rect 8131 3419 8146 3502
rect 8081 3376 8146 3419
rect 8654 3559 8719 3576
rect 8654 3554 8669 3559
rect 8654 3419 8669 3502
rect 8715 3419 8719 3559
rect 8654 3376 8719 3419
rect 8015 3282 8035 3328
rect 7969 3242 8035 3282
rect 8193 3328 8239 3368
rect 8193 3196 8239 3282
rect 8561 3328 8607 3368
rect 8561 3196 8607 3282
rect 8765 3328 8831 3614
rect 9262 3789 9273 3835
rect 9319 3789 9330 3835
rect 9262 3707 9330 3789
rect 9262 3661 9273 3707
rect 9319 3661 9330 3707
rect 9262 3579 9330 3661
rect 9262 3533 9273 3579
rect 9319 3533 9330 3579
rect 9262 3522 9330 3533
rect 9457 3793 9503 3814
rect 9457 3447 9503 3653
rect 9761 3793 9807 3860
rect 9761 3634 9807 3653
rect 9925 3801 9971 3860
rect 10498 3835 10566 3860
rect 9925 3642 9971 3661
rect 10109 3801 10175 3814
rect 10109 3666 10129 3801
rect 10109 3614 10110 3666
rect 10162 3614 10175 3661
rect 9554 3528 9568 3574
rect 9708 3528 9807 3574
rect 9457 3401 9560 3447
rect 9700 3401 9712 3447
rect 8765 3282 8785 3328
rect 8765 3242 8831 3282
rect 9262 3362 9330 3373
rect 9262 3215 9273 3362
rect 9319 3215 9330 3362
rect 9262 3196 9330 3215
rect 9457 3328 9503 3355
rect 9457 3196 9503 3282
rect 9761 3328 9807 3528
rect 9998 3559 10063 3576
rect 9998 3442 10013 3559
rect 10059 3419 10063 3559
rect 10050 3390 10063 3419
rect 9998 3376 10063 3390
rect 9761 3242 9807 3282
rect 9905 3328 9951 3368
rect 9905 3196 9951 3282
rect 10109 3328 10175 3614
rect 10498 3789 10509 3835
rect 10555 3789 10566 3835
rect 10498 3707 10566 3789
rect 10498 3661 10509 3707
rect 10555 3661 10566 3707
rect 10498 3579 10566 3661
rect 10498 3533 10509 3579
rect 10555 3533 10566 3579
rect 10498 3520 10566 3533
rect 10109 3282 10129 3328
rect 10109 3242 10175 3282
rect 10498 3362 10566 3374
rect 10498 3215 10509 3362
rect 10555 3215 10566 3362
rect 10498 3196 10566 3215
rect 1344 3162 10800 3196
rect 1344 3110 3538 3162
rect 3798 3110 5862 3162
rect 6122 3110 8186 3162
rect 8446 3110 10510 3162
rect 10770 3110 10800 3162
rect 1344 3076 10800 3110
<< via1 >>
rect 2376 8598 2636 8650
rect 4700 8598 4960 8650
rect 7024 8598 7284 8650
rect 9348 8598 9608 8650
rect 2158 8123 2173 8146
rect 2173 8123 2210 8146
rect 2158 8094 2210 8123
rect 2830 8123 2845 8146
rect 2845 8123 2882 8146
rect 2830 8094 2882 8123
rect 2270 8032 2322 8034
rect 2270 7986 2289 8032
rect 2289 7986 2322 8032
rect 2270 7982 2322 7986
rect 3502 8123 3517 8146
rect 3517 8123 3554 8146
rect 3502 8094 3554 8123
rect 3614 8094 3666 8146
rect 2942 8032 2994 8034
rect 2942 7986 2961 8032
rect 2961 7986 2994 8032
rect 2942 7982 2994 7986
rect 4174 8123 4189 8146
rect 4189 8123 4226 8146
rect 4174 8094 4226 8123
rect 4846 8123 4861 8146
rect 4861 8123 4898 8146
rect 4846 8094 4898 8123
rect 4286 8032 4338 8034
rect 4286 7986 4305 8032
rect 4305 7986 4338 8032
rect 4286 7982 4338 7986
rect 4958 8032 5010 8034
rect 4958 7986 4977 8032
rect 4977 7986 5010 8032
rect 4958 7982 5010 7986
rect 3538 7814 3798 7866
rect 5862 7814 6122 7866
rect 8186 7814 8446 7866
rect 10510 7814 10770 7866
rect 2158 7422 2173 7474
rect 2173 7422 2210 7474
rect 2830 7422 2845 7474
rect 2845 7422 2882 7474
rect 2942 7422 2994 7474
rect 2270 7198 2289 7250
rect 2289 7198 2322 7250
rect 3502 7422 3517 7474
rect 3517 7422 3554 7474
rect 4174 7422 4189 7474
rect 4189 7422 4226 7474
rect 4286 7422 4338 7474
rect 3614 7198 3633 7250
rect 3633 7198 3666 7250
rect 4846 7422 4861 7474
rect 4861 7422 4898 7474
rect 4958 7422 5010 7474
rect 5630 7422 5667 7474
rect 5667 7422 5682 7474
rect 5518 7198 5551 7250
rect 5551 7198 5570 7250
rect 6302 7422 6339 7474
rect 6339 7422 6354 7474
rect 6190 7198 6223 7250
rect 6223 7198 6242 7250
rect 10110 7422 10147 7474
rect 10147 7422 10162 7474
rect 9998 7198 10031 7250
rect 10031 7198 10050 7250
rect 2376 7030 2636 7082
rect 4700 7030 4960 7082
rect 7024 7030 7284 7082
rect 9348 7030 9608 7082
rect 1934 6555 1949 6578
rect 1949 6555 1986 6578
rect 1934 6526 1986 6555
rect 2606 6555 2621 6578
rect 2621 6555 2658 6578
rect 2606 6526 2658 6555
rect 2046 6464 2098 6466
rect 2046 6418 2065 6464
rect 2065 6418 2098 6464
rect 2046 6414 2098 6418
rect 3278 6555 3293 6578
rect 3293 6555 3330 6578
rect 3278 6526 3330 6555
rect 3390 6526 3442 6578
rect 2718 6464 2770 6466
rect 2718 6418 2737 6464
rect 2737 6418 2770 6464
rect 2718 6414 2770 6418
rect 3950 6555 3965 6578
rect 3965 6555 4002 6578
rect 3950 6526 4002 6555
rect 4622 6555 4637 6578
rect 4637 6555 4674 6578
rect 4622 6526 4674 6555
rect 4062 6464 4114 6466
rect 4062 6418 4081 6464
rect 4081 6418 4114 6464
rect 4062 6414 4114 6418
rect 5742 6555 5757 6578
rect 5757 6555 5794 6578
rect 5742 6526 5794 6555
rect 4734 6464 4786 6466
rect 4734 6418 4753 6464
rect 4753 6418 4786 6464
rect 4734 6414 4786 6418
rect 6414 6555 6429 6578
rect 6429 6555 6466 6578
rect 6414 6526 6466 6555
rect 5854 6464 5906 6466
rect 5854 6418 5873 6464
rect 5873 6418 5906 6464
rect 5854 6414 5906 6418
rect 7086 6555 7101 6578
rect 7101 6555 7138 6578
rect 7086 6526 7138 6555
rect 7198 6526 7250 6578
rect 6526 6464 6578 6466
rect 6526 6418 6545 6464
rect 6545 6418 6578 6464
rect 6526 6414 6578 6418
rect 8430 6555 8445 6578
rect 8445 6555 8482 6578
rect 8430 6526 8482 6555
rect 9774 6750 9826 6802
rect 10110 6750 10162 6802
rect 9662 6638 9714 6690
rect 8542 6464 8594 6466
rect 8542 6418 8561 6464
rect 8561 6418 8594 6464
rect 8542 6414 8594 6418
rect 3538 6246 3798 6298
rect 5862 6246 6122 6298
rect 8186 6246 8446 6298
rect 10510 6246 10770 6298
rect 1822 5989 1874 6018
rect 1822 5966 1837 5989
rect 1837 5966 1874 5989
rect 1934 5966 1986 6018
rect 2494 5989 2546 6018
rect 2494 5966 2509 5989
rect 2509 5966 2546 5989
rect 2606 5966 2658 6018
rect 3166 5989 3218 6018
rect 3166 5966 3181 5989
rect 3181 5966 3218 5989
rect 3838 5989 3890 6018
rect 3838 5966 3853 5989
rect 3853 5966 3890 5989
rect 3278 5630 3297 5682
rect 3297 5630 3330 5682
rect 4510 5854 4525 5906
rect 4525 5854 4562 5906
rect 3950 5630 3969 5682
rect 3969 5630 4002 5682
rect 5182 5854 5197 5906
rect 5197 5854 5234 5906
rect 4622 5630 4641 5682
rect 4641 5630 4674 5682
rect 5854 5989 5906 6018
rect 5854 5966 5869 5989
rect 5869 5966 5906 5989
rect 5294 5630 5313 5682
rect 5313 5630 5346 5682
rect 6526 5989 6578 6018
rect 6526 5966 6541 5989
rect 6541 5966 6578 5989
rect 6638 5966 6690 6018
rect 5966 5630 5985 5682
rect 5985 5630 6018 5682
rect 7758 5989 7810 6018
rect 7758 5966 7773 5989
rect 7773 5966 7810 5989
rect 8430 5989 8482 6018
rect 8430 5966 8445 5989
rect 8445 5966 8482 5989
rect 7870 5630 7889 5682
rect 7889 5630 7922 5682
rect 8542 5630 8561 5682
rect 8561 5630 8594 5682
rect 9998 6126 10050 6130
rect 9998 6080 10031 6126
rect 10031 6080 10050 6126
rect 9998 6078 10050 6080
rect 10110 5854 10147 5906
rect 10147 5854 10162 5906
rect 2376 5462 2636 5514
rect 4700 5462 4960 5514
rect 7024 5462 7284 5514
rect 9348 5462 9608 5514
rect 2270 5294 2289 5346
rect 2289 5294 2322 5346
rect 2158 5070 2173 5122
rect 2173 5070 2210 5122
rect 2942 5294 2961 5346
rect 2961 5294 2994 5346
rect 2830 5070 2845 5122
rect 2845 5070 2882 5122
rect 3502 5070 3517 5122
rect 3517 5070 3554 5122
rect 4286 5294 4305 5346
rect 4305 5294 4338 5346
rect 3614 5070 3666 5122
rect 4174 4987 4189 5010
rect 4189 4987 4226 5010
rect 4174 4958 4226 4987
rect 4846 4987 4861 5010
rect 4861 4987 4898 5010
rect 4846 4958 4898 4987
rect 4958 4958 5010 5010
rect 5742 4987 5757 5010
rect 5757 4987 5794 5010
rect 5742 4958 5794 4987
rect 5854 4958 5906 5010
rect 7086 5294 7105 5346
rect 7105 5294 7138 5346
rect 6974 5070 6989 5122
rect 6989 5070 7026 5122
rect 7758 5294 7777 5346
rect 7777 5294 7810 5346
rect 7646 4987 7661 5010
rect 7661 4987 7698 5010
rect 7646 4958 7698 4987
rect 8318 5070 8333 5122
rect 8333 5070 8370 5122
rect 8430 5070 8482 5122
rect 9326 4987 9341 5010
rect 9341 4987 9378 5010
rect 9326 4958 9378 4987
rect 9438 4896 9490 4898
rect 9438 4850 9457 4896
rect 9457 4850 9490 4896
rect 9438 4846 9490 4850
rect 9998 5294 10031 5346
rect 10031 5294 10050 5346
rect 10110 5070 10147 5122
rect 10147 5070 10162 5122
rect 3538 4678 3798 4730
rect 5862 4678 6122 4730
rect 8186 4678 8446 4730
rect 10510 4678 10770 4730
rect 2046 4558 2098 4562
rect 2046 4512 2065 4558
rect 2065 4512 2098 4558
rect 2046 4510 2098 4512
rect 1934 4421 1986 4450
rect 1934 4398 1949 4421
rect 1949 4398 1986 4421
rect 2606 4421 2658 4450
rect 2606 4398 2621 4421
rect 2621 4398 2658 4421
rect 3390 4558 3442 4562
rect 3390 4512 3409 4558
rect 3409 4512 3442 4558
rect 3390 4510 3442 4512
rect 3278 4286 3293 4338
rect 3293 4286 3330 4338
rect 2718 4062 2737 4114
rect 2737 4062 2770 4114
rect 3950 4421 4002 4450
rect 3950 4398 3965 4421
rect 3965 4398 4002 4421
rect 4622 4286 4637 4338
rect 4637 4286 4674 4338
rect 4062 4062 4081 4114
rect 4081 4062 4114 4114
rect 4734 4062 4753 4114
rect 4753 4062 4786 4114
rect 5742 4286 5757 4338
rect 5757 4286 5794 4338
rect 6526 4558 6578 4562
rect 6526 4512 6545 4558
rect 6545 4512 6578 4558
rect 6526 4510 6578 4512
rect 6414 4421 6466 4450
rect 6414 4398 6429 4421
rect 6429 4398 6466 4421
rect 5854 4062 5873 4114
rect 5873 4062 5906 4114
rect 7198 4558 7250 4562
rect 7198 4512 7217 4558
rect 7217 4512 7250 4558
rect 7198 4510 7250 4512
rect 7086 4421 7138 4450
rect 7086 4398 7101 4421
rect 7101 4398 7138 4421
rect 7758 4421 7810 4450
rect 7758 4398 7773 4421
rect 7773 4398 7810 4421
rect 8430 4286 8445 4338
rect 8445 4286 8482 4338
rect 7870 4062 7889 4114
rect 7889 4062 7922 4114
rect 8542 4062 8561 4114
rect 8561 4062 8594 4114
rect 9998 4286 10013 4338
rect 10013 4286 10050 4338
rect 10110 4062 10129 4114
rect 10129 4062 10162 4114
rect 2376 3894 2636 3946
rect 4700 3894 4960 3946
rect 7024 3894 7284 3946
rect 9348 3894 9608 3946
rect 1934 3390 1986 3442
rect 2046 3502 2083 3554
rect 2083 3502 2098 3554
rect 2606 3419 2621 3442
rect 2621 3419 2658 3442
rect 2606 3390 2658 3419
rect 2718 3502 2770 3554
rect 3278 3419 3293 3442
rect 3293 3419 3330 3442
rect 3278 3390 3330 3419
rect 3390 3390 3442 3442
rect 3950 3419 3965 3442
rect 3965 3419 4002 3442
rect 3950 3390 4002 3419
rect 4062 3390 4114 3442
rect 4622 3419 4637 3442
rect 4637 3419 4674 3442
rect 4622 3390 4674 3419
rect 5854 3726 5873 3778
rect 5873 3726 5906 3778
rect 4734 3390 4786 3442
rect 5742 3419 5757 3442
rect 5757 3419 5794 3442
rect 5742 3390 5794 3419
rect 6750 3726 6769 3778
rect 6769 3726 6802 3778
rect 6638 3502 6653 3554
rect 6653 3502 6690 3554
rect 7422 3726 7441 3778
rect 7441 3726 7474 3778
rect 7310 3502 7325 3554
rect 7325 3502 7362 3554
rect 7982 3726 8015 3778
rect 8015 3726 8034 3778
rect 8766 3661 8785 3666
rect 8785 3661 8818 3666
rect 8766 3614 8818 3661
rect 8094 3502 8131 3554
rect 8131 3502 8146 3554
rect 8654 3502 8669 3554
rect 8669 3502 8706 3554
rect 10110 3661 10129 3666
rect 10129 3661 10162 3666
rect 10110 3614 10162 3661
rect 9998 3419 10013 3442
rect 10013 3419 10050 3442
rect 9998 3390 10050 3419
rect 3538 3110 3798 3162
rect 5862 3110 6122 3162
rect 8186 3110 8446 3162
rect 10510 3110 10770 3162
<< metal2 >>
rect 9884 10724 9940 10734
rect 2374 8652 2638 8662
rect 2374 8586 2638 8596
rect 4698 8652 4962 8662
rect 4698 8586 4962 8596
rect 7022 8652 7286 8662
rect 7022 8586 7286 8596
rect 9346 8652 9610 8662
rect 9346 8586 9610 8596
rect 2268 8372 2324 8382
rect 2156 8148 2212 8158
rect 2268 8148 2324 8316
rect 9772 8372 9828 8382
rect 2156 8146 2324 8148
rect 2156 8094 2158 8146
rect 2210 8094 2324 8146
rect 2156 8092 2324 8094
rect 2156 8082 2212 8092
rect 2268 8034 2324 8092
rect 2828 8148 2884 8158
rect 3500 8148 3556 8158
rect 3612 8148 3668 8158
rect 2828 8146 2996 8148
rect 2828 8094 2830 8146
rect 2882 8094 2996 8146
rect 2828 8092 2996 8094
rect 2828 8082 2884 8092
rect 2268 7982 2270 8034
rect 2322 7982 2324 8034
rect 2156 7474 2212 7486
rect 2156 7422 2158 7474
rect 2210 7422 2212 7474
rect 2156 7252 2212 7422
rect 2268 7252 2324 7982
rect 2940 8034 2996 8092
rect 2940 7982 2942 8034
rect 2994 7982 2996 8034
rect 2828 7476 2884 7486
rect 2940 7476 2996 7982
rect 2156 7250 2324 7252
rect 2156 7198 2270 7250
rect 2322 7198 2324 7250
rect 2156 7196 2324 7198
rect 1932 6578 1988 6590
rect 1932 6526 1934 6578
rect 1986 6526 1988 6578
rect 1932 6468 1988 6526
rect 2044 6468 2100 6478
rect 2156 6468 2212 7196
rect 2268 7186 2324 7196
rect 2716 7474 2996 7476
rect 2716 7422 2830 7474
rect 2882 7422 2942 7474
rect 2994 7422 2996 7474
rect 2716 7420 2996 7422
rect 3388 8146 3668 8148
rect 3388 8094 3502 8146
rect 3554 8094 3614 8146
rect 3666 8094 3668 8146
rect 3388 8092 3668 8094
rect 3388 7476 3444 8092
rect 3500 8082 3556 8092
rect 3612 8082 3668 8092
rect 4172 8148 4228 8158
rect 4172 8146 4340 8148
rect 4172 8094 4174 8146
rect 4226 8094 4340 8146
rect 4172 8092 4340 8094
rect 4172 8082 4228 8092
rect 4284 8034 4340 8092
rect 4284 7982 4286 8034
rect 4338 7982 4340 8034
rect 3536 7868 3800 7878
rect 3536 7802 3800 7812
rect 3500 7476 3556 7486
rect 4172 7476 4228 7486
rect 4284 7476 4340 7982
rect 4844 8146 4900 8158
rect 4844 8094 4846 8146
rect 4898 8094 4900 8146
rect 4844 8036 4900 8094
rect 4956 8036 5012 8046
rect 4844 8034 5012 8036
rect 4844 7982 4958 8034
rect 5010 7982 5012 8034
rect 4844 7980 5012 7982
rect 4844 7476 4900 7980
rect 4956 7970 5012 7980
rect 5860 7868 6124 7878
rect 5860 7802 6124 7812
rect 8184 7868 8448 7878
rect 8184 7802 8448 7812
rect 4956 7476 5012 7486
rect 5628 7476 5684 7486
rect 6300 7476 6356 7486
rect 3388 7474 3556 7476
rect 3388 7422 3502 7474
rect 3554 7422 3556 7474
rect 3388 7420 3556 7422
rect 2374 7084 2638 7094
rect 2374 7018 2638 7028
rect 1932 6466 2212 6468
rect 1932 6414 2046 6466
rect 2098 6414 2212 6466
rect 1932 6412 2212 6414
rect 2604 6578 2660 6590
rect 2604 6526 2606 6578
rect 2658 6526 2660 6578
rect 2604 6468 2660 6526
rect 2716 6468 2772 7420
rect 2828 7410 2884 7420
rect 2940 7410 2996 7420
rect 3500 7252 3556 7420
rect 4060 7474 5012 7476
rect 4060 7422 4174 7474
rect 4226 7422 4286 7474
rect 4338 7422 4846 7474
rect 4898 7422 4958 7474
rect 5010 7422 5012 7474
rect 4060 7420 5012 7422
rect 3612 7252 3668 7262
rect 3500 7250 3668 7252
rect 3500 7198 3614 7250
rect 3666 7198 3668 7250
rect 3500 7196 3668 7198
rect 3276 6580 3332 6590
rect 3388 6580 3444 6590
rect 3500 6580 3556 7196
rect 3612 7186 3668 7196
rect 2604 6466 2772 6468
rect 2604 6414 2718 6466
rect 2770 6414 2772 6466
rect 2604 6412 2772 6414
rect 1820 6020 1876 6030
rect 1932 6020 1988 6412
rect 2044 6402 2100 6412
rect 1820 6018 1932 6020
rect 1820 5966 1822 6018
rect 1874 5966 1932 6018
rect 1820 5964 1932 5966
rect 1820 5954 1876 5964
rect 1932 5926 1988 5964
rect 2492 6020 2548 6030
rect 2604 6020 2660 6412
rect 2716 6402 2772 6412
rect 3164 6578 3556 6580
rect 3164 6526 3278 6578
rect 3330 6526 3390 6578
rect 3442 6526 3556 6578
rect 3164 6524 3556 6526
rect 3948 6578 4004 6590
rect 3948 6526 3950 6578
rect 4002 6526 4004 6578
rect 2492 6018 2604 6020
rect 2492 5966 2494 6018
rect 2546 5966 2604 6018
rect 2492 5964 2604 5966
rect 2492 5954 2548 5964
rect 2604 5926 2660 5964
rect 2940 6020 2996 6030
rect 2374 5516 2638 5526
rect 2374 5450 2638 5460
rect 2268 5348 2324 5358
rect 2044 5292 2268 5348
rect 1932 5124 1988 5134
rect 1932 4452 1988 5068
rect 1820 4450 1988 4452
rect 1820 4398 1934 4450
rect 1986 4398 1988 4450
rect 1820 4396 1988 4398
rect 1820 3444 1876 4396
rect 1932 4386 1988 4396
rect 2044 4562 2100 5292
rect 2268 5254 2324 5292
rect 2604 5348 2660 5358
rect 2156 5124 2212 5134
rect 2156 5030 2212 5068
rect 2044 4510 2046 4562
rect 2098 4510 2100 4562
rect 2044 3554 2100 4510
rect 2604 4450 2660 5292
rect 2940 5348 2996 5964
rect 3164 6020 3220 6524
rect 3276 6514 3332 6524
rect 3388 6514 3444 6524
rect 3948 6468 4004 6526
rect 4060 6468 4116 7420
rect 4172 7410 4228 7420
rect 4284 7410 4340 7420
rect 4844 7410 4900 7420
rect 4956 7410 5012 7420
rect 5516 7474 5684 7476
rect 5516 7422 5630 7474
rect 5682 7422 5684 7474
rect 5516 7420 5684 7422
rect 5516 7250 5572 7420
rect 5628 7410 5684 7420
rect 6188 7474 6356 7476
rect 6188 7422 6302 7474
rect 6354 7422 6356 7474
rect 6188 7420 6356 7422
rect 5516 7198 5518 7250
rect 5570 7198 5572 7250
rect 4698 7084 4962 7094
rect 4698 7018 4962 7028
rect 3948 6466 4116 6468
rect 3948 6414 4062 6466
rect 4114 6414 4116 6466
rect 3948 6412 4116 6414
rect 3536 6300 3800 6310
rect 3536 6234 3800 6244
rect 3164 5926 3220 5964
rect 3500 6020 3556 6030
rect 2828 5124 2884 5134
rect 2828 5030 2884 5068
rect 2604 4398 2606 4450
rect 2658 4398 2660 4450
rect 2604 4386 2660 4398
rect 2940 4228 2996 5292
rect 3276 5682 3332 5694
rect 3276 5630 3278 5682
rect 3330 5630 3332 5682
rect 3276 5124 3332 5630
rect 3500 5124 3556 5964
rect 3836 6020 3892 6030
rect 3948 6020 4004 6412
rect 4060 6402 4116 6412
rect 4620 6578 4676 6590
rect 4620 6526 4622 6578
rect 4674 6526 4676 6578
rect 4620 6468 4676 6526
rect 5516 6580 5572 7198
rect 6188 7250 6244 7420
rect 6300 7410 6356 7420
rect 6188 7198 6190 7250
rect 6242 7198 6244 7250
rect 5740 6580 5796 6590
rect 5516 6524 5740 6580
rect 4732 6468 4788 6478
rect 4620 6466 4788 6468
rect 4620 6414 4734 6466
rect 4786 6414 4788 6466
rect 4620 6412 4788 6414
rect 3892 5964 4004 6020
rect 4284 6020 4340 6030
rect 3836 5926 3892 5964
rect 3948 5684 4004 5694
rect 4060 5684 4116 5694
rect 3948 5682 4060 5684
rect 3948 5630 3950 5682
rect 4002 5630 4060 5682
rect 3948 5628 4060 5630
rect 3948 5618 4004 5628
rect 3276 5058 3332 5068
rect 3388 5122 3556 5124
rect 3388 5070 3502 5122
rect 3554 5070 3556 5122
rect 3388 5068 3556 5070
rect 3388 4564 3444 5068
rect 3500 5058 3556 5068
rect 3612 5124 3668 5134
rect 3612 5030 3668 5068
rect 4060 5012 4116 5628
rect 4284 5346 4340 5964
rect 4508 5908 4564 5918
rect 4620 5908 4676 6412
rect 4732 6402 4788 6412
rect 5740 6468 5796 6524
rect 6188 6580 6244 7198
rect 9212 7252 9268 7262
rect 7022 7084 7286 7094
rect 7022 7018 7286 7028
rect 6188 6514 6244 6524
rect 6412 6580 6468 6590
rect 5852 6468 5908 6478
rect 5740 6466 5908 6468
rect 5740 6414 5854 6466
rect 5906 6414 5908 6466
rect 5740 6412 5908 6414
rect 4508 5906 4676 5908
rect 4508 5854 4510 5906
rect 4562 5854 4676 5906
rect 4508 5852 4676 5854
rect 4508 5842 4564 5852
rect 4620 5684 4676 5852
rect 4620 5618 4676 5628
rect 5180 5906 5236 5918
rect 5180 5854 5182 5906
rect 5234 5854 5236 5906
rect 5180 5684 5236 5854
rect 5292 5684 5348 5694
rect 5236 5682 5348 5684
rect 5236 5630 5294 5682
rect 5346 5630 5348 5682
rect 5236 5628 5348 5630
rect 5180 5618 5236 5628
rect 5292 5618 5348 5628
rect 4698 5516 4962 5526
rect 4698 5450 4962 5460
rect 4284 5294 4286 5346
rect 4338 5294 4340 5346
rect 4284 5282 4340 5294
rect 4172 5012 4228 5022
rect 4844 5012 4900 5022
rect 4956 5012 5012 5022
rect 4060 5010 4228 5012
rect 4060 4958 4174 5010
rect 4226 4958 4228 5010
rect 4060 4956 4228 4958
rect 3536 4732 3800 4742
rect 3536 4666 3800 4676
rect 3388 4562 4004 4564
rect 3388 4510 3390 4562
rect 3442 4510 4004 4562
rect 3388 4508 4004 4510
rect 3388 4498 3444 4508
rect 3948 4450 4004 4508
rect 3948 4398 3950 4450
rect 4002 4398 4004 4450
rect 3948 4386 4004 4398
rect 2828 4172 2996 4228
rect 3276 4338 3332 4350
rect 3276 4286 3278 4338
rect 3330 4286 3332 4338
rect 2716 4114 2772 4126
rect 2716 4062 2718 4114
rect 2770 4062 2772 4114
rect 2374 3948 2638 3958
rect 2374 3882 2638 3892
rect 2716 3780 2772 4062
rect 2044 3502 2046 3554
rect 2098 3502 2100 3554
rect 2044 3490 2100 3502
rect 2604 3724 2772 3780
rect 1932 3444 1988 3454
rect 1820 3442 1988 3444
rect 1820 3390 1934 3442
rect 1986 3390 1988 3442
rect 1820 3388 1988 3390
rect 1932 3332 1988 3388
rect 2604 3444 2660 3724
rect 2716 3556 2772 3566
rect 2828 3556 2884 4172
rect 2716 3554 2884 3556
rect 2716 3502 2718 3554
rect 2770 3502 2884 3554
rect 2716 3500 2884 3502
rect 2716 3490 2772 3500
rect 2604 3350 2660 3388
rect 3276 3444 3332 4286
rect 4060 4114 4116 4956
rect 4172 4946 4228 4956
rect 4732 5010 5012 5012
rect 4732 4958 4846 5010
rect 4898 4958 4958 5010
rect 5010 4958 5012 5010
rect 4732 4956 5012 4958
rect 4620 4338 4676 4350
rect 4620 4286 4622 4338
rect 4674 4286 4676 4338
rect 4620 4116 4676 4286
rect 4732 4116 4788 4956
rect 4844 4946 4900 4956
rect 4956 4946 5012 4956
rect 5740 5012 5796 6412
rect 5852 6402 5908 6412
rect 6412 6468 6468 6524
rect 7084 6580 7140 6590
rect 7196 6580 7252 6590
rect 7140 6578 7252 6580
rect 7140 6526 7198 6578
rect 7250 6526 7252 6578
rect 7140 6524 7252 6526
rect 7084 6486 7140 6524
rect 7196 6514 7252 6524
rect 8428 6580 8484 6590
rect 8428 6578 8596 6580
rect 8428 6526 8430 6578
rect 8482 6526 8596 6578
rect 8428 6524 8596 6526
rect 8428 6514 8484 6524
rect 6524 6468 6580 6478
rect 6412 6466 6580 6468
rect 6412 6414 6526 6466
rect 6578 6414 6580 6466
rect 6412 6412 6580 6414
rect 5860 6300 6124 6310
rect 5860 6234 6124 6244
rect 5852 6020 5908 6030
rect 6412 6020 6468 6412
rect 6524 6402 6580 6412
rect 8540 6468 8596 6524
rect 8540 6466 8708 6468
rect 8540 6414 8542 6466
rect 8594 6414 8708 6466
rect 8540 6412 8708 6414
rect 8540 6402 8596 6412
rect 8184 6300 8448 6310
rect 8184 6234 8448 6244
rect 6524 6020 6580 6030
rect 6636 6020 6692 6030
rect 6412 6018 6692 6020
rect 6412 5966 6526 6018
rect 6578 5966 6638 6018
rect 6690 5966 6692 6018
rect 6412 5964 6692 5966
rect 5852 5926 5908 5964
rect 6524 5954 6580 5964
rect 6636 5954 6692 5964
rect 7756 6020 7812 6030
rect 7756 5926 7812 5964
rect 8316 6020 8372 6030
rect 8428 6020 8484 6030
rect 8372 6018 8484 6020
rect 8372 5966 8430 6018
rect 8482 5966 8484 6018
rect 8372 5964 8484 5966
rect 5964 5682 6020 5694
rect 5964 5630 5966 5682
rect 6018 5630 6020 5682
rect 5964 5348 6020 5630
rect 7868 5684 7924 5694
rect 7022 5516 7286 5526
rect 7022 5450 7286 5460
rect 5964 5282 6020 5292
rect 7084 5348 7140 5358
rect 6972 5124 7028 5134
rect 7084 5124 7140 5292
rect 7756 5348 7812 5358
rect 7868 5348 7924 5628
rect 7812 5292 7924 5348
rect 7756 5216 7812 5292
rect 6972 5122 7140 5124
rect 6972 5070 6974 5122
rect 7026 5070 7140 5122
rect 6972 5068 7140 5070
rect 6972 5058 7028 5068
rect 5852 5012 5908 5022
rect 5740 5010 5908 5012
rect 5740 4958 5742 5010
rect 5794 4958 5854 5010
rect 5906 4958 5908 5010
rect 5740 4956 5908 4958
rect 4060 4062 4062 4114
rect 4114 4062 4116 4114
rect 3388 3444 3444 3454
rect 3276 3442 3444 3444
rect 3276 3390 3278 3442
rect 3330 3390 3390 3442
rect 3442 3390 3444 3442
rect 3276 3388 3444 3390
rect 3276 3378 3332 3388
rect 1932 2996 1988 3276
rect 3388 3332 3444 3388
rect 3388 3266 3444 3276
rect 3948 3444 4004 3454
rect 4060 3444 4116 4062
rect 3948 3442 4116 3444
rect 3948 3390 3950 3442
rect 4002 3390 4062 3442
rect 4114 3390 4116 3442
rect 3948 3388 4116 3390
rect 4508 4114 4788 4116
rect 4508 4062 4734 4114
rect 4786 4062 4788 4114
rect 4508 4060 4788 4062
rect 4508 3444 4564 4060
rect 4732 4050 4788 4060
rect 5740 4452 5796 4956
rect 5852 4946 5908 4956
rect 5860 4732 6124 4742
rect 5860 4666 6124 4676
rect 6524 4564 6580 4574
rect 7084 4564 7140 5068
rect 8316 5122 8372 5964
rect 8428 5954 8484 5964
rect 8540 5684 8596 5694
rect 8316 5070 8318 5122
rect 8370 5070 8372 5122
rect 8316 5058 8372 5070
rect 8428 5124 8484 5134
rect 8540 5124 8596 5628
rect 8484 5068 8596 5124
rect 8428 5030 8484 5068
rect 7644 5010 7700 5022
rect 7644 4958 7646 5010
rect 7698 4958 7700 5010
rect 7196 4564 7252 4574
rect 6524 4562 7252 4564
rect 6524 4510 6526 4562
rect 6578 4510 7198 4562
rect 7250 4510 7252 4562
rect 6524 4508 7252 4510
rect 5740 4338 5796 4396
rect 6412 4452 6468 4462
rect 6524 4452 6580 4508
rect 6412 4450 6580 4452
rect 6412 4398 6414 4450
rect 6466 4398 6580 4450
rect 6412 4396 6580 4398
rect 6412 4386 6468 4396
rect 5740 4286 5742 4338
rect 5794 4286 5796 4338
rect 4698 3948 4962 3958
rect 4698 3882 4962 3892
rect 5740 3780 5796 4286
rect 5852 4116 5908 4126
rect 5852 4022 5908 4060
rect 5852 3780 5908 3790
rect 6748 3780 6804 4508
rect 7084 4450 7140 4508
rect 7196 4498 7252 4508
rect 7084 4398 7086 4450
rect 7138 4398 7140 4450
rect 7084 4386 7140 4398
rect 7420 4116 7476 4126
rect 7022 3948 7286 3958
rect 7022 3882 7286 3892
rect 5740 3778 5908 3780
rect 5740 3726 5854 3778
rect 5906 3726 5908 3778
rect 5740 3724 5908 3726
rect 4620 3444 4676 3454
rect 4732 3444 4788 3454
rect 4508 3442 4788 3444
rect 4508 3390 4622 3442
rect 4674 3390 4734 3442
rect 4786 3390 4788 3442
rect 4508 3388 4788 3390
rect 3948 3332 4004 3388
rect 4060 3378 4116 3388
rect 3948 3266 4004 3276
rect 4620 3332 4676 3388
rect 4732 3378 4788 3388
rect 5740 3444 5796 3724
rect 5852 3714 5908 3724
rect 6636 3778 7364 3780
rect 6636 3726 6750 3778
rect 6802 3726 7364 3778
rect 6636 3724 7364 3726
rect 6636 3554 6692 3724
rect 6748 3714 6804 3724
rect 6636 3502 6638 3554
rect 6690 3502 6692 3554
rect 6636 3490 6692 3502
rect 7308 3554 7364 3724
rect 7420 3778 7476 4060
rect 7644 4116 7700 4958
rect 8652 4900 8708 6412
rect 9212 5124 9268 7196
rect 9346 7084 9610 7094
rect 9346 7018 9610 7028
rect 9772 6804 9828 8316
rect 9884 7028 9940 10668
rect 10508 7868 10772 7878
rect 10508 7802 10772 7812
rect 10108 7476 10164 7486
rect 10108 7474 10276 7476
rect 10108 7422 10110 7474
rect 10162 7422 10276 7474
rect 10108 7420 10276 7422
rect 10108 7410 10164 7420
rect 9996 7252 10052 7262
rect 9996 7158 10052 7196
rect 9884 6972 10052 7028
rect 9996 6804 10052 6972
rect 10108 6804 10164 6814
rect 9772 6802 9940 6804
rect 9772 6750 9774 6802
rect 9826 6750 9940 6802
rect 9772 6748 9940 6750
rect 9996 6802 10164 6804
rect 9996 6750 10110 6802
rect 10162 6750 10164 6802
rect 9996 6748 10164 6750
rect 9772 6738 9828 6748
rect 9660 6690 9716 6702
rect 9660 6638 9662 6690
rect 9714 6638 9716 6690
rect 9660 6020 9716 6638
rect 9884 6132 9940 6748
rect 10108 6738 10164 6748
rect 9996 6132 10052 6142
rect 9884 6130 10052 6132
rect 9884 6078 9998 6130
rect 10050 6078 10052 6130
rect 9884 6076 10052 6078
rect 9996 6066 10052 6076
rect 9660 5954 9716 5964
rect 9996 5908 10052 5918
rect 9346 5516 9610 5526
rect 9346 5450 9610 5460
rect 9996 5346 10052 5852
rect 10108 5908 10164 5918
rect 10220 5908 10276 7420
rect 10508 6300 10772 6310
rect 10508 6234 10772 6244
rect 10108 5906 10276 5908
rect 10108 5854 10110 5906
rect 10162 5854 10276 5906
rect 10108 5852 10276 5854
rect 10108 5842 10164 5852
rect 9996 5294 9998 5346
rect 10050 5294 10052 5346
rect 9996 5282 10052 5294
rect 9212 5058 9268 5068
rect 9884 5124 9940 5134
rect 10108 5124 10164 5134
rect 9940 5122 10164 5124
rect 9940 5070 10110 5122
rect 10162 5070 10164 5122
rect 9940 5068 10164 5070
rect 9324 5010 9380 5022
rect 9324 4958 9326 5010
rect 9378 4958 9380 5010
rect 9324 4900 9380 4958
rect 9436 4900 9492 4910
rect 9324 4844 9436 4900
rect 8652 4834 8708 4844
rect 9436 4806 9492 4844
rect 8184 4732 8448 4742
rect 8184 4666 8448 4676
rect 7756 4452 7812 4462
rect 7756 4358 7812 4396
rect 8428 4452 8484 4462
rect 8428 4340 8484 4396
rect 8428 4338 8708 4340
rect 8428 4286 8430 4338
rect 8482 4286 8708 4338
rect 8428 4284 8708 4286
rect 8428 4274 8484 4284
rect 7644 4050 7700 4060
rect 7868 4116 7924 4126
rect 7420 3726 7422 3778
rect 7474 3726 7476 3778
rect 7420 3714 7476 3726
rect 7868 3780 7924 4060
rect 8540 4114 8596 4126
rect 8540 4062 8542 4114
rect 8594 4062 8596 4114
rect 7980 3780 8036 3790
rect 7868 3778 8036 3780
rect 7868 3726 7982 3778
rect 8034 3726 8036 3778
rect 7868 3724 8036 3726
rect 7308 3502 7310 3554
rect 7362 3502 7364 3554
rect 7308 3490 7364 3502
rect 7980 3668 8036 3724
rect 7980 3556 8036 3612
rect 8540 3668 8596 4062
rect 8540 3602 8596 3612
rect 8092 3556 8148 3566
rect 7980 3554 8148 3556
rect 7980 3502 8094 3554
rect 8146 3502 8148 3554
rect 7980 3500 8148 3502
rect 8092 3490 8148 3500
rect 8652 3554 8708 4284
rect 9346 3948 9610 3958
rect 9346 3882 9610 3892
rect 8764 3668 8820 3678
rect 8764 3574 8820 3612
rect 8652 3502 8654 3554
rect 8706 3502 8708 3554
rect 8652 3490 8708 3502
rect 9884 3444 9940 5068
rect 10108 5058 10164 5068
rect 9996 4900 10052 4910
rect 9996 4340 10052 4844
rect 10220 4900 10276 5852
rect 10220 4834 10276 4844
rect 10508 4732 10772 4742
rect 10508 4666 10772 4676
rect 9996 4338 10164 4340
rect 9996 4286 9998 4338
rect 10050 4286 10164 4338
rect 9996 4284 10164 4286
rect 9996 4274 10052 4284
rect 10108 4114 10164 4284
rect 10108 4062 10110 4114
rect 10162 4062 10164 4114
rect 10108 3668 10164 4062
rect 10108 3574 10164 3612
rect 9996 3444 10052 3454
rect 9884 3442 10052 3444
rect 9884 3390 9998 3442
rect 10050 3390 10052 3442
rect 9884 3388 10052 3390
rect 5740 3350 5796 3388
rect 4620 3266 4676 3276
rect 3536 3164 3800 3174
rect 3536 3098 3800 3108
rect 5860 3164 6124 3174
rect 5860 3098 6124 3108
rect 8184 3164 8448 3174
rect 8184 3098 8448 3108
rect 1932 2930 1988 2940
rect 9996 1316 10052 3388
rect 10508 3164 10772 3174
rect 10508 3098 10772 3108
rect 9996 1250 10052 1260
<< via2 >>
rect 9884 10668 9940 10724
rect 2374 8650 2638 8652
rect 2374 8598 2376 8650
rect 2376 8598 2636 8650
rect 2636 8598 2638 8650
rect 2374 8596 2638 8598
rect 4698 8650 4962 8652
rect 4698 8598 4700 8650
rect 4700 8598 4960 8650
rect 4960 8598 4962 8650
rect 4698 8596 4962 8598
rect 7022 8650 7286 8652
rect 7022 8598 7024 8650
rect 7024 8598 7284 8650
rect 7284 8598 7286 8650
rect 7022 8596 7286 8598
rect 9346 8650 9610 8652
rect 9346 8598 9348 8650
rect 9348 8598 9608 8650
rect 9608 8598 9610 8650
rect 9346 8596 9610 8598
rect 2268 8316 2324 8372
rect 9772 8316 9828 8372
rect 3536 7866 3800 7868
rect 3536 7814 3538 7866
rect 3538 7814 3798 7866
rect 3798 7814 3800 7866
rect 3536 7812 3800 7814
rect 5860 7866 6124 7868
rect 5860 7814 5862 7866
rect 5862 7814 6122 7866
rect 6122 7814 6124 7866
rect 5860 7812 6124 7814
rect 8184 7866 8448 7868
rect 8184 7814 8186 7866
rect 8186 7814 8446 7866
rect 8446 7814 8448 7866
rect 8184 7812 8448 7814
rect 2374 7082 2638 7084
rect 2374 7030 2376 7082
rect 2376 7030 2636 7082
rect 2636 7030 2638 7082
rect 2374 7028 2638 7030
rect 1932 6018 1988 6020
rect 1932 5966 1934 6018
rect 1934 5966 1986 6018
rect 1986 5966 1988 6018
rect 1932 5964 1988 5966
rect 2604 6018 2660 6020
rect 2604 5966 2606 6018
rect 2606 5966 2658 6018
rect 2658 5966 2660 6018
rect 2604 5964 2660 5966
rect 2940 5964 2996 6020
rect 2374 5514 2638 5516
rect 2374 5462 2376 5514
rect 2376 5462 2636 5514
rect 2636 5462 2638 5514
rect 2374 5460 2638 5462
rect 2268 5346 2324 5348
rect 2268 5294 2270 5346
rect 2270 5294 2322 5346
rect 2322 5294 2324 5346
rect 2268 5292 2324 5294
rect 1932 5068 1988 5124
rect 2604 5292 2660 5348
rect 2156 5122 2212 5124
rect 2156 5070 2158 5122
rect 2158 5070 2210 5122
rect 2210 5070 2212 5122
rect 2156 5068 2212 5070
rect 4698 7082 4962 7084
rect 4698 7030 4700 7082
rect 4700 7030 4960 7082
rect 4960 7030 4962 7082
rect 4698 7028 4962 7030
rect 3536 6298 3800 6300
rect 3536 6246 3538 6298
rect 3538 6246 3798 6298
rect 3798 6246 3800 6298
rect 3536 6244 3800 6246
rect 3164 6018 3220 6020
rect 3164 5966 3166 6018
rect 3166 5966 3218 6018
rect 3218 5966 3220 6018
rect 3164 5964 3220 5966
rect 3500 5964 3556 6020
rect 2940 5346 2996 5348
rect 2940 5294 2942 5346
rect 2942 5294 2994 5346
rect 2994 5294 2996 5346
rect 2940 5292 2996 5294
rect 2828 5122 2884 5124
rect 2828 5070 2830 5122
rect 2830 5070 2882 5122
rect 2882 5070 2884 5122
rect 2828 5068 2884 5070
rect 5740 6578 5796 6580
rect 5740 6526 5742 6578
rect 5742 6526 5794 6578
rect 5794 6526 5796 6578
rect 5740 6524 5796 6526
rect 3836 6018 3892 6020
rect 3836 5966 3838 6018
rect 3838 5966 3890 6018
rect 3890 5966 3892 6018
rect 3836 5964 3892 5966
rect 4284 5964 4340 6020
rect 4060 5628 4116 5684
rect 3276 5068 3332 5124
rect 3612 5122 3668 5124
rect 3612 5070 3614 5122
rect 3614 5070 3666 5122
rect 3666 5070 3668 5122
rect 3612 5068 3668 5070
rect 9212 7196 9268 7252
rect 7022 7082 7286 7084
rect 7022 7030 7024 7082
rect 7024 7030 7284 7082
rect 7284 7030 7286 7082
rect 7022 7028 7286 7030
rect 6188 6524 6244 6580
rect 6412 6578 6468 6580
rect 6412 6526 6414 6578
rect 6414 6526 6466 6578
rect 6466 6526 6468 6578
rect 6412 6524 6468 6526
rect 4620 5682 4676 5684
rect 4620 5630 4622 5682
rect 4622 5630 4674 5682
rect 4674 5630 4676 5682
rect 4620 5628 4676 5630
rect 5180 5628 5236 5684
rect 4698 5514 4962 5516
rect 4698 5462 4700 5514
rect 4700 5462 4960 5514
rect 4960 5462 4962 5514
rect 4698 5460 4962 5462
rect 3536 4730 3800 4732
rect 3536 4678 3538 4730
rect 3538 4678 3798 4730
rect 3798 4678 3800 4730
rect 3536 4676 3800 4678
rect 2374 3946 2638 3948
rect 2374 3894 2376 3946
rect 2376 3894 2636 3946
rect 2636 3894 2638 3946
rect 2374 3892 2638 3894
rect 2604 3442 2660 3444
rect 2604 3390 2606 3442
rect 2606 3390 2658 3442
rect 2658 3390 2660 3442
rect 2604 3388 2660 3390
rect 7084 6578 7140 6580
rect 7084 6526 7086 6578
rect 7086 6526 7138 6578
rect 7138 6526 7140 6578
rect 7084 6524 7140 6526
rect 5860 6298 6124 6300
rect 5860 6246 5862 6298
rect 5862 6246 6122 6298
rect 6122 6246 6124 6298
rect 5860 6244 6124 6246
rect 5852 6018 5908 6020
rect 5852 5966 5854 6018
rect 5854 5966 5906 6018
rect 5906 5966 5908 6018
rect 5852 5964 5908 5966
rect 8184 6298 8448 6300
rect 8184 6246 8186 6298
rect 8186 6246 8446 6298
rect 8446 6246 8448 6298
rect 8184 6244 8448 6246
rect 7756 6018 7812 6020
rect 7756 5966 7758 6018
rect 7758 5966 7810 6018
rect 7810 5966 7812 6018
rect 7756 5964 7812 5966
rect 8316 5964 8372 6020
rect 7868 5682 7924 5684
rect 7868 5630 7870 5682
rect 7870 5630 7922 5682
rect 7922 5630 7924 5682
rect 7868 5628 7924 5630
rect 7022 5514 7286 5516
rect 7022 5462 7024 5514
rect 7024 5462 7284 5514
rect 7284 5462 7286 5514
rect 7022 5460 7286 5462
rect 5964 5292 6020 5348
rect 7084 5346 7140 5348
rect 7084 5294 7086 5346
rect 7086 5294 7138 5346
rect 7138 5294 7140 5346
rect 7084 5292 7140 5294
rect 7756 5346 7812 5348
rect 7756 5294 7758 5346
rect 7758 5294 7810 5346
rect 7810 5294 7812 5346
rect 7756 5292 7812 5294
rect 1932 3276 1988 3332
rect 3388 3276 3444 3332
rect 5860 4730 6124 4732
rect 5860 4678 5862 4730
rect 5862 4678 6122 4730
rect 6122 4678 6124 4730
rect 5860 4676 6124 4678
rect 8540 5682 8596 5684
rect 8540 5630 8542 5682
rect 8542 5630 8594 5682
rect 8594 5630 8596 5682
rect 8540 5628 8596 5630
rect 8428 5122 8484 5124
rect 8428 5070 8430 5122
rect 8430 5070 8482 5122
rect 8482 5070 8484 5122
rect 8428 5068 8484 5070
rect 5740 4396 5796 4452
rect 4698 3946 4962 3948
rect 4698 3894 4700 3946
rect 4700 3894 4960 3946
rect 4960 3894 4962 3946
rect 4698 3892 4962 3894
rect 5852 4114 5908 4116
rect 5852 4062 5854 4114
rect 5854 4062 5906 4114
rect 5906 4062 5908 4114
rect 5852 4060 5908 4062
rect 7420 4060 7476 4116
rect 7022 3946 7286 3948
rect 7022 3894 7024 3946
rect 7024 3894 7284 3946
rect 7284 3894 7286 3946
rect 7022 3892 7286 3894
rect 3948 3276 4004 3332
rect 9346 7082 9610 7084
rect 9346 7030 9348 7082
rect 9348 7030 9608 7082
rect 9608 7030 9610 7082
rect 9346 7028 9610 7030
rect 10508 7866 10772 7868
rect 10508 7814 10510 7866
rect 10510 7814 10770 7866
rect 10770 7814 10772 7866
rect 10508 7812 10772 7814
rect 9996 7250 10052 7252
rect 9996 7198 9998 7250
rect 9998 7198 10050 7250
rect 10050 7198 10052 7250
rect 9996 7196 10052 7198
rect 9660 5964 9716 6020
rect 9996 5852 10052 5908
rect 9346 5514 9610 5516
rect 9346 5462 9348 5514
rect 9348 5462 9608 5514
rect 9608 5462 9610 5514
rect 9346 5460 9610 5462
rect 10508 6298 10772 6300
rect 10508 6246 10510 6298
rect 10510 6246 10770 6298
rect 10770 6246 10772 6298
rect 10508 6244 10772 6246
rect 9212 5068 9268 5124
rect 9884 5068 9940 5124
rect 8652 4844 8708 4900
rect 9436 4898 9492 4900
rect 9436 4846 9438 4898
rect 9438 4846 9490 4898
rect 9490 4846 9492 4898
rect 9436 4844 9492 4846
rect 8184 4730 8448 4732
rect 8184 4678 8186 4730
rect 8186 4678 8446 4730
rect 8446 4678 8448 4730
rect 8184 4676 8448 4678
rect 7756 4450 7812 4452
rect 7756 4398 7758 4450
rect 7758 4398 7810 4450
rect 7810 4398 7812 4450
rect 7756 4396 7812 4398
rect 8428 4396 8484 4452
rect 7644 4060 7700 4116
rect 7868 4114 7924 4116
rect 7868 4062 7870 4114
rect 7870 4062 7922 4114
rect 7922 4062 7924 4114
rect 7868 4060 7924 4062
rect 7980 3612 8036 3668
rect 8540 3612 8596 3668
rect 9346 3946 9610 3948
rect 9346 3894 9348 3946
rect 9348 3894 9608 3946
rect 9608 3894 9610 3946
rect 9346 3892 9610 3894
rect 8764 3666 8820 3668
rect 8764 3614 8766 3666
rect 8766 3614 8818 3666
rect 8818 3614 8820 3666
rect 8764 3612 8820 3614
rect 5740 3442 5796 3444
rect 5740 3390 5742 3442
rect 5742 3390 5794 3442
rect 5794 3390 5796 3442
rect 5740 3388 5796 3390
rect 9996 4844 10052 4900
rect 10220 4844 10276 4900
rect 10508 4730 10772 4732
rect 10508 4678 10510 4730
rect 10510 4678 10770 4730
rect 10770 4678 10772 4730
rect 10508 4676 10772 4678
rect 10108 3666 10164 3668
rect 10108 3614 10110 3666
rect 10110 3614 10162 3666
rect 10162 3614 10164 3666
rect 10108 3612 10164 3614
rect 4620 3276 4676 3332
rect 3536 3162 3800 3164
rect 3536 3110 3538 3162
rect 3538 3110 3798 3162
rect 3798 3110 3800 3162
rect 3536 3108 3800 3110
rect 5860 3162 6124 3164
rect 5860 3110 5862 3162
rect 5862 3110 6122 3162
rect 6122 3110 6124 3162
rect 5860 3108 6124 3110
rect 8184 3162 8448 3164
rect 8184 3110 8186 3162
rect 8186 3110 8446 3162
rect 8446 3110 8448 3162
rect 8184 3108 8448 3110
rect 1932 2940 1988 2996
rect 10508 3162 10772 3164
rect 10508 3110 10510 3162
rect 10510 3110 10770 3162
rect 10770 3110 10772 3162
rect 10508 3108 10772 3110
rect 9996 1260 10052 1316
<< metal3 >>
rect 11200 10724 12000 10752
rect 9874 10668 9884 10724
rect 9940 10668 12000 10724
rect 11200 10640 12000 10668
rect 0 8932 800 8960
rect 0 8876 1316 8932
rect 0 8848 800 8876
rect 1260 8484 1316 8876
rect 2364 8596 2374 8652
rect 2638 8596 2648 8652
rect 4688 8596 4698 8652
rect 4962 8596 4972 8652
rect 7012 8596 7022 8652
rect 7286 8596 7296 8652
rect 9336 8596 9346 8652
rect 9610 8596 9620 8652
rect 1260 8428 2324 8484
rect 2268 8372 2324 8428
rect 11200 8372 12000 8400
rect 2258 8316 2268 8372
rect 2324 8316 2334 8372
rect 9762 8316 9772 8372
rect 9828 8316 12000 8372
rect 11200 8288 12000 8316
rect 3526 7812 3536 7868
rect 3800 7812 3810 7868
rect 5850 7812 5860 7868
rect 6124 7812 6134 7868
rect 8174 7812 8184 7868
rect 8448 7812 8458 7868
rect 10498 7812 10508 7868
rect 10772 7812 10782 7868
rect 9202 7196 9212 7252
rect 9268 7196 9996 7252
rect 10052 7196 10062 7252
rect 2364 7028 2374 7084
rect 2638 7028 2648 7084
rect 4688 7028 4698 7084
rect 4962 7028 4972 7084
rect 7012 7028 7022 7084
rect 7286 7028 7296 7084
rect 9336 7028 9346 7084
rect 9610 7028 9620 7084
rect 5730 6524 5740 6580
rect 5796 6524 6188 6580
rect 6244 6524 6412 6580
rect 6468 6524 7084 6580
rect 7140 6524 7150 6580
rect 3526 6244 3536 6300
rect 3800 6244 3810 6300
rect 5850 6244 5860 6300
rect 6124 6244 6134 6300
rect 8174 6244 8184 6300
rect 8448 6244 8458 6300
rect 10498 6244 10508 6300
rect 10772 6244 10782 6300
rect 11200 6020 12000 6048
rect 1922 5964 1932 6020
rect 1988 5964 2604 6020
rect 2660 5964 2940 6020
rect 2996 5964 3164 6020
rect 3220 5964 3500 6020
rect 3556 5964 3836 6020
rect 3892 5964 4284 6020
rect 4340 5964 5852 6020
rect 5908 5964 7756 6020
rect 7812 5964 8316 6020
rect 8372 5964 8382 6020
rect 9650 5964 9660 6020
rect 9716 5964 12000 6020
rect 9996 5908 10052 5964
rect 11200 5936 12000 5964
rect 9986 5852 9996 5908
rect 10052 5852 10062 5908
rect 4050 5628 4060 5684
rect 4116 5628 4620 5684
rect 4676 5628 5180 5684
rect 5236 5628 5246 5684
rect 7858 5628 7868 5684
rect 7924 5628 8540 5684
rect 8596 5628 8606 5684
rect 2364 5460 2374 5516
rect 2638 5460 2648 5516
rect 4688 5460 4698 5516
rect 4962 5460 4972 5516
rect 7012 5460 7022 5516
rect 7286 5460 7296 5516
rect 9336 5460 9346 5516
rect 9610 5460 9620 5516
rect 2258 5292 2268 5348
rect 2324 5292 2604 5348
rect 2660 5292 2940 5348
rect 2996 5292 3006 5348
rect 5954 5292 5964 5348
rect 6020 5292 7084 5348
rect 7140 5292 7756 5348
rect 7812 5292 7822 5348
rect 1922 5068 1932 5124
rect 1988 5068 2156 5124
rect 2212 5068 2828 5124
rect 2884 5068 3276 5124
rect 3332 5068 3612 5124
rect 3668 5068 3678 5124
rect 8418 5068 8428 5124
rect 8484 5068 9212 5124
rect 9268 5068 9884 5124
rect 9940 5068 9950 5124
rect 8642 4844 8652 4900
rect 8708 4844 9436 4900
rect 9492 4844 9996 4900
rect 10052 4844 10220 4900
rect 10276 4844 10286 4900
rect 3526 4676 3536 4732
rect 3800 4676 3810 4732
rect 5850 4676 5860 4732
rect 6124 4676 6134 4732
rect 8174 4676 8184 4732
rect 8448 4676 8458 4732
rect 10498 4676 10508 4732
rect 10772 4676 10782 4732
rect 5730 4396 5740 4452
rect 5796 4396 7756 4452
rect 7812 4396 8428 4452
rect 8484 4396 8494 4452
rect 5842 4060 5852 4116
rect 5908 4060 7420 4116
rect 7476 4060 7644 4116
rect 7700 4060 7868 4116
rect 7924 4060 7934 4116
rect 2364 3892 2374 3948
rect 2638 3892 2648 3948
rect 4688 3892 4698 3948
rect 4962 3892 4972 3948
rect 7012 3892 7022 3948
rect 7286 3892 7296 3948
rect 9336 3892 9346 3948
rect 9610 3892 9620 3948
rect 11200 3668 12000 3696
rect 7970 3612 7980 3668
rect 8036 3612 8540 3668
rect 8596 3612 8764 3668
rect 8820 3612 10108 3668
rect 10164 3612 12000 3668
rect 11200 3584 12000 3612
rect 2594 3388 2604 3444
rect 2660 3388 2670 3444
rect 4956 3388 5740 3444
rect 5796 3388 5806 3444
rect 2604 3332 2660 3388
rect 4956 3332 5012 3388
rect 1922 3276 1932 3332
rect 1988 3276 3388 3332
rect 3444 3276 3948 3332
rect 4004 3276 4620 3332
rect 4676 3276 5012 3332
rect 3526 3108 3536 3164
rect 3800 3108 3810 3164
rect 5850 3108 5860 3164
rect 6124 3108 6134 3164
rect 8174 3108 8184 3164
rect 8448 3108 8458 3164
rect 10498 3108 10508 3164
rect 10772 3108 10782 3164
rect 0 2996 800 3024
rect 0 2940 1932 2996
rect 1988 2940 1998 2996
rect 0 2912 800 2940
rect 11200 1316 12000 1344
rect 9986 1260 9996 1316
rect 10052 1260 12000 1316
rect 11200 1232 12000 1260
<< via3 >>
rect 2374 8596 2638 8652
rect 4698 8596 4962 8652
rect 7022 8596 7286 8652
rect 9346 8596 9610 8652
rect 3536 7812 3800 7868
rect 5860 7812 6124 7868
rect 8184 7812 8448 7868
rect 10508 7812 10772 7868
rect 2374 7028 2638 7084
rect 4698 7028 4962 7084
rect 7022 7028 7286 7084
rect 9346 7028 9610 7084
rect 3536 6244 3800 6300
rect 5860 6244 6124 6300
rect 8184 6244 8448 6300
rect 10508 6244 10772 6300
rect 2374 5460 2638 5516
rect 4698 5460 4962 5516
rect 7022 5460 7286 5516
rect 9346 5460 9610 5516
rect 3536 4676 3800 4732
rect 5860 4676 6124 4732
rect 8184 4676 8448 4732
rect 10508 4676 10772 4732
rect 2374 3892 2638 3948
rect 4698 3892 4962 3948
rect 7022 3892 7286 3948
rect 9346 3892 9610 3948
rect 3536 3108 3800 3164
rect 5860 3108 6124 3164
rect 8184 3108 8448 3164
rect 10508 3108 10772 3164
<< metal4 >>
rect 2346 8652 2666 8684
rect 2346 8596 2374 8652
rect 2638 8596 2666 8652
rect 2346 7084 2666 8596
rect 2346 7028 2374 7084
rect 2638 7028 2666 7084
rect 2346 5516 2666 7028
rect 2346 5460 2374 5516
rect 2638 5460 2666 5516
rect 2346 3948 2666 5460
rect 2346 3892 2374 3948
rect 2638 3892 2666 3948
rect 2346 3076 2666 3892
rect 3508 7868 3828 8684
rect 3508 7812 3536 7868
rect 3800 7812 3828 7868
rect 3508 6300 3828 7812
rect 3508 6244 3536 6300
rect 3800 6244 3828 6300
rect 3508 4732 3828 6244
rect 3508 4676 3536 4732
rect 3800 4676 3828 4732
rect 3508 3164 3828 4676
rect 3508 3108 3536 3164
rect 3800 3108 3828 3164
rect 3508 3076 3828 3108
rect 4670 8652 4990 8684
rect 4670 8596 4698 8652
rect 4962 8596 4990 8652
rect 4670 7084 4990 8596
rect 4670 7028 4698 7084
rect 4962 7028 4990 7084
rect 4670 5516 4990 7028
rect 4670 5460 4698 5516
rect 4962 5460 4990 5516
rect 4670 3948 4990 5460
rect 4670 3892 4698 3948
rect 4962 3892 4990 3948
rect 4670 3076 4990 3892
rect 5832 7868 6152 8684
rect 5832 7812 5860 7868
rect 6124 7812 6152 7868
rect 5832 6300 6152 7812
rect 5832 6244 5860 6300
rect 6124 6244 6152 6300
rect 5832 4732 6152 6244
rect 5832 4676 5860 4732
rect 6124 4676 6152 4732
rect 5832 3164 6152 4676
rect 5832 3108 5860 3164
rect 6124 3108 6152 3164
rect 5832 3076 6152 3108
rect 6994 8652 7314 8684
rect 6994 8596 7022 8652
rect 7286 8596 7314 8652
rect 6994 7084 7314 8596
rect 6994 7028 7022 7084
rect 7286 7028 7314 7084
rect 6994 5516 7314 7028
rect 6994 5460 7022 5516
rect 7286 5460 7314 5516
rect 6994 3948 7314 5460
rect 6994 3892 7022 3948
rect 7286 3892 7314 3948
rect 6994 3076 7314 3892
rect 8156 7868 8476 8684
rect 8156 7812 8184 7868
rect 8448 7812 8476 7868
rect 8156 6300 8476 7812
rect 8156 6244 8184 6300
rect 8448 6244 8476 6300
rect 8156 4732 8476 6244
rect 8156 4676 8184 4732
rect 8448 4676 8476 4732
rect 8156 3164 8476 4676
rect 8156 3108 8184 3164
rect 8448 3108 8476 3164
rect 8156 3076 8476 3108
rect 9318 8652 9638 8684
rect 9318 8596 9346 8652
rect 9610 8596 9638 8652
rect 9318 7084 9638 8596
rect 9318 7028 9346 7084
rect 9610 7028 9638 7084
rect 9318 5516 9638 7028
rect 9318 5460 9346 5516
rect 9610 5460 9638 5516
rect 9318 3948 9638 5460
rect 9318 3892 9346 3948
rect 9610 3892 9638 3948
rect 9318 3076 9638 3892
rect 10480 7868 10800 8684
rect 10480 7812 10508 7868
rect 10772 7812 10800 7868
rect 10480 6300 10800 7812
rect 10480 6244 10508 6300
rect 10772 6244 10800 6300
rect 10480 4732 10800 6244
rect 10480 4676 10508 4732
rect 10772 4676 10800 4732
rect 10480 3164 10800 4676
rect 10480 3108 10508 3164
rect 10772 3108 10800 3164
rect 10480 3076 10800 3108
<< labels >>
rlabel metal1 s 5992 8624 5992 8624 4 vdd
rlabel metal2 s 6072 7840 6072 7840 4 vss
rlabel metal2 s 8344 5544 8344 5544 4 nbus
rlabel metal2 s 7448 3920 7448 3920 4 outn
rlabel metal2 s 9800 7560 9800 7560 4 outnn
rlabel metal2 s 7840 5320 7840 5320 4 outp
rlabel metal2 s 10024 5600 10024 5600 4 outpn
rlabel metal2 s 10080 6776 10080 6776 4 outxor
rlabel metal2 s 1960 3192 1960 3192 4 pbus
flabel metal3 s 0 8848 800 8960 0 FreeSans 560 0 0 0 nbus
port 1 nsew
flabel metal3 s 11200 3584 12000 3696 0 FreeSans 560 0 0 0 outn
port 2 nsew
flabel metal3 s 11200 8288 12000 8400 0 FreeSans 560 0 0 0 outnn
port 3 nsew
flabel metal3 s 11200 1232 12000 1344 0 FreeSans 560 0 0 0 outp
port 4 nsew
flabel metal3 s 11200 5936 12000 6048 0 FreeSans 560 0 0 0 outpn
port 5 nsew
flabel metal3 s 11200 10640 12000 10752 0 FreeSans 560 0 0 0 outxor
port 6 nsew
flabel metal3 s 0 2912 800 3024 0 FreeSans 560 0 0 0 pbus
port 7 nsew
flabel metal4 s 2346 3076 2666 8684 0 FreeSans 1600 90 0 0 vdd
port 8 nsew
flabel metal4 s 4670 3076 4990 8684 0 FreeSans 1600 90 0 0 vdd
port 8 nsew
flabel metal4 s 6994 3076 7314 8684 0 FreeSans 1600 90 0 0 vdd
port 8 nsew
flabel metal4 s 9318 3076 9638 8684 0 FreeSans 1600 90 0 0 vdd
port 8 nsew
flabel metal4 s 3508 3076 3828 8684 0 FreeSans 1600 90 0 0 vss
port 9 nsew
flabel metal4 s 5832 3076 6152 8684 0 FreeSans 1600 90 0 0 vss
port 9 nsew
flabel metal4 s 8156 3076 8476 8684 0 FreeSans 1600 90 0 0 vss
port 9 nsew
flabel metal4 s 10480 3076 10800 8684 0 FreeSans 1600 90 0 0 vss
port 9 nsew
<< end >>