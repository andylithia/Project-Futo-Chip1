magic
tech gf180mcuC
magscale 1 10
timestamp 1669527744
<< metal2 >>
rect 389215 -12925 389565 -12893
rect 390274 -12925 391918 -12893
rect 392622 -12925 394266 -12893
rect 394971 -12925 396615 -12893
rect 397318 -12925 398962 -12893
rect 399733 -12925 400067 -12893
rect 387840 -13041 401440 -12925
rect 387840 -13097 387986 -13041
rect 388042 -13097 388110 -13041
rect 388166 -13097 388234 -13041
rect 388290 -13097 388358 -13041
rect 388414 -13097 388482 -13041
rect 388538 -13097 388606 -13041
rect 388662 -13097 388730 -13041
rect 388786 -13097 388854 -13041
rect 388910 -13097 388978 -13041
rect 389034 -13097 389102 -13041
rect 389158 -13097 389226 -13041
rect 389282 -13097 389350 -13041
rect 389406 -13097 389474 -13041
rect 389530 -13097 389598 -13041
rect 389654 -13097 389722 -13041
rect 389778 -13097 389846 -13041
rect 389902 -13097 389970 -13041
rect 390026 -13097 390094 -13041
rect 390150 -13097 390218 -13041
rect 390274 -13097 390342 -13041
rect 390398 -13097 390466 -13041
rect 390522 -13097 390590 -13041
rect 390646 -13097 390714 -13041
rect 390770 -13097 390838 -13041
rect 390894 -13097 390962 -13041
rect 391018 -13097 391086 -13041
rect 391142 -13097 391210 -13041
rect 391266 -13097 391334 -13041
rect 391390 -13097 391458 -13041
rect 391514 -13097 391582 -13041
rect 391638 -13097 391706 -13041
rect 391762 -13097 391830 -13041
rect 391886 -13097 391954 -13041
rect 392010 -13097 392078 -13041
rect 392134 -13097 392202 -13041
rect 392258 -13097 392326 -13041
rect 392382 -13097 392450 -13041
rect 392506 -13097 392574 -13041
rect 392630 -13097 392698 -13041
rect 392754 -13097 392822 -13041
rect 392878 -13097 392946 -13041
rect 393002 -13097 393070 -13041
rect 393126 -13097 393194 -13041
rect 393250 -13097 393318 -13041
rect 393374 -13097 393442 -13041
rect 393498 -13097 393566 -13041
rect 393622 -13097 393690 -13041
rect 393746 -13097 393814 -13041
rect 393870 -13097 393938 -13041
rect 393994 -13097 394062 -13041
rect 394118 -13097 394186 -13041
rect 394242 -13097 394310 -13041
rect 394366 -13097 394434 -13041
rect 394490 -13097 394558 -13041
rect 394614 -13097 394682 -13041
rect 394738 -13097 394806 -13041
rect 394862 -13097 394930 -13041
rect 394986 -13097 395054 -13041
rect 395110 -13097 395178 -13041
rect 395234 -13097 395302 -13041
rect 395358 -13097 395426 -13041
rect 395482 -13097 395550 -13041
rect 395606 -13097 395674 -13041
rect 395730 -13097 395798 -13041
rect 395854 -13097 395922 -13041
rect 395978 -13097 396046 -13041
rect 396102 -13097 396170 -13041
rect 396226 -13097 396294 -13041
rect 396350 -13097 396418 -13041
rect 396474 -13097 396542 -13041
rect 396598 -13097 396666 -13041
rect 396722 -13097 396790 -13041
rect 396846 -13097 396914 -13041
rect 396970 -13097 397038 -13041
rect 397094 -13097 397162 -13041
rect 397218 -13097 397286 -13041
rect 397342 -13097 397410 -13041
rect 397466 -13097 397534 -13041
rect 397590 -13097 397658 -13041
rect 397714 -13097 397782 -13041
rect 397838 -13097 397906 -13041
rect 397962 -13097 398030 -13041
rect 398086 -13097 398154 -13041
rect 398210 -13097 398278 -13041
rect 398334 -13097 398402 -13041
rect 398458 -13097 398526 -13041
rect 398582 -13097 398650 -13041
rect 398706 -13097 398774 -13041
rect 398830 -13097 398898 -13041
rect 398954 -13097 399022 -13041
rect 399078 -13097 399146 -13041
rect 399202 -13097 399270 -13041
rect 399326 -13097 399394 -13041
rect 399450 -13097 399518 -13041
rect 399574 -13097 399642 -13041
rect 399698 -13097 399766 -13041
rect 399822 -13097 399890 -13041
rect 399946 -13097 400014 -13041
rect 400070 -13097 400138 -13041
rect 400194 -13097 400262 -13041
rect 400318 -13097 400386 -13041
rect 400442 -13097 400510 -13041
rect 400566 -13097 400634 -13041
rect 400690 -13097 400758 -13041
rect 400814 -13097 400882 -13041
rect 400938 -13097 401006 -13041
rect 401062 -13097 401130 -13041
rect 401186 -13097 401254 -13041
rect 401310 -13097 401440 -13041
rect 387840 -13165 401440 -13097
rect 387840 -13221 387986 -13165
rect 388042 -13221 388110 -13165
rect 388166 -13221 388234 -13165
rect 388290 -13221 388358 -13165
rect 388414 -13221 388482 -13165
rect 388538 -13221 388606 -13165
rect 388662 -13221 388730 -13165
rect 388786 -13221 388854 -13165
rect 388910 -13221 388978 -13165
rect 389034 -13221 389102 -13165
rect 389158 -13221 389226 -13165
rect 389282 -13221 389350 -13165
rect 389406 -13221 389474 -13165
rect 389530 -13221 389598 -13165
rect 389654 -13221 389722 -13165
rect 389778 -13221 389846 -13165
rect 389902 -13221 389970 -13165
rect 390026 -13221 390094 -13165
rect 390150 -13221 390218 -13165
rect 390274 -13221 390342 -13165
rect 390398 -13221 390466 -13165
rect 390522 -13221 390590 -13165
rect 390646 -13221 390714 -13165
rect 390770 -13221 390838 -13165
rect 390894 -13221 390962 -13165
rect 391018 -13221 391086 -13165
rect 391142 -13221 391210 -13165
rect 391266 -13221 391334 -13165
rect 391390 -13221 391458 -13165
rect 391514 -13221 391582 -13165
rect 391638 -13221 391706 -13165
rect 391762 -13221 391830 -13165
rect 391886 -13221 391954 -13165
rect 392010 -13221 392078 -13165
rect 392134 -13221 392202 -13165
rect 392258 -13221 392326 -13165
rect 392382 -13221 392450 -13165
rect 392506 -13221 392574 -13165
rect 392630 -13221 392698 -13165
rect 392754 -13221 392822 -13165
rect 392878 -13221 392946 -13165
rect 393002 -13221 393070 -13165
rect 393126 -13221 393194 -13165
rect 393250 -13221 393318 -13165
rect 393374 -13221 393442 -13165
rect 393498 -13221 393566 -13165
rect 393622 -13221 393690 -13165
rect 393746 -13221 393814 -13165
rect 393870 -13221 393938 -13165
rect 393994 -13221 394062 -13165
rect 394118 -13221 394186 -13165
rect 394242 -13221 394310 -13165
rect 394366 -13221 394434 -13165
rect 394490 -13221 394558 -13165
rect 394614 -13221 394682 -13165
rect 394738 -13221 394806 -13165
rect 394862 -13221 394930 -13165
rect 394986 -13221 395054 -13165
rect 395110 -13221 395178 -13165
rect 395234 -13221 395302 -13165
rect 395358 -13221 395426 -13165
rect 395482 -13221 395550 -13165
rect 395606 -13221 395674 -13165
rect 395730 -13221 395798 -13165
rect 395854 -13221 395922 -13165
rect 395978 -13221 396046 -13165
rect 396102 -13221 396170 -13165
rect 396226 -13221 396294 -13165
rect 396350 -13221 396418 -13165
rect 396474 -13221 396542 -13165
rect 396598 -13221 396666 -13165
rect 396722 -13221 396790 -13165
rect 396846 -13221 396914 -13165
rect 396970 -13221 397038 -13165
rect 397094 -13221 397162 -13165
rect 397218 -13221 397286 -13165
rect 397342 -13221 397410 -13165
rect 397466 -13221 397534 -13165
rect 397590 -13221 397658 -13165
rect 397714 -13221 397782 -13165
rect 397838 -13221 397906 -13165
rect 397962 -13221 398030 -13165
rect 398086 -13221 398154 -13165
rect 398210 -13221 398278 -13165
rect 398334 -13221 398402 -13165
rect 398458 -13221 398526 -13165
rect 398582 -13221 398650 -13165
rect 398706 -13221 398774 -13165
rect 398830 -13221 398898 -13165
rect 398954 -13221 399022 -13165
rect 399078 -13221 399146 -13165
rect 399202 -13221 399270 -13165
rect 399326 -13221 399394 -13165
rect 399450 -13221 399518 -13165
rect 399574 -13221 399642 -13165
rect 399698 -13221 399766 -13165
rect 399822 -13221 399890 -13165
rect 399946 -13221 400014 -13165
rect 400070 -13221 400138 -13165
rect 400194 -13221 400262 -13165
rect 400318 -13221 400386 -13165
rect 400442 -13221 400510 -13165
rect 400566 -13221 400634 -13165
rect 400690 -13221 400758 -13165
rect 400814 -13221 400882 -13165
rect 400938 -13221 401006 -13165
rect 401062 -13221 401130 -13165
rect 401186 -13221 401254 -13165
rect 401310 -13221 401440 -13165
rect 387840 -13289 401440 -13221
rect 387840 -13345 387986 -13289
rect 388042 -13345 388110 -13289
rect 388166 -13345 388234 -13289
rect 388290 -13345 388358 -13289
rect 388414 -13345 388482 -13289
rect 388538 -13345 388606 -13289
rect 388662 -13345 388730 -13289
rect 388786 -13345 388854 -13289
rect 388910 -13345 388978 -13289
rect 389034 -13345 389102 -13289
rect 389158 -13345 389226 -13289
rect 389282 -13345 389350 -13289
rect 389406 -13345 389474 -13289
rect 389530 -13345 389598 -13289
rect 389654 -13345 389722 -13289
rect 389778 -13345 389846 -13289
rect 389902 -13345 389970 -13289
rect 390026 -13345 390094 -13289
rect 390150 -13345 390218 -13289
rect 390274 -13345 390342 -13289
rect 390398 -13345 390466 -13289
rect 390522 -13345 390590 -13289
rect 390646 -13345 390714 -13289
rect 390770 -13345 390838 -13289
rect 390894 -13345 390962 -13289
rect 391018 -13345 391086 -13289
rect 391142 -13345 391210 -13289
rect 391266 -13345 391334 -13289
rect 391390 -13345 391458 -13289
rect 391514 -13345 391582 -13289
rect 391638 -13345 391706 -13289
rect 391762 -13345 391830 -13289
rect 391886 -13345 391954 -13289
rect 392010 -13345 392078 -13289
rect 392134 -13345 392202 -13289
rect 392258 -13345 392326 -13289
rect 392382 -13345 392450 -13289
rect 392506 -13345 392574 -13289
rect 392630 -13345 392698 -13289
rect 392754 -13345 392822 -13289
rect 392878 -13345 392946 -13289
rect 393002 -13345 393070 -13289
rect 393126 -13345 393194 -13289
rect 393250 -13345 393318 -13289
rect 393374 -13345 393442 -13289
rect 393498 -13345 393566 -13289
rect 393622 -13345 393690 -13289
rect 393746 -13345 393814 -13289
rect 393870 -13345 393938 -13289
rect 393994 -13345 394062 -13289
rect 394118 -13345 394186 -13289
rect 394242 -13345 394310 -13289
rect 394366 -13345 394434 -13289
rect 394490 -13345 394558 -13289
rect 394614 -13345 394682 -13289
rect 394738 -13345 394806 -13289
rect 394862 -13345 394930 -13289
rect 394986 -13345 395054 -13289
rect 395110 -13345 395178 -13289
rect 395234 -13345 395302 -13289
rect 395358 -13345 395426 -13289
rect 395482 -13345 395550 -13289
rect 395606 -13345 395674 -13289
rect 395730 -13345 395798 -13289
rect 395854 -13345 395922 -13289
rect 395978 -13345 396046 -13289
rect 396102 -13345 396170 -13289
rect 396226 -13345 396294 -13289
rect 396350 -13345 396418 -13289
rect 396474 -13345 396542 -13289
rect 396598 -13345 396666 -13289
rect 396722 -13345 396790 -13289
rect 396846 -13345 396914 -13289
rect 396970 -13345 397038 -13289
rect 397094 -13345 397162 -13289
rect 397218 -13345 397286 -13289
rect 397342 -13345 397410 -13289
rect 397466 -13345 397534 -13289
rect 397590 -13345 397658 -13289
rect 397714 -13345 397782 -13289
rect 397838 -13345 397906 -13289
rect 397962 -13345 398030 -13289
rect 398086 -13345 398154 -13289
rect 398210 -13345 398278 -13289
rect 398334 -13345 398402 -13289
rect 398458 -13345 398526 -13289
rect 398582 -13345 398650 -13289
rect 398706 -13345 398774 -13289
rect 398830 -13345 398898 -13289
rect 398954 -13345 399022 -13289
rect 399078 -13345 399146 -13289
rect 399202 -13345 399270 -13289
rect 399326 -13345 399394 -13289
rect 399450 -13345 399518 -13289
rect 399574 -13345 399642 -13289
rect 399698 -13345 399766 -13289
rect 399822 -13345 399890 -13289
rect 399946 -13345 400014 -13289
rect 400070 -13345 400138 -13289
rect 400194 -13345 400262 -13289
rect 400318 -13345 400386 -13289
rect 400442 -13345 400510 -13289
rect 400566 -13345 400634 -13289
rect 400690 -13345 400758 -13289
rect 400814 -13345 400882 -13289
rect 400938 -13345 401006 -13289
rect 401062 -13345 401130 -13289
rect 401186 -13345 401254 -13289
rect 401310 -13345 401440 -13289
rect 387840 -13413 401440 -13345
rect 387840 -13469 387986 -13413
rect 388042 -13469 388110 -13413
rect 388166 -13469 388234 -13413
rect 388290 -13469 388358 -13413
rect 388414 -13469 388482 -13413
rect 388538 -13469 388606 -13413
rect 388662 -13469 388730 -13413
rect 388786 -13469 388854 -13413
rect 388910 -13469 388978 -13413
rect 389034 -13469 389102 -13413
rect 389158 -13469 389226 -13413
rect 389282 -13469 389350 -13413
rect 389406 -13469 389474 -13413
rect 389530 -13469 389598 -13413
rect 389654 -13469 389722 -13413
rect 389778 -13469 389846 -13413
rect 389902 -13469 389970 -13413
rect 390026 -13469 390094 -13413
rect 390150 -13469 390218 -13413
rect 390274 -13469 390342 -13413
rect 390398 -13469 390466 -13413
rect 390522 -13469 390590 -13413
rect 390646 -13469 390714 -13413
rect 390770 -13469 390838 -13413
rect 390894 -13469 390962 -13413
rect 391018 -13469 391086 -13413
rect 391142 -13469 391210 -13413
rect 391266 -13469 391334 -13413
rect 391390 -13469 391458 -13413
rect 391514 -13469 391582 -13413
rect 391638 -13469 391706 -13413
rect 391762 -13469 391830 -13413
rect 391886 -13469 391954 -13413
rect 392010 -13469 392078 -13413
rect 392134 -13469 392202 -13413
rect 392258 -13469 392326 -13413
rect 392382 -13469 392450 -13413
rect 392506 -13469 392574 -13413
rect 392630 -13469 392698 -13413
rect 392754 -13469 392822 -13413
rect 392878 -13469 392946 -13413
rect 393002 -13469 393070 -13413
rect 393126 -13469 393194 -13413
rect 393250 -13469 393318 -13413
rect 393374 -13469 393442 -13413
rect 393498 -13469 393566 -13413
rect 393622 -13469 393690 -13413
rect 393746 -13469 393814 -13413
rect 393870 -13469 393938 -13413
rect 393994 -13469 394062 -13413
rect 394118 -13469 394186 -13413
rect 394242 -13469 394310 -13413
rect 394366 -13469 394434 -13413
rect 394490 -13469 394558 -13413
rect 394614 -13469 394682 -13413
rect 394738 -13469 394806 -13413
rect 394862 -13469 394930 -13413
rect 394986 -13469 395054 -13413
rect 395110 -13469 395178 -13413
rect 395234 -13469 395302 -13413
rect 395358 -13469 395426 -13413
rect 395482 -13469 395550 -13413
rect 395606 -13469 395674 -13413
rect 395730 -13469 395798 -13413
rect 395854 -13469 395922 -13413
rect 395978 -13469 396046 -13413
rect 396102 -13469 396170 -13413
rect 396226 -13469 396294 -13413
rect 396350 -13469 396418 -13413
rect 396474 -13469 396542 -13413
rect 396598 -13469 396666 -13413
rect 396722 -13469 396790 -13413
rect 396846 -13469 396914 -13413
rect 396970 -13469 397038 -13413
rect 397094 -13469 397162 -13413
rect 397218 -13469 397286 -13413
rect 397342 -13469 397410 -13413
rect 397466 -13469 397534 -13413
rect 397590 -13469 397658 -13413
rect 397714 -13469 397782 -13413
rect 397838 -13469 397906 -13413
rect 397962 -13469 398030 -13413
rect 398086 -13469 398154 -13413
rect 398210 -13469 398278 -13413
rect 398334 -13469 398402 -13413
rect 398458 -13469 398526 -13413
rect 398582 -13469 398650 -13413
rect 398706 -13469 398774 -13413
rect 398830 -13469 398898 -13413
rect 398954 -13469 399022 -13413
rect 399078 -13469 399146 -13413
rect 399202 -13469 399270 -13413
rect 399326 -13469 399394 -13413
rect 399450 -13469 399518 -13413
rect 399574 -13469 399642 -13413
rect 399698 -13469 399766 -13413
rect 399822 -13469 399890 -13413
rect 399946 -13469 400014 -13413
rect 400070 -13469 400138 -13413
rect 400194 -13469 400262 -13413
rect 400318 -13469 400386 -13413
rect 400442 -13469 400510 -13413
rect 400566 -13469 400634 -13413
rect 400690 -13469 400758 -13413
rect 400814 -13469 400882 -13413
rect 400938 -13469 401006 -13413
rect 401062 -13469 401130 -13413
rect 401186 -13469 401254 -13413
rect 401310 -13469 401440 -13413
rect 387840 -13590 401440 -13469
rect 387840 -13632 388640 -13590
rect 387840 -13688 387954 -13632
rect 388010 -13688 388078 -13632
rect 388134 -13688 388202 -13632
rect 388258 -13688 388326 -13632
rect 388382 -13688 388450 -13632
rect 388506 -13688 388640 -13632
rect 387840 -13756 388640 -13688
rect 387840 -13812 387954 -13756
rect 388010 -13812 388078 -13756
rect 388134 -13812 388202 -13756
rect 388258 -13812 388326 -13756
rect 388382 -13812 388450 -13756
rect 388506 -13812 388640 -13756
rect 387840 -13880 388640 -13812
rect 387840 -13936 387954 -13880
rect 388010 -13936 388078 -13880
rect 388134 -13936 388202 -13880
rect 388258 -13936 388326 -13880
rect 388382 -13936 388450 -13880
rect 388506 -13936 388640 -13880
rect 387840 -14004 388640 -13936
rect 387840 -14060 387954 -14004
rect 388010 -14060 388078 -14004
rect 388134 -14060 388202 -14004
rect 388258 -14060 388326 -14004
rect 388382 -14060 388450 -14004
rect 388506 -14060 388640 -14004
rect 387840 -14128 388640 -14060
rect 387840 -14184 387954 -14128
rect 388010 -14184 388078 -14128
rect 388134 -14184 388202 -14128
rect 388258 -14184 388326 -14128
rect 388382 -14184 388450 -14128
rect 388506 -14184 388640 -14128
rect 387840 -14252 388640 -14184
rect 387840 -14308 387954 -14252
rect 388010 -14308 388078 -14252
rect 388134 -14308 388202 -14252
rect 388258 -14308 388326 -14252
rect 388382 -14308 388450 -14252
rect 388506 -14308 388640 -14252
rect 387840 -14376 388640 -14308
rect 387840 -14432 387954 -14376
rect 388010 -14432 388078 -14376
rect 388134 -14432 388202 -14376
rect 388258 -14432 388326 -14376
rect 388382 -14432 388450 -14376
rect 388506 -14432 388640 -14376
rect 387840 -14500 388640 -14432
rect 387840 -14556 387954 -14500
rect 388010 -14556 388078 -14500
rect 388134 -14556 388202 -14500
rect 388258 -14556 388326 -14500
rect 388382 -14556 388450 -14500
rect 388506 -14556 388640 -14500
rect 387840 -14624 388640 -14556
rect 387840 -14680 387954 -14624
rect 388010 -14680 388078 -14624
rect 388134 -14680 388202 -14624
rect 388258 -14680 388326 -14624
rect 388382 -14680 388450 -14624
rect 388506 -14680 388640 -14624
rect 387840 -14748 388640 -14680
rect 387840 -14804 387954 -14748
rect 388010 -14804 388078 -14748
rect 388134 -14804 388202 -14748
rect 388258 -14804 388326 -14748
rect 388382 -14804 388450 -14748
rect 388506 -14804 388640 -14748
rect 387840 -14872 388640 -14804
rect 387840 -14928 387954 -14872
rect 388010 -14928 388078 -14872
rect 388134 -14928 388202 -14872
rect 388258 -14928 388326 -14872
rect 388382 -14928 388450 -14872
rect 388506 -14928 388640 -14872
rect 387840 -14996 388640 -14928
rect 387840 -15052 387954 -14996
rect 388010 -15052 388078 -14996
rect 388134 -15052 388202 -14996
rect 388258 -15052 388326 -14996
rect 388382 -15052 388450 -14996
rect 388506 -15052 388640 -14996
rect 387840 -15120 388640 -15052
rect 387840 -15176 387954 -15120
rect 388010 -15176 388078 -15120
rect 388134 -15176 388202 -15120
rect 388258 -15176 388326 -15120
rect 388382 -15176 388450 -15120
rect 388506 -15176 388640 -15120
rect 387840 -15244 388640 -15176
rect 387840 -15300 387954 -15244
rect 388010 -15300 388078 -15244
rect 388134 -15300 388202 -15244
rect 388258 -15300 388326 -15244
rect 388382 -15300 388450 -15244
rect 388506 -15300 388640 -15244
rect 387840 -15368 388640 -15300
rect 387840 -15424 387954 -15368
rect 388010 -15424 388078 -15368
rect 388134 -15424 388202 -15368
rect 388258 -15424 388326 -15368
rect 388382 -15424 388450 -15368
rect 388506 -15424 388640 -15368
rect 387840 -15492 388640 -15424
rect 387840 -15548 387954 -15492
rect 388010 -15548 388078 -15492
rect 388134 -15548 388202 -15492
rect 388258 -15548 388326 -15492
rect 388382 -15548 388450 -15492
rect 388506 -15548 388640 -15492
rect 387840 -15616 388640 -15548
rect 387840 -15672 387954 -15616
rect 388010 -15672 388078 -15616
rect 388134 -15672 388202 -15616
rect 388258 -15672 388326 -15616
rect 388382 -15672 388450 -15616
rect 388506 -15672 388640 -15616
rect 387840 -15740 388640 -15672
rect 387840 -15796 387954 -15740
rect 388010 -15796 388078 -15740
rect 388134 -15796 388202 -15740
rect 388258 -15796 388326 -15740
rect 388382 -15796 388450 -15740
rect 388506 -15796 388640 -15740
rect 387840 -15864 388640 -15796
rect 387840 -15920 387954 -15864
rect 388010 -15920 388078 -15864
rect 388134 -15920 388202 -15864
rect 388258 -15920 388326 -15864
rect 388382 -15920 388450 -15864
rect 388506 -15920 388640 -15864
rect 387840 -15988 388640 -15920
rect 387840 -16044 387954 -15988
rect 388010 -16044 388078 -15988
rect 388134 -16044 388202 -15988
rect 388258 -16044 388326 -15988
rect 388382 -16044 388450 -15988
rect 388506 -16044 388640 -15988
rect 387840 -16112 388640 -16044
rect 387840 -16168 387954 -16112
rect 388010 -16168 388078 -16112
rect 388134 -16168 388202 -16112
rect 388258 -16168 388326 -16112
rect 388382 -16168 388450 -16112
rect 388506 -16168 388640 -16112
rect 387840 -16236 388640 -16168
rect 387840 -16292 387954 -16236
rect 388010 -16292 388078 -16236
rect 388134 -16292 388202 -16236
rect 388258 -16292 388326 -16236
rect 388382 -16292 388450 -16236
rect 388506 -16292 388640 -16236
rect 387840 -16360 388640 -16292
rect 387840 -16416 387954 -16360
rect 388010 -16416 388078 -16360
rect 388134 -16416 388202 -16360
rect 388258 -16416 388326 -16360
rect 388382 -16416 388450 -16360
rect 388506 -16416 388640 -16360
rect 387840 -16484 388640 -16416
rect 387840 -16540 387954 -16484
rect 388010 -16540 388078 -16484
rect 388134 -16540 388202 -16484
rect 388258 -16540 388326 -16484
rect 388382 -16540 388450 -16484
rect 388506 -16540 388640 -16484
rect 387840 -16608 388640 -16540
rect 387840 -16664 387954 -16608
rect 388010 -16664 388078 -16608
rect 388134 -16664 388202 -16608
rect 388258 -16664 388326 -16608
rect 388382 -16664 388450 -16608
rect 388506 -16664 388640 -16608
rect 387840 -16732 388640 -16664
rect 387840 -16788 387954 -16732
rect 388010 -16788 388078 -16732
rect 388134 -16788 388202 -16732
rect 388258 -16788 388326 -16732
rect 388382 -16788 388450 -16732
rect 388506 -16788 388640 -16732
rect 387840 -16856 388640 -16788
rect 387840 -16912 387954 -16856
rect 388010 -16912 388078 -16856
rect 388134 -16912 388202 -16856
rect 388258 -16912 388326 -16856
rect 388382 -16912 388450 -16856
rect 388506 -16912 388640 -16856
rect 387840 -16980 388640 -16912
rect 387840 -17036 387954 -16980
rect 388010 -17036 388078 -16980
rect 388134 -17036 388202 -16980
rect 388258 -17036 388326 -16980
rect 388382 -17036 388450 -16980
rect 388506 -17036 388640 -16980
rect 387840 -17104 388640 -17036
rect 387840 -17160 387954 -17104
rect 388010 -17160 388078 -17104
rect 388134 -17160 388202 -17104
rect 388258 -17160 388326 -17104
rect 388382 -17160 388450 -17104
rect 388506 -17160 388640 -17104
rect 387840 -17228 388640 -17160
rect 387840 -17284 387954 -17228
rect 388010 -17284 388078 -17228
rect 388134 -17284 388202 -17228
rect 388258 -17284 388326 -17228
rect 388382 -17284 388450 -17228
rect 388506 -17284 388640 -17228
rect 387840 -17352 388640 -17284
rect 387840 -17408 387954 -17352
rect 388010 -17408 388078 -17352
rect 388134 -17408 388202 -17352
rect 388258 -17408 388326 -17352
rect 388382 -17408 388450 -17352
rect 388506 -17408 388640 -17352
rect 387840 -17476 388640 -17408
rect 387840 -17532 387954 -17476
rect 388010 -17532 388078 -17476
rect 388134 -17532 388202 -17476
rect 388258 -17532 388326 -17476
rect 388382 -17532 388450 -17476
rect 388506 -17532 388640 -17476
rect 387840 -17600 388640 -17532
rect 387840 -17656 387954 -17600
rect 388010 -17656 388078 -17600
rect 388134 -17656 388202 -17600
rect 388258 -17656 388326 -17600
rect 388382 -17656 388450 -17600
rect 388506 -17656 388640 -17600
rect 387840 -17724 388640 -17656
rect 387840 -17780 387954 -17724
rect 388010 -17780 388078 -17724
rect 388134 -17780 388202 -17724
rect 388258 -17780 388326 -17724
rect 388382 -17780 388450 -17724
rect 388506 -17780 388640 -17724
rect 387840 -17848 388640 -17780
rect 387840 -17904 387954 -17848
rect 388010 -17904 388078 -17848
rect 388134 -17904 388202 -17848
rect 388258 -17904 388326 -17848
rect 388382 -17904 388450 -17848
rect 388506 -17904 388640 -17848
rect 387840 -17972 388640 -17904
rect 387840 -18028 387954 -17972
rect 388010 -18028 388078 -17972
rect 388134 -18028 388202 -17972
rect 388258 -18028 388326 -17972
rect 388382 -18028 388450 -17972
rect 388506 -18028 388640 -17972
rect 387840 -18096 388640 -18028
rect 387840 -18152 387954 -18096
rect 388010 -18152 388078 -18096
rect 388134 -18152 388202 -18096
rect 388258 -18152 388326 -18096
rect 388382 -18152 388450 -18096
rect 388506 -18152 388640 -18096
rect 387840 -18220 388640 -18152
rect 387840 -18276 387954 -18220
rect 388010 -18276 388078 -18220
rect 388134 -18276 388202 -18220
rect 388258 -18276 388326 -18220
rect 388382 -18276 388450 -18220
rect 388506 -18276 388640 -18220
rect 387840 -18344 388640 -18276
rect 387840 -18400 387954 -18344
rect 388010 -18400 388078 -18344
rect 388134 -18400 388202 -18344
rect 388258 -18400 388326 -18344
rect 388382 -18400 388450 -18344
rect 388506 -18400 388640 -18344
rect 387840 -18468 388640 -18400
rect 387840 -18524 387954 -18468
rect 388010 -18524 388078 -18468
rect 388134 -18524 388202 -18468
rect 388258 -18524 388326 -18468
rect 388382 -18524 388450 -18468
rect 388506 -18524 388640 -18468
rect 387840 -18592 388640 -18524
rect 387840 -18648 387954 -18592
rect 388010 -18648 388078 -18592
rect 388134 -18648 388202 -18592
rect 388258 -18648 388326 -18592
rect 388382 -18648 388450 -18592
rect 388506 -18648 388640 -18592
rect 387840 -18716 388640 -18648
rect 387840 -18772 387954 -18716
rect 388010 -18772 388078 -18716
rect 388134 -18772 388202 -18716
rect 388258 -18772 388326 -18716
rect 388382 -18772 388450 -18716
rect 388506 -18772 388640 -18716
rect 387840 -18840 388640 -18772
rect 387840 -18896 387954 -18840
rect 388010 -18896 388078 -18840
rect 388134 -18896 388202 -18840
rect 388258 -18896 388326 -18840
rect 388382 -18896 388450 -18840
rect 388506 -18896 388640 -18840
rect 387840 -18964 388640 -18896
rect 387840 -19020 387954 -18964
rect 388010 -19020 388078 -18964
rect 388134 -19020 388202 -18964
rect 388258 -19020 388326 -18964
rect 388382 -19020 388450 -18964
rect 388506 -19020 388640 -18964
rect 387840 -19088 388640 -19020
rect 387840 -19144 387954 -19088
rect 388010 -19144 388078 -19088
rect 388134 -19144 388202 -19088
rect 388258 -19144 388326 -19088
rect 388382 -19144 388450 -19088
rect 388506 -19144 388640 -19088
rect 387840 -19212 388640 -19144
rect 387840 -19268 387954 -19212
rect 388010 -19268 388078 -19212
rect 388134 -19268 388202 -19212
rect 388258 -19268 388326 -19212
rect 388382 -19268 388450 -19212
rect 388506 -19268 388640 -19212
rect 387840 -19336 388640 -19268
rect 387840 -19392 387954 -19336
rect 388010 -19392 388078 -19336
rect 388134 -19392 388202 -19336
rect 388258 -19392 388326 -19336
rect 388382 -19392 388450 -19336
rect 388506 -19392 388640 -19336
rect 387840 -19460 388640 -19392
rect 387840 -19516 387954 -19460
rect 388010 -19516 388078 -19460
rect 388134 -19516 388202 -19460
rect 388258 -19516 388326 -19460
rect 388382 -19516 388450 -19460
rect 388506 -19516 388640 -19460
rect 387840 -19584 388640 -19516
rect 387840 -19640 387954 -19584
rect 388010 -19640 388078 -19584
rect 388134 -19640 388202 -19584
rect 388258 -19640 388326 -19584
rect 388382 -19640 388450 -19584
rect 388506 -19640 388640 -19584
rect 387840 -19708 388640 -19640
rect 387840 -19764 387954 -19708
rect 388010 -19764 388078 -19708
rect 388134 -19764 388202 -19708
rect 388258 -19764 388326 -19708
rect 388382 -19764 388450 -19708
rect 388506 -19764 388640 -19708
rect 387840 -19832 388640 -19764
rect 387840 -19888 387954 -19832
rect 388010 -19888 388078 -19832
rect 388134 -19888 388202 -19832
rect 388258 -19888 388326 -19832
rect 388382 -19888 388450 -19832
rect 388506 -19888 388640 -19832
rect 387840 -19956 388640 -19888
rect 387840 -20012 387954 -19956
rect 388010 -20012 388078 -19956
rect 388134 -20012 388202 -19956
rect 388258 -20012 388326 -19956
rect 388382 -20012 388450 -19956
rect 388506 -20012 388640 -19956
rect 387840 -20080 388640 -20012
rect 387840 -20136 387954 -20080
rect 388010 -20136 388078 -20080
rect 388134 -20136 388202 -20080
rect 388258 -20136 388326 -20080
rect 388382 -20136 388450 -20080
rect 388506 -20136 388640 -20080
rect 387840 -20204 388640 -20136
rect 387840 -20260 387954 -20204
rect 388010 -20260 388078 -20204
rect 388134 -20260 388202 -20204
rect 388258 -20260 388326 -20204
rect 388382 -20260 388450 -20204
rect 388506 -20260 388640 -20204
rect 387840 -20328 388640 -20260
rect 387840 -20384 387954 -20328
rect 388010 -20384 388078 -20328
rect 388134 -20384 388202 -20328
rect 388258 -20384 388326 -20328
rect 388382 -20384 388450 -20328
rect 388506 -20384 388640 -20328
rect 387840 -20452 388640 -20384
rect 387840 -20508 387954 -20452
rect 388010 -20508 388078 -20452
rect 388134 -20508 388202 -20452
rect 388258 -20508 388326 -20452
rect 388382 -20508 388450 -20452
rect 388506 -20508 388640 -20452
rect 387840 -20576 388640 -20508
rect 387840 -20632 387954 -20576
rect 388010 -20632 388078 -20576
rect 388134 -20632 388202 -20576
rect 388258 -20632 388326 -20576
rect 388382 -20632 388450 -20576
rect 388506 -20632 388640 -20576
rect 387840 -20700 388640 -20632
rect 387840 -20756 387954 -20700
rect 388010 -20756 388078 -20700
rect 388134 -20756 388202 -20700
rect 388258 -20756 388326 -20700
rect 388382 -20756 388450 -20700
rect 388506 -20756 388640 -20700
rect 387840 -20824 388640 -20756
rect 387840 -20880 387954 -20824
rect 388010 -20880 388078 -20824
rect 388134 -20880 388202 -20824
rect 388258 -20880 388326 -20824
rect 388382 -20880 388450 -20824
rect 388506 -20880 388640 -20824
rect 387840 -20948 388640 -20880
rect 387840 -21004 387954 -20948
rect 388010 -21004 388078 -20948
rect 388134 -21004 388202 -20948
rect 388258 -21004 388326 -20948
rect 388382 -21004 388450 -20948
rect 388506 -21004 388640 -20948
rect 387840 -21072 388640 -21004
rect 387840 -21128 387954 -21072
rect 388010 -21128 388078 -21072
rect 388134 -21128 388202 -21072
rect 388258 -21128 388326 -21072
rect 388382 -21128 388450 -21072
rect 388506 -21128 388640 -21072
rect 387840 -21196 388640 -21128
rect 387840 -21252 387954 -21196
rect 388010 -21252 388078 -21196
rect 388134 -21252 388202 -21196
rect 388258 -21252 388326 -21196
rect 388382 -21252 388450 -21196
rect 388506 -21252 388640 -21196
rect 387840 -21320 388640 -21252
rect 387840 -21376 387954 -21320
rect 388010 -21376 388078 -21320
rect 388134 -21376 388202 -21320
rect 388258 -21376 388326 -21320
rect 388382 -21376 388450 -21320
rect 388506 -21376 388640 -21320
rect 387840 -21444 388640 -21376
rect 387840 -21500 387954 -21444
rect 388010 -21500 388078 -21444
rect 388134 -21500 388202 -21444
rect 388258 -21500 388326 -21444
rect 388382 -21500 388450 -21444
rect 388506 -21500 388640 -21444
rect 387840 -21568 388640 -21500
rect 387840 -21624 387954 -21568
rect 388010 -21624 388078 -21568
rect 388134 -21624 388202 -21568
rect 388258 -21624 388326 -21568
rect 388382 -21624 388450 -21568
rect 388506 -21624 388640 -21568
rect 387840 -21692 388640 -21624
rect 387840 -21748 387954 -21692
rect 388010 -21748 388078 -21692
rect 388134 -21748 388202 -21692
rect 388258 -21748 388326 -21692
rect 388382 -21748 388450 -21692
rect 388506 -21748 388640 -21692
rect 387840 -21816 388640 -21748
rect 387840 -21872 387954 -21816
rect 388010 -21872 388078 -21816
rect 388134 -21872 388202 -21816
rect 388258 -21872 388326 -21816
rect 388382 -21872 388450 -21816
rect 388506 -21872 388640 -21816
rect 387840 -21940 388640 -21872
rect 387840 -21996 387954 -21940
rect 388010 -21996 388078 -21940
rect 388134 -21996 388202 -21940
rect 388258 -21996 388326 -21940
rect 388382 -21996 388450 -21940
rect 388506 -21996 388640 -21940
rect 387840 -22064 388640 -21996
rect 387840 -22120 387954 -22064
rect 388010 -22120 388078 -22064
rect 388134 -22120 388202 -22064
rect 388258 -22120 388326 -22064
rect 388382 -22120 388450 -22064
rect 388506 -22120 388640 -22064
rect 387840 -22188 388640 -22120
rect 387840 -22244 387954 -22188
rect 388010 -22244 388078 -22188
rect 388134 -22244 388202 -22188
rect 388258 -22244 388326 -22188
rect 388382 -22244 388450 -22188
rect 388506 -22244 388640 -22188
rect 387840 -22312 388640 -22244
rect 387840 -22368 387954 -22312
rect 388010 -22368 388078 -22312
rect 388134 -22368 388202 -22312
rect 388258 -22368 388326 -22312
rect 388382 -22368 388450 -22312
rect 388506 -22368 388640 -22312
rect 387840 -22436 388640 -22368
rect 387840 -22492 387954 -22436
rect 388010 -22492 388078 -22436
rect 388134 -22492 388202 -22436
rect 388258 -22492 388326 -22436
rect 388382 -22492 388450 -22436
rect 388506 -22492 388640 -22436
rect 387840 -22560 388640 -22492
rect 387840 -22616 387954 -22560
rect 388010 -22616 388078 -22560
rect 388134 -22616 388202 -22560
rect 388258 -22616 388326 -22560
rect 388382 -22616 388450 -22560
rect 388506 -22616 388640 -22560
rect 387840 -22684 388640 -22616
rect 387840 -22740 387954 -22684
rect 388010 -22740 388078 -22684
rect 388134 -22740 388202 -22684
rect 388258 -22740 388326 -22684
rect 388382 -22740 388450 -22684
rect 388506 -22740 388640 -22684
rect 387840 -22808 388640 -22740
rect 387840 -22864 387954 -22808
rect 388010 -22864 388078 -22808
rect 388134 -22864 388202 -22808
rect 388258 -22864 388326 -22808
rect 388382 -22864 388450 -22808
rect 388506 -22864 388640 -22808
rect 387840 -22932 388640 -22864
rect 387840 -22988 387954 -22932
rect 388010 -22988 388078 -22932
rect 388134 -22988 388202 -22932
rect 388258 -22988 388326 -22932
rect 388382 -22988 388450 -22932
rect 388506 -22988 388640 -22932
rect 387840 -23056 388640 -22988
rect 387840 -23112 387954 -23056
rect 388010 -23112 388078 -23056
rect 388134 -23112 388202 -23056
rect 388258 -23112 388326 -23056
rect 388382 -23112 388450 -23056
rect 388506 -23112 388640 -23056
rect 387840 -23180 388640 -23112
rect 387840 -23236 387954 -23180
rect 388010 -23236 388078 -23180
rect 388134 -23236 388202 -23180
rect 388258 -23236 388326 -23180
rect 388382 -23236 388450 -23180
rect 388506 -23236 388640 -23180
rect 387840 -23304 388640 -23236
rect 387840 -23360 387954 -23304
rect 388010 -23360 388078 -23304
rect 388134 -23360 388202 -23304
rect 388258 -23360 388326 -23304
rect 388382 -23360 388450 -23304
rect 388506 -23360 388640 -23304
rect 387840 -23428 388640 -23360
rect 387840 -23484 387954 -23428
rect 388010 -23484 388078 -23428
rect 388134 -23484 388202 -23428
rect 388258 -23484 388326 -23428
rect 388382 -23484 388450 -23428
rect 388506 -23484 388640 -23428
rect 387840 -23552 388640 -23484
rect 387840 -23608 387954 -23552
rect 388010 -23608 388078 -23552
rect 388134 -23608 388202 -23552
rect 388258 -23608 388326 -23552
rect 388382 -23608 388450 -23552
rect 388506 -23608 388640 -23552
rect 387840 -23676 388640 -23608
rect 387840 -23732 387954 -23676
rect 388010 -23732 388078 -23676
rect 388134 -23732 388202 -23676
rect 388258 -23732 388326 -23676
rect 388382 -23732 388450 -23676
rect 388506 -23732 388640 -23676
rect 387840 -23800 388640 -23732
rect 387840 -23856 387954 -23800
rect 388010 -23856 388078 -23800
rect 388134 -23856 388202 -23800
rect 388258 -23856 388326 -23800
rect 388382 -23856 388450 -23800
rect 388506 -23856 388640 -23800
rect 387840 -23924 388640 -23856
rect 387840 -23980 387954 -23924
rect 388010 -23980 388078 -23924
rect 388134 -23980 388202 -23924
rect 388258 -23980 388326 -23924
rect 388382 -23980 388450 -23924
rect 388506 -23980 388640 -23924
rect 387840 -24048 388640 -23980
rect 387840 -24104 387954 -24048
rect 388010 -24104 388078 -24048
rect 388134 -24104 388202 -24048
rect 388258 -24104 388326 -24048
rect 388382 -24104 388450 -24048
rect 388506 -24104 388640 -24048
rect 387840 -24172 388640 -24104
rect 387840 -24228 387954 -24172
rect 388010 -24228 388078 -24172
rect 388134 -24228 388202 -24172
rect 388258 -24228 388326 -24172
rect 388382 -24228 388450 -24172
rect 388506 -24228 388640 -24172
rect 387840 -24296 388640 -24228
rect 387840 -24352 387954 -24296
rect 388010 -24352 388078 -24296
rect 388134 -24352 388202 -24296
rect 388258 -24352 388326 -24296
rect 388382 -24352 388450 -24296
rect 388506 -24352 388640 -24296
rect 387840 -24420 388640 -24352
rect 387840 -24476 387954 -24420
rect 388010 -24476 388078 -24420
rect 388134 -24476 388202 -24420
rect 388258 -24476 388326 -24420
rect 388382 -24476 388450 -24420
rect 388506 -24476 388640 -24420
rect 387840 -24544 388640 -24476
rect 387840 -24600 387954 -24544
rect 388010 -24600 388078 -24544
rect 388134 -24600 388202 -24544
rect 388258 -24600 388326 -24544
rect 388382 -24600 388450 -24544
rect 388506 -24600 388640 -24544
rect 387840 -24668 388640 -24600
rect 387840 -24724 387954 -24668
rect 388010 -24724 388078 -24668
rect 388134 -24724 388202 -24668
rect 388258 -24724 388326 -24668
rect 388382 -24724 388450 -24668
rect 388506 -24724 388640 -24668
rect 387840 -24792 388640 -24724
rect 387840 -24848 387954 -24792
rect 388010 -24848 388078 -24792
rect 388134 -24848 388202 -24792
rect 388258 -24848 388326 -24792
rect 388382 -24848 388450 -24792
rect 388506 -24848 388640 -24792
rect 387840 -24916 388640 -24848
rect 387840 -24972 387954 -24916
rect 388010 -24972 388078 -24916
rect 388134 -24972 388202 -24916
rect 388258 -24972 388326 -24916
rect 388382 -24972 388450 -24916
rect 388506 -24972 388640 -24916
rect 387840 -25040 388640 -24972
rect 387840 -25096 387954 -25040
rect 388010 -25096 388078 -25040
rect 388134 -25096 388202 -25040
rect 388258 -25096 388326 -25040
rect 388382 -25096 388450 -25040
rect 388506 -25096 388640 -25040
rect 387840 -25164 388640 -25096
rect 387840 -25220 387954 -25164
rect 388010 -25220 388078 -25164
rect 388134 -25220 388202 -25164
rect 388258 -25220 388326 -25164
rect 388382 -25220 388450 -25164
rect 388506 -25220 388640 -25164
rect 387840 -25288 388640 -25220
rect 387840 -25344 387954 -25288
rect 388010 -25344 388078 -25288
rect 388134 -25344 388202 -25288
rect 388258 -25344 388326 -25288
rect 388382 -25344 388450 -25288
rect 388506 -25344 388640 -25288
rect 387840 -25412 388640 -25344
rect 387840 -25468 387954 -25412
rect 388010 -25468 388078 -25412
rect 388134 -25468 388202 -25412
rect 388258 -25468 388326 -25412
rect 388382 -25468 388450 -25412
rect 388506 -25468 388640 -25412
rect 387840 -25536 388640 -25468
rect 387840 -25592 387954 -25536
rect 388010 -25592 388078 -25536
rect 388134 -25592 388202 -25536
rect 388258 -25592 388326 -25536
rect 388382 -25592 388450 -25536
rect 388506 -25590 388640 -25536
rect 388908 -13680 389248 -13590
rect 388908 -13736 388981 -13680
rect 389037 -13736 389123 -13680
rect 389179 -13736 389248 -13680
rect 388908 -13822 389248 -13736
rect 388908 -13878 388981 -13822
rect 389037 -13878 389123 -13822
rect 389179 -13878 389248 -13822
rect 388908 -13964 389248 -13878
rect 388908 -14020 388981 -13964
rect 389037 -14020 389123 -13964
rect 389179 -14020 389248 -13964
rect 388908 -14106 389248 -14020
rect 388908 -14162 388981 -14106
rect 389037 -14162 389123 -14106
rect 389179 -14162 389248 -14106
rect 388908 -14248 389248 -14162
rect 388908 -14304 388981 -14248
rect 389037 -14304 389123 -14248
rect 389179 -14304 389248 -14248
rect 388908 -14390 389248 -14304
rect 388908 -14446 388981 -14390
rect 389037 -14446 389123 -14390
rect 389179 -14446 389248 -14390
rect 388908 -14532 389248 -14446
rect 388908 -14588 388981 -14532
rect 389037 -14588 389123 -14532
rect 389179 -14588 389248 -14532
rect 388908 -14674 389248 -14588
rect 388908 -14730 388981 -14674
rect 389037 -14730 389123 -14674
rect 389179 -14730 389248 -14674
rect 388908 -14816 389248 -14730
rect 388908 -14872 388981 -14816
rect 389037 -14872 389123 -14816
rect 389179 -14872 389248 -14816
rect 388908 -14958 389248 -14872
rect 388908 -15014 388981 -14958
rect 389037 -15014 389123 -14958
rect 389179 -15014 389248 -14958
rect 388908 -15100 389248 -15014
rect 388908 -15156 388981 -15100
rect 389037 -15156 389123 -15100
rect 389179 -15156 389248 -15100
rect 388908 -15242 389248 -15156
rect 388908 -15298 388981 -15242
rect 389037 -15298 389123 -15242
rect 389179 -15298 389248 -15242
rect 388908 -15384 389248 -15298
rect 388908 -15440 388981 -15384
rect 389037 -15440 389123 -15384
rect 389179 -15440 389248 -15384
rect 388908 -15526 389248 -15440
rect 388908 -15582 388981 -15526
rect 389037 -15582 389123 -15526
rect 389179 -15582 389248 -15526
rect 388908 -15668 389248 -15582
rect 388908 -15724 388981 -15668
rect 389037 -15724 389123 -15668
rect 389179 -15724 389248 -15668
rect 388908 -15810 389248 -15724
rect 388908 -15866 388981 -15810
rect 389037 -15866 389123 -15810
rect 389179 -15866 389248 -15810
rect 388908 -15952 389248 -15866
rect 388908 -16008 388981 -15952
rect 389037 -16008 389123 -15952
rect 389179 -16008 389248 -15952
rect 388908 -16094 389248 -16008
rect 388908 -16150 388981 -16094
rect 389037 -16150 389123 -16094
rect 389179 -16150 389248 -16094
rect 388908 -16236 389248 -16150
rect 388908 -16292 388981 -16236
rect 389037 -16292 389123 -16236
rect 389179 -16292 389248 -16236
rect 388908 -16378 389248 -16292
rect 388908 -16434 388981 -16378
rect 389037 -16434 389123 -16378
rect 389179 -16434 389248 -16378
rect 388908 -16520 389248 -16434
rect 388908 -16576 388981 -16520
rect 389037 -16576 389123 -16520
rect 389179 -16576 389248 -16520
rect 388908 -16662 389248 -16576
rect 388908 -16718 388981 -16662
rect 389037 -16718 389123 -16662
rect 389179 -16718 389248 -16662
rect 388908 -16804 389248 -16718
rect 388908 -16860 388981 -16804
rect 389037 -16860 389123 -16804
rect 389179 -16860 389248 -16804
rect 388908 -16946 389248 -16860
rect 388908 -17002 388981 -16946
rect 389037 -17002 389123 -16946
rect 389179 -17002 389248 -16946
rect 388908 -17088 389248 -17002
rect 388908 -17144 388981 -17088
rect 389037 -17144 389123 -17088
rect 389179 -17144 389248 -17088
rect 388908 -17230 389248 -17144
rect 388908 -17286 388981 -17230
rect 389037 -17286 389123 -17230
rect 389179 -17286 389248 -17230
rect 388908 -17372 389248 -17286
rect 388908 -17428 388981 -17372
rect 389037 -17428 389123 -17372
rect 389179 -17428 389248 -17372
rect 388908 -17514 389248 -17428
rect 388908 -17570 388981 -17514
rect 389037 -17570 389123 -17514
rect 389179 -17570 389248 -17514
rect 388908 -17656 389248 -17570
rect 388908 -17712 388981 -17656
rect 389037 -17712 389123 -17656
rect 389179 -17712 389248 -17656
rect 388908 -17798 389248 -17712
rect 388908 -17854 388981 -17798
rect 389037 -17854 389123 -17798
rect 389179 -17854 389248 -17798
rect 388908 -17940 389248 -17854
rect 388908 -17996 388981 -17940
rect 389037 -17996 389123 -17940
rect 389179 -17996 389248 -17940
rect 388908 -18082 389248 -17996
rect 388908 -18138 388981 -18082
rect 389037 -18138 389123 -18082
rect 389179 -18138 389248 -18082
rect 388908 -18224 389248 -18138
rect 388908 -18280 388981 -18224
rect 389037 -18280 389123 -18224
rect 389179 -18280 389248 -18224
rect 388908 -18366 389248 -18280
rect 388908 -18422 388981 -18366
rect 389037 -18422 389123 -18366
rect 389179 -18422 389248 -18366
rect 388908 -18508 389248 -18422
rect 388908 -18564 388981 -18508
rect 389037 -18564 389123 -18508
rect 389179 -18564 389248 -18508
rect 388908 -18650 389248 -18564
rect 388908 -18706 388981 -18650
rect 389037 -18706 389123 -18650
rect 389179 -18706 389248 -18650
rect 388908 -18792 389248 -18706
rect 388908 -18848 388981 -18792
rect 389037 -18848 389123 -18792
rect 389179 -18848 389248 -18792
rect 388908 -18934 389248 -18848
rect 388908 -18990 388981 -18934
rect 389037 -18990 389123 -18934
rect 389179 -18990 389248 -18934
rect 388908 -19076 389248 -18990
rect 388908 -19132 388981 -19076
rect 389037 -19132 389123 -19076
rect 389179 -19132 389248 -19076
rect 388908 -19218 389248 -19132
rect 388908 -19274 388981 -19218
rect 389037 -19274 389123 -19218
rect 389179 -19274 389248 -19218
rect 388908 -19360 389248 -19274
rect 388908 -19416 388981 -19360
rect 389037 -19416 389123 -19360
rect 389179 -19416 389248 -19360
rect 388908 -19502 389248 -19416
rect 388908 -19558 388981 -19502
rect 389037 -19558 389123 -19502
rect 389179 -19558 389248 -19502
rect 388908 -19644 389248 -19558
rect 388908 -19700 388981 -19644
rect 389037 -19700 389123 -19644
rect 389179 -19700 389248 -19644
rect 388908 -19786 389248 -19700
rect 388908 -19842 388981 -19786
rect 389037 -19842 389123 -19786
rect 389179 -19842 389248 -19786
rect 388908 -19928 389248 -19842
rect 388908 -19984 388981 -19928
rect 389037 -19984 389123 -19928
rect 389179 -19984 389248 -19928
rect 388908 -20070 389248 -19984
rect 388908 -20126 388981 -20070
rect 389037 -20126 389123 -20070
rect 389179 -20126 389248 -20070
rect 388908 -20212 389248 -20126
rect 388908 -20268 388981 -20212
rect 389037 -20268 389123 -20212
rect 389179 -20268 389248 -20212
rect 388908 -20354 389248 -20268
rect 388908 -20410 388981 -20354
rect 389037 -20410 389123 -20354
rect 389179 -20410 389248 -20354
rect 388908 -20496 389248 -20410
rect 388908 -20552 388981 -20496
rect 389037 -20552 389123 -20496
rect 389179 -20552 389248 -20496
rect 388908 -20638 389248 -20552
rect 388908 -20694 388981 -20638
rect 389037 -20694 389123 -20638
rect 389179 -20694 389248 -20638
rect 388908 -20780 389248 -20694
rect 388908 -20836 388981 -20780
rect 389037 -20836 389123 -20780
rect 389179 -20836 389248 -20780
rect 388908 -20922 389248 -20836
rect 388908 -20978 388981 -20922
rect 389037 -20978 389123 -20922
rect 389179 -20978 389248 -20922
rect 388908 -21064 389248 -20978
rect 388908 -21120 388981 -21064
rect 389037 -21120 389123 -21064
rect 389179 -21120 389248 -21064
rect 388908 -21206 389248 -21120
rect 388908 -21262 388981 -21206
rect 389037 -21262 389123 -21206
rect 389179 -21262 389248 -21206
rect 388908 -21348 389248 -21262
rect 388908 -21404 388981 -21348
rect 389037 -21404 389123 -21348
rect 389179 -21404 389248 -21348
rect 388908 -21490 389248 -21404
rect 388908 -21546 388981 -21490
rect 389037 -21546 389123 -21490
rect 389179 -21546 389248 -21490
rect 388908 -21632 389248 -21546
rect 388908 -21688 388981 -21632
rect 389037 -21688 389123 -21632
rect 389179 -21688 389248 -21632
rect 388908 -21774 389248 -21688
rect 388908 -21830 388981 -21774
rect 389037 -21830 389123 -21774
rect 389179 -21830 389248 -21774
rect 388908 -21916 389248 -21830
rect 388908 -21972 388981 -21916
rect 389037 -21972 389123 -21916
rect 389179 -21972 389248 -21916
rect 388908 -22058 389248 -21972
rect 388908 -22114 388981 -22058
rect 389037 -22114 389123 -22058
rect 389179 -22114 389248 -22058
rect 388908 -22200 389248 -22114
rect 388908 -22256 388981 -22200
rect 389037 -22256 389123 -22200
rect 389179 -22256 389248 -22200
rect 388908 -22342 389248 -22256
rect 388908 -22398 388981 -22342
rect 389037 -22398 389123 -22342
rect 389179 -22398 389248 -22342
rect 388908 -22484 389248 -22398
rect 388908 -22540 388981 -22484
rect 389037 -22540 389123 -22484
rect 389179 -22540 389248 -22484
rect 388908 -22626 389248 -22540
rect 388908 -22682 388981 -22626
rect 389037 -22682 389123 -22626
rect 389179 -22682 389248 -22626
rect 388908 -22768 389248 -22682
rect 388908 -22824 388981 -22768
rect 389037 -22824 389123 -22768
rect 389179 -22824 389248 -22768
rect 388908 -22910 389248 -22824
rect 388908 -22966 388981 -22910
rect 389037 -22966 389123 -22910
rect 389179 -22966 389248 -22910
rect 388908 -23052 389248 -22966
rect 388908 -23108 388981 -23052
rect 389037 -23108 389123 -23052
rect 389179 -23108 389248 -23052
rect 388908 -23194 389248 -23108
rect 388908 -23250 388981 -23194
rect 389037 -23250 389123 -23194
rect 389179 -23250 389248 -23194
rect 388908 -23336 389248 -23250
rect 388908 -23392 388981 -23336
rect 389037 -23392 389123 -23336
rect 389179 -23392 389248 -23336
rect 388908 -23478 389248 -23392
rect 388908 -23534 388981 -23478
rect 389037 -23534 389123 -23478
rect 389179 -23534 389248 -23478
rect 388908 -23620 389248 -23534
rect 388908 -23676 388981 -23620
rect 389037 -23676 389123 -23620
rect 389179 -23676 389248 -23620
rect 388908 -23762 389248 -23676
rect 388908 -23818 388981 -23762
rect 389037 -23818 389123 -23762
rect 389179 -23818 389248 -23762
rect 388908 -23904 389248 -23818
rect 388908 -23960 388981 -23904
rect 389037 -23960 389123 -23904
rect 389179 -23960 389248 -23904
rect 388908 -24046 389248 -23960
rect 388908 -24102 388981 -24046
rect 389037 -24102 389123 -24046
rect 389179 -24102 389248 -24046
rect 388908 -24188 389248 -24102
rect 388908 -24244 388981 -24188
rect 389037 -24244 389123 -24188
rect 389179 -24244 389248 -24188
rect 388908 -24330 389248 -24244
rect 388908 -24386 388981 -24330
rect 389037 -24386 389123 -24330
rect 389179 -24386 389248 -24330
rect 388908 -24472 389248 -24386
rect 388908 -24528 388981 -24472
rect 389037 -24528 389123 -24472
rect 389179 -24528 389248 -24472
rect 388908 -24614 389248 -24528
rect 388908 -24670 388981 -24614
rect 389037 -24670 389123 -24614
rect 389179 -24670 389248 -24614
rect 388908 -24756 389248 -24670
rect 388908 -24812 388981 -24756
rect 389037 -24812 389123 -24756
rect 389179 -24812 389248 -24756
rect 388908 -24898 389248 -24812
rect 388908 -24954 388981 -24898
rect 389037 -24954 389123 -24898
rect 389179 -24954 389248 -24898
rect 388908 -25040 389248 -24954
rect 388908 -25096 388981 -25040
rect 389037 -25096 389123 -25040
rect 389179 -25096 389248 -25040
rect 388908 -25182 389248 -25096
rect 388908 -25238 388981 -25182
rect 389037 -25238 389123 -25182
rect 389179 -25238 389248 -25182
rect 388908 -25324 389248 -25238
rect 388908 -25380 388981 -25324
rect 389037 -25380 389123 -25324
rect 389179 -25380 389248 -25324
rect 388908 -25466 389248 -25380
rect 388908 -25522 388981 -25466
rect 389037 -25522 389123 -25466
rect 389179 -25522 389248 -25466
rect 388908 -25590 389248 -25522
rect 389308 -13680 389648 -13590
rect 389308 -13736 389382 -13680
rect 389438 -13736 389524 -13680
rect 389580 -13736 389648 -13680
rect 389308 -13822 389648 -13736
rect 389308 -13878 389382 -13822
rect 389438 -13878 389524 -13822
rect 389580 -13878 389648 -13822
rect 389308 -13964 389648 -13878
rect 389308 -14020 389382 -13964
rect 389438 -14020 389524 -13964
rect 389580 -14020 389648 -13964
rect 389308 -14106 389648 -14020
rect 389308 -14162 389382 -14106
rect 389438 -14162 389524 -14106
rect 389580 -14162 389648 -14106
rect 389308 -14248 389648 -14162
rect 389308 -14304 389382 -14248
rect 389438 -14304 389524 -14248
rect 389580 -14304 389648 -14248
rect 389308 -14390 389648 -14304
rect 389308 -14446 389382 -14390
rect 389438 -14446 389524 -14390
rect 389580 -14446 389648 -14390
rect 389308 -14532 389648 -14446
rect 389308 -14588 389382 -14532
rect 389438 -14588 389524 -14532
rect 389580 -14588 389648 -14532
rect 389308 -14674 389648 -14588
rect 389308 -14730 389382 -14674
rect 389438 -14730 389524 -14674
rect 389580 -14730 389648 -14674
rect 389308 -14816 389648 -14730
rect 389308 -14872 389382 -14816
rect 389438 -14872 389524 -14816
rect 389580 -14872 389648 -14816
rect 389308 -14958 389648 -14872
rect 389308 -15014 389382 -14958
rect 389438 -15014 389524 -14958
rect 389580 -15014 389648 -14958
rect 389308 -15100 389648 -15014
rect 389308 -15156 389382 -15100
rect 389438 -15156 389524 -15100
rect 389580 -15156 389648 -15100
rect 389308 -15242 389648 -15156
rect 389308 -15298 389382 -15242
rect 389438 -15298 389524 -15242
rect 389580 -15298 389648 -15242
rect 389308 -15384 389648 -15298
rect 389308 -15440 389382 -15384
rect 389438 -15440 389524 -15384
rect 389580 -15440 389648 -15384
rect 389308 -15526 389648 -15440
rect 389308 -15582 389382 -15526
rect 389438 -15582 389524 -15526
rect 389580 -15582 389648 -15526
rect 389308 -15668 389648 -15582
rect 389308 -15724 389382 -15668
rect 389438 -15724 389524 -15668
rect 389580 -15724 389648 -15668
rect 389308 -15810 389648 -15724
rect 389308 -15866 389382 -15810
rect 389438 -15866 389524 -15810
rect 389580 -15866 389648 -15810
rect 389308 -15952 389648 -15866
rect 389308 -16008 389382 -15952
rect 389438 -16008 389524 -15952
rect 389580 -16008 389648 -15952
rect 389308 -16094 389648 -16008
rect 389308 -16150 389382 -16094
rect 389438 -16150 389524 -16094
rect 389580 -16150 389648 -16094
rect 389308 -16236 389648 -16150
rect 389308 -16292 389382 -16236
rect 389438 -16292 389524 -16236
rect 389580 -16292 389648 -16236
rect 389308 -16378 389648 -16292
rect 389308 -16434 389382 -16378
rect 389438 -16434 389524 -16378
rect 389580 -16434 389648 -16378
rect 389308 -16520 389648 -16434
rect 389308 -16576 389382 -16520
rect 389438 -16576 389524 -16520
rect 389580 -16576 389648 -16520
rect 389308 -16662 389648 -16576
rect 389308 -16718 389382 -16662
rect 389438 -16718 389524 -16662
rect 389580 -16718 389648 -16662
rect 389308 -16804 389648 -16718
rect 389308 -16860 389382 -16804
rect 389438 -16860 389524 -16804
rect 389580 -16860 389648 -16804
rect 389308 -16946 389648 -16860
rect 389308 -17002 389382 -16946
rect 389438 -17002 389524 -16946
rect 389580 -17002 389648 -16946
rect 389308 -17088 389648 -17002
rect 389308 -17144 389382 -17088
rect 389438 -17144 389524 -17088
rect 389580 -17144 389648 -17088
rect 389308 -17230 389648 -17144
rect 389308 -17286 389382 -17230
rect 389438 -17286 389524 -17230
rect 389580 -17286 389648 -17230
rect 389308 -17372 389648 -17286
rect 389308 -17428 389382 -17372
rect 389438 -17428 389524 -17372
rect 389580 -17428 389648 -17372
rect 389308 -17514 389648 -17428
rect 389308 -17570 389382 -17514
rect 389438 -17570 389524 -17514
rect 389580 -17570 389648 -17514
rect 389308 -17656 389648 -17570
rect 389308 -17712 389382 -17656
rect 389438 -17712 389524 -17656
rect 389580 -17712 389648 -17656
rect 389308 -17798 389648 -17712
rect 389308 -17854 389382 -17798
rect 389438 -17854 389524 -17798
rect 389580 -17854 389648 -17798
rect 389308 -17940 389648 -17854
rect 389308 -17996 389382 -17940
rect 389438 -17996 389524 -17940
rect 389580 -17996 389648 -17940
rect 389308 -18082 389648 -17996
rect 389308 -18138 389382 -18082
rect 389438 -18138 389524 -18082
rect 389580 -18138 389648 -18082
rect 389308 -18224 389648 -18138
rect 389308 -18280 389382 -18224
rect 389438 -18280 389524 -18224
rect 389580 -18280 389648 -18224
rect 389308 -18366 389648 -18280
rect 389308 -18422 389382 -18366
rect 389438 -18422 389524 -18366
rect 389580 -18422 389648 -18366
rect 389308 -18508 389648 -18422
rect 389308 -18564 389382 -18508
rect 389438 -18564 389524 -18508
rect 389580 -18564 389648 -18508
rect 389308 -18650 389648 -18564
rect 389308 -18706 389382 -18650
rect 389438 -18706 389524 -18650
rect 389580 -18706 389648 -18650
rect 389308 -18792 389648 -18706
rect 389308 -18848 389382 -18792
rect 389438 -18848 389524 -18792
rect 389580 -18848 389648 -18792
rect 389308 -18934 389648 -18848
rect 389308 -18990 389382 -18934
rect 389438 -18990 389524 -18934
rect 389580 -18990 389648 -18934
rect 389308 -19076 389648 -18990
rect 389308 -19132 389382 -19076
rect 389438 -19132 389524 -19076
rect 389580 -19132 389648 -19076
rect 389308 -19218 389648 -19132
rect 389308 -19274 389382 -19218
rect 389438 -19274 389524 -19218
rect 389580 -19274 389648 -19218
rect 389308 -19360 389648 -19274
rect 389308 -19416 389382 -19360
rect 389438 -19416 389524 -19360
rect 389580 -19416 389648 -19360
rect 389308 -19502 389648 -19416
rect 389308 -19558 389382 -19502
rect 389438 -19558 389524 -19502
rect 389580 -19558 389648 -19502
rect 389308 -19644 389648 -19558
rect 389308 -19700 389382 -19644
rect 389438 -19700 389524 -19644
rect 389580 -19700 389648 -19644
rect 389308 -19786 389648 -19700
rect 389308 -19842 389382 -19786
rect 389438 -19842 389524 -19786
rect 389580 -19842 389648 -19786
rect 389308 -19928 389648 -19842
rect 389308 -19984 389382 -19928
rect 389438 -19984 389524 -19928
rect 389580 -19984 389648 -19928
rect 389308 -20070 389648 -19984
rect 389308 -20126 389382 -20070
rect 389438 -20126 389524 -20070
rect 389580 -20126 389648 -20070
rect 389308 -20212 389648 -20126
rect 389308 -20268 389382 -20212
rect 389438 -20268 389524 -20212
rect 389580 -20268 389648 -20212
rect 389308 -20354 389648 -20268
rect 389308 -20410 389382 -20354
rect 389438 -20410 389524 -20354
rect 389580 -20410 389648 -20354
rect 389308 -20496 389648 -20410
rect 389308 -20552 389382 -20496
rect 389438 -20552 389524 -20496
rect 389580 -20552 389648 -20496
rect 389308 -20638 389648 -20552
rect 389308 -20694 389382 -20638
rect 389438 -20694 389524 -20638
rect 389580 -20694 389648 -20638
rect 389308 -20780 389648 -20694
rect 389308 -20836 389382 -20780
rect 389438 -20836 389524 -20780
rect 389580 -20836 389648 -20780
rect 389308 -20922 389648 -20836
rect 389308 -20978 389382 -20922
rect 389438 -20978 389524 -20922
rect 389580 -20978 389648 -20922
rect 389308 -21064 389648 -20978
rect 389308 -21120 389382 -21064
rect 389438 -21120 389524 -21064
rect 389580 -21120 389648 -21064
rect 389308 -21206 389648 -21120
rect 389308 -21262 389382 -21206
rect 389438 -21262 389524 -21206
rect 389580 -21262 389648 -21206
rect 389308 -21348 389648 -21262
rect 389308 -21404 389382 -21348
rect 389438 -21404 389524 -21348
rect 389580 -21404 389648 -21348
rect 389308 -21490 389648 -21404
rect 389308 -21546 389382 -21490
rect 389438 -21546 389524 -21490
rect 389580 -21546 389648 -21490
rect 389308 -21632 389648 -21546
rect 389308 -21688 389382 -21632
rect 389438 -21688 389524 -21632
rect 389580 -21688 389648 -21632
rect 389308 -21774 389648 -21688
rect 389308 -21830 389382 -21774
rect 389438 -21830 389524 -21774
rect 389580 -21830 389648 -21774
rect 389308 -21916 389648 -21830
rect 389308 -21972 389382 -21916
rect 389438 -21972 389524 -21916
rect 389580 -21972 389648 -21916
rect 389308 -22058 389648 -21972
rect 389308 -22114 389382 -22058
rect 389438 -22114 389524 -22058
rect 389580 -22114 389648 -22058
rect 389308 -22200 389648 -22114
rect 389308 -22256 389382 -22200
rect 389438 -22256 389524 -22200
rect 389580 -22256 389648 -22200
rect 389308 -22342 389648 -22256
rect 389308 -22398 389382 -22342
rect 389438 -22398 389524 -22342
rect 389580 -22398 389648 -22342
rect 389308 -22484 389648 -22398
rect 389308 -22540 389382 -22484
rect 389438 -22540 389524 -22484
rect 389580 -22540 389648 -22484
rect 389308 -22626 389648 -22540
rect 389308 -22682 389382 -22626
rect 389438 -22682 389524 -22626
rect 389580 -22682 389648 -22626
rect 389308 -22768 389648 -22682
rect 389308 -22824 389382 -22768
rect 389438 -22824 389524 -22768
rect 389580 -22824 389648 -22768
rect 389308 -22910 389648 -22824
rect 389308 -22966 389382 -22910
rect 389438 -22966 389524 -22910
rect 389580 -22966 389648 -22910
rect 389308 -23052 389648 -22966
rect 389308 -23108 389382 -23052
rect 389438 -23108 389524 -23052
rect 389580 -23108 389648 -23052
rect 389308 -23194 389648 -23108
rect 389308 -23250 389382 -23194
rect 389438 -23250 389524 -23194
rect 389580 -23250 389648 -23194
rect 389308 -23336 389648 -23250
rect 389308 -23392 389382 -23336
rect 389438 -23392 389524 -23336
rect 389580 -23392 389648 -23336
rect 389308 -23478 389648 -23392
rect 389308 -23534 389382 -23478
rect 389438 -23534 389524 -23478
rect 389580 -23534 389648 -23478
rect 389308 -23620 389648 -23534
rect 389308 -23676 389382 -23620
rect 389438 -23676 389524 -23620
rect 389580 -23676 389648 -23620
rect 389308 -23762 389648 -23676
rect 389308 -23818 389382 -23762
rect 389438 -23818 389524 -23762
rect 389580 -23818 389648 -23762
rect 389308 -23904 389648 -23818
rect 389308 -23960 389382 -23904
rect 389438 -23960 389524 -23904
rect 389580 -23960 389648 -23904
rect 389308 -24046 389648 -23960
rect 389308 -24102 389382 -24046
rect 389438 -24102 389524 -24046
rect 389580 -24102 389648 -24046
rect 389308 -24188 389648 -24102
rect 389308 -24244 389382 -24188
rect 389438 -24244 389524 -24188
rect 389580 -24244 389648 -24188
rect 389308 -24330 389648 -24244
rect 389308 -24386 389382 -24330
rect 389438 -24386 389524 -24330
rect 389580 -24386 389648 -24330
rect 389308 -24472 389648 -24386
rect 389308 -24528 389382 -24472
rect 389438 -24528 389524 -24472
rect 389580 -24528 389648 -24472
rect 389308 -24614 389648 -24528
rect 389308 -24670 389382 -24614
rect 389438 -24670 389524 -24614
rect 389580 -24670 389648 -24614
rect 389308 -24756 389648 -24670
rect 389308 -24812 389382 -24756
rect 389438 -24812 389524 -24756
rect 389580 -24812 389648 -24756
rect 389308 -24898 389648 -24812
rect 389308 -24954 389382 -24898
rect 389438 -24954 389524 -24898
rect 389580 -24954 389648 -24898
rect 389308 -25040 389648 -24954
rect 389308 -25096 389382 -25040
rect 389438 -25096 389524 -25040
rect 389580 -25096 389648 -25040
rect 389308 -25182 389648 -25096
rect 389308 -25238 389382 -25182
rect 389438 -25238 389524 -25182
rect 389580 -25238 389648 -25182
rect 389308 -25324 389648 -25238
rect 389308 -25380 389382 -25324
rect 389438 -25380 389524 -25324
rect 389580 -25380 389648 -25324
rect 389308 -25466 389648 -25380
rect 389308 -25522 389382 -25466
rect 389438 -25522 389524 -25466
rect 389580 -25522 389648 -25466
rect 389308 -25590 389648 -25522
rect 389708 -13680 390048 -13590
rect 389708 -13736 389782 -13680
rect 389838 -13736 389924 -13680
rect 389980 -13736 390048 -13680
rect 389708 -13822 390048 -13736
rect 389708 -13878 389782 -13822
rect 389838 -13878 389924 -13822
rect 389980 -13878 390048 -13822
rect 389708 -13964 390048 -13878
rect 389708 -14020 389782 -13964
rect 389838 -14020 389924 -13964
rect 389980 -14020 390048 -13964
rect 389708 -14106 390048 -14020
rect 389708 -14162 389782 -14106
rect 389838 -14162 389924 -14106
rect 389980 -14162 390048 -14106
rect 389708 -14248 390048 -14162
rect 389708 -14304 389782 -14248
rect 389838 -14304 389924 -14248
rect 389980 -14304 390048 -14248
rect 389708 -14390 390048 -14304
rect 389708 -14446 389782 -14390
rect 389838 -14446 389924 -14390
rect 389980 -14446 390048 -14390
rect 389708 -14532 390048 -14446
rect 389708 -14588 389782 -14532
rect 389838 -14588 389924 -14532
rect 389980 -14588 390048 -14532
rect 389708 -14674 390048 -14588
rect 389708 -14730 389782 -14674
rect 389838 -14730 389924 -14674
rect 389980 -14730 390048 -14674
rect 389708 -14816 390048 -14730
rect 389708 -14872 389782 -14816
rect 389838 -14872 389924 -14816
rect 389980 -14872 390048 -14816
rect 389708 -14958 390048 -14872
rect 389708 -15014 389782 -14958
rect 389838 -15014 389924 -14958
rect 389980 -15014 390048 -14958
rect 389708 -15100 390048 -15014
rect 389708 -15156 389782 -15100
rect 389838 -15156 389924 -15100
rect 389980 -15156 390048 -15100
rect 389708 -15242 390048 -15156
rect 389708 -15298 389782 -15242
rect 389838 -15298 389924 -15242
rect 389980 -15298 390048 -15242
rect 389708 -15384 390048 -15298
rect 389708 -15440 389782 -15384
rect 389838 -15440 389924 -15384
rect 389980 -15440 390048 -15384
rect 389708 -15526 390048 -15440
rect 389708 -15582 389782 -15526
rect 389838 -15582 389924 -15526
rect 389980 -15582 390048 -15526
rect 389708 -15668 390048 -15582
rect 389708 -15724 389782 -15668
rect 389838 -15724 389924 -15668
rect 389980 -15724 390048 -15668
rect 389708 -15810 390048 -15724
rect 389708 -15866 389782 -15810
rect 389838 -15866 389924 -15810
rect 389980 -15866 390048 -15810
rect 389708 -15952 390048 -15866
rect 389708 -16008 389782 -15952
rect 389838 -16008 389924 -15952
rect 389980 -16008 390048 -15952
rect 389708 -16094 390048 -16008
rect 389708 -16150 389782 -16094
rect 389838 -16150 389924 -16094
rect 389980 -16150 390048 -16094
rect 389708 -16236 390048 -16150
rect 389708 -16292 389782 -16236
rect 389838 -16292 389924 -16236
rect 389980 -16292 390048 -16236
rect 389708 -16378 390048 -16292
rect 389708 -16434 389782 -16378
rect 389838 -16434 389924 -16378
rect 389980 -16434 390048 -16378
rect 389708 -16520 390048 -16434
rect 389708 -16576 389782 -16520
rect 389838 -16576 389924 -16520
rect 389980 -16576 390048 -16520
rect 389708 -16662 390048 -16576
rect 389708 -16718 389782 -16662
rect 389838 -16718 389924 -16662
rect 389980 -16718 390048 -16662
rect 389708 -16804 390048 -16718
rect 389708 -16860 389782 -16804
rect 389838 -16860 389924 -16804
rect 389980 -16860 390048 -16804
rect 389708 -16946 390048 -16860
rect 389708 -17002 389782 -16946
rect 389838 -17002 389924 -16946
rect 389980 -17002 390048 -16946
rect 389708 -17088 390048 -17002
rect 389708 -17144 389782 -17088
rect 389838 -17144 389924 -17088
rect 389980 -17144 390048 -17088
rect 389708 -17230 390048 -17144
rect 389708 -17286 389782 -17230
rect 389838 -17286 389924 -17230
rect 389980 -17286 390048 -17230
rect 389708 -17372 390048 -17286
rect 389708 -17428 389782 -17372
rect 389838 -17428 389924 -17372
rect 389980 -17428 390048 -17372
rect 389708 -17514 390048 -17428
rect 389708 -17570 389782 -17514
rect 389838 -17570 389924 -17514
rect 389980 -17570 390048 -17514
rect 389708 -17656 390048 -17570
rect 389708 -17712 389782 -17656
rect 389838 -17712 389924 -17656
rect 389980 -17712 390048 -17656
rect 389708 -17798 390048 -17712
rect 389708 -17854 389782 -17798
rect 389838 -17854 389924 -17798
rect 389980 -17854 390048 -17798
rect 389708 -17940 390048 -17854
rect 389708 -17996 389782 -17940
rect 389838 -17996 389924 -17940
rect 389980 -17996 390048 -17940
rect 389708 -18082 390048 -17996
rect 389708 -18138 389782 -18082
rect 389838 -18138 389924 -18082
rect 389980 -18138 390048 -18082
rect 389708 -18224 390048 -18138
rect 389708 -18280 389782 -18224
rect 389838 -18280 389924 -18224
rect 389980 -18280 390048 -18224
rect 389708 -18366 390048 -18280
rect 389708 -18422 389782 -18366
rect 389838 -18422 389924 -18366
rect 389980 -18422 390048 -18366
rect 389708 -18508 390048 -18422
rect 389708 -18564 389782 -18508
rect 389838 -18564 389924 -18508
rect 389980 -18564 390048 -18508
rect 389708 -18650 390048 -18564
rect 389708 -18706 389782 -18650
rect 389838 -18706 389924 -18650
rect 389980 -18706 390048 -18650
rect 389708 -18792 390048 -18706
rect 389708 -18848 389782 -18792
rect 389838 -18848 389924 -18792
rect 389980 -18848 390048 -18792
rect 389708 -18934 390048 -18848
rect 389708 -18990 389782 -18934
rect 389838 -18990 389924 -18934
rect 389980 -18990 390048 -18934
rect 389708 -19076 390048 -18990
rect 389708 -19132 389782 -19076
rect 389838 -19132 389924 -19076
rect 389980 -19132 390048 -19076
rect 389708 -19218 390048 -19132
rect 389708 -19274 389782 -19218
rect 389838 -19274 389924 -19218
rect 389980 -19274 390048 -19218
rect 389708 -19360 390048 -19274
rect 389708 -19416 389782 -19360
rect 389838 -19416 389924 -19360
rect 389980 -19416 390048 -19360
rect 389708 -19502 390048 -19416
rect 389708 -19558 389782 -19502
rect 389838 -19558 389924 -19502
rect 389980 -19558 390048 -19502
rect 389708 -19644 390048 -19558
rect 389708 -19700 389782 -19644
rect 389838 -19700 389924 -19644
rect 389980 -19700 390048 -19644
rect 389708 -19786 390048 -19700
rect 389708 -19842 389782 -19786
rect 389838 -19842 389924 -19786
rect 389980 -19842 390048 -19786
rect 389708 -19928 390048 -19842
rect 389708 -19984 389782 -19928
rect 389838 -19984 389924 -19928
rect 389980 -19984 390048 -19928
rect 389708 -20070 390048 -19984
rect 389708 -20126 389782 -20070
rect 389838 -20126 389924 -20070
rect 389980 -20126 390048 -20070
rect 389708 -20212 390048 -20126
rect 389708 -20268 389782 -20212
rect 389838 -20268 389924 -20212
rect 389980 -20268 390048 -20212
rect 389708 -20354 390048 -20268
rect 389708 -20410 389782 -20354
rect 389838 -20410 389924 -20354
rect 389980 -20410 390048 -20354
rect 389708 -20496 390048 -20410
rect 389708 -20552 389782 -20496
rect 389838 -20552 389924 -20496
rect 389980 -20552 390048 -20496
rect 389708 -20638 390048 -20552
rect 389708 -20694 389782 -20638
rect 389838 -20694 389924 -20638
rect 389980 -20694 390048 -20638
rect 389708 -20780 390048 -20694
rect 389708 -20836 389782 -20780
rect 389838 -20836 389924 -20780
rect 389980 -20836 390048 -20780
rect 389708 -20922 390048 -20836
rect 389708 -20978 389782 -20922
rect 389838 -20978 389924 -20922
rect 389980 -20978 390048 -20922
rect 389708 -21064 390048 -20978
rect 389708 -21120 389782 -21064
rect 389838 -21120 389924 -21064
rect 389980 -21120 390048 -21064
rect 389708 -21206 390048 -21120
rect 389708 -21262 389782 -21206
rect 389838 -21262 389924 -21206
rect 389980 -21262 390048 -21206
rect 389708 -21348 390048 -21262
rect 389708 -21404 389782 -21348
rect 389838 -21404 389924 -21348
rect 389980 -21404 390048 -21348
rect 389708 -21490 390048 -21404
rect 389708 -21546 389782 -21490
rect 389838 -21546 389924 -21490
rect 389980 -21546 390048 -21490
rect 389708 -21632 390048 -21546
rect 389708 -21688 389782 -21632
rect 389838 -21688 389924 -21632
rect 389980 -21688 390048 -21632
rect 389708 -21774 390048 -21688
rect 389708 -21830 389782 -21774
rect 389838 -21830 389924 -21774
rect 389980 -21830 390048 -21774
rect 389708 -21916 390048 -21830
rect 389708 -21972 389782 -21916
rect 389838 -21972 389924 -21916
rect 389980 -21972 390048 -21916
rect 389708 -22058 390048 -21972
rect 389708 -22114 389782 -22058
rect 389838 -22114 389924 -22058
rect 389980 -22114 390048 -22058
rect 389708 -22200 390048 -22114
rect 389708 -22256 389782 -22200
rect 389838 -22256 389924 -22200
rect 389980 -22256 390048 -22200
rect 389708 -22342 390048 -22256
rect 389708 -22398 389782 -22342
rect 389838 -22398 389924 -22342
rect 389980 -22398 390048 -22342
rect 389708 -22484 390048 -22398
rect 389708 -22540 389782 -22484
rect 389838 -22540 389924 -22484
rect 389980 -22540 390048 -22484
rect 389708 -22626 390048 -22540
rect 389708 -22682 389782 -22626
rect 389838 -22682 389924 -22626
rect 389980 -22682 390048 -22626
rect 389708 -22768 390048 -22682
rect 389708 -22824 389782 -22768
rect 389838 -22824 389924 -22768
rect 389980 -22824 390048 -22768
rect 389708 -22910 390048 -22824
rect 389708 -22966 389782 -22910
rect 389838 -22966 389924 -22910
rect 389980 -22966 390048 -22910
rect 389708 -23052 390048 -22966
rect 389708 -23108 389782 -23052
rect 389838 -23108 389924 -23052
rect 389980 -23108 390048 -23052
rect 389708 -23194 390048 -23108
rect 389708 -23250 389782 -23194
rect 389838 -23250 389924 -23194
rect 389980 -23250 390048 -23194
rect 389708 -23336 390048 -23250
rect 389708 -23392 389782 -23336
rect 389838 -23392 389924 -23336
rect 389980 -23392 390048 -23336
rect 389708 -23478 390048 -23392
rect 389708 -23534 389782 -23478
rect 389838 -23534 389924 -23478
rect 389980 -23534 390048 -23478
rect 389708 -23620 390048 -23534
rect 389708 -23676 389782 -23620
rect 389838 -23676 389924 -23620
rect 389980 -23676 390048 -23620
rect 389708 -23762 390048 -23676
rect 389708 -23818 389782 -23762
rect 389838 -23818 389924 -23762
rect 389980 -23818 390048 -23762
rect 389708 -23904 390048 -23818
rect 389708 -23960 389782 -23904
rect 389838 -23960 389924 -23904
rect 389980 -23960 390048 -23904
rect 389708 -24046 390048 -23960
rect 389708 -24102 389782 -24046
rect 389838 -24102 389924 -24046
rect 389980 -24102 390048 -24046
rect 389708 -24188 390048 -24102
rect 389708 -24244 389782 -24188
rect 389838 -24244 389924 -24188
rect 389980 -24244 390048 -24188
rect 389708 -24330 390048 -24244
rect 389708 -24386 389782 -24330
rect 389838 -24386 389924 -24330
rect 389980 -24386 390048 -24330
rect 389708 -24472 390048 -24386
rect 389708 -24528 389782 -24472
rect 389838 -24528 389924 -24472
rect 389980 -24528 390048 -24472
rect 389708 -24614 390048 -24528
rect 389708 -24670 389782 -24614
rect 389838 -24670 389924 -24614
rect 389980 -24670 390048 -24614
rect 389708 -24756 390048 -24670
rect 389708 -24812 389782 -24756
rect 389838 -24812 389924 -24756
rect 389980 -24812 390048 -24756
rect 389708 -24898 390048 -24812
rect 389708 -24954 389782 -24898
rect 389838 -24954 389924 -24898
rect 389980 -24954 390048 -24898
rect 389708 -25040 390048 -24954
rect 389708 -25096 389782 -25040
rect 389838 -25096 389924 -25040
rect 389980 -25096 390048 -25040
rect 389708 -25182 390048 -25096
rect 389708 -25238 389782 -25182
rect 389838 -25238 389924 -25182
rect 389980 -25238 390048 -25182
rect 389708 -25324 390048 -25238
rect 389708 -25380 389782 -25324
rect 389838 -25380 389924 -25324
rect 389980 -25380 390048 -25324
rect 389708 -25466 390048 -25380
rect 389708 -25522 389782 -25466
rect 389838 -25522 389924 -25466
rect 389980 -25522 390048 -25466
rect 389708 -25590 390048 -25522
rect 390108 -13680 390448 -13590
rect 390108 -13736 390179 -13680
rect 390235 -13736 390321 -13680
rect 390377 -13736 390448 -13680
rect 390108 -13822 390448 -13736
rect 390108 -13878 390179 -13822
rect 390235 -13878 390321 -13822
rect 390377 -13878 390448 -13822
rect 390108 -13964 390448 -13878
rect 390108 -14020 390179 -13964
rect 390235 -14020 390321 -13964
rect 390377 -14020 390448 -13964
rect 390108 -14106 390448 -14020
rect 390108 -14162 390179 -14106
rect 390235 -14162 390321 -14106
rect 390377 -14162 390448 -14106
rect 390108 -14248 390448 -14162
rect 390108 -14304 390179 -14248
rect 390235 -14304 390321 -14248
rect 390377 -14304 390448 -14248
rect 390108 -14390 390448 -14304
rect 390108 -14446 390179 -14390
rect 390235 -14446 390321 -14390
rect 390377 -14446 390448 -14390
rect 390108 -14532 390448 -14446
rect 390108 -14588 390179 -14532
rect 390235 -14588 390321 -14532
rect 390377 -14588 390448 -14532
rect 390108 -14674 390448 -14588
rect 390108 -14730 390179 -14674
rect 390235 -14730 390321 -14674
rect 390377 -14730 390448 -14674
rect 390108 -14816 390448 -14730
rect 390108 -14872 390179 -14816
rect 390235 -14872 390321 -14816
rect 390377 -14872 390448 -14816
rect 390108 -14958 390448 -14872
rect 390108 -15014 390179 -14958
rect 390235 -15014 390321 -14958
rect 390377 -15014 390448 -14958
rect 390108 -15100 390448 -15014
rect 390108 -15156 390179 -15100
rect 390235 -15156 390321 -15100
rect 390377 -15156 390448 -15100
rect 390108 -15242 390448 -15156
rect 390108 -15298 390179 -15242
rect 390235 -15298 390321 -15242
rect 390377 -15298 390448 -15242
rect 390108 -15384 390448 -15298
rect 390108 -15440 390179 -15384
rect 390235 -15440 390321 -15384
rect 390377 -15440 390448 -15384
rect 390108 -15526 390448 -15440
rect 390108 -15582 390179 -15526
rect 390235 -15582 390321 -15526
rect 390377 -15582 390448 -15526
rect 390108 -15668 390448 -15582
rect 390108 -15724 390179 -15668
rect 390235 -15724 390321 -15668
rect 390377 -15724 390448 -15668
rect 390108 -15810 390448 -15724
rect 390108 -15866 390179 -15810
rect 390235 -15866 390321 -15810
rect 390377 -15866 390448 -15810
rect 390108 -15952 390448 -15866
rect 390108 -16008 390179 -15952
rect 390235 -16008 390321 -15952
rect 390377 -16008 390448 -15952
rect 390108 -16094 390448 -16008
rect 390108 -16150 390179 -16094
rect 390235 -16150 390321 -16094
rect 390377 -16150 390448 -16094
rect 390108 -16236 390448 -16150
rect 390108 -16292 390179 -16236
rect 390235 -16292 390321 -16236
rect 390377 -16292 390448 -16236
rect 390108 -16378 390448 -16292
rect 390108 -16434 390179 -16378
rect 390235 -16434 390321 -16378
rect 390377 -16434 390448 -16378
rect 390108 -16520 390448 -16434
rect 390108 -16576 390179 -16520
rect 390235 -16576 390321 -16520
rect 390377 -16576 390448 -16520
rect 390108 -16662 390448 -16576
rect 390108 -16718 390179 -16662
rect 390235 -16718 390321 -16662
rect 390377 -16718 390448 -16662
rect 390108 -16804 390448 -16718
rect 390108 -16860 390179 -16804
rect 390235 -16860 390321 -16804
rect 390377 -16860 390448 -16804
rect 390108 -16946 390448 -16860
rect 390108 -17002 390179 -16946
rect 390235 -17002 390321 -16946
rect 390377 -17002 390448 -16946
rect 390108 -17088 390448 -17002
rect 390108 -17144 390179 -17088
rect 390235 -17144 390321 -17088
rect 390377 -17144 390448 -17088
rect 390108 -17230 390448 -17144
rect 390108 -17286 390179 -17230
rect 390235 -17286 390321 -17230
rect 390377 -17286 390448 -17230
rect 390108 -17372 390448 -17286
rect 390108 -17428 390179 -17372
rect 390235 -17428 390321 -17372
rect 390377 -17428 390448 -17372
rect 390108 -17514 390448 -17428
rect 390108 -17570 390179 -17514
rect 390235 -17570 390321 -17514
rect 390377 -17570 390448 -17514
rect 390108 -17656 390448 -17570
rect 390108 -17712 390179 -17656
rect 390235 -17712 390321 -17656
rect 390377 -17712 390448 -17656
rect 390108 -17798 390448 -17712
rect 390108 -17854 390179 -17798
rect 390235 -17854 390321 -17798
rect 390377 -17854 390448 -17798
rect 390108 -17940 390448 -17854
rect 390108 -17996 390179 -17940
rect 390235 -17996 390321 -17940
rect 390377 -17996 390448 -17940
rect 390108 -18082 390448 -17996
rect 390108 -18138 390179 -18082
rect 390235 -18138 390321 -18082
rect 390377 -18138 390448 -18082
rect 390108 -18224 390448 -18138
rect 390108 -18280 390179 -18224
rect 390235 -18280 390321 -18224
rect 390377 -18280 390448 -18224
rect 390108 -18366 390448 -18280
rect 390108 -18422 390179 -18366
rect 390235 -18422 390321 -18366
rect 390377 -18422 390448 -18366
rect 390108 -18508 390448 -18422
rect 390108 -18564 390179 -18508
rect 390235 -18564 390321 -18508
rect 390377 -18564 390448 -18508
rect 390108 -18650 390448 -18564
rect 390108 -18706 390179 -18650
rect 390235 -18706 390321 -18650
rect 390377 -18706 390448 -18650
rect 390108 -18792 390448 -18706
rect 390108 -18848 390179 -18792
rect 390235 -18848 390321 -18792
rect 390377 -18848 390448 -18792
rect 390108 -18934 390448 -18848
rect 390108 -18990 390179 -18934
rect 390235 -18990 390321 -18934
rect 390377 -18990 390448 -18934
rect 390108 -19076 390448 -18990
rect 390108 -19132 390179 -19076
rect 390235 -19132 390321 -19076
rect 390377 -19132 390448 -19076
rect 390108 -19218 390448 -19132
rect 390108 -19274 390179 -19218
rect 390235 -19274 390321 -19218
rect 390377 -19274 390448 -19218
rect 390108 -19360 390448 -19274
rect 390108 -19416 390179 -19360
rect 390235 -19416 390321 -19360
rect 390377 -19416 390448 -19360
rect 390108 -19502 390448 -19416
rect 390108 -19558 390179 -19502
rect 390235 -19558 390321 -19502
rect 390377 -19558 390448 -19502
rect 390108 -19644 390448 -19558
rect 390108 -19700 390179 -19644
rect 390235 -19700 390321 -19644
rect 390377 -19700 390448 -19644
rect 390108 -19786 390448 -19700
rect 390108 -19842 390179 -19786
rect 390235 -19842 390321 -19786
rect 390377 -19842 390448 -19786
rect 390108 -19928 390448 -19842
rect 390108 -19984 390179 -19928
rect 390235 -19984 390321 -19928
rect 390377 -19984 390448 -19928
rect 390108 -20070 390448 -19984
rect 390108 -20126 390179 -20070
rect 390235 -20126 390321 -20070
rect 390377 -20126 390448 -20070
rect 390108 -20212 390448 -20126
rect 390108 -20268 390179 -20212
rect 390235 -20268 390321 -20212
rect 390377 -20268 390448 -20212
rect 390108 -20354 390448 -20268
rect 390108 -20410 390179 -20354
rect 390235 -20410 390321 -20354
rect 390377 -20410 390448 -20354
rect 390108 -20496 390448 -20410
rect 390108 -20552 390179 -20496
rect 390235 -20552 390321 -20496
rect 390377 -20552 390448 -20496
rect 390108 -20638 390448 -20552
rect 390108 -20694 390179 -20638
rect 390235 -20694 390321 -20638
rect 390377 -20694 390448 -20638
rect 390108 -20780 390448 -20694
rect 390108 -20836 390179 -20780
rect 390235 -20836 390321 -20780
rect 390377 -20836 390448 -20780
rect 390108 -20922 390448 -20836
rect 390108 -20978 390179 -20922
rect 390235 -20978 390321 -20922
rect 390377 -20978 390448 -20922
rect 390108 -21064 390448 -20978
rect 390108 -21120 390179 -21064
rect 390235 -21120 390321 -21064
rect 390377 -21120 390448 -21064
rect 390108 -21206 390448 -21120
rect 390108 -21262 390179 -21206
rect 390235 -21262 390321 -21206
rect 390377 -21262 390448 -21206
rect 390108 -21348 390448 -21262
rect 390108 -21404 390179 -21348
rect 390235 -21404 390321 -21348
rect 390377 -21404 390448 -21348
rect 390108 -21490 390448 -21404
rect 390108 -21546 390179 -21490
rect 390235 -21546 390321 -21490
rect 390377 -21546 390448 -21490
rect 390108 -21632 390448 -21546
rect 390108 -21688 390179 -21632
rect 390235 -21688 390321 -21632
rect 390377 -21688 390448 -21632
rect 390108 -21774 390448 -21688
rect 390108 -21830 390179 -21774
rect 390235 -21830 390321 -21774
rect 390377 -21830 390448 -21774
rect 390108 -21916 390448 -21830
rect 390108 -21972 390179 -21916
rect 390235 -21972 390321 -21916
rect 390377 -21972 390448 -21916
rect 390108 -22058 390448 -21972
rect 390108 -22114 390179 -22058
rect 390235 -22114 390321 -22058
rect 390377 -22114 390448 -22058
rect 390108 -22200 390448 -22114
rect 390108 -22256 390179 -22200
rect 390235 -22256 390321 -22200
rect 390377 -22256 390448 -22200
rect 390108 -22342 390448 -22256
rect 390108 -22398 390179 -22342
rect 390235 -22398 390321 -22342
rect 390377 -22398 390448 -22342
rect 390108 -22484 390448 -22398
rect 390108 -22540 390179 -22484
rect 390235 -22540 390321 -22484
rect 390377 -22540 390448 -22484
rect 390108 -22626 390448 -22540
rect 390108 -22682 390179 -22626
rect 390235 -22682 390321 -22626
rect 390377 -22682 390448 -22626
rect 390108 -22768 390448 -22682
rect 390108 -22824 390179 -22768
rect 390235 -22824 390321 -22768
rect 390377 -22824 390448 -22768
rect 390108 -22910 390448 -22824
rect 390108 -22966 390179 -22910
rect 390235 -22966 390321 -22910
rect 390377 -22966 390448 -22910
rect 390108 -23052 390448 -22966
rect 390108 -23108 390179 -23052
rect 390235 -23108 390321 -23052
rect 390377 -23108 390448 -23052
rect 390108 -23194 390448 -23108
rect 390108 -23250 390179 -23194
rect 390235 -23250 390321 -23194
rect 390377 -23250 390448 -23194
rect 390108 -23336 390448 -23250
rect 390108 -23392 390179 -23336
rect 390235 -23392 390321 -23336
rect 390377 -23392 390448 -23336
rect 390108 -23478 390448 -23392
rect 390108 -23534 390179 -23478
rect 390235 -23534 390321 -23478
rect 390377 -23534 390448 -23478
rect 390108 -23620 390448 -23534
rect 390108 -23676 390179 -23620
rect 390235 -23676 390321 -23620
rect 390377 -23676 390448 -23620
rect 390108 -23762 390448 -23676
rect 390108 -23818 390179 -23762
rect 390235 -23818 390321 -23762
rect 390377 -23818 390448 -23762
rect 390108 -23904 390448 -23818
rect 390108 -23960 390179 -23904
rect 390235 -23960 390321 -23904
rect 390377 -23960 390448 -23904
rect 390108 -24046 390448 -23960
rect 390108 -24102 390179 -24046
rect 390235 -24102 390321 -24046
rect 390377 -24102 390448 -24046
rect 390108 -24188 390448 -24102
rect 390108 -24244 390179 -24188
rect 390235 -24244 390321 -24188
rect 390377 -24244 390448 -24188
rect 390108 -24330 390448 -24244
rect 390108 -24386 390179 -24330
rect 390235 -24386 390321 -24330
rect 390377 -24386 390448 -24330
rect 390108 -24472 390448 -24386
rect 390108 -24528 390179 -24472
rect 390235 -24528 390321 -24472
rect 390377 -24528 390448 -24472
rect 390108 -24614 390448 -24528
rect 390108 -24670 390179 -24614
rect 390235 -24670 390321 -24614
rect 390377 -24670 390448 -24614
rect 390108 -24756 390448 -24670
rect 390108 -24812 390179 -24756
rect 390235 -24812 390321 -24756
rect 390377 -24812 390448 -24756
rect 390108 -24898 390448 -24812
rect 390108 -24954 390179 -24898
rect 390235 -24954 390321 -24898
rect 390377 -24954 390448 -24898
rect 390108 -25040 390448 -24954
rect 390108 -25096 390179 -25040
rect 390235 -25096 390321 -25040
rect 390377 -25096 390448 -25040
rect 390108 -25182 390448 -25096
rect 390108 -25238 390179 -25182
rect 390235 -25238 390321 -25182
rect 390377 -25238 390448 -25182
rect 390108 -25324 390448 -25238
rect 390108 -25380 390179 -25324
rect 390235 -25380 390321 -25324
rect 390377 -25380 390448 -25324
rect 390108 -25466 390448 -25380
rect 390108 -25522 390179 -25466
rect 390235 -25522 390321 -25466
rect 390377 -25522 390448 -25466
rect 390108 -25590 390448 -25522
rect 390508 -13680 390848 -13590
rect 390508 -13736 390576 -13680
rect 390632 -13736 390718 -13680
rect 390774 -13736 390848 -13680
rect 390508 -13822 390848 -13736
rect 390508 -13878 390576 -13822
rect 390632 -13878 390718 -13822
rect 390774 -13878 390848 -13822
rect 390508 -13964 390848 -13878
rect 390508 -14020 390576 -13964
rect 390632 -14020 390718 -13964
rect 390774 -14020 390848 -13964
rect 390508 -14106 390848 -14020
rect 390508 -14162 390576 -14106
rect 390632 -14162 390718 -14106
rect 390774 -14162 390848 -14106
rect 390508 -14248 390848 -14162
rect 390508 -14304 390576 -14248
rect 390632 -14304 390718 -14248
rect 390774 -14304 390848 -14248
rect 390508 -14390 390848 -14304
rect 390508 -14446 390576 -14390
rect 390632 -14446 390718 -14390
rect 390774 -14446 390848 -14390
rect 390508 -14532 390848 -14446
rect 390508 -14588 390576 -14532
rect 390632 -14588 390718 -14532
rect 390774 -14588 390848 -14532
rect 390508 -14674 390848 -14588
rect 390508 -14730 390576 -14674
rect 390632 -14730 390718 -14674
rect 390774 -14730 390848 -14674
rect 390508 -14816 390848 -14730
rect 390508 -14872 390576 -14816
rect 390632 -14872 390718 -14816
rect 390774 -14872 390848 -14816
rect 390508 -14958 390848 -14872
rect 390508 -15014 390576 -14958
rect 390632 -15014 390718 -14958
rect 390774 -15014 390848 -14958
rect 390508 -15100 390848 -15014
rect 390508 -15156 390576 -15100
rect 390632 -15156 390718 -15100
rect 390774 -15156 390848 -15100
rect 390508 -15242 390848 -15156
rect 390508 -15298 390576 -15242
rect 390632 -15298 390718 -15242
rect 390774 -15298 390848 -15242
rect 390508 -15384 390848 -15298
rect 390508 -15440 390576 -15384
rect 390632 -15440 390718 -15384
rect 390774 -15440 390848 -15384
rect 390508 -15526 390848 -15440
rect 390508 -15582 390576 -15526
rect 390632 -15582 390718 -15526
rect 390774 -15582 390848 -15526
rect 390508 -15668 390848 -15582
rect 390508 -15724 390576 -15668
rect 390632 -15724 390718 -15668
rect 390774 -15724 390848 -15668
rect 390508 -15810 390848 -15724
rect 390508 -15866 390576 -15810
rect 390632 -15866 390718 -15810
rect 390774 -15866 390848 -15810
rect 390508 -15952 390848 -15866
rect 390508 -16008 390576 -15952
rect 390632 -16008 390718 -15952
rect 390774 -16008 390848 -15952
rect 390508 -16094 390848 -16008
rect 390508 -16150 390576 -16094
rect 390632 -16150 390718 -16094
rect 390774 -16150 390848 -16094
rect 390508 -16236 390848 -16150
rect 390508 -16292 390576 -16236
rect 390632 -16292 390718 -16236
rect 390774 -16292 390848 -16236
rect 390508 -16378 390848 -16292
rect 390508 -16434 390576 -16378
rect 390632 -16434 390718 -16378
rect 390774 -16434 390848 -16378
rect 390508 -16520 390848 -16434
rect 390508 -16576 390576 -16520
rect 390632 -16576 390718 -16520
rect 390774 -16576 390848 -16520
rect 390508 -16662 390848 -16576
rect 390508 -16718 390576 -16662
rect 390632 -16718 390718 -16662
rect 390774 -16718 390848 -16662
rect 390508 -16804 390848 -16718
rect 390508 -16860 390576 -16804
rect 390632 -16860 390718 -16804
rect 390774 -16860 390848 -16804
rect 390508 -16946 390848 -16860
rect 390508 -17002 390576 -16946
rect 390632 -17002 390718 -16946
rect 390774 -17002 390848 -16946
rect 390508 -17088 390848 -17002
rect 390508 -17144 390576 -17088
rect 390632 -17144 390718 -17088
rect 390774 -17144 390848 -17088
rect 390508 -17230 390848 -17144
rect 390508 -17286 390576 -17230
rect 390632 -17286 390718 -17230
rect 390774 -17286 390848 -17230
rect 390508 -17372 390848 -17286
rect 390508 -17428 390576 -17372
rect 390632 -17428 390718 -17372
rect 390774 -17428 390848 -17372
rect 390508 -17514 390848 -17428
rect 390508 -17570 390576 -17514
rect 390632 -17570 390718 -17514
rect 390774 -17570 390848 -17514
rect 390508 -17656 390848 -17570
rect 390508 -17712 390576 -17656
rect 390632 -17712 390718 -17656
rect 390774 -17712 390848 -17656
rect 390508 -17798 390848 -17712
rect 390508 -17854 390576 -17798
rect 390632 -17854 390718 -17798
rect 390774 -17854 390848 -17798
rect 390508 -17940 390848 -17854
rect 390508 -17996 390576 -17940
rect 390632 -17996 390718 -17940
rect 390774 -17996 390848 -17940
rect 390508 -18082 390848 -17996
rect 390508 -18138 390576 -18082
rect 390632 -18138 390718 -18082
rect 390774 -18138 390848 -18082
rect 390508 -18224 390848 -18138
rect 390508 -18280 390576 -18224
rect 390632 -18280 390718 -18224
rect 390774 -18280 390848 -18224
rect 390508 -18366 390848 -18280
rect 390508 -18422 390576 -18366
rect 390632 -18422 390718 -18366
rect 390774 -18422 390848 -18366
rect 390508 -18508 390848 -18422
rect 390508 -18564 390576 -18508
rect 390632 -18564 390718 -18508
rect 390774 -18564 390848 -18508
rect 390508 -18650 390848 -18564
rect 390508 -18706 390576 -18650
rect 390632 -18706 390718 -18650
rect 390774 -18706 390848 -18650
rect 390508 -18792 390848 -18706
rect 390508 -18848 390576 -18792
rect 390632 -18848 390718 -18792
rect 390774 -18848 390848 -18792
rect 390508 -18934 390848 -18848
rect 390508 -18990 390576 -18934
rect 390632 -18990 390718 -18934
rect 390774 -18990 390848 -18934
rect 390508 -19076 390848 -18990
rect 390508 -19132 390576 -19076
rect 390632 -19132 390718 -19076
rect 390774 -19132 390848 -19076
rect 390508 -19218 390848 -19132
rect 390508 -19274 390576 -19218
rect 390632 -19274 390718 -19218
rect 390774 -19274 390848 -19218
rect 390508 -19360 390848 -19274
rect 390508 -19416 390576 -19360
rect 390632 -19416 390718 -19360
rect 390774 -19416 390848 -19360
rect 390508 -19502 390848 -19416
rect 390508 -19558 390576 -19502
rect 390632 -19558 390718 -19502
rect 390774 -19558 390848 -19502
rect 390508 -19644 390848 -19558
rect 390508 -19700 390576 -19644
rect 390632 -19700 390718 -19644
rect 390774 -19700 390848 -19644
rect 390508 -19786 390848 -19700
rect 390508 -19842 390576 -19786
rect 390632 -19842 390718 -19786
rect 390774 -19842 390848 -19786
rect 390508 -19928 390848 -19842
rect 390508 -19984 390576 -19928
rect 390632 -19984 390718 -19928
rect 390774 -19984 390848 -19928
rect 390508 -20070 390848 -19984
rect 390508 -20126 390576 -20070
rect 390632 -20126 390718 -20070
rect 390774 -20126 390848 -20070
rect 390508 -20212 390848 -20126
rect 390508 -20268 390576 -20212
rect 390632 -20268 390718 -20212
rect 390774 -20268 390848 -20212
rect 390508 -20354 390848 -20268
rect 390508 -20410 390576 -20354
rect 390632 -20410 390718 -20354
rect 390774 -20410 390848 -20354
rect 390508 -20496 390848 -20410
rect 390508 -20552 390576 -20496
rect 390632 -20552 390718 -20496
rect 390774 -20552 390848 -20496
rect 390508 -20638 390848 -20552
rect 390508 -20694 390576 -20638
rect 390632 -20694 390718 -20638
rect 390774 -20694 390848 -20638
rect 390508 -20780 390848 -20694
rect 390508 -20836 390576 -20780
rect 390632 -20836 390718 -20780
rect 390774 -20836 390848 -20780
rect 390508 -20922 390848 -20836
rect 390508 -20978 390576 -20922
rect 390632 -20978 390718 -20922
rect 390774 -20978 390848 -20922
rect 390508 -21064 390848 -20978
rect 390508 -21120 390576 -21064
rect 390632 -21120 390718 -21064
rect 390774 -21120 390848 -21064
rect 390508 -21206 390848 -21120
rect 390508 -21262 390576 -21206
rect 390632 -21262 390718 -21206
rect 390774 -21262 390848 -21206
rect 390508 -21348 390848 -21262
rect 390508 -21404 390576 -21348
rect 390632 -21404 390718 -21348
rect 390774 -21404 390848 -21348
rect 390508 -21490 390848 -21404
rect 390508 -21546 390576 -21490
rect 390632 -21546 390718 -21490
rect 390774 -21546 390848 -21490
rect 390508 -21632 390848 -21546
rect 390508 -21688 390576 -21632
rect 390632 -21688 390718 -21632
rect 390774 -21688 390848 -21632
rect 390508 -21774 390848 -21688
rect 390508 -21830 390576 -21774
rect 390632 -21830 390718 -21774
rect 390774 -21830 390848 -21774
rect 390508 -21916 390848 -21830
rect 390508 -21972 390576 -21916
rect 390632 -21972 390718 -21916
rect 390774 -21972 390848 -21916
rect 390508 -22058 390848 -21972
rect 390508 -22114 390576 -22058
rect 390632 -22114 390718 -22058
rect 390774 -22114 390848 -22058
rect 390508 -22200 390848 -22114
rect 390508 -22256 390576 -22200
rect 390632 -22256 390718 -22200
rect 390774 -22256 390848 -22200
rect 390508 -22342 390848 -22256
rect 390508 -22398 390576 -22342
rect 390632 -22398 390718 -22342
rect 390774 -22398 390848 -22342
rect 390508 -22484 390848 -22398
rect 390508 -22540 390576 -22484
rect 390632 -22540 390718 -22484
rect 390774 -22540 390848 -22484
rect 390508 -22626 390848 -22540
rect 390508 -22682 390576 -22626
rect 390632 -22682 390718 -22626
rect 390774 -22682 390848 -22626
rect 390508 -22768 390848 -22682
rect 390508 -22824 390576 -22768
rect 390632 -22824 390718 -22768
rect 390774 -22824 390848 -22768
rect 390508 -22910 390848 -22824
rect 390508 -22966 390576 -22910
rect 390632 -22966 390718 -22910
rect 390774 -22966 390848 -22910
rect 390508 -23052 390848 -22966
rect 390508 -23108 390576 -23052
rect 390632 -23108 390718 -23052
rect 390774 -23108 390848 -23052
rect 390508 -23194 390848 -23108
rect 390508 -23250 390576 -23194
rect 390632 -23250 390718 -23194
rect 390774 -23250 390848 -23194
rect 390508 -23336 390848 -23250
rect 390508 -23392 390576 -23336
rect 390632 -23392 390718 -23336
rect 390774 -23392 390848 -23336
rect 390508 -23478 390848 -23392
rect 390508 -23534 390576 -23478
rect 390632 -23534 390718 -23478
rect 390774 -23534 390848 -23478
rect 390508 -23620 390848 -23534
rect 390508 -23676 390576 -23620
rect 390632 -23676 390718 -23620
rect 390774 -23676 390848 -23620
rect 390508 -23762 390848 -23676
rect 390508 -23818 390576 -23762
rect 390632 -23818 390718 -23762
rect 390774 -23818 390848 -23762
rect 390508 -23904 390848 -23818
rect 390508 -23960 390576 -23904
rect 390632 -23960 390718 -23904
rect 390774 -23960 390848 -23904
rect 390508 -24046 390848 -23960
rect 390508 -24102 390576 -24046
rect 390632 -24102 390718 -24046
rect 390774 -24102 390848 -24046
rect 390508 -24188 390848 -24102
rect 390508 -24244 390576 -24188
rect 390632 -24244 390718 -24188
rect 390774 -24244 390848 -24188
rect 390508 -24330 390848 -24244
rect 390508 -24386 390576 -24330
rect 390632 -24386 390718 -24330
rect 390774 -24386 390848 -24330
rect 390508 -24472 390848 -24386
rect 390508 -24528 390576 -24472
rect 390632 -24528 390718 -24472
rect 390774 -24528 390848 -24472
rect 390508 -24614 390848 -24528
rect 390508 -24670 390576 -24614
rect 390632 -24670 390718 -24614
rect 390774 -24670 390848 -24614
rect 390508 -24756 390848 -24670
rect 390508 -24812 390576 -24756
rect 390632 -24812 390718 -24756
rect 390774 -24812 390848 -24756
rect 390508 -24898 390848 -24812
rect 390508 -24954 390576 -24898
rect 390632 -24954 390718 -24898
rect 390774 -24954 390848 -24898
rect 390508 -25040 390848 -24954
rect 390508 -25096 390576 -25040
rect 390632 -25096 390718 -25040
rect 390774 -25096 390848 -25040
rect 390508 -25182 390848 -25096
rect 390508 -25238 390576 -25182
rect 390632 -25238 390718 -25182
rect 390774 -25238 390848 -25182
rect 390508 -25324 390848 -25238
rect 390508 -25380 390576 -25324
rect 390632 -25380 390718 -25324
rect 390774 -25380 390848 -25324
rect 390508 -25466 390848 -25380
rect 390508 -25522 390576 -25466
rect 390632 -25522 390718 -25466
rect 390774 -25522 390848 -25466
rect 390508 -25590 390848 -25522
rect 390908 -13680 391248 -13590
rect 390908 -13736 390980 -13680
rect 391036 -13736 391122 -13680
rect 391178 -13736 391248 -13680
rect 390908 -13822 391248 -13736
rect 390908 -13878 390980 -13822
rect 391036 -13878 391122 -13822
rect 391178 -13878 391248 -13822
rect 390908 -13964 391248 -13878
rect 390908 -14020 390980 -13964
rect 391036 -14020 391122 -13964
rect 391178 -14020 391248 -13964
rect 390908 -14106 391248 -14020
rect 390908 -14162 390980 -14106
rect 391036 -14162 391122 -14106
rect 391178 -14162 391248 -14106
rect 390908 -14248 391248 -14162
rect 390908 -14304 390980 -14248
rect 391036 -14304 391122 -14248
rect 391178 -14304 391248 -14248
rect 390908 -14390 391248 -14304
rect 390908 -14446 390980 -14390
rect 391036 -14446 391122 -14390
rect 391178 -14446 391248 -14390
rect 390908 -14532 391248 -14446
rect 390908 -14588 390980 -14532
rect 391036 -14588 391122 -14532
rect 391178 -14588 391248 -14532
rect 390908 -14674 391248 -14588
rect 390908 -14730 390980 -14674
rect 391036 -14730 391122 -14674
rect 391178 -14730 391248 -14674
rect 390908 -14816 391248 -14730
rect 390908 -14872 390980 -14816
rect 391036 -14872 391122 -14816
rect 391178 -14872 391248 -14816
rect 390908 -14958 391248 -14872
rect 390908 -15014 390980 -14958
rect 391036 -15014 391122 -14958
rect 391178 -15014 391248 -14958
rect 390908 -15100 391248 -15014
rect 390908 -15156 390980 -15100
rect 391036 -15156 391122 -15100
rect 391178 -15156 391248 -15100
rect 390908 -15242 391248 -15156
rect 390908 -15298 390980 -15242
rect 391036 -15298 391122 -15242
rect 391178 -15298 391248 -15242
rect 390908 -15384 391248 -15298
rect 390908 -15440 390980 -15384
rect 391036 -15440 391122 -15384
rect 391178 -15440 391248 -15384
rect 390908 -15526 391248 -15440
rect 390908 -15582 390980 -15526
rect 391036 -15582 391122 -15526
rect 391178 -15582 391248 -15526
rect 390908 -15668 391248 -15582
rect 390908 -15724 390980 -15668
rect 391036 -15724 391122 -15668
rect 391178 -15724 391248 -15668
rect 390908 -15810 391248 -15724
rect 390908 -15866 390980 -15810
rect 391036 -15866 391122 -15810
rect 391178 -15866 391248 -15810
rect 390908 -15952 391248 -15866
rect 390908 -16008 390980 -15952
rect 391036 -16008 391122 -15952
rect 391178 -16008 391248 -15952
rect 390908 -16094 391248 -16008
rect 390908 -16150 390980 -16094
rect 391036 -16150 391122 -16094
rect 391178 -16150 391248 -16094
rect 390908 -16236 391248 -16150
rect 390908 -16292 390980 -16236
rect 391036 -16292 391122 -16236
rect 391178 -16292 391248 -16236
rect 390908 -16378 391248 -16292
rect 390908 -16434 390980 -16378
rect 391036 -16434 391122 -16378
rect 391178 -16434 391248 -16378
rect 390908 -16520 391248 -16434
rect 390908 -16576 390980 -16520
rect 391036 -16576 391122 -16520
rect 391178 -16576 391248 -16520
rect 390908 -16662 391248 -16576
rect 390908 -16718 390980 -16662
rect 391036 -16718 391122 -16662
rect 391178 -16718 391248 -16662
rect 390908 -16804 391248 -16718
rect 390908 -16860 390980 -16804
rect 391036 -16860 391122 -16804
rect 391178 -16860 391248 -16804
rect 390908 -16946 391248 -16860
rect 390908 -17002 390980 -16946
rect 391036 -17002 391122 -16946
rect 391178 -17002 391248 -16946
rect 390908 -17088 391248 -17002
rect 390908 -17144 390980 -17088
rect 391036 -17144 391122 -17088
rect 391178 -17144 391248 -17088
rect 390908 -17230 391248 -17144
rect 390908 -17286 390980 -17230
rect 391036 -17286 391122 -17230
rect 391178 -17286 391248 -17230
rect 390908 -17372 391248 -17286
rect 390908 -17428 390980 -17372
rect 391036 -17428 391122 -17372
rect 391178 -17428 391248 -17372
rect 390908 -17514 391248 -17428
rect 390908 -17570 390980 -17514
rect 391036 -17570 391122 -17514
rect 391178 -17570 391248 -17514
rect 390908 -17656 391248 -17570
rect 390908 -17712 390980 -17656
rect 391036 -17712 391122 -17656
rect 391178 -17712 391248 -17656
rect 390908 -17798 391248 -17712
rect 390908 -17854 390980 -17798
rect 391036 -17854 391122 -17798
rect 391178 -17854 391248 -17798
rect 390908 -17940 391248 -17854
rect 390908 -17996 390980 -17940
rect 391036 -17996 391122 -17940
rect 391178 -17996 391248 -17940
rect 390908 -18082 391248 -17996
rect 390908 -18138 390980 -18082
rect 391036 -18138 391122 -18082
rect 391178 -18138 391248 -18082
rect 390908 -18224 391248 -18138
rect 390908 -18280 390980 -18224
rect 391036 -18280 391122 -18224
rect 391178 -18280 391248 -18224
rect 390908 -18366 391248 -18280
rect 390908 -18422 390980 -18366
rect 391036 -18422 391122 -18366
rect 391178 -18422 391248 -18366
rect 390908 -18508 391248 -18422
rect 390908 -18564 390980 -18508
rect 391036 -18564 391122 -18508
rect 391178 -18564 391248 -18508
rect 390908 -18650 391248 -18564
rect 390908 -18706 390980 -18650
rect 391036 -18706 391122 -18650
rect 391178 -18706 391248 -18650
rect 390908 -18792 391248 -18706
rect 390908 -18848 390980 -18792
rect 391036 -18848 391122 -18792
rect 391178 -18848 391248 -18792
rect 390908 -18934 391248 -18848
rect 390908 -18990 390980 -18934
rect 391036 -18990 391122 -18934
rect 391178 -18990 391248 -18934
rect 390908 -19076 391248 -18990
rect 390908 -19132 390980 -19076
rect 391036 -19132 391122 -19076
rect 391178 -19132 391248 -19076
rect 390908 -19218 391248 -19132
rect 390908 -19274 390980 -19218
rect 391036 -19274 391122 -19218
rect 391178 -19274 391248 -19218
rect 390908 -19360 391248 -19274
rect 390908 -19416 390980 -19360
rect 391036 -19416 391122 -19360
rect 391178 -19416 391248 -19360
rect 390908 -19502 391248 -19416
rect 390908 -19558 390980 -19502
rect 391036 -19558 391122 -19502
rect 391178 -19558 391248 -19502
rect 390908 -19644 391248 -19558
rect 390908 -19700 390980 -19644
rect 391036 -19700 391122 -19644
rect 391178 -19700 391248 -19644
rect 390908 -19786 391248 -19700
rect 390908 -19842 390980 -19786
rect 391036 -19842 391122 -19786
rect 391178 -19842 391248 -19786
rect 390908 -19928 391248 -19842
rect 390908 -19984 390980 -19928
rect 391036 -19984 391122 -19928
rect 391178 -19984 391248 -19928
rect 390908 -20070 391248 -19984
rect 390908 -20126 390980 -20070
rect 391036 -20126 391122 -20070
rect 391178 -20126 391248 -20070
rect 390908 -20212 391248 -20126
rect 390908 -20268 390980 -20212
rect 391036 -20268 391122 -20212
rect 391178 -20268 391248 -20212
rect 390908 -20354 391248 -20268
rect 390908 -20410 390980 -20354
rect 391036 -20410 391122 -20354
rect 391178 -20410 391248 -20354
rect 390908 -20496 391248 -20410
rect 390908 -20552 390980 -20496
rect 391036 -20552 391122 -20496
rect 391178 -20552 391248 -20496
rect 390908 -20638 391248 -20552
rect 390908 -20694 390980 -20638
rect 391036 -20694 391122 -20638
rect 391178 -20694 391248 -20638
rect 390908 -20780 391248 -20694
rect 390908 -20836 390980 -20780
rect 391036 -20836 391122 -20780
rect 391178 -20836 391248 -20780
rect 390908 -20922 391248 -20836
rect 390908 -20978 390980 -20922
rect 391036 -20978 391122 -20922
rect 391178 -20978 391248 -20922
rect 390908 -21064 391248 -20978
rect 390908 -21120 390980 -21064
rect 391036 -21120 391122 -21064
rect 391178 -21120 391248 -21064
rect 390908 -21206 391248 -21120
rect 390908 -21262 390980 -21206
rect 391036 -21262 391122 -21206
rect 391178 -21262 391248 -21206
rect 390908 -21348 391248 -21262
rect 390908 -21404 390980 -21348
rect 391036 -21404 391122 -21348
rect 391178 -21404 391248 -21348
rect 390908 -21490 391248 -21404
rect 390908 -21546 390980 -21490
rect 391036 -21546 391122 -21490
rect 391178 -21546 391248 -21490
rect 390908 -21632 391248 -21546
rect 390908 -21688 390980 -21632
rect 391036 -21688 391122 -21632
rect 391178 -21688 391248 -21632
rect 390908 -21774 391248 -21688
rect 390908 -21830 390980 -21774
rect 391036 -21830 391122 -21774
rect 391178 -21830 391248 -21774
rect 390908 -21916 391248 -21830
rect 390908 -21972 390980 -21916
rect 391036 -21972 391122 -21916
rect 391178 -21972 391248 -21916
rect 390908 -22058 391248 -21972
rect 390908 -22114 390980 -22058
rect 391036 -22114 391122 -22058
rect 391178 -22114 391248 -22058
rect 390908 -22200 391248 -22114
rect 390908 -22256 390980 -22200
rect 391036 -22256 391122 -22200
rect 391178 -22256 391248 -22200
rect 390908 -22342 391248 -22256
rect 390908 -22398 390980 -22342
rect 391036 -22398 391122 -22342
rect 391178 -22398 391248 -22342
rect 390908 -22484 391248 -22398
rect 390908 -22540 390980 -22484
rect 391036 -22540 391122 -22484
rect 391178 -22540 391248 -22484
rect 390908 -22626 391248 -22540
rect 390908 -22682 390980 -22626
rect 391036 -22682 391122 -22626
rect 391178 -22682 391248 -22626
rect 390908 -22768 391248 -22682
rect 390908 -22824 390980 -22768
rect 391036 -22824 391122 -22768
rect 391178 -22824 391248 -22768
rect 390908 -22910 391248 -22824
rect 390908 -22966 390980 -22910
rect 391036 -22966 391122 -22910
rect 391178 -22966 391248 -22910
rect 390908 -23052 391248 -22966
rect 390908 -23108 390980 -23052
rect 391036 -23108 391122 -23052
rect 391178 -23108 391248 -23052
rect 390908 -23194 391248 -23108
rect 390908 -23250 390980 -23194
rect 391036 -23250 391122 -23194
rect 391178 -23250 391248 -23194
rect 390908 -23336 391248 -23250
rect 390908 -23392 390980 -23336
rect 391036 -23392 391122 -23336
rect 391178 -23392 391248 -23336
rect 390908 -23478 391248 -23392
rect 390908 -23534 390980 -23478
rect 391036 -23534 391122 -23478
rect 391178 -23534 391248 -23478
rect 390908 -23620 391248 -23534
rect 390908 -23676 390980 -23620
rect 391036 -23676 391122 -23620
rect 391178 -23676 391248 -23620
rect 390908 -23762 391248 -23676
rect 390908 -23818 390980 -23762
rect 391036 -23818 391122 -23762
rect 391178 -23818 391248 -23762
rect 390908 -23904 391248 -23818
rect 390908 -23960 390980 -23904
rect 391036 -23960 391122 -23904
rect 391178 -23960 391248 -23904
rect 390908 -24046 391248 -23960
rect 390908 -24102 390980 -24046
rect 391036 -24102 391122 -24046
rect 391178 -24102 391248 -24046
rect 390908 -24188 391248 -24102
rect 390908 -24244 390980 -24188
rect 391036 -24244 391122 -24188
rect 391178 -24244 391248 -24188
rect 390908 -24330 391248 -24244
rect 390908 -24386 390980 -24330
rect 391036 -24386 391122 -24330
rect 391178 -24386 391248 -24330
rect 390908 -24472 391248 -24386
rect 390908 -24528 390980 -24472
rect 391036 -24528 391122 -24472
rect 391178 -24528 391248 -24472
rect 390908 -24614 391248 -24528
rect 390908 -24670 390980 -24614
rect 391036 -24670 391122 -24614
rect 391178 -24670 391248 -24614
rect 390908 -24756 391248 -24670
rect 390908 -24812 390980 -24756
rect 391036 -24812 391122 -24756
rect 391178 -24812 391248 -24756
rect 390908 -24898 391248 -24812
rect 390908 -24954 390980 -24898
rect 391036 -24954 391122 -24898
rect 391178 -24954 391248 -24898
rect 390908 -25040 391248 -24954
rect 390908 -25096 390980 -25040
rect 391036 -25096 391122 -25040
rect 391178 -25096 391248 -25040
rect 390908 -25182 391248 -25096
rect 390908 -25238 390980 -25182
rect 391036 -25238 391122 -25182
rect 391178 -25238 391248 -25182
rect 390908 -25324 391248 -25238
rect 390908 -25380 390980 -25324
rect 391036 -25380 391122 -25324
rect 391178 -25380 391248 -25324
rect 390908 -25466 391248 -25380
rect 390908 -25522 390980 -25466
rect 391036 -25522 391122 -25466
rect 391178 -25522 391248 -25466
rect 390908 -25590 391248 -25522
rect 391308 -13680 391648 -13590
rect 391308 -13736 391376 -13680
rect 391432 -13736 391518 -13680
rect 391574 -13736 391648 -13680
rect 391308 -13822 391648 -13736
rect 391308 -13878 391376 -13822
rect 391432 -13878 391518 -13822
rect 391574 -13878 391648 -13822
rect 391308 -13964 391648 -13878
rect 391308 -14020 391376 -13964
rect 391432 -14020 391518 -13964
rect 391574 -14020 391648 -13964
rect 391308 -14106 391648 -14020
rect 391308 -14162 391376 -14106
rect 391432 -14162 391518 -14106
rect 391574 -14162 391648 -14106
rect 391308 -14248 391648 -14162
rect 391308 -14304 391376 -14248
rect 391432 -14304 391518 -14248
rect 391574 -14304 391648 -14248
rect 391308 -14390 391648 -14304
rect 391308 -14446 391376 -14390
rect 391432 -14446 391518 -14390
rect 391574 -14446 391648 -14390
rect 391308 -14532 391648 -14446
rect 391308 -14588 391376 -14532
rect 391432 -14588 391518 -14532
rect 391574 -14588 391648 -14532
rect 391308 -14674 391648 -14588
rect 391308 -14730 391376 -14674
rect 391432 -14730 391518 -14674
rect 391574 -14730 391648 -14674
rect 391308 -14816 391648 -14730
rect 391308 -14872 391376 -14816
rect 391432 -14872 391518 -14816
rect 391574 -14872 391648 -14816
rect 391308 -14958 391648 -14872
rect 391308 -15014 391376 -14958
rect 391432 -15014 391518 -14958
rect 391574 -15014 391648 -14958
rect 391308 -15100 391648 -15014
rect 391308 -15156 391376 -15100
rect 391432 -15156 391518 -15100
rect 391574 -15156 391648 -15100
rect 391308 -15242 391648 -15156
rect 391308 -15298 391376 -15242
rect 391432 -15298 391518 -15242
rect 391574 -15298 391648 -15242
rect 391308 -15384 391648 -15298
rect 391308 -15440 391376 -15384
rect 391432 -15440 391518 -15384
rect 391574 -15440 391648 -15384
rect 391308 -15526 391648 -15440
rect 391308 -15582 391376 -15526
rect 391432 -15582 391518 -15526
rect 391574 -15582 391648 -15526
rect 391308 -15668 391648 -15582
rect 391308 -15724 391376 -15668
rect 391432 -15724 391518 -15668
rect 391574 -15724 391648 -15668
rect 391308 -15810 391648 -15724
rect 391308 -15866 391376 -15810
rect 391432 -15866 391518 -15810
rect 391574 -15866 391648 -15810
rect 391308 -15952 391648 -15866
rect 391308 -16008 391376 -15952
rect 391432 -16008 391518 -15952
rect 391574 -16008 391648 -15952
rect 391308 -16094 391648 -16008
rect 391308 -16150 391376 -16094
rect 391432 -16150 391518 -16094
rect 391574 -16150 391648 -16094
rect 391308 -16236 391648 -16150
rect 391308 -16292 391376 -16236
rect 391432 -16292 391518 -16236
rect 391574 -16292 391648 -16236
rect 391308 -16378 391648 -16292
rect 391308 -16434 391376 -16378
rect 391432 -16434 391518 -16378
rect 391574 -16434 391648 -16378
rect 391308 -16520 391648 -16434
rect 391308 -16576 391376 -16520
rect 391432 -16576 391518 -16520
rect 391574 -16576 391648 -16520
rect 391308 -16662 391648 -16576
rect 391308 -16718 391376 -16662
rect 391432 -16718 391518 -16662
rect 391574 -16718 391648 -16662
rect 391308 -16804 391648 -16718
rect 391308 -16860 391376 -16804
rect 391432 -16860 391518 -16804
rect 391574 -16860 391648 -16804
rect 391308 -16946 391648 -16860
rect 391308 -17002 391376 -16946
rect 391432 -17002 391518 -16946
rect 391574 -17002 391648 -16946
rect 391308 -17088 391648 -17002
rect 391308 -17144 391376 -17088
rect 391432 -17144 391518 -17088
rect 391574 -17144 391648 -17088
rect 391308 -17230 391648 -17144
rect 391308 -17286 391376 -17230
rect 391432 -17286 391518 -17230
rect 391574 -17286 391648 -17230
rect 391308 -17372 391648 -17286
rect 391308 -17428 391376 -17372
rect 391432 -17428 391518 -17372
rect 391574 -17428 391648 -17372
rect 391308 -17514 391648 -17428
rect 391308 -17570 391376 -17514
rect 391432 -17570 391518 -17514
rect 391574 -17570 391648 -17514
rect 391308 -17656 391648 -17570
rect 391308 -17712 391376 -17656
rect 391432 -17712 391518 -17656
rect 391574 -17712 391648 -17656
rect 391308 -17798 391648 -17712
rect 391308 -17854 391376 -17798
rect 391432 -17854 391518 -17798
rect 391574 -17854 391648 -17798
rect 391308 -17940 391648 -17854
rect 391308 -17996 391376 -17940
rect 391432 -17996 391518 -17940
rect 391574 -17996 391648 -17940
rect 391308 -18082 391648 -17996
rect 391308 -18138 391376 -18082
rect 391432 -18138 391518 -18082
rect 391574 -18138 391648 -18082
rect 391308 -18224 391648 -18138
rect 391308 -18280 391376 -18224
rect 391432 -18280 391518 -18224
rect 391574 -18280 391648 -18224
rect 391308 -18366 391648 -18280
rect 391308 -18422 391376 -18366
rect 391432 -18422 391518 -18366
rect 391574 -18422 391648 -18366
rect 391308 -18508 391648 -18422
rect 391308 -18564 391376 -18508
rect 391432 -18564 391518 -18508
rect 391574 -18564 391648 -18508
rect 391308 -18650 391648 -18564
rect 391308 -18706 391376 -18650
rect 391432 -18706 391518 -18650
rect 391574 -18706 391648 -18650
rect 391308 -18792 391648 -18706
rect 391308 -18848 391376 -18792
rect 391432 -18848 391518 -18792
rect 391574 -18848 391648 -18792
rect 391308 -18934 391648 -18848
rect 391308 -18990 391376 -18934
rect 391432 -18990 391518 -18934
rect 391574 -18990 391648 -18934
rect 391308 -19076 391648 -18990
rect 391308 -19132 391376 -19076
rect 391432 -19132 391518 -19076
rect 391574 -19132 391648 -19076
rect 391308 -19218 391648 -19132
rect 391308 -19274 391376 -19218
rect 391432 -19274 391518 -19218
rect 391574 -19274 391648 -19218
rect 391308 -19360 391648 -19274
rect 391308 -19416 391376 -19360
rect 391432 -19416 391518 -19360
rect 391574 -19416 391648 -19360
rect 391308 -19502 391648 -19416
rect 391308 -19558 391376 -19502
rect 391432 -19558 391518 -19502
rect 391574 -19558 391648 -19502
rect 391308 -19644 391648 -19558
rect 391308 -19700 391376 -19644
rect 391432 -19700 391518 -19644
rect 391574 -19700 391648 -19644
rect 391308 -19786 391648 -19700
rect 391308 -19842 391376 -19786
rect 391432 -19842 391518 -19786
rect 391574 -19842 391648 -19786
rect 391308 -19928 391648 -19842
rect 391308 -19984 391376 -19928
rect 391432 -19984 391518 -19928
rect 391574 -19984 391648 -19928
rect 391308 -20070 391648 -19984
rect 391308 -20126 391376 -20070
rect 391432 -20126 391518 -20070
rect 391574 -20126 391648 -20070
rect 391308 -20212 391648 -20126
rect 391308 -20268 391376 -20212
rect 391432 -20268 391518 -20212
rect 391574 -20268 391648 -20212
rect 391308 -20354 391648 -20268
rect 391308 -20410 391376 -20354
rect 391432 -20410 391518 -20354
rect 391574 -20410 391648 -20354
rect 391308 -20496 391648 -20410
rect 391308 -20552 391376 -20496
rect 391432 -20552 391518 -20496
rect 391574 -20552 391648 -20496
rect 391308 -20638 391648 -20552
rect 391308 -20694 391376 -20638
rect 391432 -20694 391518 -20638
rect 391574 -20694 391648 -20638
rect 391308 -20780 391648 -20694
rect 391308 -20836 391376 -20780
rect 391432 -20836 391518 -20780
rect 391574 -20836 391648 -20780
rect 391308 -20922 391648 -20836
rect 391308 -20978 391376 -20922
rect 391432 -20978 391518 -20922
rect 391574 -20978 391648 -20922
rect 391308 -21064 391648 -20978
rect 391308 -21120 391376 -21064
rect 391432 -21120 391518 -21064
rect 391574 -21120 391648 -21064
rect 391308 -21206 391648 -21120
rect 391308 -21262 391376 -21206
rect 391432 -21262 391518 -21206
rect 391574 -21262 391648 -21206
rect 391308 -21348 391648 -21262
rect 391308 -21404 391376 -21348
rect 391432 -21404 391518 -21348
rect 391574 -21404 391648 -21348
rect 391308 -21490 391648 -21404
rect 391308 -21546 391376 -21490
rect 391432 -21546 391518 -21490
rect 391574 -21546 391648 -21490
rect 391308 -21632 391648 -21546
rect 391308 -21688 391376 -21632
rect 391432 -21688 391518 -21632
rect 391574 -21688 391648 -21632
rect 391308 -21774 391648 -21688
rect 391308 -21830 391376 -21774
rect 391432 -21830 391518 -21774
rect 391574 -21830 391648 -21774
rect 391308 -21916 391648 -21830
rect 391308 -21972 391376 -21916
rect 391432 -21972 391518 -21916
rect 391574 -21972 391648 -21916
rect 391308 -22058 391648 -21972
rect 391308 -22114 391376 -22058
rect 391432 -22114 391518 -22058
rect 391574 -22114 391648 -22058
rect 391308 -22200 391648 -22114
rect 391308 -22256 391376 -22200
rect 391432 -22256 391518 -22200
rect 391574 -22256 391648 -22200
rect 391308 -22342 391648 -22256
rect 391308 -22398 391376 -22342
rect 391432 -22398 391518 -22342
rect 391574 -22398 391648 -22342
rect 391308 -22484 391648 -22398
rect 391308 -22540 391376 -22484
rect 391432 -22540 391518 -22484
rect 391574 -22540 391648 -22484
rect 391308 -22626 391648 -22540
rect 391308 -22682 391376 -22626
rect 391432 -22682 391518 -22626
rect 391574 -22682 391648 -22626
rect 391308 -22768 391648 -22682
rect 391308 -22824 391376 -22768
rect 391432 -22824 391518 -22768
rect 391574 -22824 391648 -22768
rect 391308 -22910 391648 -22824
rect 391308 -22966 391376 -22910
rect 391432 -22966 391518 -22910
rect 391574 -22966 391648 -22910
rect 391308 -23052 391648 -22966
rect 391308 -23108 391376 -23052
rect 391432 -23108 391518 -23052
rect 391574 -23108 391648 -23052
rect 391308 -23194 391648 -23108
rect 391308 -23250 391376 -23194
rect 391432 -23250 391518 -23194
rect 391574 -23250 391648 -23194
rect 391308 -23336 391648 -23250
rect 391308 -23392 391376 -23336
rect 391432 -23392 391518 -23336
rect 391574 -23392 391648 -23336
rect 391308 -23478 391648 -23392
rect 391308 -23534 391376 -23478
rect 391432 -23534 391518 -23478
rect 391574 -23534 391648 -23478
rect 391308 -23620 391648 -23534
rect 391308 -23676 391376 -23620
rect 391432 -23676 391518 -23620
rect 391574 -23676 391648 -23620
rect 391308 -23762 391648 -23676
rect 391308 -23818 391376 -23762
rect 391432 -23818 391518 -23762
rect 391574 -23818 391648 -23762
rect 391308 -23904 391648 -23818
rect 391308 -23960 391376 -23904
rect 391432 -23960 391518 -23904
rect 391574 -23960 391648 -23904
rect 391308 -24046 391648 -23960
rect 391308 -24102 391376 -24046
rect 391432 -24102 391518 -24046
rect 391574 -24102 391648 -24046
rect 391308 -24188 391648 -24102
rect 391308 -24244 391376 -24188
rect 391432 -24244 391518 -24188
rect 391574 -24244 391648 -24188
rect 391308 -24330 391648 -24244
rect 391308 -24386 391376 -24330
rect 391432 -24386 391518 -24330
rect 391574 -24386 391648 -24330
rect 391308 -24472 391648 -24386
rect 391308 -24528 391376 -24472
rect 391432 -24528 391518 -24472
rect 391574 -24528 391648 -24472
rect 391308 -24614 391648 -24528
rect 391308 -24670 391376 -24614
rect 391432 -24670 391518 -24614
rect 391574 -24670 391648 -24614
rect 391308 -24756 391648 -24670
rect 391308 -24812 391376 -24756
rect 391432 -24812 391518 -24756
rect 391574 -24812 391648 -24756
rect 391308 -24898 391648 -24812
rect 391308 -24954 391376 -24898
rect 391432 -24954 391518 -24898
rect 391574 -24954 391648 -24898
rect 391308 -25040 391648 -24954
rect 391308 -25096 391376 -25040
rect 391432 -25096 391518 -25040
rect 391574 -25096 391648 -25040
rect 391308 -25182 391648 -25096
rect 391308 -25238 391376 -25182
rect 391432 -25238 391518 -25182
rect 391574 -25238 391648 -25182
rect 391308 -25324 391648 -25238
rect 391308 -25380 391376 -25324
rect 391432 -25380 391518 -25324
rect 391574 -25380 391648 -25324
rect 391308 -25466 391648 -25380
rect 391308 -25522 391376 -25466
rect 391432 -25522 391518 -25466
rect 391574 -25522 391648 -25466
rect 391308 -25590 391648 -25522
rect 391708 -13680 392048 -13590
rect 391708 -13736 391776 -13680
rect 391832 -13736 391918 -13680
rect 391974 -13736 392048 -13680
rect 391708 -13822 392048 -13736
rect 391708 -13878 391776 -13822
rect 391832 -13878 391918 -13822
rect 391974 -13878 392048 -13822
rect 391708 -13964 392048 -13878
rect 391708 -14020 391776 -13964
rect 391832 -14020 391918 -13964
rect 391974 -14020 392048 -13964
rect 391708 -14106 392048 -14020
rect 391708 -14162 391776 -14106
rect 391832 -14162 391918 -14106
rect 391974 -14162 392048 -14106
rect 391708 -14248 392048 -14162
rect 391708 -14304 391776 -14248
rect 391832 -14304 391918 -14248
rect 391974 -14304 392048 -14248
rect 391708 -14390 392048 -14304
rect 391708 -14446 391776 -14390
rect 391832 -14446 391918 -14390
rect 391974 -14446 392048 -14390
rect 391708 -14532 392048 -14446
rect 391708 -14588 391776 -14532
rect 391832 -14588 391918 -14532
rect 391974 -14588 392048 -14532
rect 391708 -14674 392048 -14588
rect 391708 -14730 391776 -14674
rect 391832 -14730 391918 -14674
rect 391974 -14730 392048 -14674
rect 391708 -14816 392048 -14730
rect 391708 -14872 391776 -14816
rect 391832 -14872 391918 -14816
rect 391974 -14872 392048 -14816
rect 391708 -14958 392048 -14872
rect 391708 -15014 391776 -14958
rect 391832 -15014 391918 -14958
rect 391974 -15014 392048 -14958
rect 391708 -15100 392048 -15014
rect 391708 -15156 391776 -15100
rect 391832 -15156 391918 -15100
rect 391974 -15156 392048 -15100
rect 391708 -15242 392048 -15156
rect 391708 -15298 391776 -15242
rect 391832 -15298 391918 -15242
rect 391974 -15298 392048 -15242
rect 391708 -15384 392048 -15298
rect 391708 -15440 391776 -15384
rect 391832 -15440 391918 -15384
rect 391974 -15440 392048 -15384
rect 391708 -15526 392048 -15440
rect 391708 -15582 391776 -15526
rect 391832 -15582 391918 -15526
rect 391974 -15582 392048 -15526
rect 391708 -15668 392048 -15582
rect 391708 -15724 391776 -15668
rect 391832 -15724 391918 -15668
rect 391974 -15724 392048 -15668
rect 391708 -15810 392048 -15724
rect 391708 -15866 391776 -15810
rect 391832 -15866 391918 -15810
rect 391974 -15866 392048 -15810
rect 391708 -15952 392048 -15866
rect 391708 -16008 391776 -15952
rect 391832 -16008 391918 -15952
rect 391974 -16008 392048 -15952
rect 391708 -16094 392048 -16008
rect 391708 -16150 391776 -16094
rect 391832 -16150 391918 -16094
rect 391974 -16150 392048 -16094
rect 391708 -16236 392048 -16150
rect 391708 -16292 391776 -16236
rect 391832 -16292 391918 -16236
rect 391974 -16292 392048 -16236
rect 391708 -16378 392048 -16292
rect 391708 -16434 391776 -16378
rect 391832 -16434 391918 -16378
rect 391974 -16434 392048 -16378
rect 391708 -16520 392048 -16434
rect 391708 -16576 391776 -16520
rect 391832 -16576 391918 -16520
rect 391974 -16576 392048 -16520
rect 391708 -16662 392048 -16576
rect 391708 -16718 391776 -16662
rect 391832 -16718 391918 -16662
rect 391974 -16718 392048 -16662
rect 391708 -16804 392048 -16718
rect 391708 -16860 391776 -16804
rect 391832 -16860 391918 -16804
rect 391974 -16860 392048 -16804
rect 391708 -16946 392048 -16860
rect 391708 -17002 391776 -16946
rect 391832 -17002 391918 -16946
rect 391974 -17002 392048 -16946
rect 391708 -17088 392048 -17002
rect 391708 -17144 391776 -17088
rect 391832 -17144 391918 -17088
rect 391974 -17144 392048 -17088
rect 391708 -17230 392048 -17144
rect 391708 -17286 391776 -17230
rect 391832 -17286 391918 -17230
rect 391974 -17286 392048 -17230
rect 391708 -17372 392048 -17286
rect 391708 -17428 391776 -17372
rect 391832 -17428 391918 -17372
rect 391974 -17428 392048 -17372
rect 391708 -17514 392048 -17428
rect 391708 -17570 391776 -17514
rect 391832 -17570 391918 -17514
rect 391974 -17570 392048 -17514
rect 391708 -17656 392048 -17570
rect 391708 -17712 391776 -17656
rect 391832 -17712 391918 -17656
rect 391974 -17712 392048 -17656
rect 391708 -17798 392048 -17712
rect 391708 -17854 391776 -17798
rect 391832 -17854 391918 -17798
rect 391974 -17854 392048 -17798
rect 391708 -17940 392048 -17854
rect 391708 -17996 391776 -17940
rect 391832 -17996 391918 -17940
rect 391974 -17996 392048 -17940
rect 391708 -18082 392048 -17996
rect 391708 -18138 391776 -18082
rect 391832 -18138 391918 -18082
rect 391974 -18138 392048 -18082
rect 391708 -18224 392048 -18138
rect 391708 -18280 391776 -18224
rect 391832 -18280 391918 -18224
rect 391974 -18280 392048 -18224
rect 391708 -18366 392048 -18280
rect 391708 -18422 391776 -18366
rect 391832 -18422 391918 -18366
rect 391974 -18422 392048 -18366
rect 391708 -18508 392048 -18422
rect 391708 -18564 391776 -18508
rect 391832 -18564 391918 -18508
rect 391974 -18564 392048 -18508
rect 391708 -18650 392048 -18564
rect 391708 -18706 391776 -18650
rect 391832 -18706 391918 -18650
rect 391974 -18706 392048 -18650
rect 391708 -18792 392048 -18706
rect 391708 -18848 391776 -18792
rect 391832 -18848 391918 -18792
rect 391974 -18848 392048 -18792
rect 391708 -18934 392048 -18848
rect 391708 -18990 391776 -18934
rect 391832 -18990 391918 -18934
rect 391974 -18990 392048 -18934
rect 391708 -19076 392048 -18990
rect 391708 -19132 391776 -19076
rect 391832 -19132 391918 -19076
rect 391974 -19132 392048 -19076
rect 391708 -19218 392048 -19132
rect 391708 -19274 391776 -19218
rect 391832 -19274 391918 -19218
rect 391974 -19274 392048 -19218
rect 391708 -19360 392048 -19274
rect 391708 -19416 391776 -19360
rect 391832 -19416 391918 -19360
rect 391974 -19416 392048 -19360
rect 391708 -19502 392048 -19416
rect 391708 -19558 391776 -19502
rect 391832 -19558 391918 -19502
rect 391974 -19558 392048 -19502
rect 391708 -19644 392048 -19558
rect 391708 -19700 391776 -19644
rect 391832 -19700 391918 -19644
rect 391974 -19700 392048 -19644
rect 391708 -19786 392048 -19700
rect 391708 -19842 391776 -19786
rect 391832 -19842 391918 -19786
rect 391974 -19842 392048 -19786
rect 391708 -19928 392048 -19842
rect 391708 -19984 391776 -19928
rect 391832 -19984 391918 -19928
rect 391974 -19984 392048 -19928
rect 391708 -20070 392048 -19984
rect 391708 -20126 391776 -20070
rect 391832 -20126 391918 -20070
rect 391974 -20126 392048 -20070
rect 391708 -20212 392048 -20126
rect 391708 -20268 391776 -20212
rect 391832 -20268 391918 -20212
rect 391974 -20268 392048 -20212
rect 391708 -20354 392048 -20268
rect 391708 -20410 391776 -20354
rect 391832 -20410 391918 -20354
rect 391974 -20410 392048 -20354
rect 391708 -20496 392048 -20410
rect 391708 -20552 391776 -20496
rect 391832 -20552 391918 -20496
rect 391974 -20552 392048 -20496
rect 391708 -20638 392048 -20552
rect 391708 -20694 391776 -20638
rect 391832 -20694 391918 -20638
rect 391974 -20694 392048 -20638
rect 391708 -20780 392048 -20694
rect 391708 -20836 391776 -20780
rect 391832 -20836 391918 -20780
rect 391974 -20836 392048 -20780
rect 391708 -20922 392048 -20836
rect 391708 -20978 391776 -20922
rect 391832 -20978 391918 -20922
rect 391974 -20978 392048 -20922
rect 391708 -21064 392048 -20978
rect 391708 -21120 391776 -21064
rect 391832 -21120 391918 -21064
rect 391974 -21120 392048 -21064
rect 391708 -21206 392048 -21120
rect 391708 -21262 391776 -21206
rect 391832 -21262 391918 -21206
rect 391974 -21262 392048 -21206
rect 391708 -21348 392048 -21262
rect 391708 -21404 391776 -21348
rect 391832 -21404 391918 -21348
rect 391974 -21404 392048 -21348
rect 391708 -21490 392048 -21404
rect 391708 -21546 391776 -21490
rect 391832 -21546 391918 -21490
rect 391974 -21546 392048 -21490
rect 391708 -21632 392048 -21546
rect 391708 -21688 391776 -21632
rect 391832 -21688 391918 -21632
rect 391974 -21688 392048 -21632
rect 391708 -21774 392048 -21688
rect 391708 -21830 391776 -21774
rect 391832 -21830 391918 -21774
rect 391974 -21830 392048 -21774
rect 391708 -21916 392048 -21830
rect 391708 -21972 391776 -21916
rect 391832 -21972 391918 -21916
rect 391974 -21972 392048 -21916
rect 391708 -22058 392048 -21972
rect 391708 -22114 391776 -22058
rect 391832 -22114 391918 -22058
rect 391974 -22114 392048 -22058
rect 391708 -22200 392048 -22114
rect 391708 -22256 391776 -22200
rect 391832 -22256 391918 -22200
rect 391974 -22256 392048 -22200
rect 391708 -22342 392048 -22256
rect 391708 -22398 391776 -22342
rect 391832 -22398 391918 -22342
rect 391974 -22398 392048 -22342
rect 391708 -22484 392048 -22398
rect 391708 -22540 391776 -22484
rect 391832 -22540 391918 -22484
rect 391974 -22540 392048 -22484
rect 391708 -22626 392048 -22540
rect 391708 -22682 391776 -22626
rect 391832 -22682 391918 -22626
rect 391974 -22682 392048 -22626
rect 391708 -22768 392048 -22682
rect 391708 -22824 391776 -22768
rect 391832 -22824 391918 -22768
rect 391974 -22824 392048 -22768
rect 391708 -22910 392048 -22824
rect 391708 -22966 391776 -22910
rect 391832 -22966 391918 -22910
rect 391974 -22966 392048 -22910
rect 391708 -23052 392048 -22966
rect 391708 -23108 391776 -23052
rect 391832 -23108 391918 -23052
rect 391974 -23108 392048 -23052
rect 391708 -23194 392048 -23108
rect 391708 -23250 391776 -23194
rect 391832 -23250 391918 -23194
rect 391974 -23250 392048 -23194
rect 391708 -23336 392048 -23250
rect 391708 -23392 391776 -23336
rect 391832 -23392 391918 -23336
rect 391974 -23392 392048 -23336
rect 391708 -23478 392048 -23392
rect 391708 -23534 391776 -23478
rect 391832 -23534 391918 -23478
rect 391974 -23534 392048 -23478
rect 391708 -23620 392048 -23534
rect 391708 -23676 391776 -23620
rect 391832 -23676 391918 -23620
rect 391974 -23676 392048 -23620
rect 391708 -23762 392048 -23676
rect 391708 -23818 391776 -23762
rect 391832 -23818 391918 -23762
rect 391974 -23818 392048 -23762
rect 391708 -23904 392048 -23818
rect 391708 -23960 391776 -23904
rect 391832 -23960 391918 -23904
rect 391974 -23960 392048 -23904
rect 391708 -24046 392048 -23960
rect 391708 -24102 391776 -24046
rect 391832 -24102 391918 -24046
rect 391974 -24102 392048 -24046
rect 391708 -24188 392048 -24102
rect 391708 -24244 391776 -24188
rect 391832 -24244 391918 -24188
rect 391974 -24244 392048 -24188
rect 391708 -24330 392048 -24244
rect 391708 -24386 391776 -24330
rect 391832 -24386 391918 -24330
rect 391974 -24386 392048 -24330
rect 391708 -24472 392048 -24386
rect 391708 -24528 391776 -24472
rect 391832 -24528 391918 -24472
rect 391974 -24528 392048 -24472
rect 391708 -24614 392048 -24528
rect 391708 -24670 391776 -24614
rect 391832 -24670 391918 -24614
rect 391974 -24670 392048 -24614
rect 391708 -24756 392048 -24670
rect 391708 -24812 391776 -24756
rect 391832 -24812 391918 -24756
rect 391974 -24812 392048 -24756
rect 391708 -24898 392048 -24812
rect 391708 -24954 391776 -24898
rect 391832 -24954 391918 -24898
rect 391974 -24954 392048 -24898
rect 391708 -25040 392048 -24954
rect 391708 -25096 391776 -25040
rect 391832 -25096 391918 -25040
rect 391974 -25096 392048 -25040
rect 391708 -25182 392048 -25096
rect 391708 -25238 391776 -25182
rect 391832 -25238 391918 -25182
rect 391974 -25238 392048 -25182
rect 391708 -25324 392048 -25238
rect 391708 -25380 391776 -25324
rect 391832 -25380 391918 -25324
rect 391974 -25380 392048 -25324
rect 391708 -25466 392048 -25380
rect 391708 -25522 391776 -25466
rect 391832 -25522 391918 -25466
rect 391974 -25522 392048 -25466
rect 391708 -25590 392048 -25522
rect 392108 -13680 392448 -13590
rect 392108 -13736 392173 -13680
rect 392229 -13736 392315 -13680
rect 392371 -13736 392448 -13680
rect 392108 -13822 392448 -13736
rect 392108 -13878 392173 -13822
rect 392229 -13878 392315 -13822
rect 392371 -13878 392448 -13822
rect 392108 -13964 392448 -13878
rect 392108 -14020 392173 -13964
rect 392229 -14020 392315 -13964
rect 392371 -14020 392448 -13964
rect 392108 -14106 392448 -14020
rect 392108 -14162 392173 -14106
rect 392229 -14162 392315 -14106
rect 392371 -14162 392448 -14106
rect 392108 -14248 392448 -14162
rect 392108 -14304 392173 -14248
rect 392229 -14304 392315 -14248
rect 392371 -14304 392448 -14248
rect 392108 -14390 392448 -14304
rect 392108 -14446 392173 -14390
rect 392229 -14446 392315 -14390
rect 392371 -14446 392448 -14390
rect 392108 -14532 392448 -14446
rect 392108 -14588 392173 -14532
rect 392229 -14588 392315 -14532
rect 392371 -14588 392448 -14532
rect 392108 -14674 392448 -14588
rect 392108 -14730 392173 -14674
rect 392229 -14730 392315 -14674
rect 392371 -14730 392448 -14674
rect 392108 -14816 392448 -14730
rect 392108 -14872 392173 -14816
rect 392229 -14872 392315 -14816
rect 392371 -14872 392448 -14816
rect 392108 -14958 392448 -14872
rect 392108 -15014 392173 -14958
rect 392229 -15014 392315 -14958
rect 392371 -15014 392448 -14958
rect 392108 -15100 392448 -15014
rect 392108 -15156 392173 -15100
rect 392229 -15156 392315 -15100
rect 392371 -15156 392448 -15100
rect 392108 -15242 392448 -15156
rect 392108 -15298 392173 -15242
rect 392229 -15298 392315 -15242
rect 392371 -15298 392448 -15242
rect 392108 -15384 392448 -15298
rect 392108 -15440 392173 -15384
rect 392229 -15440 392315 -15384
rect 392371 -15440 392448 -15384
rect 392108 -15526 392448 -15440
rect 392108 -15582 392173 -15526
rect 392229 -15582 392315 -15526
rect 392371 -15582 392448 -15526
rect 392108 -15668 392448 -15582
rect 392108 -15724 392173 -15668
rect 392229 -15724 392315 -15668
rect 392371 -15724 392448 -15668
rect 392108 -15810 392448 -15724
rect 392108 -15866 392173 -15810
rect 392229 -15866 392315 -15810
rect 392371 -15866 392448 -15810
rect 392108 -15952 392448 -15866
rect 392108 -16008 392173 -15952
rect 392229 -16008 392315 -15952
rect 392371 -16008 392448 -15952
rect 392108 -16094 392448 -16008
rect 392108 -16150 392173 -16094
rect 392229 -16150 392315 -16094
rect 392371 -16150 392448 -16094
rect 392108 -16236 392448 -16150
rect 392108 -16292 392173 -16236
rect 392229 -16292 392315 -16236
rect 392371 -16292 392448 -16236
rect 392108 -16378 392448 -16292
rect 392108 -16434 392173 -16378
rect 392229 -16434 392315 -16378
rect 392371 -16434 392448 -16378
rect 392108 -16520 392448 -16434
rect 392108 -16576 392173 -16520
rect 392229 -16576 392315 -16520
rect 392371 -16576 392448 -16520
rect 392108 -16662 392448 -16576
rect 392108 -16718 392173 -16662
rect 392229 -16718 392315 -16662
rect 392371 -16718 392448 -16662
rect 392108 -16804 392448 -16718
rect 392108 -16860 392173 -16804
rect 392229 -16860 392315 -16804
rect 392371 -16860 392448 -16804
rect 392108 -16946 392448 -16860
rect 392108 -17002 392173 -16946
rect 392229 -17002 392315 -16946
rect 392371 -17002 392448 -16946
rect 392108 -17088 392448 -17002
rect 392108 -17144 392173 -17088
rect 392229 -17144 392315 -17088
rect 392371 -17144 392448 -17088
rect 392108 -17230 392448 -17144
rect 392108 -17286 392173 -17230
rect 392229 -17286 392315 -17230
rect 392371 -17286 392448 -17230
rect 392108 -17372 392448 -17286
rect 392108 -17428 392173 -17372
rect 392229 -17428 392315 -17372
rect 392371 -17428 392448 -17372
rect 392108 -17514 392448 -17428
rect 392108 -17570 392173 -17514
rect 392229 -17570 392315 -17514
rect 392371 -17570 392448 -17514
rect 392108 -17656 392448 -17570
rect 392108 -17712 392173 -17656
rect 392229 -17712 392315 -17656
rect 392371 -17712 392448 -17656
rect 392108 -17798 392448 -17712
rect 392108 -17854 392173 -17798
rect 392229 -17854 392315 -17798
rect 392371 -17854 392448 -17798
rect 392108 -17940 392448 -17854
rect 392108 -17996 392173 -17940
rect 392229 -17996 392315 -17940
rect 392371 -17996 392448 -17940
rect 392108 -18082 392448 -17996
rect 392108 -18138 392173 -18082
rect 392229 -18138 392315 -18082
rect 392371 -18138 392448 -18082
rect 392108 -18224 392448 -18138
rect 392108 -18280 392173 -18224
rect 392229 -18280 392315 -18224
rect 392371 -18280 392448 -18224
rect 392108 -18366 392448 -18280
rect 392108 -18422 392173 -18366
rect 392229 -18422 392315 -18366
rect 392371 -18422 392448 -18366
rect 392108 -18508 392448 -18422
rect 392108 -18564 392173 -18508
rect 392229 -18564 392315 -18508
rect 392371 -18564 392448 -18508
rect 392108 -18650 392448 -18564
rect 392108 -18706 392173 -18650
rect 392229 -18706 392315 -18650
rect 392371 -18706 392448 -18650
rect 392108 -18792 392448 -18706
rect 392108 -18848 392173 -18792
rect 392229 -18848 392315 -18792
rect 392371 -18848 392448 -18792
rect 392108 -18934 392448 -18848
rect 392108 -18990 392173 -18934
rect 392229 -18990 392315 -18934
rect 392371 -18990 392448 -18934
rect 392108 -19076 392448 -18990
rect 392108 -19132 392173 -19076
rect 392229 -19132 392315 -19076
rect 392371 -19132 392448 -19076
rect 392108 -19218 392448 -19132
rect 392108 -19274 392173 -19218
rect 392229 -19274 392315 -19218
rect 392371 -19274 392448 -19218
rect 392108 -19360 392448 -19274
rect 392108 -19416 392173 -19360
rect 392229 -19416 392315 -19360
rect 392371 -19416 392448 -19360
rect 392108 -19502 392448 -19416
rect 392108 -19558 392173 -19502
rect 392229 -19558 392315 -19502
rect 392371 -19558 392448 -19502
rect 392108 -19644 392448 -19558
rect 392108 -19700 392173 -19644
rect 392229 -19700 392315 -19644
rect 392371 -19700 392448 -19644
rect 392108 -19786 392448 -19700
rect 392108 -19842 392173 -19786
rect 392229 -19842 392315 -19786
rect 392371 -19842 392448 -19786
rect 392108 -19928 392448 -19842
rect 392108 -19984 392173 -19928
rect 392229 -19984 392315 -19928
rect 392371 -19984 392448 -19928
rect 392108 -20070 392448 -19984
rect 392108 -20126 392173 -20070
rect 392229 -20126 392315 -20070
rect 392371 -20126 392448 -20070
rect 392108 -20212 392448 -20126
rect 392108 -20268 392173 -20212
rect 392229 -20268 392315 -20212
rect 392371 -20268 392448 -20212
rect 392108 -20354 392448 -20268
rect 392108 -20410 392173 -20354
rect 392229 -20410 392315 -20354
rect 392371 -20410 392448 -20354
rect 392108 -20496 392448 -20410
rect 392108 -20552 392173 -20496
rect 392229 -20552 392315 -20496
rect 392371 -20552 392448 -20496
rect 392108 -20638 392448 -20552
rect 392108 -20694 392173 -20638
rect 392229 -20694 392315 -20638
rect 392371 -20694 392448 -20638
rect 392108 -20780 392448 -20694
rect 392108 -20836 392173 -20780
rect 392229 -20836 392315 -20780
rect 392371 -20836 392448 -20780
rect 392108 -20922 392448 -20836
rect 392108 -20978 392173 -20922
rect 392229 -20978 392315 -20922
rect 392371 -20978 392448 -20922
rect 392108 -21064 392448 -20978
rect 392108 -21120 392173 -21064
rect 392229 -21120 392315 -21064
rect 392371 -21120 392448 -21064
rect 392108 -21206 392448 -21120
rect 392108 -21262 392173 -21206
rect 392229 -21262 392315 -21206
rect 392371 -21262 392448 -21206
rect 392108 -21348 392448 -21262
rect 392108 -21404 392173 -21348
rect 392229 -21404 392315 -21348
rect 392371 -21404 392448 -21348
rect 392108 -21490 392448 -21404
rect 392108 -21546 392173 -21490
rect 392229 -21546 392315 -21490
rect 392371 -21546 392448 -21490
rect 392108 -21632 392448 -21546
rect 392108 -21688 392173 -21632
rect 392229 -21688 392315 -21632
rect 392371 -21688 392448 -21632
rect 392108 -21774 392448 -21688
rect 392108 -21830 392173 -21774
rect 392229 -21830 392315 -21774
rect 392371 -21830 392448 -21774
rect 392108 -21916 392448 -21830
rect 392108 -21972 392173 -21916
rect 392229 -21972 392315 -21916
rect 392371 -21972 392448 -21916
rect 392108 -22058 392448 -21972
rect 392108 -22114 392173 -22058
rect 392229 -22114 392315 -22058
rect 392371 -22114 392448 -22058
rect 392108 -22200 392448 -22114
rect 392108 -22256 392173 -22200
rect 392229 -22256 392315 -22200
rect 392371 -22256 392448 -22200
rect 392108 -22342 392448 -22256
rect 392108 -22398 392173 -22342
rect 392229 -22398 392315 -22342
rect 392371 -22398 392448 -22342
rect 392108 -22484 392448 -22398
rect 392108 -22540 392173 -22484
rect 392229 -22540 392315 -22484
rect 392371 -22540 392448 -22484
rect 392108 -22626 392448 -22540
rect 392108 -22682 392173 -22626
rect 392229 -22682 392315 -22626
rect 392371 -22682 392448 -22626
rect 392108 -22768 392448 -22682
rect 392108 -22824 392173 -22768
rect 392229 -22824 392315 -22768
rect 392371 -22824 392448 -22768
rect 392108 -22910 392448 -22824
rect 392108 -22966 392173 -22910
rect 392229 -22966 392315 -22910
rect 392371 -22966 392448 -22910
rect 392108 -23052 392448 -22966
rect 392108 -23108 392173 -23052
rect 392229 -23108 392315 -23052
rect 392371 -23108 392448 -23052
rect 392108 -23194 392448 -23108
rect 392108 -23250 392173 -23194
rect 392229 -23250 392315 -23194
rect 392371 -23250 392448 -23194
rect 392108 -23336 392448 -23250
rect 392108 -23392 392173 -23336
rect 392229 -23392 392315 -23336
rect 392371 -23392 392448 -23336
rect 392108 -23478 392448 -23392
rect 392108 -23534 392173 -23478
rect 392229 -23534 392315 -23478
rect 392371 -23534 392448 -23478
rect 392108 -23620 392448 -23534
rect 392108 -23676 392173 -23620
rect 392229 -23676 392315 -23620
rect 392371 -23676 392448 -23620
rect 392108 -23762 392448 -23676
rect 392108 -23818 392173 -23762
rect 392229 -23818 392315 -23762
rect 392371 -23818 392448 -23762
rect 392108 -23904 392448 -23818
rect 392108 -23960 392173 -23904
rect 392229 -23960 392315 -23904
rect 392371 -23960 392448 -23904
rect 392108 -24046 392448 -23960
rect 392108 -24102 392173 -24046
rect 392229 -24102 392315 -24046
rect 392371 -24102 392448 -24046
rect 392108 -24188 392448 -24102
rect 392108 -24244 392173 -24188
rect 392229 -24244 392315 -24188
rect 392371 -24244 392448 -24188
rect 392108 -24330 392448 -24244
rect 392108 -24386 392173 -24330
rect 392229 -24386 392315 -24330
rect 392371 -24386 392448 -24330
rect 392108 -24472 392448 -24386
rect 392108 -24528 392173 -24472
rect 392229 -24528 392315 -24472
rect 392371 -24528 392448 -24472
rect 392108 -24614 392448 -24528
rect 392108 -24670 392173 -24614
rect 392229 -24670 392315 -24614
rect 392371 -24670 392448 -24614
rect 392108 -24756 392448 -24670
rect 392108 -24812 392173 -24756
rect 392229 -24812 392315 -24756
rect 392371 -24812 392448 -24756
rect 392108 -24898 392448 -24812
rect 392108 -24954 392173 -24898
rect 392229 -24954 392315 -24898
rect 392371 -24954 392448 -24898
rect 392108 -25040 392448 -24954
rect 392108 -25096 392173 -25040
rect 392229 -25096 392315 -25040
rect 392371 -25096 392448 -25040
rect 392108 -25182 392448 -25096
rect 392108 -25238 392173 -25182
rect 392229 -25238 392315 -25182
rect 392371 -25238 392448 -25182
rect 392108 -25324 392448 -25238
rect 392108 -25380 392173 -25324
rect 392229 -25380 392315 -25324
rect 392371 -25380 392448 -25324
rect 392108 -25466 392448 -25380
rect 392108 -25522 392173 -25466
rect 392229 -25522 392315 -25466
rect 392371 -25522 392448 -25466
rect 392108 -25590 392448 -25522
rect 392508 -13680 392848 -13590
rect 392508 -13736 392578 -13680
rect 392634 -13736 392720 -13680
rect 392776 -13736 392848 -13680
rect 392508 -13822 392848 -13736
rect 392508 -13878 392578 -13822
rect 392634 -13878 392720 -13822
rect 392776 -13878 392848 -13822
rect 392508 -13964 392848 -13878
rect 392508 -14020 392578 -13964
rect 392634 -14020 392720 -13964
rect 392776 -14020 392848 -13964
rect 392508 -14106 392848 -14020
rect 392508 -14162 392578 -14106
rect 392634 -14162 392720 -14106
rect 392776 -14162 392848 -14106
rect 392508 -14248 392848 -14162
rect 392508 -14304 392578 -14248
rect 392634 -14304 392720 -14248
rect 392776 -14304 392848 -14248
rect 392508 -14390 392848 -14304
rect 392508 -14446 392578 -14390
rect 392634 -14446 392720 -14390
rect 392776 -14446 392848 -14390
rect 392508 -14532 392848 -14446
rect 392508 -14588 392578 -14532
rect 392634 -14588 392720 -14532
rect 392776 -14588 392848 -14532
rect 392508 -14674 392848 -14588
rect 392508 -14730 392578 -14674
rect 392634 -14730 392720 -14674
rect 392776 -14730 392848 -14674
rect 392508 -14816 392848 -14730
rect 392508 -14872 392578 -14816
rect 392634 -14872 392720 -14816
rect 392776 -14872 392848 -14816
rect 392508 -14958 392848 -14872
rect 392508 -15014 392578 -14958
rect 392634 -15014 392720 -14958
rect 392776 -15014 392848 -14958
rect 392508 -15100 392848 -15014
rect 392508 -15156 392578 -15100
rect 392634 -15156 392720 -15100
rect 392776 -15156 392848 -15100
rect 392508 -15242 392848 -15156
rect 392508 -15298 392578 -15242
rect 392634 -15298 392720 -15242
rect 392776 -15298 392848 -15242
rect 392508 -15384 392848 -15298
rect 392508 -15440 392578 -15384
rect 392634 -15440 392720 -15384
rect 392776 -15440 392848 -15384
rect 392508 -15526 392848 -15440
rect 392508 -15582 392578 -15526
rect 392634 -15582 392720 -15526
rect 392776 -15582 392848 -15526
rect 392508 -15668 392848 -15582
rect 392508 -15724 392578 -15668
rect 392634 -15724 392720 -15668
rect 392776 -15724 392848 -15668
rect 392508 -15810 392848 -15724
rect 392508 -15866 392578 -15810
rect 392634 -15866 392720 -15810
rect 392776 -15866 392848 -15810
rect 392508 -15952 392848 -15866
rect 392508 -16008 392578 -15952
rect 392634 -16008 392720 -15952
rect 392776 -16008 392848 -15952
rect 392508 -16094 392848 -16008
rect 392508 -16150 392578 -16094
rect 392634 -16150 392720 -16094
rect 392776 -16150 392848 -16094
rect 392508 -16236 392848 -16150
rect 392508 -16292 392578 -16236
rect 392634 -16292 392720 -16236
rect 392776 -16292 392848 -16236
rect 392508 -16378 392848 -16292
rect 392508 -16434 392578 -16378
rect 392634 -16434 392720 -16378
rect 392776 -16434 392848 -16378
rect 392508 -16520 392848 -16434
rect 392508 -16576 392578 -16520
rect 392634 -16576 392720 -16520
rect 392776 -16576 392848 -16520
rect 392508 -16662 392848 -16576
rect 392508 -16718 392578 -16662
rect 392634 -16718 392720 -16662
rect 392776 -16718 392848 -16662
rect 392508 -16804 392848 -16718
rect 392508 -16860 392578 -16804
rect 392634 -16860 392720 -16804
rect 392776 -16860 392848 -16804
rect 392508 -16946 392848 -16860
rect 392508 -17002 392578 -16946
rect 392634 -17002 392720 -16946
rect 392776 -17002 392848 -16946
rect 392508 -17088 392848 -17002
rect 392508 -17144 392578 -17088
rect 392634 -17144 392720 -17088
rect 392776 -17144 392848 -17088
rect 392508 -17230 392848 -17144
rect 392508 -17286 392578 -17230
rect 392634 -17286 392720 -17230
rect 392776 -17286 392848 -17230
rect 392508 -17372 392848 -17286
rect 392508 -17428 392578 -17372
rect 392634 -17428 392720 -17372
rect 392776 -17428 392848 -17372
rect 392508 -17514 392848 -17428
rect 392508 -17570 392578 -17514
rect 392634 -17570 392720 -17514
rect 392776 -17570 392848 -17514
rect 392508 -17656 392848 -17570
rect 392508 -17712 392578 -17656
rect 392634 -17712 392720 -17656
rect 392776 -17712 392848 -17656
rect 392508 -17798 392848 -17712
rect 392508 -17854 392578 -17798
rect 392634 -17854 392720 -17798
rect 392776 -17854 392848 -17798
rect 392508 -17940 392848 -17854
rect 392508 -17996 392578 -17940
rect 392634 -17996 392720 -17940
rect 392776 -17996 392848 -17940
rect 392508 -18082 392848 -17996
rect 392508 -18138 392578 -18082
rect 392634 -18138 392720 -18082
rect 392776 -18138 392848 -18082
rect 392508 -18224 392848 -18138
rect 392508 -18280 392578 -18224
rect 392634 -18280 392720 -18224
rect 392776 -18280 392848 -18224
rect 392508 -18366 392848 -18280
rect 392508 -18422 392578 -18366
rect 392634 -18422 392720 -18366
rect 392776 -18422 392848 -18366
rect 392508 -18508 392848 -18422
rect 392508 -18564 392578 -18508
rect 392634 -18564 392720 -18508
rect 392776 -18564 392848 -18508
rect 392508 -18650 392848 -18564
rect 392508 -18706 392578 -18650
rect 392634 -18706 392720 -18650
rect 392776 -18706 392848 -18650
rect 392508 -18792 392848 -18706
rect 392508 -18848 392578 -18792
rect 392634 -18848 392720 -18792
rect 392776 -18848 392848 -18792
rect 392508 -18934 392848 -18848
rect 392508 -18990 392578 -18934
rect 392634 -18990 392720 -18934
rect 392776 -18990 392848 -18934
rect 392508 -19076 392848 -18990
rect 392508 -19132 392578 -19076
rect 392634 -19132 392720 -19076
rect 392776 -19132 392848 -19076
rect 392508 -19218 392848 -19132
rect 392508 -19274 392578 -19218
rect 392634 -19274 392720 -19218
rect 392776 -19274 392848 -19218
rect 392508 -19360 392848 -19274
rect 392508 -19416 392578 -19360
rect 392634 -19416 392720 -19360
rect 392776 -19416 392848 -19360
rect 392508 -19502 392848 -19416
rect 392508 -19558 392578 -19502
rect 392634 -19558 392720 -19502
rect 392776 -19558 392848 -19502
rect 392508 -19644 392848 -19558
rect 392508 -19700 392578 -19644
rect 392634 -19700 392720 -19644
rect 392776 -19700 392848 -19644
rect 392508 -19786 392848 -19700
rect 392508 -19842 392578 -19786
rect 392634 -19842 392720 -19786
rect 392776 -19842 392848 -19786
rect 392508 -19928 392848 -19842
rect 392508 -19984 392578 -19928
rect 392634 -19984 392720 -19928
rect 392776 -19984 392848 -19928
rect 392508 -20070 392848 -19984
rect 392508 -20126 392578 -20070
rect 392634 -20126 392720 -20070
rect 392776 -20126 392848 -20070
rect 392508 -20212 392848 -20126
rect 392508 -20268 392578 -20212
rect 392634 -20268 392720 -20212
rect 392776 -20268 392848 -20212
rect 392508 -20354 392848 -20268
rect 392508 -20410 392578 -20354
rect 392634 -20410 392720 -20354
rect 392776 -20410 392848 -20354
rect 392508 -20496 392848 -20410
rect 392508 -20552 392578 -20496
rect 392634 -20552 392720 -20496
rect 392776 -20552 392848 -20496
rect 392508 -20638 392848 -20552
rect 392508 -20694 392578 -20638
rect 392634 -20694 392720 -20638
rect 392776 -20694 392848 -20638
rect 392508 -20780 392848 -20694
rect 392508 -20836 392578 -20780
rect 392634 -20836 392720 -20780
rect 392776 -20836 392848 -20780
rect 392508 -20922 392848 -20836
rect 392508 -20978 392578 -20922
rect 392634 -20978 392720 -20922
rect 392776 -20978 392848 -20922
rect 392508 -21064 392848 -20978
rect 392508 -21120 392578 -21064
rect 392634 -21120 392720 -21064
rect 392776 -21120 392848 -21064
rect 392508 -21206 392848 -21120
rect 392508 -21262 392578 -21206
rect 392634 -21262 392720 -21206
rect 392776 -21262 392848 -21206
rect 392508 -21348 392848 -21262
rect 392508 -21404 392578 -21348
rect 392634 -21404 392720 -21348
rect 392776 -21404 392848 -21348
rect 392508 -21490 392848 -21404
rect 392508 -21546 392578 -21490
rect 392634 -21546 392720 -21490
rect 392776 -21546 392848 -21490
rect 392508 -21632 392848 -21546
rect 392508 -21688 392578 -21632
rect 392634 -21688 392720 -21632
rect 392776 -21688 392848 -21632
rect 392508 -21774 392848 -21688
rect 392508 -21830 392578 -21774
rect 392634 -21830 392720 -21774
rect 392776 -21830 392848 -21774
rect 392508 -21916 392848 -21830
rect 392508 -21972 392578 -21916
rect 392634 -21972 392720 -21916
rect 392776 -21972 392848 -21916
rect 392508 -22058 392848 -21972
rect 392508 -22114 392578 -22058
rect 392634 -22114 392720 -22058
rect 392776 -22114 392848 -22058
rect 392508 -22200 392848 -22114
rect 392508 -22256 392578 -22200
rect 392634 -22256 392720 -22200
rect 392776 -22256 392848 -22200
rect 392508 -22342 392848 -22256
rect 392508 -22398 392578 -22342
rect 392634 -22398 392720 -22342
rect 392776 -22398 392848 -22342
rect 392508 -22484 392848 -22398
rect 392508 -22540 392578 -22484
rect 392634 -22540 392720 -22484
rect 392776 -22540 392848 -22484
rect 392508 -22626 392848 -22540
rect 392508 -22682 392578 -22626
rect 392634 -22682 392720 -22626
rect 392776 -22682 392848 -22626
rect 392508 -22768 392848 -22682
rect 392508 -22824 392578 -22768
rect 392634 -22824 392720 -22768
rect 392776 -22824 392848 -22768
rect 392508 -22910 392848 -22824
rect 392508 -22966 392578 -22910
rect 392634 -22966 392720 -22910
rect 392776 -22966 392848 -22910
rect 392508 -23052 392848 -22966
rect 392508 -23108 392578 -23052
rect 392634 -23108 392720 -23052
rect 392776 -23108 392848 -23052
rect 392508 -23194 392848 -23108
rect 392508 -23250 392578 -23194
rect 392634 -23250 392720 -23194
rect 392776 -23250 392848 -23194
rect 392508 -23336 392848 -23250
rect 392508 -23392 392578 -23336
rect 392634 -23392 392720 -23336
rect 392776 -23392 392848 -23336
rect 392508 -23478 392848 -23392
rect 392508 -23534 392578 -23478
rect 392634 -23534 392720 -23478
rect 392776 -23534 392848 -23478
rect 392508 -23620 392848 -23534
rect 392508 -23676 392578 -23620
rect 392634 -23676 392720 -23620
rect 392776 -23676 392848 -23620
rect 392508 -23762 392848 -23676
rect 392508 -23818 392578 -23762
rect 392634 -23818 392720 -23762
rect 392776 -23818 392848 -23762
rect 392508 -23904 392848 -23818
rect 392508 -23960 392578 -23904
rect 392634 -23960 392720 -23904
rect 392776 -23960 392848 -23904
rect 392508 -24046 392848 -23960
rect 392508 -24102 392578 -24046
rect 392634 -24102 392720 -24046
rect 392776 -24102 392848 -24046
rect 392508 -24188 392848 -24102
rect 392508 -24244 392578 -24188
rect 392634 -24244 392720 -24188
rect 392776 -24244 392848 -24188
rect 392508 -24330 392848 -24244
rect 392508 -24386 392578 -24330
rect 392634 -24386 392720 -24330
rect 392776 -24386 392848 -24330
rect 392508 -24472 392848 -24386
rect 392508 -24528 392578 -24472
rect 392634 -24528 392720 -24472
rect 392776 -24528 392848 -24472
rect 392508 -24614 392848 -24528
rect 392508 -24670 392578 -24614
rect 392634 -24670 392720 -24614
rect 392776 -24670 392848 -24614
rect 392508 -24756 392848 -24670
rect 392508 -24812 392578 -24756
rect 392634 -24812 392720 -24756
rect 392776 -24812 392848 -24756
rect 392508 -24898 392848 -24812
rect 392508 -24954 392578 -24898
rect 392634 -24954 392720 -24898
rect 392776 -24954 392848 -24898
rect 392508 -25040 392848 -24954
rect 392508 -25096 392578 -25040
rect 392634 -25096 392720 -25040
rect 392776 -25096 392848 -25040
rect 392508 -25182 392848 -25096
rect 392508 -25238 392578 -25182
rect 392634 -25238 392720 -25182
rect 392776 -25238 392848 -25182
rect 392508 -25324 392848 -25238
rect 392508 -25380 392578 -25324
rect 392634 -25380 392720 -25324
rect 392776 -25380 392848 -25324
rect 392508 -25466 392848 -25380
rect 392508 -25522 392578 -25466
rect 392634 -25522 392720 -25466
rect 392776 -25522 392848 -25466
rect 392508 -25590 392848 -25522
rect 392908 -13680 393248 -13590
rect 392908 -13736 392978 -13680
rect 393034 -13736 393120 -13680
rect 393176 -13736 393248 -13680
rect 392908 -13822 393248 -13736
rect 392908 -13878 392978 -13822
rect 393034 -13878 393120 -13822
rect 393176 -13878 393248 -13822
rect 392908 -13964 393248 -13878
rect 392908 -14020 392978 -13964
rect 393034 -14020 393120 -13964
rect 393176 -14020 393248 -13964
rect 392908 -14106 393248 -14020
rect 392908 -14162 392978 -14106
rect 393034 -14162 393120 -14106
rect 393176 -14162 393248 -14106
rect 392908 -14248 393248 -14162
rect 392908 -14304 392978 -14248
rect 393034 -14304 393120 -14248
rect 393176 -14304 393248 -14248
rect 392908 -14390 393248 -14304
rect 392908 -14446 392978 -14390
rect 393034 -14446 393120 -14390
rect 393176 -14446 393248 -14390
rect 392908 -14532 393248 -14446
rect 392908 -14588 392978 -14532
rect 393034 -14588 393120 -14532
rect 393176 -14588 393248 -14532
rect 392908 -14674 393248 -14588
rect 392908 -14730 392978 -14674
rect 393034 -14730 393120 -14674
rect 393176 -14730 393248 -14674
rect 392908 -14816 393248 -14730
rect 392908 -14872 392978 -14816
rect 393034 -14872 393120 -14816
rect 393176 -14872 393248 -14816
rect 392908 -14958 393248 -14872
rect 392908 -15014 392978 -14958
rect 393034 -15014 393120 -14958
rect 393176 -15014 393248 -14958
rect 392908 -15100 393248 -15014
rect 392908 -15156 392978 -15100
rect 393034 -15156 393120 -15100
rect 393176 -15156 393248 -15100
rect 392908 -15242 393248 -15156
rect 392908 -15298 392978 -15242
rect 393034 -15298 393120 -15242
rect 393176 -15298 393248 -15242
rect 392908 -15384 393248 -15298
rect 392908 -15440 392978 -15384
rect 393034 -15440 393120 -15384
rect 393176 -15440 393248 -15384
rect 392908 -15526 393248 -15440
rect 392908 -15582 392978 -15526
rect 393034 -15582 393120 -15526
rect 393176 -15582 393248 -15526
rect 392908 -15668 393248 -15582
rect 392908 -15724 392978 -15668
rect 393034 -15724 393120 -15668
rect 393176 -15724 393248 -15668
rect 392908 -15810 393248 -15724
rect 392908 -15866 392978 -15810
rect 393034 -15866 393120 -15810
rect 393176 -15866 393248 -15810
rect 392908 -15952 393248 -15866
rect 392908 -16008 392978 -15952
rect 393034 -16008 393120 -15952
rect 393176 -16008 393248 -15952
rect 392908 -16094 393248 -16008
rect 392908 -16150 392978 -16094
rect 393034 -16150 393120 -16094
rect 393176 -16150 393248 -16094
rect 392908 -16236 393248 -16150
rect 392908 -16292 392978 -16236
rect 393034 -16292 393120 -16236
rect 393176 -16292 393248 -16236
rect 392908 -16378 393248 -16292
rect 392908 -16434 392978 -16378
rect 393034 -16434 393120 -16378
rect 393176 -16434 393248 -16378
rect 392908 -16520 393248 -16434
rect 392908 -16576 392978 -16520
rect 393034 -16576 393120 -16520
rect 393176 -16576 393248 -16520
rect 392908 -16662 393248 -16576
rect 392908 -16718 392978 -16662
rect 393034 -16718 393120 -16662
rect 393176 -16718 393248 -16662
rect 392908 -16804 393248 -16718
rect 392908 -16860 392978 -16804
rect 393034 -16860 393120 -16804
rect 393176 -16860 393248 -16804
rect 392908 -16946 393248 -16860
rect 392908 -17002 392978 -16946
rect 393034 -17002 393120 -16946
rect 393176 -17002 393248 -16946
rect 392908 -17088 393248 -17002
rect 392908 -17144 392978 -17088
rect 393034 -17144 393120 -17088
rect 393176 -17144 393248 -17088
rect 392908 -17230 393248 -17144
rect 392908 -17286 392978 -17230
rect 393034 -17286 393120 -17230
rect 393176 -17286 393248 -17230
rect 392908 -17372 393248 -17286
rect 392908 -17428 392978 -17372
rect 393034 -17428 393120 -17372
rect 393176 -17428 393248 -17372
rect 392908 -17514 393248 -17428
rect 392908 -17570 392978 -17514
rect 393034 -17570 393120 -17514
rect 393176 -17570 393248 -17514
rect 392908 -17656 393248 -17570
rect 392908 -17712 392978 -17656
rect 393034 -17712 393120 -17656
rect 393176 -17712 393248 -17656
rect 392908 -17798 393248 -17712
rect 392908 -17854 392978 -17798
rect 393034 -17854 393120 -17798
rect 393176 -17854 393248 -17798
rect 392908 -17940 393248 -17854
rect 392908 -17996 392978 -17940
rect 393034 -17996 393120 -17940
rect 393176 -17996 393248 -17940
rect 392908 -18082 393248 -17996
rect 392908 -18138 392978 -18082
rect 393034 -18138 393120 -18082
rect 393176 -18138 393248 -18082
rect 392908 -18224 393248 -18138
rect 392908 -18280 392978 -18224
rect 393034 -18280 393120 -18224
rect 393176 -18280 393248 -18224
rect 392908 -18366 393248 -18280
rect 392908 -18422 392978 -18366
rect 393034 -18422 393120 -18366
rect 393176 -18422 393248 -18366
rect 392908 -18508 393248 -18422
rect 392908 -18564 392978 -18508
rect 393034 -18564 393120 -18508
rect 393176 -18564 393248 -18508
rect 392908 -18650 393248 -18564
rect 392908 -18706 392978 -18650
rect 393034 -18706 393120 -18650
rect 393176 -18706 393248 -18650
rect 392908 -18792 393248 -18706
rect 392908 -18848 392978 -18792
rect 393034 -18848 393120 -18792
rect 393176 -18848 393248 -18792
rect 392908 -18934 393248 -18848
rect 392908 -18990 392978 -18934
rect 393034 -18990 393120 -18934
rect 393176 -18990 393248 -18934
rect 392908 -19076 393248 -18990
rect 392908 -19132 392978 -19076
rect 393034 -19132 393120 -19076
rect 393176 -19132 393248 -19076
rect 392908 -19218 393248 -19132
rect 392908 -19274 392978 -19218
rect 393034 -19274 393120 -19218
rect 393176 -19274 393248 -19218
rect 392908 -19360 393248 -19274
rect 392908 -19416 392978 -19360
rect 393034 -19416 393120 -19360
rect 393176 -19416 393248 -19360
rect 392908 -19502 393248 -19416
rect 392908 -19558 392978 -19502
rect 393034 -19558 393120 -19502
rect 393176 -19558 393248 -19502
rect 392908 -19644 393248 -19558
rect 392908 -19700 392978 -19644
rect 393034 -19700 393120 -19644
rect 393176 -19700 393248 -19644
rect 392908 -19786 393248 -19700
rect 392908 -19842 392978 -19786
rect 393034 -19842 393120 -19786
rect 393176 -19842 393248 -19786
rect 392908 -19928 393248 -19842
rect 392908 -19984 392978 -19928
rect 393034 -19984 393120 -19928
rect 393176 -19984 393248 -19928
rect 392908 -20070 393248 -19984
rect 392908 -20126 392978 -20070
rect 393034 -20126 393120 -20070
rect 393176 -20126 393248 -20070
rect 392908 -20212 393248 -20126
rect 392908 -20268 392978 -20212
rect 393034 -20268 393120 -20212
rect 393176 -20268 393248 -20212
rect 392908 -20354 393248 -20268
rect 392908 -20410 392978 -20354
rect 393034 -20410 393120 -20354
rect 393176 -20410 393248 -20354
rect 392908 -20496 393248 -20410
rect 392908 -20552 392978 -20496
rect 393034 -20552 393120 -20496
rect 393176 -20552 393248 -20496
rect 392908 -20638 393248 -20552
rect 392908 -20694 392978 -20638
rect 393034 -20694 393120 -20638
rect 393176 -20694 393248 -20638
rect 392908 -20780 393248 -20694
rect 392908 -20836 392978 -20780
rect 393034 -20836 393120 -20780
rect 393176 -20836 393248 -20780
rect 392908 -20922 393248 -20836
rect 392908 -20978 392978 -20922
rect 393034 -20978 393120 -20922
rect 393176 -20978 393248 -20922
rect 392908 -21064 393248 -20978
rect 392908 -21120 392978 -21064
rect 393034 -21120 393120 -21064
rect 393176 -21120 393248 -21064
rect 392908 -21206 393248 -21120
rect 392908 -21262 392978 -21206
rect 393034 -21262 393120 -21206
rect 393176 -21262 393248 -21206
rect 392908 -21348 393248 -21262
rect 392908 -21404 392978 -21348
rect 393034 -21404 393120 -21348
rect 393176 -21404 393248 -21348
rect 392908 -21490 393248 -21404
rect 392908 -21546 392978 -21490
rect 393034 -21546 393120 -21490
rect 393176 -21546 393248 -21490
rect 392908 -21632 393248 -21546
rect 392908 -21688 392978 -21632
rect 393034 -21688 393120 -21632
rect 393176 -21688 393248 -21632
rect 392908 -21774 393248 -21688
rect 392908 -21830 392978 -21774
rect 393034 -21830 393120 -21774
rect 393176 -21830 393248 -21774
rect 392908 -21916 393248 -21830
rect 392908 -21972 392978 -21916
rect 393034 -21972 393120 -21916
rect 393176 -21972 393248 -21916
rect 392908 -22058 393248 -21972
rect 392908 -22114 392978 -22058
rect 393034 -22114 393120 -22058
rect 393176 -22114 393248 -22058
rect 392908 -22200 393248 -22114
rect 392908 -22256 392978 -22200
rect 393034 -22256 393120 -22200
rect 393176 -22256 393248 -22200
rect 392908 -22342 393248 -22256
rect 392908 -22398 392978 -22342
rect 393034 -22398 393120 -22342
rect 393176 -22398 393248 -22342
rect 392908 -22484 393248 -22398
rect 392908 -22540 392978 -22484
rect 393034 -22540 393120 -22484
rect 393176 -22540 393248 -22484
rect 392908 -22626 393248 -22540
rect 392908 -22682 392978 -22626
rect 393034 -22682 393120 -22626
rect 393176 -22682 393248 -22626
rect 392908 -22768 393248 -22682
rect 392908 -22824 392978 -22768
rect 393034 -22824 393120 -22768
rect 393176 -22824 393248 -22768
rect 392908 -22910 393248 -22824
rect 392908 -22966 392978 -22910
rect 393034 -22966 393120 -22910
rect 393176 -22966 393248 -22910
rect 392908 -23052 393248 -22966
rect 392908 -23108 392978 -23052
rect 393034 -23108 393120 -23052
rect 393176 -23108 393248 -23052
rect 392908 -23194 393248 -23108
rect 392908 -23250 392978 -23194
rect 393034 -23250 393120 -23194
rect 393176 -23250 393248 -23194
rect 392908 -23336 393248 -23250
rect 392908 -23392 392978 -23336
rect 393034 -23392 393120 -23336
rect 393176 -23392 393248 -23336
rect 392908 -23478 393248 -23392
rect 392908 -23534 392978 -23478
rect 393034 -23534 393120 -23478
rect 393176 -23534 393248 -23478
rect 392908 -23620 393248 -23534
rect 392908 -23676 392978 -23620
rect 393034 -23676 393120 -23620
rect 393176 -23676 393248 -23620
rect 392908 -23762 393248 -23676
rect 392908 -23818 392978 -23762
rect 393034 -23818 393120 -23762
rect 393176 -23818 393248 -23762
rect 392908 -23904 393248 -23818
rect 392908 -23960 392978 -23904
rect 393034 -23960 393120 -23904
rect 393176 -23960 393248 -23904
rect 392908 -24046 393248 -23960
rect 392908 -24102 392978 -24046
rect 393034 -24102 393120 -24046
rect 393176 -24102 393248 -24046
rect 392908 -24188 393248 -24102
rect 392908 -24244 392978 -24188
rect 393034 -24244 393120 -24188
rect 393176 -24244 393248 -24188
rect 392908 -24330 393248 -24244
rect 392908 -24386 392978 -24330
rect 393034 -24386 393120 -24330
rect 393176 -24386 393248 -24330
rect 392908 -24472 393248 -24386
rect 392908 -24528 392978 -24472
rect 393034 -24528 393120 -24472
rect 393176 -24528 393248 -24472
rect 392908 -24614 393248 -24528
rect 392908 -24670 392978 -24614
rect 393034 -24670 393120 -24614
rect 393176 -24670 393248 -24614
rect 392908 -24756 393248 -24670
rect 392908 -24812 392978 -24756
rect 393034 -24812 393120 -24756
rect 393176 -24812 393248 -24756
rect 392908 -24898 393248 -24812
rect 392908 -24954 392978 -24898
rect 393034 -24954 393120 -24898
rect 393176 -24954 393248 -24898
rect 392908 -25040 393248 -24954
rect 392908 -25096 392978 -25040
rect 393034 -25096 393120 -25040
rect 393176 -25096 393248 -25040
rect 392908 -25182 393248 -25096
rect 392908 -25238 392978 -25182
rect 393034 -25238 393120 -25182
rect 393176 -25238 393248 -25182
rect 392908 -25324 393248 -25238
rect 392908 -25380 392978 -25324
rect 393034 -25380 393120 -25324
rect 393176 -25380 393248 -25324
rect 392908 -25466 393248 -25380
rect 392908 -25522 392978 -25466
rect 393034 -25522 393120 -25466
rect 393176 -25522 393248 -25466
rect 392908 -25590 393248 -25522
rect 393308 -13680 393648 -13590
rect 393308 -13736 393383 -13680
rect 393439 -13736 393525 -13680
rect 393581 -13736 393648 -13680
rect 393308 -13822 393648 -13736
rect 393308 -13878 393383 -13822
rect 393439 -13878 393525 -13822
rect 393581 -13878 393648 -13822
rect 393308 -13964 393648 -13878
rect 393308 -14020 393383 -13964
rect 393439 -14020 393525 -13964
rect 393581 -14020 393648 -13964
rect 393308 -14106 393648 -14020
rect 393308 -14162 393383 -14106
rect 393439 -14162 393525 -14106
rect 393581 -14162 393648 -14106
rect 393308 -14248 393648 -14162
rect 393308 -14304 393383 -14248
rect 393439 -14304 393525 -14248
rect 393581 -14304 393648 -14248
rect 393308 -14390 393648 -14304
rect 393308 -14446 393383 -14390
rect 393439 -14446 393525 -14390
rect 393581 -14446 393648 -14390
rect 393308 -14532 393648 -14446
rect 393308 -14588 393383 -14532
rect 393439 -14588 393525 -14532
rect 393581 -14588 393648 -14532
rect 393308 -14674 393648 -14588
rect 393308 -14730 393383 -14674
rect 393439 -14730 393525 -14674
rect 393581 -14730 393648 -14674
rect 393308 -14816 393648 -14730
rect 393308 -14872 393383 -14816
rect 393439 -14872 393525 -14816
rect 393581 -14872 393648 -14816
rect 393308 -14958 393648 -14872
rect 393308 -15014 393383 -14958
rect 393439 -15014 393525 -14958
rect 393581 -15014 393648 -14958
rect 393308 -15100 393648 -15014
rect 393308 -15156 393383 -15100
rect 393439 -15156 393525 -15100
rect 393581 -15156 393648 -15100
rect 393308 -15242 393648 -15156
rect 393308 -15298 393383 -15242
rect 393439 -15298 393525 -15242
rect 393581 -15298 393648 -15242
rect 393308 -15384 393648 -15298
rect 393308 -15440 393383 -15384
rect 393439 -15440 393525 -15384
rect 393581 -15440 393648 -15384
rect 393308 -15526 393648 -15440
rect 393308 -15582 393383 -15526
rect 393439 -15582 393525 -15526
rect 393581 -15582 393648 -15526
rect 393308 -15668 393648 -15582
rect 393308 -15724 393383 -15668
rect 393439 -15724 393525 -15668
rect 393581 -15724 393648 -15668
rect 393308 -15810 393648 -15724
rect 393308 -15866 393383 -15810
rect 393439 -15866 393525 -15810
rect 393581 -15866 393648 -15810
rect 393308 -15952 393648 -15866
rect 393308 -16008 393383 -15952
rect 393439 -16008 393525 -15952
rect 393581 -16008 393648 -15952
rect 393308 -16094 393648 -16008
rect 393308 -16150 393383 -16094
rect 393439 -16150 393525 -16094
rect 393581 -16150 393648 -16094
rect 393308 -16236 393648 -16150
rect 393308 -16292 393383 -16236
rect 393439 -16292 393525 -16236
rect 393581 -16292 393648 -16236
rect 393308 -16378 393648 -16292
rect 393308 -16434 393383 -16378
rect 393439 -16434 393525 -16378
rect 393581 -16434 393648 -16378
rect 393308 -16520 393648 -16434
rect 393308 -16576 393383 -16520
rect 393439 -16576 393525 -16520
rect 393581 -16576 393648 -16520
rect 393308 -16662 393648 -16576
rect 393308 -16718 393383 -16662
rect 393439 -16718 393525 -16662
rect 393581 -16718 393648 -16662
rect 393308 -16804 393648 -16718
rect 393308 -16860 393383 -16804
rect 393439 -16860 393525 -16804
rect 393581 -16860 393648 -16804
rect 393308 -16946 393648 -16860
rect 393308 -17002 393383 -16946
rect 393439 -17002 393525 -16946
rect 393581 -17002 393648 -16946
rect 393308 -17088 393648 -17002
rect 393308 -17144 393383 -17088
rect 393439 -17144 393525 -17088
rect 393581 -17144 393648 -17088
rect 393308 -17230 393648 -17144
rect 393308 -17286 393383 -17230
rect 393439 -17286 393525 -17230
rect 393581 -17286 393648 -17230
rect 393308 -17372 393648 -17286
rect 393308 -17428 393383 -17372
rect 393439 -17428 393525 -17372
rect 393581 -17428 393648 -17372
rect 393308 -17514 393648 -17428
rect 393308 -17570 393383 -17514
rect 393439 -17570 393525 -17514
rect 393581 -17570 393648 -17514
rect 393308 -17656 393648 -17570
rect 393308 -17712 393383 -17656
rect 393439 -17712 393525 -17656
rect 393581 -17712 393648 -17656
rect 393308 -17798 393648 -17712
rect 393308 -17854 393383 -17798
rect 393439 -17854 393525 -17798
rect 393581 -17854 393648 -17798
rect 393308 -17940 393648 -17854
rect 393308 -17996 393383 -17940
rect 393439 -17996 393525 -17940
rect 393581 -17996 393648 -17940
rect 393308 -18082 393648 -17996
rect 393308 -18138 393383 -18082
rect 393439 -18138 393525 -18082
rect 393581 -18138 393648 -18082
rect 393308 -18224 393648 -18138
rect 393308 -18280 393383 -18224
rect 393439 -18280 393525 -18224
rect 393581 -18280 393648 -18224
rect 393308 -18366 393648 -18280
rect 393308 -18422 393383 -18366
rect 393439 -18422 393525 -18366
rect 393581 -18422 393648 -18366
rect 393308 -18508 393648 -18422
rect 393308 -18564 393383 -18508
rect 393439 -18564 393525 -18508
rect 393581 -18564 393648 -18508
rect 393308 -18650 393648 -18564
rect 393308 -18706 393383 -18650
rect 393439 -18706 393525 -18650
rect 393581 -18706 393648 -18650
rect 393308 -18792 393648 -18706
rect 393308 -18848 393383 -18792
rect 393439 -18848 393525 -18792
rect 393581 -18848 393648 -18792
rect 393308 -18934 393648 -18848
rect 393308 -18990 393383 -18934
rect 393439 -18990 393525 -18934
rect 393581 -18990 393648 -18934
rect 393308 -19076 393648 -18990
rect 393308 -19132 393383 -19076
rect 393439 -19132 393525 -19076
rect 393581 -19132 393648 -19076
rect 393308 -19218 393648 -19132
rect 393308 -19274 393383 -19218
rect 393439 -19274 393525 -19218
rect 393581 -19274 393648 -19218
rect 393308 -19360 393648 -19274
rect 393308 -19416 393383 -19360
rect 393439 -19416 393525 -19360
rect 393581 -19416 393648 -19360
rect 393308 -19502 393648 -19416
rect 393308 -19558 393383 -19502
rect 393439 -19558 393525 -19502
rect 393581 -19558 393648 -19502
rect 393308 -19644 393648 -19558
rect 393308 -19700 393383 -19644
rect 393439 -19700 393525 -19644
rect 393581 -19700 393648 -19644
rect 393308 -19786 393648 -19700
rect 393308 -19842 393383 -19786
rect 393439 -19842 393525 -19786
rect 393581 -19842 393648 -19786
rect 393308 -19928 393648 -19842
rect 393308 -19984 393383 -19928
rect 393439 -19984 393525 -19928
rect 393581 -19984 393648 -19928
rect 393308 -20070 393648 -19984
rect 393308 -20126 393383 -20070
rect 393439 -20126 393525 -20070
rect 393581 -20126 393648 -20070
rect 393308 -20212 393648 -20126
rect 393308 -20268 393383 -20212
rect 393439 -20268 393525 -20212
rect 393581 -20268 393648 -20212
rect 393308 -20354 393648 -20268
rect 393308 -20410 393383 -20354
rect 393439 -20410 393525 -20354
rect 393581 -20410 393648 -20354
rect 393308 -20496 393648 -20410
rect 393308 -20552 393383 -20496
rect 393439 -20552 393525 -20496
rect 393581 -20552 393648 -20496
rect 393308 -20638 393648 -20552
rect 393308 -20694 393383 -20638
rect 393439 -20694 393525 -20638
rect 393581 -20694 393648 -20638
rect 393308 -20780 393648 -20694
rect 393308 -20836 393383 -20780
rect 393439 -20836 393525 -20780
rect 393581 -20836 393648 -20780
rect 393308 -20922 393648 -20836
rect 393308 -20978 393383 -20922
rect 393439 -20978 393525 -20922
rect 393581 -20978 393648 -20922
rect 393308 -21064 393648 -20978
rect 393308 -21120 393383 -21064
rect 393439 -21120 393525 -21064
rect 393581 -21120 393648 -21064
rect 393308 -21206 393648 -21120
rect 393308 -21262 393383 -21206
rect 393439 -21262 393525 -21206
rect 393581 -21262 393648 -21206
rect 393308 -21348 393648 -21262
rect 393308 -21404 393383 -21348
rect 393439 -21404 393525 -21348
rect 393581 -21404 393648 -21348
rect 393308 -21490 393648 -21404
rect 393308 -21546 393383 -21490
rect 393439 -21546 393525 -21490
rect 393581 -21546 393648 -21490
rect 393308 -21632 393648 -21546
rect 393308 -21688 393383 -21632
rect 393439 -21688 393525 -21632
rect 393581 -21688 393648 -21632
rect 393308 -21774 393648 -21688
rect 393308 -21830 393383 -21774
rect 393439 -21830 393525 -21774
rect 393581 -21830 393648 -21774
rect 393308 -21916 393648 -21830
rect 393308 -21972 393383 -21916
rect 393439 -21972 393525 -21916
rect 393581 -21972 393648 -21916
rect 393308 -22058 393648 -21972
rect 393308 -22114 393383 -22058
rect 393439 -22114 393525 -22058
rect 393581 -22114 393648 -22058
rect 393308 -22200 393648 -22114
rect 393308 -22256 393383 -22200
rect 393439 -22256 393525 -22200
rect 393581 -22256 393648 -22200
rect 393308 -22342 393648 -22256
rect 393308 -22398 393383 -22342
rect 393439 -22398 393525 -22342
rect 393581 -22398 393648 -22342
rect 393308 -22484 393648 -22398
rect 393308 -22540 393383 -22484
rect 393439 -22540 393525 -22484
rect 393581 -22540 393648 -22484
rect 393308 -22626 393648 -22540
rect 393308 -22682 393383 -22626
rect 393439 -22682 393525 -22626
rect 393581 -22682 393648 -22626
rect 393308 -22768 393648 -22682
rect 393308 -22824 393383 -22768
rect 393439 -22824 393525 -22768
rect 393581 -22824 393648 -22768
rect 393308 -22910 393648 -22824
rect 393308 -22966 393383 -22910
rect 393439 -22966 393525 -22910
rect 393581 -22966 393648 -22910
rect 393308 -23052 393648 -22966
rect 393308 -23108 393383 -23052
rect 393439 -23108 393525 -23052
rect 393581 -23108 393648 -23052
rect 393308 -23194 393648 -23108
rect 393308 -23250 393383 -23194
rect 393439 -23250 393525 -23194
rect 393581 -23250 393648 -23194
rect 393308 -23336 393648 -23250
rect 393308 -23392 393383 -23336
rect 393439 -23392 393525 -23336
rect 393581 -23392 393648 -23336
rect 393308 -23478 393648 -23392
rect 393308 -23534 393383 -23478
rect 393439 -23534 393525 -23478
rect 393581 -23534 393648 -23478
rect 393308 -23620 393648 -23534
rect 393308 -23676 393383 -23620
rect 393439 -23676 393525 -23620
rect 393581 -23676 393648 -23620
rect 393308 -23762 393648 -23676
rect 393308 -23818 393383 -23762
rect 393439 -23818 393525 -23762
rect 393581 -23818 393648 -23762
rect 393308 -23904 393648 -23818
rect 393308 -23960 393383 -23904
rect 393439 -23960 393525 -23904
rect 393581 -23960 393648 -23904
rect 393308 -24046 393648 -23960
rect 393308 -24102 393383 -24046
rect 393439 -24102 393525 -24046
rect 393581 -24102 393648 -24046
rect 393308 -24188 393648 -24102
rect 393308 -24244 393383 -24188
rect 393439 -24244 393525 -24188
rect 393581 -24244 393648 -24188
rect 393308 -24330 393648 -24244
rect 393308 -24386 393383 -24330
rect 393439 -24386 393525 -24330
rect 393581 -24386 393648 -24330
rect 393308 -24472 393648 -24386
rect 393308 -24528 393383 -24472
rect 393439 -24528 393525 -24472
rect 393581 -24528 393648 -24472
rect 393308 -24614 393648 -24528
rect 393308 -24670 393383 -24614
rect 393439 -24670 393525 -24614
rect 393581 -24670 393648 -24614
rect 393308 -24756 393648 -24670
rect 393308 -24812 393383 -24756
rect 393439 -24812 393525 -24756
rect 393581 -24812 393648 -24756
rect 393308 -24898 393648 -24812
rect 393308 -24954 393383 -24898
rect 393439 -24954 393525 -24898
rect 393581 -24954 393648 -24898
rect 393308 -25040 393648 -24954
rect 393308 -25096 393383 -25040
rect 393439 -25096 393525 -25040
rect 393581 -25096 393648 -25040
rect 393308 -25182 393648 -25096
rect 393308 -25238 393383 -25182
rect 393439 -25238 393525 -25182
rect 393581 -25238 393648 -25182
rect 393308 -25324 393648 -25238
rect 393308 -25380 393383 -25324
rect 393439 -25380 393525 -25324
rect 393581 -25380 393648 -25324
rect 393308 -25466 393648 -25380
rect 393308 -25522 393383 -25466
rect 393439 -25522 393525 -25466
rect 393581 -25522 393648 -25466
rect 393308 -25590 393648 -25522
rect 393708 -13680 394048 -13590
rect 393708 -13736 393780 -13680
rect 393836 -13736 393922 -13680
rect 393978 -13736 394048 -13680
rect 393708 -13822 394048 -13736
rect 393708 -13878 393780 -13822
rect 393836 -13878 393922 -13822
rect 393978 -13878 394048 -13822
rect 393708 -13964 394048 -13878
rect 393708 -14020 393780 -13964
rect 393836 -14020 393922 -13964
rect 393978 -14020 394048 -13964
rect 393708 -14106 394048 -14020
rect 393708 -14162 393780 -14106
rect 393836 -14162 393922 -14106
rect 393978 -14162 394048 -14106
rect 393708 -14248 394048 -14162
rect 393708 -14304 393780 -14248
rect 393836 -14304 393922 -14248
rect 393978 -14304 394048 -14248
rect 393708 -14390 394048 -14304
rect 393708 -14446 393780 -14390
rect 393836 -14446 393922 -14390
rect 393978 -14446 394048 -14390
rect 393708 -14532 394048 -14446
rect 393708 -14588 393780 -14532
rect 393836 -14588 393922 -14532
rect 393978 -14588 394048 -14532
rect 393708 -14674 394048 -14588
rect 393708 -14730 393780 -14674
rect 393836 -14730 393922 -14674
rect 393978 -14730 394048 -14674
rect 393708 -14816 394048 -14730
rect 393708 -14872 393780 -14816
rect 393836 -14872 393922 -14816
rect 393978 -14872 394048 -14816
rect 393708 -14958 394048 -14872
rect 393708 -15014 393780 -14958
rect 393836 -15014 393922 -14958
rect 393978 -15014 394048 -14958
rect 393708 -15100 394048 -15014
rect 393708 -15156 393780 -15100
rect 393836 -15156 393922 -15100
rect 393978 -15156 394048 -15100
rect 393708 -15242 394048 -15156
rect 393708 -15298 393780 -15242
rect 393836 -15298 393922 -15242
rect 393978 -15298 394048 -15242
rect 393708 -15384 394048 -15298
rect 393708 -15440 393780 -15384
rect 393836 -15440 393922 -15384
rect 393978 -15440 394048 -15384
rect 393708 -15526 394048 -15440
rect 393708 -15582 393780 -15526
rect 393836 -15582 393922 -15526
rect 393978 -15582 394048 -15526
rect 393708 -15668 394048 -15582
rect 393708 -15724 393780 -15668
rect 393836 -15724 393922 -15668
rect 393978 -15724 394048 -15668
rect 393708 -15810 394048 -15724
rect 393708 -15866 393780 -15810
rect 393836 -15866 393922 -15810
rect 393978 -15866 394048 -15810
rect 393708 -15952 394048 -15866
rect 393708 -16008 393780 -15952
rect 393836 -16008 393922 -15952
rect 393978 -16008 394048 -15952
rect 393708 -16094 394048 -16008
rect 393708 -16150 393780 -16094
rect 393836 -16150 393922 -16094
rect 393978 -16150 394048 -16094
rect 393708 -16236 394048 -16150
rect 393708 -16292 393780 -16236
rect 393836 -16292 393922 -16236
rect 393978 -16292 394048 -16236
rect 393708 -16378 394048 -16292
rect 393708 -16434 393780 -16378
rect 393836 -16434 393922 -16378
rect 393978 -16434 394048 -16378
rect 393708 -16520 394048 -16434
rect 393708 -16576 393780 -16520
rect 393836 -16576 393922 -16520
rect 393978 -16576 394048 -16520
rect 393708 -16662 394048 -16576
rect 393708 -16718 393780 -16662
rect 393836 -16718 393922 -16662
rect 393978 -16718 394048 -16662
rect 393708 -16804 394048 -16718
rect 393708 -16860 393780 -16804
rect 393836 -16860 393922 -16804
rect 393978 -16860 394048 -16804
rect 393708 -16946 394048 -16860
rect 393708 -17002 393780 -16946
rect 393836 -17002 393922 -16946
rect 393978 -17002 394048 -16946
rect 393708 -17088 394048 -17002
rect 393708 -17144 393780 -17088
rect 393836 -17144 393922 -17088
rect 393978 -17144 394048 -17088
rect 393708 -17230 394048 -17144
rect 393708 -17286 393780 -17230
rect 393836 -17286 393922 -17230
rect 393978 -17286 394048 -17230
rect 393708 -17372 394048 -17286
rect 393708 -17428 393780 -17372
rect 393836 -17428 393922 -17372
rect 393978 -17428 394048 -17372
rect 393708 -17514 394048 -17428
rect 393708 -17570 393780 -17514
rect 393836 -17570 393922 -17514
rect 393978 -17570 394048 -17514
rect 393708 -17656 394048 -17570
rect 393708 -17712 393780 -17656
rect 393836 -17712 393922 -17656
rect 393978 -17712 394048 -17656
rect 393708 -17798 394048 -17712
rect 393708 -17854 393780 -17798
rect 393836 -17854 393922 -17798
rect 393978 -17854 394048 -17798
rect 393708 -17940 394048 -17854
rect 393708 -17996 393780 -17940
rect 393836 -17996 393922 -17940
rect 393978 -17996 394048 -17940
rect 393708 -18082 394048 -17996
rect 393708 -18138 393780 -18082
rect 393836 -18138 393922 -18082
rect 393978 -18138 394048 -18082
rect 393708 -18224 394048 -18138
rect 393708 -18280 393780 -18224
rect 393836 -18280 393922 -18224
rect 393978 -18280 394048 -18224
rect 393708 -18366 394048 -18280
rect 393708 -18422 393780 -18366
rect 393836 -18422 393922 -18366
rect 393978 -18422 394048 -18366
rect 393708 -18508 394048 -18422
rect 393708 -18564 393780 -18508
rect 393836 -18564 393922 -18508
rect 393978 -18564 394048 -18508
rect 393708 -18650 394048 -18564
rect 393708 -18706 393780 -18650
rect 393836 -18706 393922 -18650
rect 393978 -18706 394048 -18650
rect 393708 -18792 394048 -18706
rect 393708 -18848 393780 -18792
rect 393836 -18848 393922 -18792
rect 393978 -18848 394048 -18792
rect 393708 -18934 394048 -18848
rect 393708 -18990 393780 -18934
rect 393836 -18990 393922 -18934
rect 393978 -18990 394048 -18934
rect 393708 -19076 394048 -18990
rect 393708 -19132 393780 -19076
rect 393836 -19132 393922 -19076
rect 393978 -19132 394048 -19076
rect 393708 -19218 394048 -19132
rect 393708 -19274 393780 -19218
rect 393836 -19274 393922 -19218
rect 393978 -19274 394048 -19218
rect 393708 -19360 394048 -19274
rect 393708 -19416 393780 -19360
rect 393836 -19416 393922 -19360
rect 393978 -19416 394048 -19360
rect 393708 -19502 394048 -19416
rect 393708 -19558 393780 -19502
rect 393836 -19558 393922 -19502
rect 393978 -19558 394048 -19502
rect 393708 -19644 394048 -19558
rect 393708 -19700 393780 -19644
rect 393836 -19700 393922 -19644
rect 393978 -19700 394048 -19644
rect 393708 -19786 394048 -19700
rect 393708 -19842 393780 -19786
rect 393836 -19842 393922 -19786
rect 393978 -19842 394048 -19786
rect 393708 -19928 394048 -19842
rect 393708 -19984 393780 -19928
rect 393836 -19984 393922 -19928
rect 393978 -19984 394048 -19928
rect 393708 -20070 394048 -19984
rect 393708 -20126 393780 -20070
rect 393836 -20126 393922 -20070
rect 393978 -20126 394048 -20070
rect 393708 -20212 394048 -20126
rect 393708 -20268 393780 -20212
rect 393836 -20268 393922 -20212
rect 393978 -20268 394048 -20212
rect 393708 -20354 394048 -20268
rect 393708 -20410 393780 -20354
rect 393836 -20410 393922 -20354
rect 393978 -20410 394048 -20354
rect 393708 -20496 394048 -20410
rect 393708 -20552 393780 -20496
rect 393836 -20552 393922 -20496
rect 393978 -20552 394048 -20496
rect 393708 -20638 394048 -20552
rect 393708 -20694 393780 -20638
rect 393836 -20694 393922 -20638
rect 393978 -20694 394048 -20638
rect 393708 -20780 394048 -20694
rect 393708 -20836 393780 -20780
rect 393836 -20836 393922 -20780
rect 393978 -20836 394048 -20780
rect 393708 -20922 394048 -20836
rect 393708 -20978 393780 -20922
rect 393836 -20978 393922 -20922
rect 393978 -20978 394048 -20922
rect 393708 -21064 394048 -20978
rect 393708 -21120 393780 -21064
rect 393836 -21120 393922 -21064
rect 393978 -21120 394048 -21064
rect 393708 -21206 394048 -21120
rect 393708 -21262 393780 -21206
rect 393836 -21262 393922 -21206
rect 393978 -21262 394048 -21206
rect 393708 -21348 394048 -21262
rect 393708 -21404 393780 -21348
rect 393836 -21404 393922 -21348
rect 393978 -21404 394048 -21348
rect 393708 -21490 394048 -21404
rect 393708 -21546 393780 -21490
rect 393836 -21546 393922 -21490
rect 393978 -21546 394048 -21490
rect 393708 -21632 394048 -21546
rect 393708 -21688 393780 -21632
rect 393836 -21688 393922 -21632
rect 393978 -21688 394048 -21632
rect 393708 -21774 394048 -21688
rect 393708 -21830 393780 -21774
rect 393836 -21830 393922 -21774
rect 393978 -21830 394048 -21774
rect 393708 -21916 394048 -21830
rect 393708 -21972 393780 -21916
rect 393836 -21972 393922 -21916
rect 393978 -21972 394048 -21916
rect 393708 -22058 394048 -21972
rect 393708 -22114 393780 -22058
rect 393836 -22114 393922 -22058
rect 393978 -22114 394048 -22058
rect 393708 -22200 394048 -22114
rect 393708 -22256 393780 -22200
rect 393836 -22256 393922 -22200
rect 393978 -22256 394048 -22200
rect 393708 -22342 394048 -22256
rect 393708 -22398 393780 -22342
rect 393836 -22398 393922 -22342
rect 393978 -22398 394048 -22342
rect 393708 -22484 394048 -22398
rect 393708 -22540 393780 -22484
rect 393836 -22540 393922 -22484
rect 393978 -22540 394048 -22484
rect 393708 -22626 394048 -22540
rect 393708 -22682 393780 -22626
rect 393836 -22682 393922 -22626
rect 393978 -22682 394048 -22626
rect 393708 -22768 394048 -22682
rect 393708 -22824 393780 -22768
rect 393836 -22824 393922 -22768
rect 393978 -22824 394048 -22768
rect 393708 -22910 394048 -22824
rect 393708 -22966 393780 -22910
rect 393836 -22966 393922 -22910
rect 393978 -22966 394048 -22910
rect 393708 -23052 394048 -22966
rect 393708 -23108 393780 -23052
rect 393836 -23108 393922 -23052
rect 393978 -23108 394048 -23052
rect 393708 -23194 394048 -23108
rect 393708 -23250 393780 -23194
rect 393836 -23250 393922 -23194
rect 393978 -23250 394048 -23194
rect 393708 -23336 394048 -23250
rect 393708 -23392 393780 -23336
rect 393836 -23392 393922 -23336
rect 393978 -23392 394048 -23336
rect 393708 -23478 394048 -23392
rect 393708 -23534 393780 -23478
rect 393836 -23534 393922 -23478
rect 393978 -23534 394048 -23478
rect 393708 -23620 394048 -23534
rect 393708 -23676 393780 -23620
rect 393836 -23676 393922 -23620
rect 393978 -23676 394048 -23620
rect 393708 -23762 394048 -23676
rect 393708 -23818 393780 -23762
rect 393836 -23818 393922 -23762
rect 393978 -23818 394048 -23762
rect 393708 -23904 394048 -23818
rect 393708 -23960 393780 -23904
rect 393836 -23960 393922 -23904
rect 393978 -23960 394048 -23904
rect 393708 -24046 394048 -23960
rect 393708 -24102 393780 -24046
rect 393836 -24102 393922 -24046
rect 393978 -24102 394048 -24046
rect 393708 -24188 394048 -24102
rect 393708 -24244 393780 -24188
rect 393836 -24244 393922 -24188
rect 393978 -24244 394048 -24188
rect 393708 -24330 394048 -24244
rect 393708 -24386 393780 -24330
rect 393836 -24386 393922 -24330
rect 393978 -24386 394048 -24330
rect 393708 -24472 394048 -24386
rect 393708 -24528 393780 -24472
rect 393836 -24528 393922 -24472
rect 393978 -24528 394048 -24472
rect 393708 -24614 394048 -24528
rect 393708 -24670 393780 -24614
rect 393836 -24670 393922 -24614
rect 393978 -24670 394048 -24614
rect 393708 -24756 394048 -24670
rect 393708 -24812 393780 -24756
rect 393836 -24812 393922 -24756
rect 393978 -24812 394048 -24756
rect 393708 -24898 394048 -24812
rect 393708 -24954 393780 -24898
rect 393836 -24954 393922 -24898
rect 393978 -24954 394048 -24898
rect 393708 -25040 394048 -24954
rect 393708 -25096 393780 -25040
rect 393836 -25096 393922 -25040
rect 393978 -25096 394048 -25040
rect 393708 -25182 394048 -25096
rect 393708 -25238 393780 -25182
rect 393836 -25238 393922 -25182
rect 393978 -25238 394048 -25182
rect 393708 -25324 394048 -25238
rect 393708 -25380 393780 -25324
rect 393836 -25380 393922 -25324
rect 393978 -25380 394048 -25324
rect 393708 -25466 394048 -25380
rect 393708 -25522 393780 -25466
rect 393836 -25522 393922 -25466
rect 393978 -25522 394048 -25466
rect 393708 -25590 394048 -25522
rect 394108 -13680 394448 -13590
rect 394108 -13736 394177 -13680
rect 394233 -13736 394319 -13680
rect 394375 -13736 394448 -13680
rect 394108 -13822 394448 -13736
rect 394108 -13878 394177 -13822
rect 394233 -13878 394319 -13822
rect 394375 -13878 394448 -13822
rect 394108 -13964 394448 -13878
rect 394108 -14020 394177 -13964
rect 394233 -14020 394319 -13964
rect 394375 -14020 394448 -13964
rect 394108 -14106 394448 -14020
rect 394108 -14162 394177 -14106
rect 394233 -14162 394319 -14106
rect 394375 -14162 394448 -14106
rect 394108 -14248 394448 -14162
rect 394108 -14304 394177 -14248
rect 394233 -14304 394319 -14248
rect 394375 -14304 394448 -14248
rect 394108 -14390 394448 -14304
rect 394108 -14446 394177 -14390
rect 394233 -14446 394319 -14390
rect 394375 -14446 394448 -14390
rect 394108 -14532 394448 -14446
rect 394108 -14588 394177 -14532
rect 394233 -14588 394319 -14532
rect 394375 -14588 394448 -14532
rect 394108 -14674 394448 -14588
rect 394108 -14730 394177 -14674
rect 394233 -14730 394319 -14674
rect 394375 -14730 394448 -14674
rect 394108 -14816 394448 -14730
rect 394108 -14872 394177 -14816
rect 394233 -14872 394319 -14816
rect 394375 -14872 394448 -14816
rect 394108 -14958 394448 -14872
rect 394108 -15014 394177 -14958
rect 394233 -15014 394319 -14958
rect 394375 -15014 394448 -14958
rect 394108 -15100 394448 -15014
rect 394108 -15156 394177 -15100
rect 394233 -15156 394319 -15100
rect 394375 -15156 394448 -15100
rect 394108 -15242 394448 -15156
rect 394108 -15298 394177 -15242
rect 394233 -15298 394319 -15242
rect 394375 -15298 394448 -15242
rect 394108 -15384 394448 -15298
rect 394108 -15440 394177 -15384
rect 394233 -15440 394319 -15384
rect 394375 -15440 394448 -15384
rect 394108 -15526 394448 -15440
rect 394108 -15582 394177 -15526
rect 394233 -15582 394319 -15526
rect 394375 -15582 394448 -15526
rect 394108 -15668 394448 -15582
rect 394108 -15724 394177 -15668
rect 394233 -15724 394319 -15668
rect 394375 -15724 394448 -15668
rect 394108 -15810 394448 -15724
rect 394108 -15866 394177 -15810
rect 394233 -15866 394319 -15810
rect 394375 -15866 394448 -15810
rect 394108 -15952 394448 -15866
rect 394108 -16008 394177 -15952
rect 394233 -16008 394319 -15952
rect 394375 -16008 394448 -15952
rect 394108 -16094 394448 -16008
rect 394108 -16150 394177 -16094
rect 394233 -16150 394319 -16094
rect 394375 -16150 394448 -16094
rect 394108 -16236 394448 -16150
rect 394108 -16292 394177 -16236
rect 394233 -16292 394319 -16236
rect 394375 -16292 394448 -16236
rect 394108 -16378 394448 -16292
rect 394108 -16434 394177 -16378
rect 394233 -16434 394319 -16378
rect 394375 -16434 394448 -16378
rect 394108 -16520 394448 -16434
rect 394108 -16576 394177 -16520
rect 394233 -16576 394319 -16520
rect 394375 -16576 394448 -16520
rect 394108 -16662 394448 -16576
rect 394108 -16718 394177 -16662
rect 394233 -16718 394319 -16662
rect 394375 -16718 394448 -16662
rect 394108 -16804 394448 -16718
rect 394108 -16860 394177 -16804
rect 394233 -16860 394319 -16804
rect 394375 -16860 394448 -16804
rect 394108 -16946 394448 -16860
rect 394108 -17002 394177 -16946
rect 394233 -17002 394319 -16946
rect 394375 -17002 394448 -16946
rect 394108 -17088 394448 -17002
rect 394108 -17144 394177 -17088
rect 394233 -17144 394319 -17088
rect 394375 -17144 394448 -17088
rect 394108 -17230 394448 -17144
rect 394108 -17286 394177 -17230
rect 394233 -17286 394319 -17230
rect 394375 -17286 394448 -17230
rect 394108 -17372 394448 -17286
rect 394108 -17428 394177 -17372
rect 394233 -17428 394319 -17372
rect 394375 -17428 394448 -17372
rect 394108 -17514 394448 -17428
rect 394108 -17570 394177 -17514
rect 394233 -17570 394319 -17514
rect 394375 -17570 394448 -17514
rect 394108 -17656 394448 -17570
rect 394108 -17712 394177 -17656
rect 394233 -17712 394319 -17656
rect 394375 -17712 394448 -17656
rect 394108 -17798 394448 -17712
rect 394108 -17854 394177 -17798
rect 394233 -17854 394319 -17798
rect 394375 -17854 394448 -17798
rect 394108 -17940 394448 -17854
rect 394108 -17996 394177 -17940
rect 394233 -17996 394319 -17940
rect 394375 -17996 394448 -17940
rect 394108 -18082 394448 -17996
rect 394108 -18138 394177 -18082
rect 394233 -18138 394319 -18082
rect 394375 -18138 394448 -18082
rect 394108 -18224 394448 -18138
rect 394108 -18280 394177 -18224
rect 394233 -18280 394319 -18224
rect 394375 -18280 394448 -18224
rect 394108 -18366 394448 -18280
rect 394108 -18422 394177 -18366
rect 394233 -18422 394319 -18366
rect 394375 -18422 394448 -18366
rect 394108 -18508 394448 -18422
rect 394108 -18564 394177 -18508
rect 394233 -18564 394319 -18508
rect 394375 -18564 394448 -18508
rect 394108 -18650 394448 -18564
rect 394108 -18706 394177 -18650
rect 394233 -18706 394319 -18650
rect 394375 -18706 394448 -18650
rect 394108 -18792 394448 -18706
rect 394108 -18848 394177 -18792
rect 394233 -18848 394319 -18792
rect 394375 -18848 394448 -18792
rect 394108 -18934 394448 -18848
rect 394108 -18990 394177 -18934
rect 394233 -18990 394319 -18934
rect 394375 -18990 394448 -18934
rect 394108 -19076 394448 -18990
rect 394108 -19132 394177 -19076
rect 394233 -19132 394319 -19076
rect 394375 -19132 394448 -19076
rect 394108 -19218 394448 -19132
rect 394108 -19274 394177 -19218
rect 394233 -19274 394319 -19218
rect 394375 -19274 394448 -19218
rect 394108 -19360 394448 -19274
rect 394108 -19416 394177 -19360
rect 394233 -19416 394319 -19360
rect 394375 -19416 394448 -19360
rect 394108 -19502 394448 -19416
rect 394108 -19558 394177 -19502
rect 394233 -19558 394319 -19502
rect 394375 -19558 394448 -19502
rect 394108 -19644 394448 -19558
rect 394108 -19700 394177 -19644
rect 394233 -19700 394319 -19644
rect 394375 -19700 394448 -19644
rect 394108 -19786 394448 -19700
rect 394108 -19842 394177 -19786
rect 394233 -19842 394319 -19786
rect 394375 -19842 394448 -19786
rect 394108 -19928 394448 -19842
rect 394108 -19984 394177 -19928
rect 394233 -19984 394319 -19928
rect 394375 -19984 394448 -19928
rect 394108 -20070 394448 -19984
rect 394108 -20126 394177 -20070
rect 394233 -20126 394319 -20070
rect 394375 -20126 394448 -20070
rect 394108 -20212 394448 -20126
rect 394108 -20268 394177 -20212
rect 394233 -20268 394319 -20212
rect 394375 -20268 394448 -20212
rect 394108 -20354 394448 -20268
rect 394108 -20410 394177 -20354
rect 394233 -20410 394319 -20354
rect 394375 -20410 394448 -20354
rect 394108 -20496 394448 -20410
rect 394108 -20552 394177 -20496
rect 394233 -20552 394319 -20496
rect 394375 -20552 394448 -20496
rect 394108 -20638 394448 -20552
rect 394108 -20694 394177 -20638
rect 394233 -20694 394319 -20638
rect 394375 -20694 394448 -20638
rect 394108 -20780 394448 -20694
rect 394108 -20836 394177 -20780
rect 394233 -20836 394319 -20780
rect 394375 -20836 394448 -20780
rect 394108 -20922 394448 -20836
rect 394108 -20978 394177 -20922
rect 394233 -20978 394319 -20922
rect 394375 -20978 394448 -20922
rect 394108 -21064 394448 -20978
rect 394108 -21120 394177 -21064
rect 394233 -21120 394319 -21064
rect 394375 -21120 394448 -21064
rect 394108 -21206 394448 -21120
rect 394108 -21262 394177 -21206
rect 394233 -21262 394319 -21206
rect 394375 -21262 394448 -21206
rect 394108 -21348 394448 -21262
rect 394108 -21404 394177 -21348
rect 394233 -21404 394319 -21348
rect 394375 -21404 394448 -21348
rect 394108 -21490 394448 -21404
rect 394108 -21546 394177 -21490
rect 394233 -21546 394319 -21490
rect 394375 -21546 394448 -21490
rect 394108 -21632 394448 -21546
rect 394108 -21688 394177 -21632
rect 394233 -21688 394319 -21632
rect 394375 -21688 394448 -21632
rect 394108 -21774 394448 -21688
rect 394108 -21830 394177 -21774
rect 394233 -21830 394319 -21774
rect 394375 -21830 394448 -21774
rect 394108 -21916 394448 -21830
rect 394108 -21972 394177 -21916
rect 394233 -21972 394319 -21916
rect 394375 -21972 394448 -21916
rect 394108 -22058 394448 -21972
rect 394108 -22114 394177 -22058
rect 394233 -22114 394319 -22058
rect 394375 -22114 394448 -22058
rect 394108 -22200 394448 -22114
rect 394108 -22256 394177 -22200
rect 394233 -22256 394319 -22200
rect 394375 -22256 394448 -22200
rect 394108 -22342 394448 -22256
rect 394108 -22398 394177 -22342
rect 394233 -22398 394319 -22342
rect 394375 -22398 394448 -22342
rect 394108 -22484 394448 -22398
rect 394108 -22540 394177 -22484
rect 394233 -22540 394319 -22484
rect 394375 -22540 394448 -22484
rect 394108 -22626 394448 -22540
rect 394108 -22682 394177 -22626
rect 394233 -22682 394319 -22626
rect 394375 -22682 394448 -22626
rect 394108 -22768 394448 -22682
rect 394108 -22824 394177 -22768
rect 394233 -22824 394319 -22768
rect 394375 -22824 394448 -22768
rect 394108 -22910 394448 -22824
rect 394108 -22966 394177 -22910
rect 394233 -22966 394319 -22910
rect 394375 -22966 394448 -22910
rect 394108 -23052 394448 -22966
rect 394108 -23108 394177 -23052
rect 394233 -23108 394319 -23052
rect 394375 -23108 394448 -23052
rect 394108 -23194 394448 -23108
rect 394108 -23250 394177 -23194
rect 394233 -23250 394319 -23194
rect 394375 -23250 394448 -23194
rect 394108 -23336 394448 -23250
rect 394108 -23392 394177 -23336
rect 394233 -23392 394319 -23336
rect 394375 -23392 394448 -23336
rect 394108 -23478 394448 -23392
rect 394108 -23534 394177 -23478
rect 394233 -23534 394319 -23478
rect 394375 -23534 394448 -23478
rect 394108 -23620 394448 -23534
rect 394108 -23676 394177 -23620
rect 394233 -23676 394319 -23620
rect 394375 -23676 394448 -23620
rect 394108 -23762 394448 -23676
rect 394108 -23818 394177 -23762
rect 394233 -23818 394319 -23762
rect 394375 -23818 394448 -23762
rect 394108 -23904 394448 -23818
rect 394108 -23960 394177 -23904
rect 394233 -23960 394319 -23904
rect 394375 -23960 394448 -23904
rect 394108 -24046 394448 -23960
rect 394108 -24102 394177 -24046
rect 394233 -24102 394319 -24046
rect 394375 -24102 394448 -24046
rect 394108 -24188 394448 -24102
rect 394108 -24244 394177 -24188
rect 394233 -24244 394319 -24188
rect 394375 -24244 394448 -24188
rect 394108 -24330 394448 -24244
rect 394108 -24386 394177 -24330
rect 394233 -24386 394319 -24330
rect 394375 -24386 394448 -24330
rect 394108 -24472 394448 -24386
rect 394108 -24528 394177 -24472
rect 394233 -24528 394319 -24472
rect 394375 -24528 394448 -24472
rect 394108 -24614 394448 -24528
rect 394108 -24670 394177 -24614
rect 394233 -24670 394319 -24614
rect 394375 -24670 394448 -24614
rect 394108 -24756 394448 -24670
rect 394108 -24812 394177 -24756
rect 394233 -24812 394319 -24756
rect 394375 -24812 394448 -24756
rect 394108 -24898 394448 -24812
rect 394108 -24954 394177 -24898
rect 394233 -24954 394319 -24898
rect 394375 -24954 394448 -24898
rect 394108 -25040 394448 -24954
rect 394108 -25096 394177 -25040
rect 394233 -25096 394319 -25040
rect 394375 -25096 394448 -25040
rect 394108 -25182 394448 -25096
rect 394108 -25238 394177 -25182
rect 394233 -25238 394319 -25182
rect 394375 -25238 394448 -25182
rect 394108 -25324 394448 -25238
rect 394108 -25380 394177 -25324
rect 394233 -25380 394319 -25324
rect 394375 -25380 394448 -25324
rect 394108 -25466 394448 -25380
rect 394108 -25522 394177 -25466
rect 394233 -25522 394319 -25466
rect 394375 -25522 394448 -25466
rect 394108 -25590 394448 -25522
rect 394508 -13680 394848 -13590
rect 394508 -13736 394580 -13680
rect 394636 -13736 394722 -13680
rect 394778 -13736 394848 -13680
rect 394508 -13822 394848 -13736
rect 394508 -13878 394580 -13822
rect 394636 -13878 394722 -13822
rect 394778 -13878 394848 -13822
rect 394508 -13964 394848 -13878
rect 394508 -14020 394580 -13964
rect 394636 -14020 394722 -13964
rect 394778 -14020 394848 -13964
rect 394508 -14106 394848 -14020
rect 394508 -14162 394580 -14106
rect 394636 -14162 394722 -14106
rect 394778 -14162 394848 -14106
rect 394508 -14248 394848 -14162
rect 394508 -14304 394580 -14248
rect 394636 -14304 394722 -14248
rect 394778 -14304 394848 -14248
rect 394508 -14390 394848 -14304
rect 394508 -14446 394580 -14390
rect 394636 -14446 394722 -14390
rect 394778 -14446 394848 -14390
rect 394508 -14532 394848 -14446
rect 394508 -14588 394580 -14532
rect 394636 -14588 394722 -14532
rect 394778 -14588 394848 -14532
rect 394508 -14674 394848 -14588
rect 394508 -14730 394580 -14674
rect 394636 -14730 394722 -14674
rect 394778 -14730 394848 -14674
rect 394508 -14816 394848 -14730
rect 394508 -14872 394580 -14816
rect 394636 -14872 394722 -14816
rect 394778 -14872 394848 -14816
rect 394508 -14958 394848 -14872
rect 394508 -15014 394580 -14958
rect 394636 -15014 394722 -14958
rect 394778 -15014 394848 -14958
rect 394508 -15100 394848 -15014
rect 394508 -15156 394580 -15100
rect 394636 -15156 394722 -15100
rect 394778 -15156 394848 -15100
rect 394508 -15242 394848 -15156
rect 394508 -15298 394580 -15242
rect 394636 -15298 394722 -15242
rect 394778 -15298 394848 -15242
rect 394508 -15384 394848 -15298
rect 394508 -15440 394580 -15384
rect 394636 -15440 394722 -15384
rect 394778 -15440 394848 -15384
rect 394508 -15526 394848 -15440
rect 394508 -15582 394580 -15526
rect 394636 -15582 394722 -15526
rect 394778 -15582 394848 -15526
rect 394508 -15668 394848 -15582
rect 394508 -15724 394580 -15668
rect 394636 -15724 394722 -15668
rect 394778 -15724 394848 -15668
rect 394508 -15810 394848 -15724
rect 394508 -15866 394580 -15810
rect 394636 -15866 394722 -15810
rect 394778 -15866 394848 -15810
rect 394508 -15952 394848 -15866
rect 394508 -16008 394580 -15952
rect 394636 -16008 394722 -15952
rect 394778 -16008 394848 -15952
rect 394508 -16094 394848 -16008
rect 394508 -16150 394580 -16094
rect 394636 -16150 394722 -16094
rect 394778 -16150 394848 -16094
rect 394508 -16236 394848 -16150
rect 394508 -16292 394580 -16236
rect 394636 -16292 394722 -16236
rect 394778 -16292 394848 -16236
rect 394508 -16378 394848 -16292
rect 394508 -16434 394580 -16378
rect 394636 -16434 394722 -16378
rect 394778 -16434 394848 -16378
rect 394508 -16520 394848 -16434
rect 394508 -16576 394580 -16520
rect 394636 -16576 394722 -16520
rect 394778 -16576 394848 -16520
rect 394508 -16662 394848 -16576
rect 394508 -16718 394580 -16662
rect 394636 -16718 394722 -16662
rect 394778 -16718 394848 -16662
rect 394508 -16804 394848 -16718
rect 394508 -16860 394580 -16804
rect 394636 -16860 394722 -16804
rect 394778 -16860 394848 -16804
rect 394508 -16946 394848 -16860
rect 394508 -17002 394580 -16946
rect 394636 -17002 394722 -16946
rect 394778 -17002 394848 -16946
rect 394508 -17088 394848 -17002
rect 394508 -17144 394580 -17088
rect 394636 -17144 394722 -17088
rect 394778 -17144 394848 -17088
rect 394508 -17230 394848 -17144
rect 394508 -17286 394580 -17230
rect 394636 -17286 394722 -17230
rect 394778 -17286 394848 -17230
rect 394508 -17372 394848 -17286
rect 394508 -17428 394580 -17372
rect 394636 -17428 394722 -17372
rect 394778 -17428 394848 -17372
rect 394508 -17514 394848 -17428
rect 394508 -17570 394580 -17514
rect 394636 -17570 394722 -17514
rect 394778 -17570 394848 -17514
rect 394508 -17656 394848 -17570
rect 394508 -17712 394580 -17656
rect 394636 -17712 394722 -17656
rect 394778 -17712 394848 -17656
rect 394508 -17798 394848 -17712
rect 394508 -17854 394580 -17798
rect 394636 -17854 394722 -17798
rect 394778 -17854 394848 -17798
rect 394508 -17940 394848 -17854
rect 394508 -17996 394580 -17940
rect 394636 -17996 394722 -17940
rect 394778 -17996 394848 -17940
rect 394508 -18082 394848 -17996
rect 394508 -18138 394580 -18082
rect 394636 -18138 394722 -18082
rect 394778 -18138 394848 -18082
rect 394508 -18224 394848 -18138
rect 394508 -18280 394580 -18224
rect 394636 -18280 394722 -18224
rect 394778 -18280 394848 -18224
rect 394508 -18366 394848 -18280
rect 394508 -18422 394580 -18366
rect 394636 -18422 394722 -18366
rect 394778 -18422 394848 -18366
rect 394508 -18508 394848 -18422
rect 394508 -18564 394580 -18508
rect 394636 -18564 394722 -18508
rect 394778 -18564 394848 -18508
rect 394508 -18650 394848 -18564
rect 394508 -18706 394580 -18650
rect 394636 -18706 394722 -18650
rect 394778 -18706 394848 -18650
rect 394508 -18792 394848 -18706
rect 394508 -18848 394580 -18792
rect 394636 -18848 394722 -18792
rect 394778 -18848 394848 -18792
rect 394508 -18934 394848 -18848
rect 394508 -18990 394580 -18934
rect 394636 -18990 394722 -18934
rect 394778 -18990 394848 -18934
rect 394508 -19076 394848 -18990
rect 394508 -19132 394580 -19076
rect 394636 -19132 394722 -19076
rect 394778 -19132 394848 -19076
rect 394508 -19218 394848 -19132
rect 394508 -19274 394580 -19218
rect 394636 -19274 394722 -19218
rect 394778 -19274 394848 -19218
rect 394508 -19360 394848 -19274
rect 394508 -19416 394580 -19360
rect 394636 -19416 394722 -19360
rect 394778 -19416 394848 -19360
rect 394508 -19502 394848 -19416
rect 394508 -19558 394580 -19502
rect 394636 -19558 394722 -19502
rect 394778 -19558 394848 -19502
rect 394508 -19644 394848 -19558
rect 394508 -19700 394580 -19644
rect 394636 -19700 394722 -19644
rect 394778 -19700 394848 -19644
rect 394508 -19786 394848 -19700
rect 394508 -19842 394580 -19786
rect 394636 -19842 394722 -19786
rect 394778 -19842 394848 -19786
rect 394508 -19928 394848 -19842
rect 394508 -19984 394580 -19928
rect 394636 -19984 394722 -19928
rect 394778 -19984 394848 -19928
rect 394508 -20070 394848 -19984
rect 394508 -20126 394580 -20070
rect 394636 -20126 394722 -20070
rect 394778 -20126 394848 -20070
rect 394508 -20212 394848 -20126
rect 394508 -20268 394580 -20212
rect 394636 -20268 394722 -20212
rect 394778 -20268 394848 -20212
rect 394508 -20354 394848 -20268
rect 394508 -20410 394580 -20354
rect 394636 -20410 394722 -20354
rect 394778 -20410 394848 -20354
rect 394508 -20496 394848 -20410
rect 394508 -20552 394580 -20496
rect 394636 -20552 394722 -20496
rect 394778 -20552 394848 -20496
rect 394508 -20638 394848 -20552
rect 394508 -20694 394580 -20638
rect 394636 -20694 394722 -20638
rect 394778 -20694 394848 -20638
rect 394508 -20780 394848 -20694
rect 394508 -20836 394580 -20780
rect 394636 -20836 394722 -20780
rect 394778 -20836 394848 -20780
rect 394508 -20922 394848 -20836
rect 394508 -20978 394580 -20922
rect 394636 -20978 394722 -20922
rect 394778 -20978 394848 -20922
rect 394508 -21064 394848 -20978
rect 394508 -21120 394580 -21064
rect 394636 -21120 394722 -21064
rect 394778 -21120 394848 -21064
rect 394508 -21206 394848 -21120
rect 394508 -21262 394580 -21206
rect 394636 -21262 394722 -21206
rect 394778 -21262 394848 -21206
rect 394508 -21348 394848 -21262
rect 394508 -21404 394580 -21348
rect 394636 -21404 394722 -21348
rect 394778 -21404 394848 -21348
rect 394508 -21490 394848 -21404
rect 394508 -21546 394580 -21490
rect 394636 -21546 394722 -21490
rect 394778 -21546 394848 -21490
rect 394508 -21632 394848 -21546
rect 394508 -21688 394580 -21632
rect 394636 -21688 394722 -21632
rect 394778 -21688 394848 -21632
rect 394508 -21774 394848 -21688
rect 394508 -21830 394580 -21774
rect 394636 -21830 394722 -21774
rect 394778 -21830 394848 -21774
rect 394508 -21916 394848 -21830
rect 394508 -21972 394580 -21916
rect 394636 -21972 394722 -21916
rect 394778 -21972 394848 -21916
rect 394508 -22058 394848 -21972
rect 394508 -22114 394580 -22058
rect 394636 -22114 394722 -22058
rect 394778 -22114 394848 -22058
rect 394508 -22200 394848 -22114
rect 394508 -22256 394580 -22200
rect 394636 -22256 394722 -22200
rect 394778 -22256 394848 -22200
rect 394508 -22342 394848 -22256
rect 394508 -22398 394580 -22342
rect 394636 -22398 394722 -22342
rect 394778 -22398 394848 -22342
rect 394508 -22484 394848 -22398
rect 394508 -22540 394580 -22484
rect 394636 -22540 394722 -22484
rect 394778 -22540 394848 -22484
rect 394508 -22626 394848 -22540
rect 394508 -22682 394580 -22626
rect 394636 -22682 394722 -22626
rect 394778 -22682 394848 -22626
rect 394508 -22768 394848 -22682
rect 394508 -22824 394580 -22768
rect 394636 -22824 394722 -22768
rect 394778 -22824 394848 -22768
rect 394508 -22910 394848 -22824
rect 394508 -22966 394580 -22910
rect 394636 -22966 394722 -22910
rect 394778 -22966 394848 -22910
rect 394508 -23052 394848 -22966
rect 394508 -23108 394580 -23052
rect 394636 -23108 394722 -23052
rect 394778 -23108 394848 -23052
rect 394508 -23194 394848 -23108
rect 394508 -23250 394580 -23194
rect 394636 -23250 394722 -23194
rect 394778 -23250 394848 -23194
rect 394508 -23336 394848 -23250
rect 394508 -23392 394580 -23336
rect 394636 -23392 394722 -23336
rect 394778 -23392 394848 -23336
rect 394508 -23478 394848 -23392
rect 394508 -23534 394580 -23478
rect 394636 -23534 394722 -23478
rect 394778 -23534 394848 -23478
rect 394508 -23620 394848 -23534
rect 394508 -23676 394580 -23620
rect 394636 -23676 394722 -23620
rect 394778 -23676 394848 -23620
rect 394508 -23762 394848 -23676
rect 394508 -23818 394580 -23762
rect 394636 -23818 394722 -23762
rect 394778 -23818 394848 -23762
rect 394508 -23904 394848 -23818
rect 394508 -23960 394580 -23904
rect 394636 -23960 394722 -23904
rect 394778 -23960 394848 -23904
rect 394508 -24046 394848 -23960
rect 394508 -24102 394580 -24046
rect 394636 -24102 394722 -24046
rect 394778 -24102 394848 -24046
rect 394508 -24188 394848 -24102
rect 394508 -24244 394580 -24188
rect 394636 -24244 394722 -24188
rect 394778 -24244 394848 -24188
rect 394508 -24330 394848 -24244
rect 394508 -24386 394580 -24330
rect 394636 -24386 394722 -24330
rect 394778 -24386 394848 -24330
rect 394508 -24472 394848 -24386
rect 394508 -24528 394580 -24472
rect 394636 -24528 394722 -24472
rect 394778 -24528 394848 -24472
rect 394508 -24614 394848 -24528
rect 394508 -24670 394580 -24614
rect 394636 -24670 394722 -24614
rect 394778 -24670 394848 -24614
rect 394508 -24756 394848 -24670
rect 394508 -24812 394580 -24756
rect 394636 -24812 394722 -24756
rect 394778 -24812 394848 -24756
rect 394508 -24898 394848 -24812
rect 394508 -24954 394580 -24898
rect 394636 -24954 394722 -24898
rect 394778 -24954 394848 -24898
rect 394508 -25040 394848 -24954
rect 394508 -25096 394580 -25040
rect 394636 -25096 394722 -25040
rect 394778 -25096 394848 -25040
rect 394508 -25182 394848 -25096
rect 394508 -25238 394580 -25182
rect 394636 -25238 394722 -25182
rect 394778 -25238 394848 -25182
rect 394508 -25324 394848 -25238
rect 394508 -25380 394580 -25324
rect 394636 -25380 394722 -25324
rect 394778 -25380 394848 -25324
rect 394508 -25466 394848 -25380
rect 394508 -25522 394580 -25466
rect 394636 -25522 394722 -25466
rect 394778 -25522 394848 -25466
rect 394508 -25590 394848 -25522
rect 394908 -13680 395248 -13590
rect 394908 -13736 394982 -13680
rect 395038 -13736 395124 -13680
rect 395180 -13736 395248 -13680
rect 394908 -13822 395248 -13736
rect 394908 -13878 394982 -13822
rect 395038 -13878 395124 -13822
rect 395180 -13878 395248 -13822
rect 394908 -13964 395248 -13878
rect 394908 -14020 394982 -13964
rect 395038 -14020 395124 -13964
rect 395180 -14020 395248 -13964
rect 394908 -14106 395248 -14020
rect 394908 -14162 394982 -14106
rect 395038 -14162 395124 -14106
rect 395180 -14162 395248 -14106
rect 394908 -14248 395248 -14162
rect 394908 -14304 394982 -14248
rect 395038 -14304 395124 -14248
rect 395180 -14304 395248 -14248
rect 394908 -14390 395248 -14304
rect 394908 -14446 394982 -14390
rect 395038 -14446 395124 -14390
rect 395180 -14446 395248 -14390
rect 394908 -14532 395248 -14446
rect 394908 -14588 394982 -14532
rect 395038 -14588 395124 -14532
rect 395180 -14588 395248 -14532
rect 394908 -14674 395248 -14588
rect 394908 -14730 394982 -14674
rect 395038 -14730 395124 -14674
rect 395180 -14730 395248 -14674
rect 394908 -14816 395248 -14730
rect 394908 -14872 394982 -14816
rect 395038 -14872 395124 -14816
rect 395180 -14872 395248 -14816
rect 394908 -14958 395248 -14872
rect 394908 -15014 394982 -14958
rect 395038 -15014 395124 -14958
rect 395180 -15014 395248 -14958
rect 394908 -15100 395248 -15014
rect 394908 -15156 394982 -15100
rect 395038 -15156 395124 -15100
rect 395180 -15156 395248 -15100
rect 394908 -15242 395248 -15156
rect 394908 -15298 394982 -15242
rect 395038 -15298 395124 -15242
rect 395180 -15298 395248 -15242
rect 394908 -15384 395248 -15298
rect 394908 -15440 394982 -15384
rect 395038 -15440 395124 -15384
rect 395180 -15440 395248 -15384
rect 394908 -15526 395248 -15440
rect 394908 -15582 394982 -15526
rect 395038 -15582 395124 -15526
rect 395180 -15582 395248 -15526
rect 394908 -15668 395248 -15582
rect 394908 -15724 394982 -15668
rect 395038 -15724 395124 -15668
rect 395180 -15724 395248 -15668
rect 394908 -15810 395248 -15724
rect 394908 -15866 394982 -15810
rect 395038 -15866 395124 -15810
rect 395180 -15866 395248 -15810
rect 394908 -15952 395248 -15866
rect 394908 -16008 394982 -15952
rect 395038 -16008 395124 -15952
rect 395180 -16008 395248 -15952
rect 394908 -16094 395248 -16008
rect 394908 -16150 394982 -16094
rect 395038 -16150 395124 -16094
rect 395180 -16150 395248 -16094
rect 394908 -16236 395248 -16150
rect 394908 -16292 394982 -16236
rect 395038 -16292 395124 -16236
rect 395180 -16292 395248 -16236
rect 394908 -16378 395248 -16292
rect 394908 -16434 394982 -16378
rect 395038 -16434 395124 -16378
rect 395180 -16434 395248 -16378
rect 394908 -16520 395248 -16434
rect 394908 -16576 394982 -16520
rect 395038 -16576 395124 -16520
rect 395180 -16576 395248 -16520
rect 394908 -16662 395248 -16576
rect 394908 -16718 394982 -16662
rect 395038 -16718 395124 -16662
rect 395180 -16718 395248 -16662
rect 394908 -16804 395248 -16718
rect 394908 -16860 394982 -16804
rect 395038 -16860 395124 -16804
rect 395180 -16860 395248 -16804
rect 394908 -16946 395248 -16860
rect 394908 -17002 394982 -16946
rect 395038 -17002 395124 -16946
rect 395180 -17002 395248 -16946
rect 394908 -17088 395248 -17002
rect 394908 -17144 394982 -17088
rect 395038 -17144 395124 -17088
rect 395180 -17144 395248 -17088
rect 394908 -17230 395248 -17144
rect 394908 -17286 394982 -17230
rect 395038 -17286 395124 -17230
rect 395180 -17286 395248 -17230
rect 394908 -17372 395248 -17286
rect 394908 -17428 394982 -17372
rect 395038 -17428 395124 -17372
rect 395180 -17428 395248 -17372
rect 394908 -17514 395248 -17428
rect 394908 -17570 394982 -17514
rect 395038 -17570 395124 -17514
rect 395180 -17570 395248 -17514
rect 394908 -17656 395248 -17570
rect 394908 -17712 394982 -17656
rect 395038 -17712 395124 -17656
rect 395180 -17712 395248 -17656
rect 394908 -17798 395248 -17712
rect 394908 -17854 394982 -17798
rect 395038 -17854 395124 -17798
rect 395180 -17854 395248 -17798
rect 394908 -17940 395248 -17854
rect 394908 -17996 394982 -17940
rect 395038 -17996 395124 -17940
rect 395180 -17996 395248 -17940
rect 394908 -18082 395248 -17996
rect 394908 -18138 394982 -18082
rect 395038 -18138 395124 -18082
rect 395180 -18138 395248 -18082
rect 394908 -18224 395248 -18138
rect 394908 -18280 394982 -18224
rect 395038 -18280 395124 -18224
rect 395180 -18280 395248 -18224
rect 394908 -18366 395248 -18280
rect 394908 -18422 394982 -18366
rect 395038 -18422 395124 -18366
rect 395180 -18422 395248 -18366
rect 394908 -18508 395248 -18422
rect 394908 -18564 394982 -18508
rect 395038 -18564 395124 -18508
rect 395180 -18564 395248 -18508
rect 394908 -18650 395248 -18564
rect 394908 -18706 394982 -18650
rect 395038 -18706 395124 -18650
rect 395180 -18706 395248 -18650
rect 394908 -18792 395248 -18706
rect 394908 -18848 394982 -18792
rect 395038 -18848 395124 -18792
rect 395180 -18848 395248 -18792
rect 394908 -18934 395248 -18848
rect 394908 -18990 394982 -18934
rect 395038 -18990 395124 -18934
rect 395180 -18990 395248 -18934
rect 394908 -19076 395248 -18990
rect 394908 -19132 394982 -19076
rect 395038 -19132 395124 -19076
rect 395180 -19132 395248 -19076
rect 394908 -19218 395248 -19132
rect 394908 -19274 394982 -19218
rect 395038 -19274 395124 -19218
rect 395180 -19274 395248 -19218
rect 394908 -19360 395248 -19274
rect 394908 -19416 394982 -19360
rect 395038 -19416 395124 -19360
rect 395180 -19416 395248 -19360
rect 394908 -19502 395248 -19416
rect 394908 -19558 394982 -19502
rect 395038 -19558 395124 -19502
rect 395180 -19558 395248 -19502
rect 394908 -19644 395248 -19558
rect 394908 -19700 394982 -19644
rect 395038 -19700 395124 -19644
rect 395180 -19700 395248 -19644
rect 394908 -19786 395248 -19700
rect 394908 -19842 394982 -19786
rect 395038 -19842 395124 -19786
rect 395180 -19842 395248 -19786
rect 394908 -19928 395248 -19842
rect 394908 -19984 394982 -19928
rect 395038 -19984 395124 -19928
rect 395180 -19984 395248 -19928
rect 394908 -20070 395248 -19984
rect 394908 -20126 394982 -20070
rect 395038 -20126 395124 -20070
rect 395180 -20126 395248 -20070
rect 394908 -20212 395248 -20126
rect 394908 -20268 394982 -20212
rect 395038 -20268 395124 -20212
rect 395180 -20268 395248 -20212
rect 394908 -20354 395248 -20268
rect 394908 -20410 394982 -20354
rect 395038 -20410 395124 -20354
rect 395180 -20410 395248 -20354
rect 394908 -20496 395248 -20410
rect 394908 -20552 394982 -20496
rect 395038 -20552 395124 -20496
rect 395180 -20552 395248 -20496
rect 394908 -20638 395248 -20552
rect 394908 -20694 394982 -20638
rect 395038 -20694 395124 -20638
rect 395180 -20694 395248 -20638
rect 394908 -20780 395248 -20694
rect 394908 -20836 394982 -20780
rect 395038 -20836 395124 -20780
rect 395180 -20836 395248 -20780
rect 394908 -20922 395248 -20836
rect 394908 -20978 394982 -20922
rect 395038 -20978 395124 -20922
rect 395180 -20978 395248 -20922
rect 394908 -21064 395248 -20978
rect 394908 -21120 394982 -21064
rect 395038 -21120 395124 -21064
rect 395180 -21120 395248 -21064
rect 394908 -21206 395248 -21120
rect 394908 -21262 394982 -21206
rect 395038 -21262 395124 -21206
rect 395180 -21262 395248 -21206
rect 394908 -21348 395248 -21262
rect 394908 -21404 394982 -21348
rect 395038 -21404 395124 -21348
rect 395180 -21404 395248 -21348
rect 394908 -21490 395248 -21404
rect 394908 -21546 394982 -21490
rect 395038 -21546 395124 -21490
rect 395180 -21546 395248 -21490
rect 394908 -21632 395248 -21546
rect 394908 -21688 394982 -21632
rect 395038 -21688 395124 -21632
rect 395180 -21688 395248 -21632
rect 394908 -21774 395248 -21688
rect 394908 -21830 394982 -21774
rect 395038 -21830 395124 -21774
rect 395180 -21830 395248 -21774
rect 394908 -21916 395248 -21830
rect 394908 -21972 394982 -21916
rect 395038 -21972 395124 -21916
rect 395180 -21972 395248 -21916
rect 394908 -22058 395248 -21972
rect 394908 -22114 394982 -22058
rect 395038 -22114 395124 -22058
rect 395180 -22114 395248 -22058
rect 394908 -22200 395248 -22114
rect 394908 -22256 394982 -22200
rect 395038 -22256 395124 -22200
rect 395180 -22256 395248 -22200
rect 394908 -22342 395248 -22256
rect 394908 -22398 394982 -22342
rect 395038 -22398 395124 -22342
rect 395180 -22398 395248 -22342
rect 394908 -22484 395248 -22398
rect 394908 -22540 394982 -22484
rect 395038 -22540 395124 -22484
rect 395180 -22540 395248 -22484
rect 394908 -22626 395248 -22540
rect 394908 -22682 394982 -22626
rect 395038 -22682 395124 -22626
rect 395180 -22682 395248 -22626
rect 394908 -22768 395248 -22682
rect 394908 -22824 394982 -22768
rect 395038 -22824 395124 -22768
rect 395180 -22824 395248 -22768
rect 394908 -22910 395248 -22824
rect 394908 -22966 394982 -22910
rect 395038 -22966 395124 -22910
rect 395180 -22966 395248 -22910
rect 394908 -23052 395248 -22966
rect 394908 -23108 394982 -23052
rect 395038 -23108 395124 -23052
rect 395180 -23108 395248 -23052
rect 394908 -23194 395248 -23108
rect 394908 -23250 394982 -23194
rect 395038 -23250 395124 -23194
rect 395180 -23250 395248 -23194
rect 394908 -23336 395248 -23250
rect 394908 -23392 394982 -23336
rect 395038 -23392 395124 -23336
rect 395180 -23392 395248 -23336
rect 394908 -23478 395248 -23392
rect 394908 -23534 394982 -23478
rect 395038 -23534 395124 -23478
rect 395180 -23534 395248 -23478
rect 394908 -23620 395248 -23534
rect 394908 -23676 394982 -23620
rect 395038 -23676 395124 -23620
rect 395180 -23676 395248 -23620
rect 394908 -23762 395248 -23676
rect 394908 -23818 394982 -23762
rect 395038 -23818 395124 -23762
rect 395180 -23818 395248 -23762
rect 394908 -23904 395248 -23818
rect 394908 -23960 394982 -23904
rect 395038 -23960 395124 -23904
rect 395180 -23960 395248 -23904
rect 394908 -24046 395248 -23960
rect 394908 -24102 394982 -24046
rect 395038 -24102 395124 -24046
rect 395180 -24102 395248 -24046
rect 394908 -24188 395248 -24102
rect 394908 -24244 394982 -24188
rect 395038 -24244 395124 -24188
rect 395180 -24244 395248 -24188
rect 394908 -24330 395248 -24244
rect 394908 -24386 394982 -24330
rect 395038 -24386 395124 -24330
rect 395180 -24386 395248 -24330
rect 394908 -24472 395248 -24386
rect 394908 -24528 394982 -24472
rect 395038 -24528 395124 -24472
rect 395180 -24528 395248 -24472
rect 394908 -24614 395248 -24528
rect 394908 -24670 394982 -24614
rect 395038 -24670 395124 -24614
rect 395180 -24670 395248 -24614
rect 394908 -24756 395248 -24670
rect 394908 -24812 394982 -24756
rect 395038 -24812 395124 -24756
rect 395180 -24812 395248 -24756
rect 394908 -24898 395248 -24812
rect 394908 -24954 394982 -24898
rect 395038 -24954 395124 -24898
rect 395180 -24954 395248 -24898
rect 394908 -25040 395248 -24954
rect 394908 -25096 394982 -25040
rect 395038 -25096 395124 -25040
rect 395180 -25096 395248 -25040
rect 394908 -25182 395248 -25096
rect 394908 -25238 394982 -25182
rect 395038 -25238 395124 -25182
rect 395180 -25238 395248 -25182
rect 394908 -25324 395248 -25238
rect 394908 -25380 394982 -25324
rect 395038 -25380 395124 -25324
rect 395180 -25380 395248 -25324
rect 394908 -25466 395248 -25380
rect 394908 -25522 394982 -25466
rect 395038 -25522 395124 -25466
rect 395180 -25522 395248 -25466
rect 394908 -25590 395248 -25522
rect 395308 -13680 395648 -13590
rect 395308 -13736 395385 -13680
rect 395441 -13736 395527 -13680
rect 395583 -13736 395648 -13680
rect 395308 -13822 395648 -13736
rect 395308 -13878 395385 -13822
rect 395441 -13878 395527 -13822
rect 395583 -13878 395648 -13822
rect 395308 -13964 395648 -13878
rect 395308 -14020 395385 -13964
rect 395441 -14020 395527 -13964
rect 395583 -14020 395648 -13964
rect 395308 -14106 395648 -14020
rect 395308 -14162 395385 -14106
rect 395441 -14162 395527 -14106
rect 395583 -14162 395648 -14106
rect 395308 -14248 395648 -14162
rect 395308 -14304 395385 -14248
rect 395441 -14304 395527 -14248
rect 395583 -14304 395648 -14248
rect 395308 -14390 395648 -14304
rect 395308 -14446 395385 -14390
rect 395441 -14446 395527 -14390
rect 395583 -14446 395648 -14390
rect 395308 -14532 395648 -14446
rect 395308 -14588 395385 -14532
rect 395441 -14588 395527 -14532
rect 395583 -14588 395648 -14532
rect 395308 -14674 395648 -14588
rect 395308 -14730 395385 -14674
rect 395441 -14730 395527 -14674
rect 395583 -14730 395648 -14674
rect 395308 -14816 395648 -14730
rect 395308 -14872 395385 -14816
rect 395441 -14872 395527 -14816
rect 395583 -14872 395648 -14816
rect 395308 -14958 395648 -14872
rect 395308 -15014 395385 -14958
rect 395441 -15014 395527 -14958
rect 395583 -15014 395648 -14958
rect 395308 -15100 395648 -15014
rect 395308 -15156 395385 -15100
rect 395441 -15156 395527 -15100
rect 395583 -15156 395648 -15100
rect 395308 -15242 395648 -15156
rect 395308 -15298 395385 -15242
rect 395441 -15298 395527 -15242
rect 395583 -15298 395648 -15242
rect 395308 -15384 395648 -15298
rect 395308 -15440 395385 -15384
rect 395441 -15440 395527 -15384
rect 395583 -15440 395648 -15384
rect 395308 -15526 395648 -15440
rect 395308 -15582 395385 -15526
rect 395441 -15582 395527 -15526
rect 395583 -15582 395648 -15526
rect 395308 -15668 395648 -15582
rect 395308 -15724 395385 -15668
rect 395441 -15724 395527 -15668
rect 395583 -15724 395648 -15668
rect 395308 -15810 395648 -15724
rect 395308 -15866 395385 -15810
rect 395441 -15866 395527 -15810
rect 395583 -15866 395648 -15810
rect 395308 -15952 395648 -15866
rect 395308 -16008 395385 -15952
rect 395441 -16008 395527 -15952
rect 395583 -16008 395648 -15952
rect 395308 -16094 395648 -16008
rect 395308 -16150 395385 -16094
rect 395441 -16150 395527 -16094
rect 395583 -16150 395648 -16094
rect 395308 -16236 395648 -16150
rect 395308 -16292 395385 -16236
rect 395441 -16292 395527 -16236
rect 395583 -16292 395648 -16236
rect 395308 -16378 395648 -16292
rect 395308 -16434 395385 -16378
rect 395441 -16434 395527 -16378
rect 395583 -16434 395648 -16378
rect 395308 -16520 395648 -16434
rect 395308 -16576 395385 -16520
rect 395441 -16576 395527 -16520
rect 395583 -16576 395648 -16520
rect 395308 -16662 395648 -16576
rect 395308 -16718 395385 -16662
rect 395441 -16718 395527 -16662
rect 395583 -16718 395648 -16662
rect 395308 -16804 395648 -16718
rect 395308 -16860 395385 -16804
rect 395441 -16860 395527 -16804
rect 395583 -16860 395648 -16804
rect 395308 -16946 395648 -16860
rect 395308 -17002 395385 -16946
rect 395441 -17002 395527 -16946
rect 395583 -17002 395648 -16946
rect 395308 -17088 395648 -17002
rect 395308 -17144 395385 -17088
rect 395441 -17144 395527 -17088
rect 395583 -17144 395648 -17088
rect 395308 -17230 395648 -17144
rect 395308 -17286 395385 -17230
rect 395441 -17286 395527 -17230
rect 395583 -17286 395648 -17230
rect 395308 -17372 395648 -17286
rect 395308 -17428 395385 -17372
rect 395441 -17428 395527 -17372
rect 395583 -17428 395648 -17372
rect 395308 -17514 395648 -17428
rect 395308 -17570 395385 -17514
rect 395441 -17570 395527 -17514
rect 395583 -17570 395648 -17514
rect 395308 -17656 395648 -17570
rect 395308 -17712 395385 -17656
rect 395441 -17712 395527 -17656
rect 395583 -17712 395648 -17656
rect 395308 -17798 395648 -17712
rect 395308 -17854 395385 -17798
rect 395441 -17854 395527 -17798
rect 395583 -17854 395648 -17798
rect 395308 -17940 395648 -17854
rect 395308 -17996 395385 -17940
rect 395441 -17996 395527 -17940
rect 395583 -17996 395648 -17940
rect 395308 -18082 395648 -17996
rect 395308 -18138 395385 -18082
rect 395441 -18138 395527 -18082
rect 395583 -18138 395648 -18082
rect 395308 -18224 395648 -18138
rect 395308 -18280 395385 -18224
rect 395441 -18280 395527 -18224
rect 395583 -18280 395648 -18224
rect 395308 -18366 395648 -18280
rect 395308 -18422 395385 -18366
rect 395441 -18422 395527 -18366
rect 395583 -18422 395648 -18366
rect 395308 -18508 395648 -18422
rect 395308 -18564 395385 -18508
rect 395441 -18564 395527 -18508
rect 395583 -18564 395648 -18508
rect 395308 -18650 395648 -18564
rect 395308 -18706 395385 -18650
rect 395441 -18706 395527 -18650
rect 395583 -18706 395648 -18650
rect 395308 -18792 395648 -18706
rect 395308 -18848 395385 -18792
rect 395441 -18848 395527 -18792
rect 395583 -18848 395648 -18792
rect 395308 -18934 395648 -18848
rect 395308 -18990 395385 -18934
rect 395441 -18990 395527 -18934
rect 395583 -18990 395648 -18934
rect 395308 -19076 395648 -18990
rect 395308 -19132 395385 -19076
rect 395441 -19132 395527 -19076
rect 395583 -19132 395648 -19076
rect 395308 -19218 395648 -19132
rect 395308 -19274 395385 -19218
rect 395441 -19274 395527 -19218
rect 395583 -19274 395648 -19218
rect 395308 -19360 395648 -19274
rect 395308 -19416 395385 -19360
rect 395441 -19416 395527 -19360
rect 395583 -19416 395648 -19360
rect 395308 -19502 395648 -19416
rect 395308 -19558 395385 -19502
rect 395441 -19558 395527 -19502
rect 395583 -19558 395648 -19502
rect 395308 -19644 395648 -19558
rect 395308 -19700 395385 -19644
rect 395441 -19700 395527 -19644
rect 395583 -19700 395648 -19644
rect 395308 -19786 395648 -19700
rect 395308 -19842 395385 -19786
rect 395441 -19842 395527 -19786
rect 395583 -19842 395648 -19786
rect 395308 -19928 395648 -19842
rect 395308 -19984 395385 -19928
rect 395441 -19984 395527 -19928
rect 395583 -19984 395648 -19928
rect 395308 -20070 395648 -19984
rect 395308 -20126 395385 -20070
rect 395441 -20126 395527 -20070
rect 395583 -20126 395648 -20070
rect 395308 -20212 395648 -20126
rect 395308 -20268 395385 -20212
rect 395441 -20268 395527 -20212
rect 395583 -20268 395648 -20212
rect 395308 -20354 395648 -20268
rect 395308 -20410 395385 -20354
rect 395441 -20410 395527 -20354
rect 395583 -20410 395648 -20354
rect 395308 -20496 395648 -20410
rect 395308 -20552 395385 -20496
rect 395441 -20552 395527 -20496
rect 395583 -20552 395648 -20496
rect 395308 -20638 395648 -20552
rect 395308 -20694 395385 -20638
rect 395441 -20694 395527 -20638
rect 395583 -20694 395648 -20638
rect 395308 -20780 395648 -20694
rect 395308 -20836 395385 -20780
rect 395441 -20836 395527 -20780
rect 395583 -20836 395648 -20780
rect 395308 -20922 395648 -20836
rect 395308 -20978 395385 -20922
rect 395441 -20978 395527 -20922
rect 395583 -20978 395648 -20922
rect 395308 -21064 395648 -20978
rect 395308 -21120 395385 -21064
rect 395441 -21120 395527 -21064
rect 395583 -21120 395648 -21064
rect 395308 -21206 395648 -21120
rect 395308 -21262 395385 -21206
rect 395441 -21262 395527 -21206
rect 395583 -21262 395648 -21206
rect 395308 -21348 395648 -21262
rect 395308 -21404 395385 -21348
rect 395441 -21404 395527 -21348
rect 395583 -21404 395648 -21348
rect 395308 -21490 395648 -21404
rect 395308 -21546 395385 -21490
rect 395441 -21546 395527 -21490
rect 395583 -21546 395648 -21490
rect 395308 -21632 395648 -21546
rect 395308 -21688 395385 -21632
rect 395441 -21688 395527 -21632
rect 395583 -21688 395648 -21632
rect 395308 -21774 395648 -21688
rect 395308 -21830 395385 -21774
rect 395441 -21830 395527 -21774
rect 395583 -21830 395648 -21774
rect 395308 -21916 395648 -21830
rect 395308 -21972 395385 -21916
rect 395441 -21972 395527 -21916
rect 395583 -21972 395648 -21916
rect 395308 -22058 395648 -21972
rect 395308 -22114 395385 -22058
rect 395441 -22114 395527 -22058
rect 395583 -22114 395648 -22058
rect 395308 -22200 395648 -22114
rect 395308 -22256 395385 -22200
rect 395441 -22256 395527 -22200
rect 395583 -22256 395648 -22200
rect 395308 -22342 395648 -22256
rect 395308 -22398 395385 -22342
rect 395441 -22398 395527 -22342
rect 395583 -22398 395648 -22342
rect 395308 -22484 395648 -22398
rect 395308 -22540 395385 -22484
rect 395441 -22540 395527 -22484
rect 395583 -22540 395648 -22484
rect 395308 -22626 395648 -22540
rect 395308 -22682 395385 -22626
rect 395441 -22682 395527 -22626
rect 395583 -22682 395648 -22626
rect 395308 -22768 395648 -22682
rect 395308 -22824 395385 -22768
rect 395441 -22824 395527 -22768
rect 395583 -22824 395648 -22768
rect 395308 -22910 395648 -22824
rect 395308 -22966 395385 -22910
rect 395441 -22966 395527 -22910
rect 395583 -22966 395648 -22910
rect 395308 -23052 395648 -22966
rect 395308 -23108 395385 -23052
rect 395441 -23108 395527 -23052
rect 395583 -23108 395648 -23052
rect 395308 -23194 395648 -23108
rect 395308 -23250 395385 -23194
rect 395441 -23250 395527 -23194
rect 395583 -23250 395648 -23194
rect 395308 -23336 395648 -23250
rect 395308 -23392 395385 -23336
rect 395441 -23392 395527 -23336
rect 395583 -23392 395648 -23336
rect 395308 -23478 395648 -23392
rect 395308 -23534 395385 -23478
rect 395441 -23534 395527 -23478
rect 395583 -23534 395648 -23478
rect 395308 -23620 395648 -23534
rect 395308 -23676 395385 -23620
rect 395441 -23676 395527 -23620
rect 395583 -23676 395648 -23620
rect 395308 -23762 395648 -23676
rect 395308 -23818 395385 -23762
rect 395441 -23818 395527 -23762
rect 395583 -23818 395648 -23762
rect 395308 -23904 395648 -23818
rect 395308 -23960 395385 -23904
rect 395441 -23960 395527 -23904
rect 395583 -23960 395648 -23904
rect 395308 -24046 395648 -23960
rect 395308 -24102 395385 -24046
rect 395441 -24102 395527 -24046
rect 395583 -24102 395648 -24046
rect 395308 -24188 395648 -24102
rect 395308 -24244 395385 -24188
rect 395441 -24244 395527 -24188
rect 395583 -24244 395648 -24188
rect 395308 -24330 395648 -24244
rect 395308 -24386 395385 -24330
rect 395441 -24386 395527 -24330
rect 395583 -24386 395648 -24330
rect 395308 -24472 395648 -24386
rect 395308 -24528 395385 -24472
rect 395441 -24528 395527 -24472
rect 395583 -24528 395648 -24472
rect 395308 -24614 395648 -24528
rect 395308 -24670 395385 -24614
rect 395441 -24670 395527 -24614
rect 395583 -24670 395648 -24614
rect 395308 -24756 395648 -24670
rect 395308 -24812 395385 -24756
rect 395441 -24812 395527 -24756
rect 395583 -24812 395648 -24756
rect 395308 -24898 395648 -24812
rect 395308 -24954 395385 -24898
rect 395441 -24954 395527 -24898
rect 395583 -24954 395648 -24898
rect 395308 -25040 395648 -24954
rect 395308 -25096 395385 -25040
rect 395441 -25096 395527 -25040
rect 395583 -25096 395648 -25040
rect 395308 -25182 395648 -25096
rect 395308 -25238 395385 -25182
rect 395441 -25238 395527 -25182
rect 395583 -25238 395648 -25182
rect 395308 -25324 395648 -25238
rect 395308 -25380 395385 -25324
rect 395441 -25380 395527 -25324
rect 395583 -25380 395648 -25324
rect 395308 -25466 395648 -25380
rect 395308 -25522 395385 -25466
rect 395441 -25522 395527 -25466
rect 395583 -25522 395648 -25466
rect 395308 -25590 395648 -25522
rect 395708 -13680 396048 -13590
rect 395708 -13736 395779 -13680
rect 395835 -13736 395921 -13680
rect 395977 -13736 396048 -13680
rect 395708 -13822 396048 -13736
rect 395708 -13878 395779 -13822
rect 395835 -13878 395921 -13822
rect 395977 -13878 396048 -13822
rect 395708 -13964 396048 -13878
rect 395708 -14020 395779 -13964
rect 395835 -14020 395921 -13964
rect 395977 -14020 396048 -13964
rect 395708 -14106 396048 -14020
rect 395708 -14162 395779 -14106
rect 395835 -14162 395921 -14106
rect 395977 -14162 396048 -14106
rect 395708 -14248 396048 -14162
rect 395708 -14304 395779 -14248
rect 395835 -14304 395921 -14248
rect 395977 -14304 396048 -14248
rect 395708 -14390 396048 -14304
rect 395708 -14446 395779 -14390
rect 395835 -14446 395921 -14390
rect 395977 -14446 396048 -14390
rect 395708 -14532 396048 -14446
rect 395708 -14588 395779 -14532
rect 395835 -14588 395921 -14532
rect 395977 -14588 396048 -14532
rect 395708 -14674 396048 -14588
rect 395708 -14730 395779 -14674
rect 395835 -14730 395921 -14674
rect 395977 -14730 396048 -14674
rect 395708 -14816 396048 -14730
rect 395708 -14872 395779 -14816
rect 395835 -14872 395921 -14816
rect 395977 -14872 396048 -14816
rect 395708 -14958 396048 -14872
rect 395708 -15014 395779 -14958
rect 395835 -15014 395921 -14958
rect 395977 -15014 396048 -14958
rect 395708 -15100 396048 -15014
rect 395708 -15156 395779 -15100
rect 395835 -15156 395921 -15100
rect 395977 -15156 396048 -15100
rect 395708 -15242 396048 -15156
rect 395708 -15298 395779 -15242
rect 395835 -15298 395921 -15242
rect 395977 -15298 396048 -15242
rect 395708 -15384 396048 -15298
rect 395708 -15440 395779 -15384
rect 395835 -15440 395921 -15384
rect 395977 -15440 396048 -15384
rect 395708 -15526 396048 -15440
rect 395708 -15582 395779 -15526
rect 395835 -15582 395921 -15526
rect 395977 -15582 396048 -15526
rect 395708 -15668 396048 -15582
rect 395708 -15724 395779 -15668
rect 395835 -15724 395921 -15668
rect 395977 -15724 396048 -15668
rect 395708 -15810 396048 -15724
rect 395708 -15866 395779 -15810
rect 395835 -15866 395921 -15810
rect 395977 -15866 396048 -15810
rect 395708 -15952 396048 -15866
rect 395708 -16008 395779 -15952
rect 395835 -16008 395921 -15952
rect 395977 -16008 396048 -15952
rect 395708 -16094 396048 -16008
rect 395708 -16150 395779 -16094
rect 395835 -16150 395921 -16094
rect 395977 -16150 396048 -16094
rect 395708 -16236 396048 -16150
rect 395708 -16292 395779 -16236
rect 395835 -16292 395921 -16236
rect 395977 -16292 396048 -16236
rect 395708 -16378 396048 -16292
rect 395708 -16434 395779 -16378
rect 395835 -16434 395921 -16378
rect 395977 -16434 396048 -16378
rect 395708 -16520 396048 -16434
rect 395708 -16576 395779 -16520
rect 395835 -16576 395921 -16520
rect 395977 -16576 396048 -16520
rect 395708 -16662 396048 -16576
rect 395708 -16718 395779 -16662
rect 395835 -16718 395921 -16662
rect 395977 -16718 396048 -16662
rect 395708 -16804 396048 -16718
rect 395708 -16860 395779 -16804
rect 395835 -16860 395921 -16804
rect 395977 -16860 396048 -16804
rect 395708 -16946 396048 -16860
rect 395708 -17002 395779 -16946
rect 395835 -17002 395921 -16946
rect 395977 -17002 396048 -16946
rect 395708 -17088 396048 -17002
rect 395708 -17144 395779 -17088
rect 395835 -17144 395921 -17088
rect 395977 -17144 396048 -17088
rect 395708 -17230 396048 -17144
rect 395708 -17286 395779 -17230
rect 395835 -17286 395921 -17230
rect 395977 -17286 396048 -17230
rect 395708 -17372 396048 -17286
rect 395708 -17428 395779 -17372
rect 395835 -17428 395921 -17372
rect 395977 -17428 396048 -17372
rect 395708 -17514 396048 -17428
rect 395708 -17570 395779 -17514
rect 395835 -17570 395921 -17514
rect 395977 -17570 396048 -17514
rect 395708 -17656 396048 -17570
rect 395708 -17712 395779 -17656
rect 395835 -17712 395921 -17656
rect 395977 -17712 396048 -17656
rect 395708 -17798 396048 -17712
rect 395708 -17854 395779 -17798
rect 395835 -17854 395921 -17798
rect 395977 -17854 396048 -17798
rect 395708 -17940 396048 -17854
rect 395708 -17996 395779 -17940
rect 395835 -17996 395921 -17940
rect 395977 -17996 396048 -17940
rect 395708 -18082 396048 -17996
rect 395708 -18138 395779 -18082
rect 395835 -18138 395921 -18082
rect 395977 -18138 396048 -18082
rect 395708 -18224 396048 -18138
rect 395708 -18280 395779 -18224
rect 395835 -18280 395921 -18224
rect 395977 -18280 396048 -18224
rect 395708 -18366 396048 -18280
rect 395708 -18422 395779 -18366
rect 395835 -18422 395921 -18366
rect 395977 -18422 396048 -18366
rect 395708 -18508 396048 -18422
rect 395708 -18564 395779 -18508
rect 395835 -18564 395921 -18508
rect 395977 -18564 396048 -18508
rect 395708 -18650 396048 -18564
rect 395708 -18706 395779 -18650
rect 395835 -18706 395921 -18650
rect 395977 -18706 396048 -18650
rect 395708 -18792 396048 -18706
rect 395708 -18848 395779 -18792
rect 395835 -18848 395921 -18792
rect 395977 -18848 396048 -18792
rect 395708 -18934 396048 -18848
rect 395708 -18990 395779 -18934
rect 395835 -18990 395921 -18934
rect 395977 -18990 396048 -18934
rect 395708 -19076 396048 -18990
rect 395708 -19132 395779 -19076
rect 395835 -19132 395921 -19076
rect 395977 -19132 396048 -19076
rect 395708 -19218 396048 -19132
rect 395708 -19274 395779 -19218
rect 395835 -19274 395921 -19218
rect 395977 -19274 396048 -19218
rect 395708 -19360 396048 -19274
rect 395708 -19416 395779 -19360
rect 395835 -19416 395921 -19360
rect 395977 -19416 396048 -19360
rect 395708 -19502 396048 -19416
rect 395708 -19558 395779 -19502
rect 395835 -19558 395921 -19502
rect 395977 -19558 396048 -19502
rect 395708 -19644 396048 -19558
rect 395708 -19700 395779 -19644
rect 395835 -19700 395921 -19644
rect 395977 -19700 396048 -19644
rect 395708 -19786 396048 -19700
rect 395708 -19842 395779 -19786
rect 395835 -19842 395921 -19786
rect 395977 -19842 396048 -19786
rect 395708 -19928 396048 -19842
rect 395708 -19984 395779 -19928
rect 395835 -19984 395921 -19928
rect 395977 -19984 396048 -19928
rect 395708 -20070 396048 -19984
rect 395708 -20126 395779 -20070
rect 395835 -20126 395921 -20070
rect 395977 -20126 396048 -20070
rect 395708 -20212 396048 -20126
rect 395708 -20268 395779 -20212
rect 395835 -20268 395921 -20212
rect 395977 -20268 396048 -20212
rect 395708 -20354 396048 -20268
rect 395708 -20410 395779 -20354
rect 395835 -20410 395921 -20354
rect 395977 -20410 396048 -20354
rect 395708 -20496 396048 -20410
rect 395708 -20552 395779 -20496
rect 395835 -20552 395921 -20496
rect 395977 -20552 396048 -20496
rect 395708 -20638 396048 -20552
rect 395708 -20694 395779 -20638
rect 395835 -20694 395921 -20638
rect 395977 -20694 396048 -20638
rect 395708 -20780 396048 -20694
rect 395708 -20836 395779 -20780
rect 395835 -20836 395921 -20780
rect 395977 -20836 396048 -20780
rect 395708 -20922 396048 -20836
rect 395708 -20978 395779 -20922
rect 395835 -20978 395921 -20922
rect 395977 -20978 396048 -20922
rect 395708 -21064 396048 -20978
rect 395708 -21120 395779 -21064
rect 395835 -21120 395921 -21064
rect 395977 -21120 396048 -21064
rect 395708 -21206 396048 -21120
rect 395708 -21262 395779 -21206
rect 395835 -21262 395921 -21206
rect 395977 -21262 396048 -21206
rect 395708 -21348 396048 -21262
rect 395708 -21404 395779 -21348
rect 395835 -21404 395921 -21348
rect 395977 -21404 396048 -21348
rect 395708 -21490 396048 -21404
rect 395708 -21546 395779 -21490
rect 395835 -21546 395921 -21490
rect 395977 -21546 396048 -21490
rect 395708 -21632 396048 -21546
rect 395708 -21688 395779 -21632
rect 395835 -21688 395921 -21632
rect 395977 -21688 396048 -21632
rect 395708 -21774 396048 -21688
rect 395708 -21830 395779 -21774
rect 395835 -21830 395921 -21774
rect 395977 -21830 396048 -21774
rect 395708 -21916 396048 -21830
rect 395708 -21972 395779 -21916
rect 395835 -21972 395921 -21916
rect 395977 -21972 396048 -21916
rect 395708 -22058 396048 -21972
rect 395708 -22114 395779 -22058
rect 395835 -22114 395921 -22058
rect 395977 -22114 396048 -22058
rect 395708 -22200 396048 -22114
rect 395708 -22256 395779 -22200
rect 395835 -22256 395921 -22200
rect 395977 -22256 396048 -22200
rect 395708 -22342 396048 -22256
rect 395708 -22398 395779 -22342
rect 395835 -22398 395921 -22342
rect 395977 -22398 396048 -22342
rect 395708 -22484 396048 -22398
rect 395708 -22540 395779 -22484
rect 395835 -22540 395921 -22484
rect 395977 -22540 396048 -22484
rect 395708 -22626 396048 -22540
rect 395708 -22682 395779 -22626
rect 395835 -22682 395921 -22626
rect 395977 -22682 396048 -22626
rect 395708 -22768 396048 -22682
rect 395708 -22824 395779 -22768
rect 395835 -22824 395921 -22768
rect 395977 -22824 396048 -22768
rect 395708 -22910 396048 -22824
rect 395708 -22966 395779 -22910
rect 395835 -22966 395921 -22910
rect 395977 -22966 396048 -22910
rect 395708 -23052 396048 -22966
rect 395708 -23108 395779 -23052
rect 395835 -23108 395921 -23052
rect 395977 -23108 396048 -23052
rect 395708 -23194 396048 -23108
rect 395708 -23250 395779 -23194
rect 395835 -23250 395921 -23194
rect 395977 -23250 396048 -23194
rect 395708 -23336 396048 -23250
rect 395708 -23392 395779 -23336
rect 395835 -23392 395921 -23336
rect 395977 -23392 396048 -23336
rect 395708 -23478 396048 -23392
rect 395708 -23534 395779 -23478
rect 395835 -23534 395921 -23478
rect 395977 -23534 396048 -23478
rect 395708 -23620 396048 -23534
rect 395708 -23676 395779 -23620
rect 395835 -23676 395921 -23620
rect 395977 -23676 396048 -23620
rect 395708 -23762 396048 -23676
rect 395708 -23818 395779 -23762
rect 395835 -23818 395921 -23762
rect 395977 -23818 396048 -23762
rect 395708 -23904 396048 -23818
rect 395708 -23960 395779 -23904
rect 395835 -23960 395921 -23904
rect 395977 -23960 396048 -23904
rect 395708 -24046 396048 -23960
rect 395708 -24102 395779 -24046
rect 395835 -24102 395921 -24046
rect 395977 -24102 396048 -24046
rect 395708 -24188 396048 -24102
rect 395708 -24244 395779 -24188
rect 395835 -24244 395921 -24188
rect 395977 -24244 396048 -24188
rect 395708 -24330 396048 -24244
rect 395708 -24386 395779 -24330
rect 395835 -24386 395921 -24330
rect 395977 -24386 396048 -24330
rect 395708 -24472 396048 -24386
rect 395708 -24528 395779 -24472
rect 395835 -24528 395921 -24472
rect 395977 -24528 396048 -24472
rect 395708 -24614 396048 -24528
rect 395708 -24670 395779 -24614
rect 395835 -24670 395921 -24614
rect 395977 -24670 396048 -24614
rect 395708 -24756 396048 -24670
rect 395708 -24812 395779 -24756
rect 395835 -24812 395921 -24756
rect 395977 -24812 396048 -24756
rect 395708 -24898 396048 -24812
rect 395708 -24954 395779 -24898
rect 395835 -24954 395921 -24898
rect 395977 -24954 396048 -24898
rect 395708 -25040 396048 -24954
rect 395708 -25096 395779 -25040
rect 395835 -25096 395921 -25040
rect 395977 -25096 396048 -25040
rect 395708 -25182 396048 -25096
rect 395708 -25238 395779 -25182
rect 395835 -25238 395921 -25182
rect 395977 -25238 396048 -25182
rect 395708 -25324 396048 -25238
rect 395708 -25380 395779 -25324
rect 395835 -25380 395921 -25324
rect 395977 -25380 396048 -25324
rect 395708 -25466 396048 -25380
rect 395708 -25522 395779 -25466
rect 395835 -25522 395921 -25466
rect 395977 -25522 396048 -25466
rect 395708 -25590 396048 -25522
rect 396108 -13680 396448 -13590
rect 396108 -13736 396180 -13680
rect 396236 -13736 396322 -13680
rect 396378 -13736 396448 -13680
rect 396108 -13822 396448 -13736
rect 396108 -13878 396180 -13822
rect 396236 -13878 396322 -13822
rect 396378 -13878 396448 -13822
rect 396108 -13964 396448 -13878
rect 396108 -14020 396180 -13964
rect 396236 -14020 396322 -13964
rect 396378 -14020 396448 -13964
rect 396108 -14106 396448 -14020
rect 396108 -14162 396180 -14106
rect 396236 -14162 396322 -14106
rect 396378 -14162 396448 -14106
rect 396108 -14248 396448 -14162
rect 396108 -14304 396180 -14248
rect 396236 -14304 396322 -14248
rect 396378 -14304 396448 -14248
rect 396108 -14390 396448 -14304
rect 396108 -14446 396180 -14390
rect 396236 -14446 396322 -14390
rect 396378 -14446 396448 -14390
rect 396108 -14532 396448 -14446
rect 396108 -14588 396180 -14532
rect 396236 -14588 396322 -14532
rect 396378 -14588 396448 -14532
rect 396108 -14674 396448 -14588
rect 396108 -14730 396180 -14674
rect 396236 -14730 396322 -14674
rect 396378 -14730 396448 -14674
rect 396108 -14816 396448 -14730
rect 396108 -14872 396180 -14816
rect 396236 -14872 396322 -14816
rect 396378 -14872 396448 -14816
rect 396108 -14958 396448 -14872
rect 396108 -15014 396180 -14958
rect 396236 -15014 396322 -14958
rect 396378 -15014 396448 -14958
rect 396108 -15100 396448 -15014
rect 396108 -15156 396180 -15100
rect 396236 -15156 396322 -15100
rect 396378 -15156 396448 -15100
rect 396108 -15242 396448 -15156
rect 396108 -15298 396180 -15242
rect 396236 -15298 396322 -15242
rect 396378 -15298 396448 -15242
rect 396108 -15384 396448 -15298
rect 396108 -15440 396180 -15384
rect 396236 -15440 396322 -15384
rect 396378 -15440 396448 -15384
rect 396108 -15526 396448 -15440
rect 396108 -15582 396180 -15526
rect 396236 -15582 396322 -15526
rect 396378 -15582 396448 -15526
rect 396108 -15668 396448 -15582
rect 396108 -15724 396180 -15668
rect 396236 -15724 396322 -15668
rect 396378 -15724 396448 -15668
rect 396108 -15810 396448 -15724
rect 396108 -15866 396180 -15810
rect 396236 -15866 396322 -15810
rect 396378 -15866 396448 -15810
rect 396108 -15952 396448 -15866
rect 396108 -16008 396180 -15952
rect 396236 -16008 396322 -15952
rect 396378 -16008 396448 -15952
rect 396108 -16094 396448 -16008
rect 396108 -16150 396180 -16094
rect 396236 -16150 396322 -16094
rect 396378 -16150 396448 -16094
rect 396108 -16236 396448 -16150
rect 396108 -16292 396180 -16236
rect 396236 -16292 396322 -16236
rect 396378 -16292 396448 -16236
rect 396108 -16378 396448 -16292
rect 396108 -16434 396180 -16378
rect 396236 -16434 396322 -16378
rect 396378 -16434 396448 -16378
rect 396108 -16520 396448 -16434
rect 396108 -16576 396180 -16520
rect 396236 -16576 396322 -16520
rect 396378 -16576 396448 -16520
rect 396108 -16662 396448 -16576
rect 396108 -16718 396180 -16662
rect 396236 -16718 396322 -16662
rect 396378 -16718 396448 -16662
rect 396108 -16804 396448 -16718
rect 396108 -16860 396180 -16804
rect 396236 -16860 396322 -16804
rect 396378 -16860 396448 -16804
rect 396108 -16946 396448 -16860
rect 396108 -17002 396180 -16946
rect 396236 -17002 396322 -16946
rect 396378 -17002 396448 -16946
rect 396108 -17088 396448 -17002
rect 396108 -17144 396180 -17088
rect 396236 -17144 396322 -17088
rect 396378 -17144 396448 -17088
rect 396108 -17230 396448 -17144
rect 396108 -17286 396180 -17230
rect 396236 -17286 396322 -17230
rect 396378 -17286 396448 -17230
rect 396108 -17372 396448 -17286
rect 396108 -17428 396180 -17372
rect 396236 -17428 396322 -17372
rect 396378 -17428 396448 -17372
rect 396108 -17514 396448 -17428
rect 396108 -17570 396180 -17514
rect 396236 -17570 396322 -17514
rect 396378 -17570 396448 -17514
rect 396108 -17656 396448 -17570
rect 396108 -17712 396180 -17656
rect 396236 -17712 396322 -17656
rect 396378 -17712 396448 -17656
rect 396108 -17798 396448 -17712
rect 396108 -17854 396180 -17798
rect 396236 -17854 396322 -17798
rect 396378 -17854 396448 -17798
rect 396108 -17940 396448 -17854
rect 396108 -17996 396180 -17940
rect 396236 -17996 396322 -17940
rect 396378 -17996 396448 -17940
rect 396108 -18082 396448 -17996
rect 396108 -18138 396180 -18082
rect 396236 -18138 396322 -18082
rect 396378 -18138 396448 -18082
rect 396108 -18224 396448 -18138
rect 396108 -18280 396180 -18224
rect 396236 -18280 396322 -18224
rect 396378 -18280 396448 -18224
rect 396108 -18366 396448 -18280
rect 396108 -18422 396180 -18366
rect 396236 -18422 396322 -18366
rect 396378 -18422 396448 -18366
rect 396108 -18508 396448 -18422
rect 396108 -18564 396180 -18508
rect 396236 -18564 396322 -18508
rect 396378 -18564 396448 -18508
rect 396108 -18650 396448 -18564
rect 396108 -18706 396180 -18650
rect 396236 -18706 396322 -18650
rect 396378 -18706 396448 -18650
rect 396108 -18792 396448 -18706
rect 396108 -18848 396180 -18792
rect 396236 -18848 396322 -18792
rect 396378 -18848 396448 -18792
rect 396108 -18934 396448 -18848
rect 396108 -18990 396180 -18934
rect 396236 -18990 396322 -18934
rect 396378 -18990 396448 -18934
rect 396108 -19076 396448 -18990
rect 396108 -19132 396180 -19076
rect 396236 -19132 396322 -19076
rect 396378 -19132 396448 -19076
rect 396108 -19218 396448 -19132
rect 396108 -19274 396180 -19218
rect 396236 -19274 396322 -19218
rect 396378 -19274 396448 -19218
rect 396108 -19360 396448 -19274
rect 396108 -19416 396180 -19360
rect 396236 -19416 396322 -19360
rect 396378 -19416 396448 -19360
rect 396108 -19502 396448 -19416
rect 396108 -19558 396180 -19502
rect 396236 -19558 396322 -19502
rect 396378 -19558 396448 -19502
rect 396108 -19644 396448 -19558
rect 396108 -19700 396180 -19644
rect 396236 -19700 396322 -19644
rect 396378 -19700 396448 -19644
rect 396108 -19786 396448 -19700
rect 396108 -19842 396180 -19786
rect 396236 -19842 396322 -19786
rect 396378 -19842 396448 -19786
rect 396108 -19928 396448 -19842
rect 396108 -19984 396180 -19928
rect 396236 -19984 396322 -19928
rect 396378 -19984 396448 -19928
rect 396108 -20070 396448 -19984
rect 396108 -20126 396180 -20070
rect 396236 -20126 396322 -20070
rect 396378 -20126 396448 -20070
rect 396108 -20212 396448 -20126
rect 396108 -20268 396180 -20212
rect 396236 -20268 396322 -20212
rect 396378 -20268 396448 -20212
rect 396108 -20354 396448 -20268
rect 396108 -20410 396180 -20354
rect 396236 -20410 396322 -20354
rect 396378 -20410 396448 -20354
rect 396108 -20496 396448 -20410
rect 396108 -20552 396180 -20496
rect 396236 -20552 396322 -20496
rect 396378 -20552 396448 -20496
rect 396108 -20638 396448 -20552
rect 396108 -20694 396180 -20638
rect 396236 -20694 396322 -20638
rect 396378 -20694 396448 -20638
rect 396108 -20780 396448 -20694
rect 396108 -20836 396180 -20780
rect 396236 -20836 396322 -20780
rect 396378 -20836 396448 -20780
rect 396108 -20922 396448 -20836
rect 396108 -20978 396180 -20922
rect 396236 -20978 396322 -20922
rect 396378 -20978 396448 -20922
rect 396108 -21064 396448 -20978
rect 396108 -21120 396180 -21064
rect 396236 -21120 396322 -21064
rect 396378 -21120 396448 -21064
rect 396108 -21206 396448 -21120
rect 396108 -21262 396180 -21206
rect 396236 -21262 396322 -21206
rect 396378 -21262 396448 -21206
rect 396108 -21348 396448 -21262
rect 396108 -21404 396180 -21348
rect 396236 -21404 396322 -21348
rect 396378 -21404 396448 -21348
rect 396108 -21490 396448 -21404
rect 396108 -21546 396180 -21490
rect 396236 -21546 396322 -21490
rect 396378 -21546 396448 -21490
rect 396108 -21632 396448 -21546
rect 396108 -21688 396180 -21632
rect 396236 -21688 396322 -21632
rect 396378 -21688 396448 -21632
rect 396108 -21774 396448 -21688
rect 396108 -21830 396180 -21774
rect 396236 -21830 396322 -21774
rect 396378 -21830 396448 -21774
rect 396108 -21916 396448 -21830
rect 396108 -21972 396180 -21916
rect 396236 -21972 396322 -21916
rect 396378 -21972 396448 -21916
rect 396108 -22058 396448 -21972
rect 396108 -22114 396180 -22058
rect 396236 -22114 396322 -22058
rect 396378 -22114 396448 -22058
rect 396108 -22200 396448 -22114
rect 396108 -22256 396180 -22200
rect 396236 -22256 396322 -22200
rect 396378 -22256 396448 -22200
rect 396108 -22342 396448 -22256
rect 396108 -22398 396180 -22342
rect 396236 -22398 396322 -22342
rect 396378 -22398 396448 -22342
rect 396108 -22484 396448 -22398
rect 396108 -22540 396180 -22484
rect 396236 -22540 396322 -22484
rect 396378 -22540 396448 -22484
rect 396108 -22626 396448 -22540
rect 396108 -22682 396180 -22626
rect 396236 -22682 396322 -22626
rect 396378 -22682 396448 -22626
rect 396108 -22768 396448 -22682
rect 396108 -22824 396180 -22768
rect 396236 -22824 396322 -22768
rect 396378 -22824 396448 -22768
rect 396108 -22910 396448 -22824
rect 396108 -22966 396180 -22910
rect 396236 -22966 396322 -22910
rect 396378 -22966 396448 -22910
rect 396108 -23052 396448 -22966
rect 396108 -23108 396180 -23052
rect 396236 -23108 396322 -23052
rect 396378 -23108 396448 -23052
rect 396108 -23194 396448 -23108
rect 396108 -23250 396180 -23194
rect 396236 -23250 396322 -23194
rect 396378 -23250 396448 -23194
rect 396108 -23336 396448 -23250
rect 396108 -23392 396180 -23336
rect 396236 -23392 396322 -23336
rect 396378 -23392 396448 -23336
rect 396108 -23478 396448 -23392
rect 396108 -23534 396180 -23478
rect 396236 -23534 396322 -23478
rect 396378 -23534 396448 -23478
rect 396108 -23620 396448 -23534
rect 396108 -23676 396180 -23620
rect 396236 -23676 396322 -23620
rect 396378 -23676 396448 -23620
rect 396108 -23762 396448 -23676
rect 396108 -23818 396180 -23762
rect 396236 -23818 396322 -23762
rect 396378 -23818 396448 -23762
rect 396108 -23904 396448 -23818
rect 396108 -23960 396180 -23904
rect 396236 -23960 396322 -23904
rect 396378 -23960 396448 -23904
rect 396108 -24046 396448 -23960
rect 396108 -24102 396180 -24046
rect 396236 -24102 396322 -24046
rect 396378 -24102 396448 -24046
rect 396108 -24188 396448 -24102
rect 396108 -24244 396180 -24188
rect 396236 -24244 396322 -24188
rect 396378 -24244 396448 -24188
rect 396108 -24330 396448 -24244
rect 396108 -24386 396180 -24330
rect 396236 -24386 396322 -24330
rect 396378 -24386 396448 -24330
rect 396108 -24472 396448 -24386
rect 396108 -24528 396180 -24472
rect 396236 -24528 396322 -24472
rect 396378 -24528 396448 -24472
rect 396108 -24614 396448 -24528
rect 396108 -24670 396180 -24614
rect 396236 -24670 396322 -24614
rect 396378 -24670 396448 -24614
rect 396108 -24756 396448 -24670
rect 396108 -24812 396180 -24756
rect 396236 -24812 396322 -24756
rect 396378 -24812 396448 -24756
rect 396108 -24898 396448 -24812
rect 396108 -24954 396180 -24898
rect 396236 -24954 396322 -24898
rect 396378 -24954 396448 -24898
rect 396108 -25040 396448 -24954
rect 396108 -25096 396180 -25040
rect 396236 -25096 396322 -25040
rect 396378 -25096 396448 -25040
rect 396108 -25182 396448 -25096
rect 396108 -25238 396180 -25182
rect 396236 -25238 396322 -25182
rect 396378 -25238 396448 -25182
rect 396108 -25324 396448 -25238
rect 396108 -25380 396180 -25324
rect 396236 -25380 396322 -25324
rect 396378 -25380 396448 -25324
rect 396108 -25466 396448 -25380
rect 396108 -25522 396180 -25466
rect 396236 -25522 396322 -25466
rect 396378 -25522 396448 -25466
rect 396108 -25590 396448 -25522
rect 396508 -13680 396848 -13590
rect 396508 -13736 396580 -13680
rect 396636 -13736 396722 -13680
rect 396778 -13736 396848 -13680
rect 396508 -13822 396848 -13736
rect 396508 -13878 396580 -13822
rect 396636 -13878 396722 -13822
rect 396778 -13878 396848 -13822
rect 396508 -13964 396848 -13878
rect 396508 -14020 396580 -13964
rect 396636 -14020 396722 -13964
rect 396778 -14020 396848 -13964
rect 396508 -14106 396848 -14020
rect 396508 -14162 396580 -14106
rect 396636 -14162 396722 -14106
rect 396778 -14162 396848 -14106
rect 396508 -14248 396848 -14162
rect 396508 -14304 396580 -14248
rect 396636 -14304 396722 -14248
rect 396778 -14304 396848 -14248
rect 396508 -14390 396848 -14304
rect 396508 -14446 396580 -14390
rect 396636 -14446 396722 -14390
rect 396778 -14446 396848 -14390
rect 396508 -14532 396848 -14446
rect 396508 -14588 396580 -14532
rect 396636 -14588 396722 -14532
rect 396778 -14588 396848 -14532
rect 396508 -14674 396848 -14588
rect 396508 -14730 396580 -14674
rect 396636 -14730 396722 -14674
rect 396778 -14730 396848 -14674
rect 396508 -14816 396848 -14730
rect 396508 -14872 396580 -14816
rect 396636 -14872 396722 -14816
rect 396778 -14872 396848 -14816
rect 396508 -14958 396848 -14872
rect 396508 -15014 396580 -14958
rect 396636 -15014 396722 -14958
rect 396778 -15014 396848 -14958
rect 396508 -15100 396848 -15014
rect 396508 -15156 396580 -15100
rect 396636 -15156 396722 -15100
rect 396778 -15156 396848 -15100
rect 396508 -15242 396848 -15156
rect 396508 -15298 396580 -15242
rect 396636 -15298 396722 -15242
rect 396778 -15298 396848 -15242
rect 396508 -15384 396848 -15298
rect 396508 -15440 396580 -15384
rect 396636 -15440 396722 -15384
rect 396778 -15440 396848 -15384
rect 396508 -15526 396848 -15440
rect 396508 -15582 396580 -15526
rect 396636 -15582 396722 -15526
rect 396778 -15582 396848 -15526
rect 396508 -15668 396848 -15582
rect 396508 -15724 396580 -15668
rect 396636 -15724 396722 -15668
rect 396778 -15724 396848 -15668
rect 396508 -15810 396848 -15724
rect 396508 -15866 396580 -15810
rect 396636 -15866 396722 -15810
rect 396778 -15866 396848 -15810
rect 396508 -15952 396848 -15866
rect 396508 -16008 396580 -15952
rect 396636 -16008 396722 -15952
rect 396778 -16008 396848 -15952
rect 396508 -16094 396848 -16008
rect 396508 -16150 396580 -16094
rect 396636 -16150 396722 -16094
rect 396778 -16150 396848 -16094
rect 396508 -16236 396848 -16150
rect 396508 -16292 396580 -16236
rect 396636 -16292 396722 -16236
rect 396778 -16292 396848 -16236
rect 396508 -16378 396848 -16292
rect 396508 -16434 396580 -16378
rect 396636 -16434 396722 -16378
rect 396778 -16434 396848 -16378
rect 396508 -16520 396848 -16434
rect 396508 -16576 396580 -16520
rect 396636 -16576 396722 -16520
rect 396778 -16576 396848 -16520
rect 396508 -16662 396848 -16576
rect 396508 -16718 396580 -16662
rect 396636 -16718 396722 -16662
rect 396778 -16718 396848 -16662
rect 396508 -16804 396848 -16718
rect 396508 -16860 396580 -16804
rect 396636 -16860 396722 -16804
rect 396778 -16860 396848 -16804
rect 396508 -16946 396848 -16860
rect 396508 -17002 396580 -16946
rect 396636 -17002 396722 -16946
rect 396778 -17002 396848 -16946
rect 396508 -17088 396848 -17002
rect 396508 -17144 396580 -17088
rect 396636 -17144 396722 -17088
rect 396778 -17144 396848 -17088
rect 396508 -17230 396848 -17144
rect 396508 -17286 396580 -17230
rect 396636 -17286 396722 -17230
rect 396778 -17286 396848 -17230
rect 396508 -17372 396848 -17286
rect 396508 -17428 396580 -17372
rect 396636 -17428 396722 -17372
rect 396778 -17428 396848 -17372
rect 396508 -17514 396848 -17428
rect 396508 -17570 396580 -17514
rect 396636 -17570 396722 -17514
rect 396778 -17570 396848 -17514
rect 396508 -17656 396848 -17570
rect 396508 -17712 396580 -17656
rect 396636 -17712 396722 -17656
rect 396778 -17712 396848 -17656
rect 396508 -17798 396848 -17712
rect 396508 -17854 396580 -17798
rect 396636 -17854 396722 -17798
rect 396778 -17854 396848 -17798
rect 396508 -17940 396848 -17854
rect 396508 -17996 396580 -17940
rect 396636 -17996 396722 -17940
rect 396778 -17996 396848 -17940
rect 396508 -18082 396848 -17996
rect 396508 -18138 396580 -18082
rect 396636 -18138 396722 -18082
rect 396778 -18138 396848 -18082
rect 396508 -18224 396848 -18138
rect 396508 -18280 396580 -18224
rect 396636 -18280 396722 -18224
rect 396778 -18280 396848 -18224
rect 396508 -18366 396848 -18280
rect 396508 -18422 396580 -18366
rect 396636 -18422 396722 -18366
rect 396778 -18422 396848 -18366
rect 396508 -18508 396848 -18422
rect 396508 -18564 396580 -18508
rect 396636 -18564 396722 -18508
rect 396778 -18564 396848 -18508
rect 396508 -18650 396848 -18564
rect 396508 -18706 396580 -18650
rect 396636 -18706 396722 -18650
rect 396778 -18706 396848 -18650
rect 396508 -18792 396848 -18706
rect 396508 -18848 396580 -18792
rect 396636 -18848 396722 -18792
rect 396778 -18848 396848 -18792
rect 396508 -18934 396848 -18848
rect 396508 -18990 396580 -18934
rect 396636 -18990 396722 -18934
rect 396778 -18990 396848 -18934
rect 396508 -19076 396848 -18990
rect 396508 -19132 396580 -19076
rect 396636 -19132 396722 -19076
rect 396778 -19132 396848 -19076
rect 396508 -19218 396848 -19132
rect 396508 -19274 396580 -19218
rect 396636 -19274 396722 -19218
rect 396778 -19274 396848 -19218
rect 396508 -19360 396848 -19274
rect 396508 -19416 396580 -19360
rect 396636 -19416 396722 -19360
rect 396778 -19416 396848 -19360
rect 396508 -19502 396848 -19416
rect 396508 -19558 396580 -19502
rect 396636 -19558 396722 -19502
rect 396778 -19558 396848 -19502
rect 396508 -19644 396848 -19558
rect 396508 -19700 396580 -19644
rect 396636 -19700 396722 -19644
rect 396778 -19700 396848 -19644
rect 396508 -19786 396848 -19700
rect 396508 -19842 396580 -19786
rect 396636 -19842 396722 -19786
rect 396778 -19842 396848 -19786
rect 396508 -19928 396848 -19842
rect 396508 -19984 396580 -19928
rect 396636 -19984 396722 -19928
rect 396778 -19984 396848 -19928
rect 396508 -20070 396848 -19984
rect 396508 -20126 396580 -20070
rect 396636 -20126 396722 -20070
rect 396778 -20126 396848 -20070
rect 396508 -20212 396848 -20126
rect 396508 -20268 396580 -20212
rect 396636 -20268 396722 -20212
rect 396778 -20268 396848 -20212
rect 396508 -20354 396848 -20268
rect 396508 -20410 396580 -20354
rect 396636 -20410 396722 -20354
rect 396778 -20410 396848 -20354
rect 396508 -20496 396848 -20410
rect 396508 -20552 396580 -20496
rect 396636 -20552 396722 -20496
rect 396778 -20552 396848 -20496
rect 396508 -20638 396848 -20552
rect 396508 -20694 396580 -20638
rect 396636 -20694 396722 -20638
rect 396778 -20694 396848 -20638
rect 396508 -20780 396848 -20694
rect 396508 -20836 396580 -20780
rect 396636 -20836 396722 -20780
rect 396778 -20836 396848 -20780
rect 396508 -20922 396848 -20836
rect 396508 -20978 396580 -20922
rect 396636 -20978 396722 -20922
rect 396778 -20978 396848 -20922
rect 396508 -21064 396848 -20978
rect 396508 -21120 396580 -21064
rect 396636 -21120 396722 -21064
rect 396778 -21120 396848 -21064
rect 396508 -21206 396848 -21120
rect 396508 -21262 396580 -21206
rect 396636 -21262 396722 -21206
rect 396778 -21262 396848 -21206
rect 396508 -21348 396848 -21262
rect 396508 -21404 396580 -21348
rect 396636 -21404 396722 -21348
rect 396778 -21404 396848 -21348
rect 396508 -21490 396848 -21404
rect 396508 -21546 396580 -21490
rect 396636 -21546 396722 -21490
rect 396778 -21546 396848 -21490
rect 396508 -21632 396848 -21546
rect 396508 -21688 396580 -21632
rect 396636 -21688 396722 -21632
rect 396778 -21688 396848 -21632
rect 396508 -21774 396848 -21688
rect 396508 -21830 396580 -21774
rect 396636 -21830 396722 -21774
rect 396778 -21830 396848 -21774
rect 396508 -21916 396848 -21830
rect 396508 -21972 396580 -21916
rect 396636 -21972 396722 -21916
rect 396778 -21972 396848 -21916
rect 396508 -22058 396848 -21972
rect 396508 -22114 396580 -22058
rect 396636 -22114 396722 -22058
rect 396778 -22114 396848 -22058
rect 396508 -22200 396848 -22114
rect 396508 -22256 396580 -22200
rect 396636 -22256 396722 -22200
rect 396778 -22256 396848 -22200
rect 396508 -22342 396848 -22256
rect 396508 -22398 396580 -22342
rect 396636 -22398 396722 -22342
rect 396778 -22398 396848 -22342
rect 396508 -22484 396848 -22398
rect 396508 -22540 396580 -22484
rect 396636 -22540 396722 -22484
rect 396778 -22540 396848 -22484
rect 396508 -22626 396848 -22540
rect 396508 -22682 396580 -22626
rect 396636 -22682 396722 -22626
rect 396778 -22682 396848 -22626
rect 396508 -22768 396848 -22682
rect 396508 -22824 396580 -22768
rect 396636 -22824 396722 -22768
rect 396778 -22824 396848 -22768
rect 396508 -22910 396848 -22824
rect 396508 -22966 396580 -22910
rect 396636 -22966 396722 -22910
rect 396778 -22966 396848 -22910
rect 396508 -23052 396848 -22966
rect 396508 -23108 396580 -23052
rect 396636 -23108 396722 -23052
rect 396778 -23108 396848 -23052
rect 396508 -23194 396848 -23108
rect 396508 -23250 396580 -23194
rect 396636 -23250 396722 -23194
rect 396778 -23250 396848 -23194
rect 396508 -23336 396848 -23250
rect 396508 -23392 396580 -23336
rect 396636 -23392 396722 -23336
rect 396778 -23392 396848 -23336
rect 396508 -23478 396848 -23392
rect 396508 -23534 396580 -23478
rect 396636 -23534 396722 -23478
rect 396778 -23534 396848 -23478
rect 396508 -23620 396848 -23534
rect 396508 -23676 396580 -23620
rect 396636 -23676 396722 -23620
rect 396778 -23676 396848 -23620
rect 396508 -23762 396848 -23676
rect 396508 -23818 396580 -23762
rect 396636 -23818 396722 -23762
rect 396778 -23818 396848 -23762
rect 396508 -23904 396848 -23818
rect 396508 -23960 396580 -23904
rect 396636 -23960 396722 -23904
rect 396778 -23960 396848 -23904
rect 396508 -24046 396848 -23960
rect 396508 -24102 396580 -24046
rect 396636 -24102 396722 -24046
rect 396778 -24102 396848 -24046
rect 396508 -24188 396848 -24102
rect 396508 -24244 396580 -24188
rect 396636 -24244 396722 -24188
rect 396778 -24244 396848 -24188
rect 396508 -24330 396848 -24244
rect 396508 -24386 396580 -24330
rect 396636 -24386 396722 -24330
rect 396778 -24386 396848 -24330
rect 396508 -24472 396848 -24386
rect 396508 -24528 396580 -24472
rect 396636 -24528 396722 -24472
rect 396778 -24528 396848 -24472
rect 396508 -24614 396848 -24528
rect 396508 -24670 396580 -24614
rect 396636 -24670 396722 -24614
rect 396778 -24670 396848 -24614
rect 396508 -24756 396848 -24670
rect 396508 -24812 396580 -24756
rect 396636 -24812 396722 -24756
rect 396778 -24812 396848 -24756
rect 396508 -24898 396848 -24812
rect 396508 -24954 396580 -24898
rect 396636 -24954 396722 -24898
rect 396778 -24954 396848 -24898
rect 396508 -25040 396848 -24954
rect 396508 -25096 396580 -25040
rect 396636 -25096 396722 -25040
rect 396778 -25096 396848 -25040
rect 396508 -25182 396848 -25096
rect 396508 -25238 396580 -25182
rect 396636 -25238 396722 -25182
rect 396778 -25238 396848 -25182
rect 396508 -25324 396848 -25238
rect 396508 -25380 396580 -25324
rect 396636 -25380 396722 -25324
rect 396778 -25380 396848 -25324
rect 396508 -25466 396848 -25380
rect 396508 -25522 396580 -25466
rect 396636 -25522 396722 -25466
rect 396778 -25522 396848 -25466
rect 396508 -25590 396848 -25522
rect 396908 -13680 397248 -13590
rect 396908 -13736 396977 -13680
rect 397033 -13736 397119 -13680
rect 397175 -13736 397248 -13680
rect 396908 -13822 397248 -13736
rect 396908 -13878 396977 -13822
rect 397033 -13878 397119 -13822
rect 397175 -13878 397248 -13822
rect 396908 -13964 397248 -13878
rect 396908 -14020 396977 -13964
rect 397033 -14020 397119 -13964
rect 397175 -14020 397248 -13964
rect 396908 -14106 397248 -14020
rect 396908 -14162 396977 -14106
rect 397033 -14162 397119 -14106
rect 397175 -14162 397248 -14106
rect 396908 -14248 397248 -14162
rect 396908 -14304 396977 -14248
rect 397033 -14304 397119 -14248
rect 397175 -14304 397248 -14248
rect 396908 -14390 397248 -14304
rect 396908 -14446 396977 -14390
rect 397033 -14446 397119 -14390
rect 397175 -14446 397248 -14390
rect 396908 -14532 397248 -14446
rect 396908 -14588 396977 -14532
rect 397033 -14588 397119 -14532
rect 397175 -14588 397248 -14532
rect 396908 -14674 397248 -14588
rect 396908 -14730 396977 -14674
rect 397033 -14730 397119 -14674
rect 397175 -14730 397248 -14674
rect 396908 -14816 397248 -14730
rect 396908 -14872 396977 -14816
rect 397033 -14872 397119 -14816
rect 397175 -14872 397248 -14816
rect 396908 -14958 397248 -14872
rect 396908 -15014 396977 -14958
rect 397033 -15014 397119 -14958
rect 397175 -15014 397248 -14958
rect 396908 -15100 397248 -15014
rect 396908 -15156 396977 -15100
rect 397033 -15156 397119 -15100
rect 397175 -15156 397248 -15100
rect 396908 -15242 397248 -15156
rect 396908 -15298 396977 -15242
rect 397033 -15298 397119 -15242
rect 397175 -15298 397248 -15242
rect 396908 -15384 397248 -15298
rect 396908 -15440 396977 -15384
rect 397033 -15440 397119 -15384
rect 397175 -15440 397248 -15384
rect 396908 -15526 397248 -15440
rect 396908 -15582 396977 -15526
rect 397033 -15582 397119 -15526
rect 397175 -15582 397248 -15526
rect 396908 -15668 397248 -15582
rect 396908 -15724 396977 -15668
rect 397033 -15724 397119 -15668
rect 397175 -15724 397248 -15668
rect 396908 -15810 397248 -15724
rect 396908 -15866 396977 -15810
rect 397033 -15866 397119 -15810
rect 397175 -15866 397248 -15810
rect 396908 -15952 397248 -15866
rect 396908 -16008 396977 -15952
rect 397033 -16008 397119 -15952
rect 397175 -16008 397248 -15952
rect 396908 -16094 397248 -16008
rect 396908 -16150 396977 -16094
rect 397033 -16150 397119 -16094
rect 397175 -16150 397248 -16094
rect 396908 -16236 397248 -16150
rect 396908 -16292 396977 -16236
rect 397033 -16292 397119 -16236
rect 397175 -16292 397248 -16236
rect 396908 -16378 397248 -16292
rect 396908 -16434 396977 -16378
rect 397033 -16434 397119 -16378
rect 397175 -16434 397248 -16378
rect 396908 -16520 397248 -16434
rect 396908 -16576 396977 -16520
rect 397033 -16576 397119 -16520
rect 397175 -16576 397248 -16520
rect 396908 -16662 397248 -16576
rect 396908 -16718 396977 -16662
rect 397033 -16718 397119 -16662
rect 397175 -16718 397248 -16662
rect 396908 -16804 397248 -16718
rect 396908 -16860 396977 -16804
rect 397033 -16860 397119 -16804
rect 397175 -16860 397248 -16804
rect 396908 -16946 397248 -16860
rect 396908 -17002 396977 -16946
rect 397033 -17002 397119 -16946
rect 397175 -17002 397248 -16946
rect 396908 -17088 397248 -17002
rect 396908 -17144 396977 -17088
rect 397033 -17144 397119 -17088
rect 397175 -17144 397248 -17088
rect 396908 -17230 397248 -17144
rect 396908 -17286 396977 -17230
rect 397033 -17286 397119 -17230
rect 397175 -17286 397248 -17230
rect 396908 -17372 397248 -17286
rect 396908 -17428 396977 -17372
rect 397033 -17428 397119 -17372
rect 397175 -17428 397248 -17372
rect 396908 -17514 397248 -17428
rect 396908 -17570 396977 -17514
rect 397033 -17570 397119 -17514
rect 397175 -17570 397248 -17514
rect 396908 -17656 397248 -17570
rect 396908 -17712 396977 -17656
rect 397033 -17712 397119 -17656
rect 397175 -17712 397248 -17656
rect 396908 -17798 397248 -17712
rect 396908 -17854 396977 -17798
rect 397033 -17854 397119 -17798
rect 397175 -17854 397248 -17798
rect 396908 -17940 397248 -17854
rect 396908 -17996 396977 -17940
rect 397033 -17996 397119 -17940
rect 397175 -17996 397248 -17940
rect 396908 -18082 397248 -17996
rect 396908 -18138 396977 -18082
rect 397033 -18138 397119 -18082
rect 397175 -18138 397248 -18082
rect 396908 -18224 397248 -18138
rect 396908 -18280 396977 -18224
rect 397033 -18280 397119 -18224
rect 397175 -18280 397248 -18224
rect 396908 -18366 397248 -18280
rect 396908 -18422 396977 -18366
rect 397033 -18422 397119 -18366
rect 397175 -18422 397248 -18366
rect 396908 -18508 397248 -18422
rect 396908 -18564 396977 -18508
rect 397033 -18564 397119 -18508
rect 397175 -18564 397248 -18508
rect 396908 -18650 397248 -18564
rect 396908 -18706 396977 -18650
rect 397033 -18706 397119 -18650
rect 397175 -18706 397248 -18650
rect 396908 -18792 397248 -18706
rect 396908 -18848 396977 -18792
rect 397033 -18848 397119 -18792
rect 397175 -18848 397248 -18792
rect 396908 -18934 397248 -18848
rect 396908 -18990 396977 -18934
rect 397033 -18990 397119 -18934
rect 397175 -18990 397248 -18934
rect 396908 -19076 397248 -18990
rect 396908 -19132 396977 -19076
rect 397033 -19132 397119 -19076
rect 397175 -19132 397248 -19076
rect 396908 -19218 397248 -19132
rect 396908 -19274 396977 -19218
rect 397033 -19274 397119 -19218
rect 397175 -19274 397248 -19218
rect 396908 -19360 397248 -19274
rect 396908 -19416 396977 -19360
rect 397033 -19416 397119 -19360
rect 397175 -19416 397248 -19360
rect 396908 -19502 397248 -19416
rect 396908 -19558 396977 -19502
rect 397033 -19558 397119 -19502
rect 397175 -19558 397248 -19502
rect 396908 -19644 397248 -19558
rect 396908 -19700 396977 -19644
rect 397033 -19700 397119 -19644
rect 397175 -19700 397248 -19644
rect 396908 -19786 397248 -19700
rect 396908 -19842 396977 -19786
rect 397033 -19842 397119 -19786
rect 397175 -19842 397248 -19786
rect 396908 -19928 397248 -19842
rect 396908 -19984 396977 -19928
rect 397033 -19984 397119 -19928
rect 397175 -19984 397248 -19928
rect 396908 -20070 397248 -19984
rect 396908 -20126 396977 -20070
rect 397033 -20126 397119 -20070
rect 397175 -20126 397248 -20070
rect 396908 -20212 397248 -20126
rect 396908 -20268 396977 -20212
rect 397033 -20268 397119 -20212
rect 397175 -20268 397248 -20212
rect 396908 -20354 397248 -20268
rect 396908 -20410 396977 -20354
rect 397033 -20410 397119 -20354
rect 397175 -20410 397248 -20354
rect 396908 -20496 397248 -20410
rect 396908 -20552 396977 -20496
rect 397033 -20552 397119 -20496
rect 397175 -20552 397248 -20496
rect 396908 -20638 397248 -20552
rect 396908 -20694 396977 -20638
rect 397033 -20694 397119 -20638
rect 397175 -20694 397248 -20638
rect 396908 -20780 397248 -20694
rect 396908 -20836 396977 -20780
rect 397033 -20836 397119 -20780
rect 397175 -20836 397248 -20780
rect 396908 -20922 397248 -20836
rect 396908 -20978 396977 -20922
rect 397033 -20978 397119 -20922
rect 397175 -20978 397248 -20922
rect 396908 -21064 397248 -20978
rect 396908 -21120 396977 -21064
rect 397033 -21120 397119 -21064
rect 397175 -21120 397248 -21064
rect 396908 -21206 397248 -21120
rect 396908 -21262 396977 -21206
rect 397033 -21262 397119 -21206
rect 397175 -21262 397248 -21206
rect 396908 -21348 397248 -21262
rect 396908 -21404 396977 -21348
rect 397033 -21404 397119 -21348
rect 397175 -21404 397248 -21348
rect 396908 -21490 397248 -21404
rect 396908 -21546 396977 -21490
rect 397033 -21546 397119 -21490
rect 397175 -21546 397248 -21490
rect 396908 -21632 397248 -21546
rect 396908 -21688 396977 -21632
rect 397033 -21688 397119 -21632
rect 397175 -21688 397248 -21632
rect 396908 -21774 397248 -21688
rect 396908 -21830 396977 -21774
rect 397033 -21830 397119 -21774
rect 397175 -21830 397248 -21774
rect 396908 -21916 397248 -21830
rect 396908 -21972 396977 -21916
rect 397033 -21972 397119 -21916
rect 397175 -21972 397248 -21916
rect 396908 -22058 397248 -21972
rect 396908 -22114 396977 -22058
rect 397033 -22114 397119 -22058
rect 397175 -22114 397248 -22058
rect 396908 -22200 397248 -22114
rect 396908 -22256 396977 -22200
rect 397033 -22256 397119 -22200
rect 397175 -22256 397248 -22200
rect 396908 -22342 397248 -22256
rect 396908 -22398 396977 -22342
rect 397033 -22398 397119 -22342
rect 397175 -22398 397248 -22342
rect 396908 -22484 397248 -22398
rect 396908 -22540 396977 -22484
rect 397033 -22540 397119 -22484
rect 397175 -22540 397248 -22484
rect 396908 -22626 397248 -22540
rect 396908 -22682 396977 -22626
rect 397033 -22682 397119 -22626
rect 397175 -22682 397248 -22626
rect 396908 -22768 397248 -22682
rect 396908 -22824 396977 -22768
rect 397033 -22824 397119 -22768
rect 397175 -22824 397248 -22768
rect 396908 -22910 397248 -22824
rect 396908 -22966 396977 -22910
rect 397033 -22966 397119 -22910
rect 397175 -22966 397248 -22910
rect 396908 -23052 397248 -22966
rect 396908 -23108 396977 -23052
rect 397033 -23108 397119 -23052
rect 397175 -23108 397248 -23052
rect 396908 -23194 397248 -23108
rect 396908 -23250 396977 -23194
rect 397033 -23250 397119 -23194
rect 397175 -23250 397248 -23194
rect 396908 -23336 397248 -23250
rect 396908 -23392 396977 -23336
rect 397033 -23392 397119 -23336
rect 397175 -23392 397248 -23336
rect 396908 -23478 397248 -23392
rect 396908 -23534 396977 -23478
rect 397033 -23534 397119 -23478
rect 397175 -23534 397248 -23478
rect 396908 -23620 397248 -23534
rect 396908 -23676 396977 -23620
rect 397033 -23676 397119 -23620
rect 397175 -23676 397248 -23620
rect 396908 -23762 397248 -23676
rect 396908 -23818 396977 -23762
rect 397033 -23818 397119 -23762
rect 397175 -23818 397248 -23762
rect 396908 -23904 397248 -23818
rect 396908 -23960 396977 -23904
rect 397033 -23960 397119 -23904
rect 397175 -23960 397248 -23904
rect 396908 -24046 397248 -23960
rect 396908 -24102 396977 -24046
rect 397033 -24102 397119 -24046
rect 397175 -24102 397248 -24046
rect 396908 -24188 397248 -24102
rect 396908 -24244 396977 -24188
rect 397033 -24244 397119 -24188
rect 397175 -24244 397248 -24188
rect 396908 -24330 397248 -24244
rect 396908 -24386 396977 -24330
rect 397033 -24386 397119 -24330
rect 397175 -24386 397248 -24330
rect 396908 -24472 397248 -24386
rect 396908 -24528 396977 -24472
rect 397033 -24528 397119 -24472
rect 397175 -24528 397248 -24472
rect 396908 -24614 397248 -24528
rect 396908 -24670 396977 -24614
rect 397033 -24670 397119 -24614
rect 397175 -24670 397248 -24614
rect 396908 -24756 397248 -24670
rect 396908 -24812 396977 -24756
rect 397033 -24812 397119 -24756
rect 397175 -24812 397248 -24756
rect 396908 -24898 397248 -24812
rect 396908 -24954 396977 -24898
rect 397033 -24954 397119 -24898
rect 397175 -24954 397248 -24898
rect 396908 -25040 397248 -24954
rect 396908 -25096 396977 -25040
rect 397033 -25096 397119 -25040
rect 397175 -25096 397248 -25040
rect 396908 -25182 397248 -25096
rect 396908 -25238 396977 -25182
rect 397033 -25238 397119 -25182
rect 397175 -25238 397248 -25182
rect 396908 -25324 397248 -25238
rect 396908 -25380 396977 -25324
rect 397033 -25380 397119 -25324
rect 397175 -25380 397248 -25324
rect 396908 -25466 397248 -25380
rect 396908 -25522 396977 -25466
rect 397033 -25522 397119 -25466
rect 397175 -25522 397248 -25466
rect 396908 -25590 397248 -25522
rect 397308 -13680 397648 -13590
rect 397308 -13736 397374 -13680
rect 397430 -13736 397516 -13680
rect 397572 -13736 397648 -13680
rect 397308 -13822 397648 -13736
rect 397308 -13878 397374 -13822
rect 397430 -13878 397516 -13822
rect 397572 -13878 397648 -13822
rect 397308 -13964 397648 -13878
rect 397308 -14020 397374 -13964
rect 397430 -14020 397516 -13964
rect 397572 -14020 397648 -13964
rect 397308 -14106 397648 -14020
rect 397308 -14162 397374 -14106
rect 397430 -14162 397516 -14106
rect 397572 -14162 397648 -14106
rect 397308 -14248 397648 -14162
rect 397308 -14304 397374 -14248
rect 397430 -14304 397516 -14248
rect 397572 -14304 397648 -14248
rect 397308 -14390 397648 -14304
rect 397308 -14446 397374 -14390
rect 397430 -14446 397516 -14390
rect 397572 -14446 397648 -14390
rect 397308 -14532 397648 -14446
rect 397308 -14588 397374 -14532
rect 397430 -14588 397516 -14532
rect 397572 -14588 397648 -14532
rect 397308 -14674 397648 -14588
rect 397308 -14730 397374 -14674
rect 397430 -14730 397516 -14674
rect 397572 -14730 397648 -14674
rect 397308 -14816 397648 -14730
rect 397308 -14872 397374 -14816
rect 397430 -14872 397516 -14816
rect 397572 -14872 397648 -14816
rect 397308 -14958 397648 -14872
rect 397308 -15014 397374 -14958
rect 397430 -15014 397516 -14958
rect 397572 -15014 397648 -14958
rect 397308 -15100 397648 -15014
rect 397308 -15156 397374 -15100
rect 397430 -15156 397516 -15100
rect 397572 -15156 397648 -15100
rect 397308 -15242 397648 -15156
rect 397308 -15298 397374 -15242
rect 397430 -15298 397516 -15242
rect 397572 -15298 397648 -15242
rect 397308 -15384 397648 -15298
rect 397308 -15440 397374 -15384
rect 397430 -15440 397516 -15384
rect 397572 -15440 397648 -15384
rect 397308 -15526 397648 -15440
rect 397308 -15582 397374 -15526
rect 397430 -15582 397516 -15526
rect 397572 -15582 397648 -15526
rect 397308 -15668 397648 -15582
rect 397308 -15724 397374 -15668
rect 397430 -15724 397516 -15668
rect 397572 -15724 397648 -15668
rect 397308 -15810 397648 -15724
rect 397308 -15866 397374 -15810
rect 397430 -15866 397516 -15810
rect 397572 -15866 397648 -15810
rect 397308 -15952 397648 -15866
rect 397308 -16008 397374 -15952
rect 397430 -16008 397516 -15952
rect 397572 -16008 397648 -15952
rect 397308 -16094 397648 -16008
rect 397308 -16150 397374 -16094
rect 397430 -16150 397516 -16094
rect 397572 -16150 397648 -16094
rect 397308 -16236 397648 -16150
rect 397308 -16292 397374 -16236
rect 397430 -16292 397516 -16236
rect 397572 -16292 397648 -16236
rect 397308 -16378 397648 -16292
rect 397308 -16434 397374 -16378
rect 397430 -16434 397516 -16378
rect 397572 -16434 397648 -16378
rect 397308 -16520 397648 -16434
rect 397308 -16576 397374 -16520
rect 397430 -16576 397516 -16520
rect 397572 -16576 397648 -16520
rect 397308 -16662 397648 -16576
rect 397308 -16718 397374 -16662
rect 397430 -16718 397516 -16662
rect 397572 -16718 397648 -16662
rect 397308 -16804 397648 -16718
rect 397308 -16860 397374 -16804
rect 397430 -16860 397516 -16804
rect 397572 -16860 397648 -16804
rect 397308 -16946 397648 -16860
rect 397308 -17002 397374 -16946
rect 397430 -17002 397516 -16946
rect 397572 -17002 397648 -16946
rect 397308 -17088 397648 -17002
rect 397308 -17144 397374 -17088
rect 397430 -17144 397516 -17088
rect 397572 -17144 397648 -17088
rect 397308 -17230 397648 -17144
rect 397308 -17286 397374 -17230
rect 397430 -17286 397516 -17230
rect 397572 -17286 397648 -17230
rect 397308 -17372 397648 -17286
rect 397308 -17428 397374 -17372
rect 397430 -17428 397516 -17372
rect 397572 -17428 397648 -17372
rect 397308 -17514 397648 -17428
rect 397308 -17570 397374 -17514
rect 397430 -17570 397516 -17514
rect 397572 -17570 397648 -17514
rect 397308 -17656 397648 -17570
rect 397308 -17712 397374 -17656
rect 397430 -17712 397516 -17656
rect 397572 -17712 397648 -17656
rect 397308 -17798 397648 -17712
rect 397308 -17854 397374 -17798
rect 397430 -17854 397516 -17798
rect 397572 -17854 397648 -17798
rect 397308 -17940 397648 -17854
rect 397308 -17996 397374 -17940
rect 397430 -17996 397516 -17940
rect 397572 -17996 397648 -17940
rect 397308 -18082 397648 -17996
rect 397308 -18138 397374 -18082
rect 397430 -18138 397516 -18082
rect 397572 -18138 397648 -18082
rect 397308 -18224 397648 -18138
rect 397308 -18280 397374 -18224
rect 397430 -18280 397516 -18224
rect 397572 -18280 397648 -18224
rect 397308 -18366 397648 -18280
rect 397308 -18422 397374 -18366
rect 397430 -18422 397516 -18366
rect 397572 -18422 397648 -18366
rect 397308 -18508 397648 -18422
rect 397308 -18564 397374 -18508
rect 397430 -18564 397516 -18508
rect 397572 -18564 397648 -18508
rect 397308 -18650 397648 -18564
rect 397308 -18706 397374 -18650
rect 397430 -18706 397516 -18650
rect 397572 -18706 397648 -18650
rect 397308 -18792 397648 -18706
rect 397308 -18848 397374 -18792
rect 397430 -18848 397516 -18792
rect 397572 -18848 397648 -18792
rect 397308 -18934 397648 -18848
rect 397308 -18990 397374 -18934
rect 397430 -18990 397516 -18934
rect 397572 -18990 397648 -18934
rect 397308 -19076 397648 -18990
rect 397308 -19132 397374 -19076
rect 397430 -19132 397516 -19076
rect 397572 -19132 397648 -19076
rect 397308 -19218 397648 -19132
rect 397308 -19274 397374 -19218
rect 397430 -19274 397516 -19218
rect 397572 -19274 397648 -19218
rect 397308 -19360 397648 -19274
rect 397308 -19416 397374 -19360
rect 397430 -19416 397516 -19360
rect 397572 -19416 397648 -19360
rect 397308 -19502 397648 -19416
rect 397308 -19558 397374 -19502
rect 397430 -19558 397516 -19502
rect 397572 -19558 397648 -19502
rect 397308 -19644 397648 -19558
rect 397308 -19700 397374 -19644
rect 397430 -19700 397516 -19644
rect 397572 -19700 397648 -19644
rect 397308 -19786 397648 -19700
rect 397308 -19842 397374 -19786
rect 397430 -19842 397516 -19786
rect 397572 -19842 397648 -19786
rect 397308 -19928 397648 -19842
rect 397308 -19984 397374 -19928
rect 397430 -19984 397516 -19928
rect 397572 -19984 397648 -19928
rect 397308 -20070 397648 -19984
rect 397308 -20126 397374 -20070
rect 397430 -20126 397516 -20070
rect 397572 -20126 397648 -20070
rect 397308 -20212 397648 -20126
rect 397308 -20268 397374 -20212
rect 397430 -20268 397516 -20212
rect 397572 -20268 397648 -20212
rect 397308 -20354 397648 -20268
rect 397308 -20410 397374 -20354
rect 397430 -20410 397516 -20354
rect 397572 -20410 397648 -20354
rect 397308 -20496 397648 -20410
rect 397308 -20552 397374 -20496
rect 397430 -20552 397516 -20496
rect 397572 -20552 397648 -20496
rect 397308 -20638 397648 -20552
rect 397308 -20694 397374 -20638
rect 397430 -20694 397516 -20638
rect 397572 -20694 397648 -20638
rect 397308 -20780 397648 -20694
rect 397308 -20836 397374 -20780
rect 397430 -20836 397516 -20780
rect 397572 -20836 397648 -20780
rect 397308 -20922 397648 -20836
rect 397308 -20978 397374 -20922
rect 397430 -20978 397516 -20922
rect 397572 -20978 397648 -20922
rect 397308 -21064 397648 -20978
rect 397308 -21120 397374 -21064
rect 397430 -21120 397516 -21064
rect 397572 -21120 397648 -21064
rect 397308 -21206 397648 -21120
rect 397308 -21262 397374 -21206
rect 397430 -21262 397516 -21206
rect 397572 -21262 397648 -21206
rect 397308 -21348 397648 -21262
rect 397308 -21404 397374 -21348
rect 397430 -21404 397516 -21348
rect 397572 -21404 397648 -21348
rect 397308 -21490 397648 -21404
rect 397308 -21546 397374 -21490
rect 397430 -21546 397516 -21490
rect 397572 -21546 397648 -21490
rect 397308 -21632 397648 -21546
rect 397308 -21688 397374 -21632
rect 397430 -21688 397516 -21632
rect 397572 -21688 397648 -21632
rect 397308 -21774 397648 -21688
rect 397308 -21830 397374 -21774
rect 397430 -21830 397516 -21774
rect 397572 -21830 397648 -21774
rect 397308 -21916 397648 -21830
rect 397308 -21972 397374 -21916
rect 397430 -21972 397516 -21916
rect 397572 -21972 397648 -21916
rect 397308 -22058 397648 -21972
rect 397308 -22114 397374 -22058
rect 397430 -22114 397516 -22058
rect 397572 -22114 397648 -22058
rect 397308 -22200 397648 -22114
rect 397308 -22256 397374 -22200
rect 397430 -22256 397516 -22200
rect 397572 -22256 397648 -22200
rect 397308 -22342 397648 -22256
rect 397308 -22398 397374 -22342
rect 397430 -22398 397516 -22342
rect 397572 -22398 397648 -22342
rect 397308 -22484 397648 -22398
rect 397308 -22540 397374 -22484
rect 397430 -22540 397516 -22484
rect 397572 -22540 397648 -22484
rect 397308 -22626 397648 -22540
rect 397308 -22682 397374 -22626
rect 397430 -22682 397516 -22626
rect 397572 -22682 397648 -22626
rect 397308 -22768 397648 -22682
rect 397308 -22824 397374 -22768
rect 397430 -22824 397516 -22768
rect 397572 -22824 397648 -22768
rect 397308 -22910 397648 -22824
rect 397308 -22966 397374 -22910
rect 397430 -22966 397516 -22910
rect 397572 -22966 397648 -22910
rect 397308 -23052 397648 -22966
rect 397308 -23108 397374 -23052
rect 397430 -23108 397516 -23052
rect 397572 -23108 397648 -23052
rect 397308 -23194 397648 -23108
rect 397308 -23250 397374 -23194
rect 397430 -23250 397516 -23194
rect 397572 -23250 397648 -23194
rect 397308 -23336 397648 -23250
rect 397308 -23392 397374 -23336
rect 397430 -23392 397516 -23336
rect 397572 -23392 397648 -23336
rect 397308 -23478 397648 -23392
rect 397308 -23534 397374 -23478
rect 397430 -23534 397516 -23478
rect 397572 -23534 397648 -23478
rect 397308 -23620 397648 -23534
rect 397308 -23676 397374 -23620
rect 397430 -23676 397516 -23620
rect 397572 -23676 397648 -23620
rect 397308 -23762 397648 -23676
rect 397308 -23818 397374 -23762
rect 397430 -23818 397516 -23762
rect 397572 -23818 397648 -23762
rect 397308 -23904 397648 -23818
rect 397308 -23960 397374 -23904
rect 397430 -23960 397516 -23904
rect 397572 -23960 397648 -23904
rect 397308 -24046 397648 -23960
rect 397308 -24102 397374 -24046
rect 397430 -24102 397516 -24046
rect 397572 -24102 397648 -24046
rect 397308 -24188 397648 -24102
rect 397308 -24244 397374 -24188
rect 397430 -24244 397516 -24188
rect 397572 -24244 397648 -24188
rect 397308 -24330 397648 -24244
rect 397308 -24386 397374 -24330
rect 397430 -24386 397516 -24330
rect 397572 -24386 397648 -24330
rect 397308 -24472 397648 -24386
rect 397308 -24528 397374 -24472
rect 397430 -24528 397516 -24472
rect 397572 -24528 397648 -24472
rect 397308 -24614 397648 -24528
rect 397308 -24670 397374 -24614
rect 397430 -24670 397516 -24614
rect 397572 -24670 397648 -24614
rect 397308 -24756 397648 -24670
rect 397308 -24812 397374 -24756
rect 397430 -24812 397516 -24756
rect 397572 -24812 397648 -24756
rect 397308 -24898 397648 -24812
rect 397308 -24954 397374 -24898
rect 397430 -24954 397516 -24898
rect 397572 -24954 397648 -24898
rect 397308 -25040 397648 -24954
rect 397308 -25096 397374 -25040
rect 397430 -25096 397516 -25040
rect 397572 -25096 397648 -25040
rect 397308 -25182 397648 -25096
rect 397308 -25238 397374 -25182
rect 397430 -25238 397516 -25182
rect 397572 -25238 397648 -25182
rect 397308 -25324 397648 -25238
rect 397308 -25380 397374 -25324
rect 397430 -25380 397516 -25324
rect 397572 -25380 397648 -25324
rect 397308 -25466 397648 -25380
rect 397308 -25522 397374 -25466
rect 397430 -25522 397516 -25466
rect 397572 -25522 397648 -25466
rect 397308 -25590 397648 -25522
rect 397708 -13680 398048 -13590
rect 397708 -13736 397778 -13680
rect 397834 -13736 397920 -13680
rect 397976 -13736 398048 -13680
rect 397708 -13822 398048 -13736
rect 397708 -13878 397778 -13822
rect 397834 -13878 397920 -13822
rect 397976 -13878 398048 -13822
rect 397708 -13964 398048 -13878
rect 397708 -14020 397778 -13964
rect 397834 -14020 397920 -13964
rect 397976 -14020 398048 -13964
rect 397708 -14106 398048 -14020
rect 397708 -14162 397778 -14106
rect 397834 -14162 397920 -14106
rect 397976 -14162 398048 -14106
rect 397708 -14248 398048 -14162
rect 397708 -14304 397778 -14248
rect 397834 -14304 397920 -14248
rect 397976 -14304 398048 -14248
rect 397708 -14390 398048 -14304
rect 397708 -14446 397778 -14390
rect 397834 -14446 397920 -14390
rect 397976 -14446 398048 -14390
rect 397708 -14532 398048 -14446
rect 397708 -14588 397778 -14532
rect 397834 -14588 397920 -14532
rect 397976 -14588 398048 -14532
rect 397708 -14674 398048 -14588
rect 397708 -14730 397778 -14674
rect 397834 -14730 397920 -14674
rect 397976 -14730 398048 -14674
rect 397708 -14816 398048 -14730
rect 397708 -14872 397778 -14816
rect 397834 -14872 397920 -14816
rect 397976 -14872 398048 -14816
rect 397708 -14958 398048 -14872
rect 397708 -15014 397778 -14958
rect 397834 -15014 397920 -14958
rect 397976 -15014 398048 -14958
rect 397708 -15100 398048 -15014
rect 397708 -15156 397778 -15100
rect 397834 -15156 397920 -15100
rect 397976 -15156 398048 -15100
rect 397708 -15242 398048 -15156
rect 397708 -15298 397778 -15242
rect 397834 -15298 397920 -15242
rect 397976 -15298 398048 -15242
rect 397708 -15384 398048 -15298
rect 397708 -15440 397778 -15384
rect 397834 -15440 397920 -15384
rect 397976 -15440 398048 -15384
rect 397708 -15526 398048 -15440
rect 397708 -15582 397778 -15526
rect 397834 -15582 397920 -15526
rect 397976 -15582 398048 -15526
rect 397708 -15668 398048 -15582
rect 397708 -15724 397778 -15668
rect 397834 -15724 397920 -15668
rect 397976 -15724 398048 -15668
rect 397708 -15810 398048 -15724
rect 397708 -15866 397778 -15810
rect 397834 -15866 397920 -15810
rect 397976 -15866 398048 -15810
rect 397708 -15952 398048 -15866
rect 397708 -16008 397778 -15952
rect 397834 -16008 397920 -15952
rect 397976 -16008 398048 -15952
rect 397708 -16094 398048 -16008
rect 397708 -16150 397778 -16094
rect 397834 -16150 397920 -16094
rect 397976 -16150 398048 -16094
rect 397708 -16236 398048 -16150
rect 397708 -16292 397778 -16236
rect 397834 -16292 397920 -16236
rect 397976 -16292 398048 -16236
rect 397708 -16378 398048 -16292
rect 397708 -16434 397778 -16378
rect 397834 -16434 397920 -16378
rect 397976 -16434 398048 -16378
rect 397708 -16520 398048 -16434
rect 397708 -16576 397778 -16520
rect 397834 -16576 397920 -16520
rect 397976 -16576 398048 -16520
rect 397708 -16662 398048 -16576
rect 397708 -16718 397778 -16662
rect 397834 -16718 397920 -16662
rect 397976 -16718 398048 -16662
rect 397708 -16804 398048 -16718
rect 397708 -16860 397778 -16804
rect 397834 -16860 397920 -16804
rect 397976 -16860 398048 -16804
rect 397708 -16946 398048 -16860
rect 397708 -17002 397778 -16946
rect 397834 -17002 397920 -16946
rect 397976 -17002 398048 -16946
rect 397708 -17088 398048 -17002
rect 397708 -17144 397778 -17088
rect 397834 -17144 397920 -17088
rect 397976 -17144 398048 -17088
rect 397708 -17230 398048 -17144
rect 397708 -17286 397778 -17230
rect 397834 -17286 397920 -17230
rect 397976 -17286 398048 -17230
rect 397708 -17372 398048 -17286
rect 397708 -17428 397778 -17372
rect 397834 -17428 397920 -17372
rect 397976 -17428 398048 -17372
rect 397708 -17514 398048 -17428
rect 397708 -17570 397778 -17514
rect 397834 -17570 397920 -17514
rect 397976 -17570 398048 -17514
rect 397708 -17656 398048 -17570
rect 397708 -17712 397778 -17656
rect 397834 -17712 397920 -17656
rect 397976 -17712 398048 -17656
rect 397708 -17798 398048 -17712
rect 397708 -17854 397778 -17798
rect 397834 -17854 397920 -17798
rect 397976 -17854 398048 -17798
rect 397708 -17940 398048 -17854
rect 397708 -17996 397778 -17940
rect 397834 -17996 397920 -17940
rect 397976 -17996 398048 -17940
rect 397708 -18082 398048 -17996
rect 397708 -18138 397778 -18082
rect 397834 -18138 397920 -18082
rect 397976 -18138 398048 -18082
rect 397708 -18224 398048 -18138
rect 397708 -18280 397778 -18224
rect 397834 -18280 397920 -18224
rect 397976 -18280 398048 -18224
rect 397708 -18366 398048 -18280
rect 397708 -18422 397778 -18366
rect 397834 -18422 397920 -18366
rect 397976 -18422 398048 -18366
rect 397708 -18508 398048 -18422
rect 397708 -18564 397778 -18508
rect 397834 -18564 397920 -18508
rect 397976 -18564 398048 -18508
rect 397708 -18650 398048 -18564
rect 397708 -18706 397778 -18650
rect 397834 -18706 397920 -18650
rect 397976 -18706 398048 -18650
rect 397708 -18792 398048 -18706
rect 397708 -18848 397778 -18792
rect 397834 -18848 397920 -18792
rect 397976 -18848 398048 -18792
rect 397708 -18934 398048 -18848
rect 397708 -18990 397778 -18934
rect 397834 -18990 397920 -18934
rect 397976 -18990 398048 -18934
rect 397708 -19076 398048 -18990
rect 397708 -19132 397778 -19076
rect 397834 -19132 397920 -19076
rect 397976 -19132 398048 -19076
rect 397708 -19218 398048 -19132
rect 397708 -19274 397778 -19218
rect 397834 -19274 397920 -19218
rect 397976 -19274 398048 -19218
rect 397708 -19360 398048 -19274
rect 397708 -19416 397778 -19360
rect 397834 -19416 397920 -19360
rect 397976 -19416 398048 -19360
rect 397708 -19502 398048 -19416
rect 397708 -19558 397778 -19502
rect 397834 -19558 397920 -19502
rect 397976 -19558 398048 -19502
rect 397708 -19644 398048 -19558
rect 397708 -19700 397778 -19644
rect 397834 -19700 397920 -19644
rect 397976 -19700 398048 -19644
rect 397708 -19786 398048 -19700
rect 397708 -19842 397778 -19786
rect 397834 -19842 397920 -19786
rect 397976 -19842 398048 -19786
rect 397708 -19928 398048 -19842
rect 397708 -19984 397778 -19928
rect 397834 -19984 397920 -19928
rect 397976 -19984 398048 -19928
rect 397708 -20070 398048 -19984
rect 397708 -20126 397778 -20070
rect 397834 -20126 397920 -20070
rect 397976 -20126 398048 -20070
rect 397708 -20212 398048 -20126
rect 397708 -20268 397778 -20212
rect 397834 -20268 397920 -20212
rect 397976 -20268 398048 -20212
rect 397708 -20354 398048 -20268
rect 397708 -20410 397778 -20354
rect 397834 -20410 397920 -20354
rect 397976 -20410 398048 -20354
rect 397708 -20496 398048 -20410
rect 397708 -20552 397778 -20496
rect 397834 -20552 397920 -20496
rect 397976 -20552 398048 -20496
rect 397708 -20638 398048 -20552
rect 397708 -20694 397778 -20638
rect 397834 -20694 397920 -20638
rect 397976 -20694 398048 -20638
rect 397708 -20780 398048 -20694
rect 397708 -20836 397778 -20780
rect 397834 -20836 397920 -20780
rect 397976 -20836 398048 -20780
rect 397708 -20922 398048 -20836
rect 397708 -20978 397778 -20922
rect 397834 -20978 397920 -20922
rect 397976 -20978 398048 -20922
rect 397708 -21064 398048 -20978
rect 397708 -21120 397778 -21064
rect 397834 -21120 397920 -21064
rect 397976 -21120 398048 -21064
rect 397708 -21206 398048 -21120
rect 397708 -21262 397778 -21206
rect 397834 -21262 397920 -21206
rect 397976 -21262 398048 -21206
rect 397708 -21348 398048 -21262
rect 397708 -21404 397778 -21348
rect 397834 -21404 397920 -21348
rect 397976 -21404 398048 -21348
rect 397708 -21490 398048 -21404
rect 397708 -21546 397778 -21490
rect 397834 -21546 397920 -21490
rect 397976 -21546 398048 -21490
rect 397708 -21632 398048 -21546
rect 397708 -21688 397778 -21632
rect 397834 -21688 397920 -21632
rect 397976 -21688 398048 -21632
rect 397708 -21774 398048 -21688
rect 397708 -21830 397778 -21774
rect 397834 -21830 397920 -21774
rect 397976 -21830 398048 -21774
rect 397708 -21916 398048 -21830
rect 397708 -21972 397778 -21916
rect 397834 -21972 397920 -21916
rect 397976 -21972 398048 -21916
rect 397708 -22058 398048 -21972
rect 397708 -22114 397778 -22058
rect 397834 -22114 397920 -22058
rect 397976 -22114 398048 -22058
rect 397708 -22200 398048 -22114
rect 397708 -22256 397778 -22200
rect 397834 -22256 397920 -22200
rect 397976 -22256 398048 -22200
rect 397708 -22342 398048 -22256
rect 397708 -22398 397778 -22342
rect 397834 -22398 397920 -22342
rect 397976 -22398 398048 -22342
rect 397708 -22484 398048 -22398
rect 397708 -22540 397778 -22484
rect 397834 -22540 397920 -22484
rect 397976 -22540 398048 -22484
rect 397708 -22626 398048 -22540
rect 397708 -22682 397778 -22626
rect 397834 -22682 397920 -22626
rect 397976 -22682 398048 -22626
rect 397708 -22768 398048 -22682
rect 397708 -22824 397778 -22768
rect 397834 -22824 397920 -22768
rect 397976 -22824 398048 -22768
rect 397708 -22910 398048 -22824
rect 397708 -22966 397778 -22910
rect 397834 -22966 397920 -22910
rect 397976 -22966 398048 -22910
rect 397708 -23052 398048 -22966
rect 397708 -23108 397778 -23052
rect 397834 -23108 397920 -23052
rect 397976 -23108 398048 -23052
rect 397708 -23194 398048 -23108
rect 397708 -23250 397778 -23194
rect 397834 -23250 397920 -23194
rect 397976 -23250 398048 -23194
rect 397708 -23336 398048 -23250
rect 397708 -23392 397778 -23336
rect 397834 -23392 397920 -23336
rect 397976 -23392 398048 -23336
rect 397708 -23478 398048 -23392
rect 397708 -23534 397778 -23478
rect 397834 -23534 397920 -23478
rect 397976 -23534 398048 -23478
rect 397708 -23620 398048 -23534
rect 397708 -23676 397778 -23620
rect 397834 -23676 397920 -23620
rect 397976 -23676 398048 -23620
rect 397708 -23762 398048 -23676
rect 397708 -23818 397778 -23762
rect 397834 -23818 397920 -23762
rect 397976 -23818 398048 -23762
rect 397708 -23904 398048 -23818
rect 397708 -23960 397778 -23904
rect 397834 -23960 397920 -23904
rect 397976 -23960 398048 -23904
rect 397708 -24046 398048 -23960
rect 397708 -24102 397778 -24046
rect 397834 -24102 397920 -24046
rect 397976 -24102 398048 -24046
rect 397708 -24188 398048 -24102
rect 397708 -24244 397778 -24188
rect 397834 -24244 397920 -24188
rect 397976 -24244 398048 -24188
rect 397708 -24330 398048 -24244
rect 397708 -24386 397778 -24330
rect 397834 -24386 397920 -24330
rect 397976 -24386 398048 -24330
rect 397708 -24472 398048 -24386
rect 397708 -24528 397778 -24472
rect 397834 -24528 397920 -24472
rect 397976 -24528 398048 -24472
rect 397708 -24614 398048 -24528
rect 397708 -24670 397778 -24614
rect 397834 -24670 397920 -24614
rect 397976 -24670 398048 -24614
rect 397708 -24756 398048 -24670
rect 397708 -24812 397778 -24756
rect 397834 -24812 397920 -24756
rect 397976 -24812 398048 -24756
rect 397708 -24898 398048 -24812
rect 397708 -24954 397778 -24898
rect 397834 -24954 397920 -24898
rect 397976 -24954 398048 -24898
rect 397708 -25040 398048 -24954
rect 397708 -25096 397778 -25040
rect 397834 -25096 397920 -25040
rect 397976 -25096 398048 -25040
rect 397708 -25182 398048 -25096
rect 397708 -25238 397778 -25182
rect 397834 -25238 397920 -25182
rect 397976 -25238 398048 -25182
rect 397708 -25324 398048 -25238
rect 397708 -25380 397778 -25324
rect 397834 -25380 397920 -25324
rect 397976 -25380 398048 -25324
rect 397708 -25466 398048 -25380
rect 397708 -25522 397778 -25466
rect 397834 -25522 397920 -25466
rect 397976 -25522 398048 -25466
rect 397708 -25590 398048 -25522
rect 398108 -13680 398448 -13590
rect 398108 -13736 398174 -13680
rect 398230 -13736 398316 -13680
rect 398372 -13736 398448 -13680
rect 398108 -13822 398448 -13736
rect 398108 -13878 398174 -13822
rect 398230 -13878 398316 -13822
rect 398372 -13878 398448 -13822
rect 398108 -13964 398448 -13878
rect 398108 -14020 398174 -13964
rect 398230 -14020 398316 -13964
rect 398372 -14020 398448 -13964
rect 398108 -14106 398448 -14020
rect 398108 -14162 398174 -14106
rect 398230 -14162 398316 -14106
rect 398372 -14162 398448 -14106
rect 398108 -14248 398448 -14162
rect 398108 -14304 398174 -14248
rect 398230 -14304 398316 -14248
rect 398372 -14304 398448 -14248
rect 398108 -14390 398448 -14304
rect 398108 -14446 398174 -14390
rect 398230 -14446 398316 -14390
rect 398372 -14446 398448 -14390
rect 398108 -14532 398448 -14446
rect 398108 -14588 398174 -14532
rect 398230 -14588 398316 -14532
rect 398372 -14588 398448 -14532
rect 398108 -14674 398448 -14588
rect 398108 -14730 398174 -14674
rect 398230 -14730 398316 -14674
rect 398372 -14730 398448 -14674
rect 398108 -14816 398448 -14730
rect 398108 -14872 398174 -14816
rect 398230 -14872 398316 -14816
rect 398372 -14872 398448 -14816
rect 398108 -14958 398448 -14872
rect 398108 -15014 398174 -14958
rect 398230 -15014 398316 -14958
rect 398372 -15014 398448 -14958
rect 398108 -15100 398448 -15014
rect 398108 -15156 398174 -15100
rect 398230 -15156 398316 -15100
rect 398372 -15156 398448 -15100
rect 398108 -15242 398448 -15156
rect 398108 -15298 398174 -15242
rect 398230 -15298 398316 -15242
rect 398372 -15298 398448 -15242
rect 398108 -15384 398448 -15298
rect 398108 -15440 398174 -15384
rect 398230 -15440 398316 -15384
rect 398372 -15440 398448 -15384
rect 398108 -15526 398448 -15440
rect 398108 -15582 398174 -15526
rect 398230 -15582 398316 -15526
rect 398372 -15582 398448 -15526
rect 398108 -15668 398448 -15582
rect 398108 -15724 398174 -15668
rect 398230 -15724 398316 -15668
rect 398372 -15724 398448 -15668
rect 398108 -15810 398448 -15724
rect 398108 -15866 398174 -15810
rect 398230 -15866 398316 -15810
rect 398372 -15866 398448 -15810
rect 398108 -15952 398448 -15866
rect 398108 -16008 398174 -15952
rect 398230 -16008 398316 -15952
rect 398372 -16008 398448 -15952
rect 398108 -16094 398448 -16008
rect 398108 -16150 398174 -16094
rect 398230 -16150 398316 -16094
rect 398372 -16150 398448 -16094
rect 398108 -16236 398448 -16150
rect 398108 -16292 398174 -16236
rect 398230 -16292 398316 -16236
rect 398372 -16292 398448 -16236
rect 398108 -16378 398448 -16292
rect 398108 -16434 398174 -16378
rect 398230 -16434 398316 -16378
rect 398372 -16434 398448 -16378
rect 398108 -16520 398448 -16434
rect 398108 -16576 398174 -16520
rect 398230 -16576 398316 -16520
rect 398372 -16576 398448 -16520
rect 398108 -16662 398448 -16576
rect 398108 -16718 398174 -16662
rect 398230 -16718 398316 -16662
rect 398372 -16718 398448 -16662
rect 398108 -16804 398448 -16718
rect 398108 -16860 398174 -16804
rect 398230 -16860 398316 -16804
rect 398372 -16860 398448 -16804
rect 398108 -16946 398448 -16860
rect 398108 -17002 398174 -16946
rect 398230 -17002 398316 -16946
rect 398372 -17002 398448 -16946
rect 398108 -17088 398448 -17002
rect 398108 -17144 398174 -17088
rect 398230 -17144 398316 -17088
rect 398372 -17144 398448 -17088
rect 398108 -17230 398448 -17144
rect 398108 -17286 398174 -17230
rect 398230 -17286 398316 -17230
rect 398372 -17286 398448 -17230
rect 398108 -17372 398448 -17286
rect 398108 -17428 398174 -17372
rect 398230 -17428 398316 -17372
rect 398372 -17428 398448 -17372
rect 398108 -17514 398448 -17428
rect 398108 -17570 398174 -17514
rect 398230 -17570 398316 -17514
rect 398372 -17570 398448 -17514
rect 398108 -17656 398448 -17570
rect 398108 -17712 398174 -17656
rect 398230 -17712 398316 -17656
rect 398372 -17712 398448 -17656
rect 398108 -17798 398448 -17712
rect 398108 -17854 398174 -17798
rect 398230 -17854 398316 -17798
rect 398372 -17854 398448 -17798
rect 398108 -17940 398448 -17854
rect 398108 -17996 398174 -17940
rect 398230 -17996 398316 -17940
rect 398372 -17996 398448 -17940
rect 398108 -18082 398448 -17996
rect 398108 -18138 398174 -18082
rect 398230 -18138 398316 -18082
rect 398372 -18138 398448 -18082
rect 398108 -18224 398448 -18138
rect 398108 -18280 398174 -18224
rect 398230 -18280 398316 -18224
rect 398372 -18280 398448 -18224
rect 398108 -18366 398448 -18280
rect 398108 -18422 398174 -18366
rect 398230 -18422 398316 -18366
rect 398372 -18422 398448 -18366
rect 398108 -18508 398448 -18422
rect 398108 -18564 398174 -18508
rect 398230 -18564 398316 -18508
rect 398372 -18564 398448 -18508
rect 398108 -18650 398448 -18564
rect 398108 -18706 398174 -18650
rect 398230 -18706 398316 -18650
rect 398372 -18706 398448 -18650
rect 398108 -18792 398448 -18706
rect 398108 -18848 398174 -18792
rect 398230 -18848 398316 -18792
rect 398372 -18848 398448 -18792
rect 398108 -18934 398448 -18848
rect 398108 -18990 398174 -18934
rect 398230 -18990 398316 -18934
rect 398372 -18990 398448 -18934
rect 398108 -19076 398448 -18990
rect 398108 -19132 398174 -19076
rect 398230 -19132 398316 -19076
rect 398372 -19132 398448 -19076
rect 398108 -19218 398448 -19132
rect 398108 -19274 398174 -19218
rect 398230 -19274 398316 -19218
rect 398372 -19274 398448 -19218
rect 398108 -19360 398448 -19274
rect 398108 -19416 398174 -19360
rect 398230 -19416 398316 -19360
rect 398372 -19416 398448 -19360
rect 398108 -19502 398448 -19416
rect 398108 -19558 398174 -19502
rect 398230 -19558 398316 -19502
rect 398372 -19558 398448 -19502
rect 398108 -19644 398448 -19558
rect 398108 -19700 398174 -19644
rect 398230 -19700 398316 -19644
rect 398372 -19700 398448 -19644
rect 398108 -19786 398448 -19700
rect 398108 -19842 398174 -19786
rect 398230 -19842 398316 -19786
rect 398372 -19842 398448 -19786
rect 398108 -19928 398448 -19842
rect 398108 -19984 398174 -19928
rect 398230 -19984 398316 -19928
rect 398372 -19984 398448 -19928
rect 398108 -20070 398448 -19984
rect 398108 -20126 398174 -20070
rect 398230 -20126 398316 -20070
rect 398372 -20126 398448 -20070
rect 398108 -20212 398448 -20126
rect 398108 -20268 398174 -20212
rect 398230 -20268 398316 -20212
rect 398372 -20268 398448 -20212
rect 398108 -20354 398448 -20268
rect 398108 -20410 398174 -20354
rect 398230 -20410 398316 -20354
rect 398372 -20410 398448 -20354
rect 398108 -20496 398448 -20410
rect 398108 -20552 398174 -20496
rect 398230 -20552 398316 -20496
rect 398372 -20552 398448 -20496
rect 398108 -20638 398448 -20552
rect 398108 -20694 398174 -20638
rect 398230 -20694 398316 -20638
rect 398372 -20694 398448 -20638
rect 398108 -20780 398448 -20694
rect 398108 -20836 398174 -20780
rect 398230 -20836 398316 -20780
rect 398372 -20836 398448 -20780
rect 398108 -20922 398448 -20836
rect 398108 -20978 398174 -20922
rect 398230 -20978 398316 -20922
rect 398372 -20978 398448 -20922
rect 398108 -21064 398448 -20978
rect 398108 -21120 398174 -21064
rect 398230 -21120 398316 -21064
rect 398372 -21120 398448 -21064
rect 398108 -21206 398448 -21120
rect 398108 -21262 398174 -21206
rect 398230 -21262 398316 -21206
rect 398372 -21262 398448 -21206
rect 398108 -21348 398448 -21262
rect 398108 -21404 398174 -21348
rect 398230 -21404 398316 -21348
rect 398372 -21404 398448 -21348
rect 398108 -21490 398448 -21404
rect 398108 -21546 398174 -21490
rect 398230 -21546 398316 -21490
rect 398372 -21546 398448 -21490
rect 398108 -21632 398448 -21546
rect 398108 -21688 398174 -21632
rect 398230 -21688 398316 -21632
rect 398372 -21688 398448 -21632
rect 398108 -21774 398448 -21688
rect 398108 -21830 398174 -21774
rect 398230 -21830 398316 -21774
rect 398372 -21830 398448 -21774
rect 398108 -21916 398448 -21830
rect 398108 -21972 398174 -21916
rect 398230 -21972 398316 -21916
rect 398372 -21972 398448 -21916
rect 398108 -22058 398448 -21972
rect 398108 -22114 398174 -22058
rect 398230 -22114 398316 -22058
rect 398372 -22114 398448 -22058
rect 398108 -22200 398448 -22114
rect 398108 -22256 398174 -22200
rect 398230 -22256 398316 -22200
rect 398372 -22256 398448 -22200
rect 398108 -22342 398448 -22256
rect 398108 -22398 398174 -22342
rect 398230 -22398 398316 -22342
rect 398372 -22398 398448 -22342
rect 398108 -22484 398448 -22398
rect 398108 -22540 398174 -22484
rect 398230 -22540 398316 -22484
rect 398372 -22540 398448 -22484
rect 398108 -22626 398448 -22540
rect 398108 -22682 398174 -22626
rect 398230 -22682 398316 -22626
rect 398372 -22682 398448 -22626
rect 398108 -22768 398448 -22682
rect 398108 -22824 398174 -22768
rect 398230 -22824 398316 -22768
rect 398372 -22824 398448 -22768
rect 398108 -22910 398448 -22824
rect 398108 -22966 398174 -22910
rect 398230 -22966 398316 -22910
rect 398372 -22966 398448 -22910
rect 398108 -23052 398448 -22966
rect 398108 -23108 398174 -23052
rect 398230 -23108 398316 -23052
rect 398372 -23108 398448 -23052
rect 398108 -23194 398448 -23108
rect 398108 -23250 398174 -23194
rect 398230 -23250 398316 -23194
rect 398372 -23250 398448 -23194
rect 398108 -23336 398448 -23250
rect 398108 -23392 398174 -23336
rect 398230 -23392 398316 -23336
rect 398372 -23392 398448 -23336
rect 398108 -23478 398448 -23392
rect 398108 -23534 398174 -23478
rect 398230 -23534 398316 -23478
rect 398372 -23534 398448 -23478
rect 398108 -23620 398448 -23534
rect 398108 -23676 398174 -23620
rect 398230 -23676 398316 -23620
rect 398372 -23676 398448 -23620
rect 398108 -23762 398448 -23676
rect 398108 -23818 398174 -23762
rect 398230 -23818 398316 -23762
rect 398372 -23818 398448 -23762
rect 398108 -23904 398448 -23818
rect 398108 -23960 398174 -23904
rect 398230 -23960 398316 -23904
rect 398372 -23960 398448 -23904
rect 398108 -24046 398448 -23960
rect 398108 -24102 398174 -24046
rect 398230 -24102 398316 -24046
rect 398372 -24102 398448 -24046
rect 398108 -24188 398448 -24102
rect 398108 -24244 398174 -24188
rect 398230 -24244 398316 -24188
rect 398372 -24244 398448 -24188
rect 398108 -24330 398448 -24244
rect 398108 -24386 398174 -24330
rect 398230 -24386 398316 -24330
rect 398372 -24386 398448 -24330
rect 398108 -24472 398448 -24386
rect 398108 -24528 398174 -24472
rect 398230 -24528 398316 -24472
rect 398372 -24528 398448 -24472
rect 398108 -24614 398448 -24528
rect 398108 -24670 398174 -24614
rect 398230 -24670 398316 -24614
rect 398372 -24670 398448 -24614
rect 398108 -24756 398448 -24670
rect 398108 -24812 398174 -24756
rect 398230 -24812 398316 -24756
rect 398372 -24812 398448 -24756
rect 398108 -24898 398448 -24812
rect 398108 -24954 398174 -24898
rect 398230 -24954 398316 -24898
rect 398372 -24954 398448 -24898
rect 398108 -25040 398448 -24954
rect 398108 -25096 398174 -25040
rect 398230 -25096 398316 -25040
rect 398372 -25096 398448 -25040
rect 398108 -25182 398448 -25096
rect 398108 -25238 398174 -25182
rect 398230 -25238 398316 -25182
rect 398372 -25238 398448 -25182
rect 398108 -25324 398448 -25238
rect 398108 -25380 398174 -25324
rect 398230 -25380 398316 -25324
rect 398372 -25380 398448 -25324
rect 398108 -25466 398448 -25380
rect 398108 -25522 398174 -25466
rect 398230 -25522 398316 -25466
rect 398372 -25522 398448 -25466
rect 398108 -25590 398448 -25522
rect 398508 -13680 398848 -13590
rect 398508 -13736 398574 -13680
rect 398630 -13736 398716 -13680
rect 398772 -13736 398848 -13680
rect 398508 -13822 398848 -13736
rect 398508 -13878 398574 -13822
rect 398630 -13878 398716 -13822
rect 398772 -13878 398848 -13822
rect 398508 -13964 398848 -13878
rect 398508 -14020 398574 -13964
rect 398630 -14020 398716 -13964
rect 398772 -14020 398848 -13964
rect 398508 -14106 398848 -14020
rect 398508 -14162 398574 -14106
rect 398630 -14162 398716 -14106
rect 398772 -14162 398848 -14106
rect 398508 -14248 398848 -14162
rect 398508 -14304 398574 -14248
rect 398630 -14304 398716 -14248
rect 398772 -14304 398848 -14248
rect 398508 -14390 398848 -14304
rect 398508 -14446 398574 -14390
rect 398630 -14446 398716 -14390
rect 398772 -14446 398848 -14390
rect 398508 -14532 398848 -14446
rect 398508 -14588 398574 -14532
rect 398630 -14588 398716 -14532
rect 398772 -14588 398848 -14532
rect 398508 -14674 398848 -14588
rect 398508 -14730 398574 -14674
rect 398630 -14730 398716 -14674
rect 398772 -14730 398848 -14674
rect 398508 -14816 398848 -14730
rect 398508 -14872 398574 -14816
rect 398630 -14872 398716 -14816
rect 398772 -14872 398848 -14816
rect 398508 -14958 398848 -14872
rect 398508 -15014 398574 -14958
rect 398630 -15014 398716 -14958
rect 398772 -15014 398848 -14958
rect 398508 -15100 398848 -15014
rect 398508 -15156 398574 -15100
rect 398630 -15156 398716 -15100
rect 398772 -15156 398848 -15100
rect 398508 -15242 398848 -15156
rect 398508 -15298 398574 -15242
rect 398630 -15298 398716 -15242
rect 398772 -15298 398848 -15242
rect 398508 -15384 398848 -15298
rect 398508 -15440 398574 -15384
rect 398630 -15440 398716 -15384
rect 398772 -15440 398848 -15384
rect 398508 -15526 398848 -15440
rect 398508 -15582 398574 -15526
rect 398630 -15582 398716 -15526
rect 398772 -15582 398848 -15526
rect 398508 -15668 398848 -15582
rect 398508 -15724 398574 -15668
rect 398630 -15724 398716 -15668
rect 398772 -15724 398848 -15668
rect 398508 -15810 398848 -15724
rect 398508 -15866 398574 -15810
rect 398630 -15866 398716 -15810
rect 398772 -15866 398848 -15810
rect 398508 -15952 398848 -15866
rect 398508 -16008 398574 -15952
rect 398630 -16008 398716 -15952
rect 398772 -16008 398848 -15952
rect 398508 -16094 398848 -16008
rect 398508 -16150 398574 -16094
rect 398630 -16150 398716 -16094
rect 398772 -16150 398848 -16094
rect 398508 -16236 398848 -16150
rect 398508 -16292 398574 -16236
rect 398630 -16292 398716 -16236
rect 398772 -16292 398848 -16236
rect 398508 -16378 398848 -16292
rect 398508 -16434 398574 -16378
rect 398630 -16434 398716 -16378
rect 398772 -16434 398848 -16378
rect 398508 -16520 398848 -16434
rect 398508 -16576 398574 -16520
rect 398630 -16576 398716 -16520
rect 398772 -16576 398848 -16520
rect 398508 -16662 398848 -16576
rect 398508 -16718 398574 -16662
rect 398630 -16718 398716 -16662
rect 398772 -16718 398848 -16662
rect 398508 -16804 398848 -16718
rect 398508 -16860 398574 -16804
rect 398630 -16860 398716 -16804
rect 398772 -16860 398848 -16804
rect 398508 -16946 398848 -16860
rect 398508 -17002 398574 -16946
rect 398630 -17002 398716 -16946
rect 398772 -17002 398848 -16946
rect 398508 -17088 398848 -17002
rect 398508 -17144 398574 -17088
rect 398630 -17144 398716 -17088
rect 398772 -17144 398848 -17088
rect 398508 -17230 398848 -17144
rect 398508 -17286 398574 -17230
rect 398630 -17286 398716 -17230
rect 398772 -17286 398848 -17230
rect 398508 -17372 398848 -17286
rect 398508 -17428 398574 -17372
rect 398630 -17428 398716 -17372
rect 398772 -17428 398848 -17372
rect 398508 -17514 398848 -17428
rect 398508 -17570 398574 -17514
rect 398630 -17570 398716 -17514
rect 398772 -17570 398848 -17514
rect 398508 -17656 398848 -17570
rect 398508 -17712 398574 -17656
rect 398630 -17712 398716 -17656
rect 398772 -17712 398848 -17656
rect 398508 -17798 398848 -17712
rect 398508 -17854 398574 -17798
rect 398630 -17854 398716 -17798
rect 398772 -17854 398848 -17798
rect 398508 -17940 398848 -17854
rect 398508 -17996 398574 -17940
rect 398630 -17996 398716 -17940
rect 398772 -17996 398848 -17940
rect 398508 -18082 398848 -17996
rect 398508 -18138 398574 -18082
rect 398630 -18138 398716 -18082
rect 398772 -18138 398848 -18082
rect 398508 -18224 398848 -18138
rect 398508 -18280 398574 -18224
rect 398630 -18280 398716 -18224
rect 398772 -18280 398848 -18224
rect 398508 -18366 398848 -18280
rect 398508 -18422 398574 -18366
rect 398630 -18422 398716 -18366
rect 398772 -18422 398848 -18366
rect 398508 -18508 398848 -18422
rect 398508 -18564 398574 -18508
rect 398630 -18564 398716 -18508
rect 398772 -18564 398848 -18508
rect 398508 -18650 398848 -18564
rect 398508 -18706 398574 -18650
rect 398630 -18706 398716 -18650
rect 398772 -18706 398848 -18650
rect 398508 -18792 398848 -18706
rect 398508 -18848 398574 -18792
rect 398630 -18848 398716 -18792
rect 398772 -18848 398848 -18792
rect 398508 -18934 398848 -18848
rect 398508 -18990 398574 -18934
rect 398630 -18990 398716 -18934
rect 398772 -18990 398848 -18934
rect 398508 -19076 398848 -18990
rect 398508 -19132 398574 -19076
rect 398630 -19132 398716 -19076
rect 398772 -19132 398848 -19076
rect 398508 -19218 398848 -19132
rect 398508 -19274 398574 -19218
rect 398630 -19274 398716 -19218
rect 398772 -19274 398848 -19218
rect 398508 -19360 398848 -19274
rect 398508 -19416 398574 -19360
rect 398630 -19416 398716 -19360
rect 398772 -19416 398848 -19360
rect 398508 -19502 398848 -19416
rect 398508 -19558 398574 -19502
rect 398630 -19558 398716 -19502
rect 398772 -19558 398848 -19502
rect 398508 -19644 398848 -19558
rect 398508 -19700 398574 -19644
rect 398630 -19700 398716 -19644
rect 398772 -19700 398848 -19644
rect 398508 -19786 398848 -19700
rect 398508 -19842 398574 -19786
rect 398630 -19842 398716 -19786
rect 398772 -19842 398848 -19786
rect 398508 -19928 398848 -19842
rect 398508 -19984 398574 -19928
rect 398630 -19984 398716 -19928
rect 398772 -19984 398848 -19928
rect 398508 -20070 398848 -19984
rect 398508 -20126 398574 -20070
rect 398630 -20126 398716 -20070
rect 398772 -20126 398848 -20070
rect 398508 -20212 398848 -20126
rect 398508 -20268 398574 -20212
rect 398630 -20268 398716 -20212
rect 398772 -20268 398848 -20212
rect 398508 -20354 398848 -20268
rect 398508 -20410 398574 -20354
rect 398630 -20410 398716 -20354
rect 398772 -20410 398848 -20354
rect 398508 -20496 398848 -20410
rect 398508 -20552 398574 -20496
rect 398630 -20552 398716 -20496
rect 398772 -20552 398848 -20496
rect 398508 -20638 398848 -20552
rect 398508 -20694 398574 -20638
rect 398630 -20694 398716 -20638
rect 398772 -20694 398848 -20638
rect 398508 -20780 398848 -20694
rect 398508 -20836 398574 -20780
rect 398630 -20836 398716 -20780
rect 398772 -20836 398848 -20780
rect 398508 -20922 398848 -20836
rect 398508 -20978 398574 -20922
rect 398630 -20978 398716 -20922
rect 398772 -20978 398848 -20922
rect 398508 -21064 398848 -20978
rect 398508 -21120 398574 -21064
rect 398630 -21120 398716 -21064
rect 398772 -21120 398848 -21064
rect 398508 -21206 398848 -21120
rect 398508 -21262 398574 -21206
rect 398630 -21262 398716 -21206
rect 398772 -21262 398848 -21206
rect 398508 -21348 398848 -21262
rect 398508 -21404 398574 -21348
rect 398630 -21404 398716 -21348
rect 398772 -21404 398848 -21348
rect 398508 -21490 398848 -21404
rect 398508 -21546 398574 -21490
rect 398630 -21546 398716 -21490
rect 398772 -21546 398848 -21490
rect 398508 -21632 398848 -21546
rect 398508 -21688 398574 -21632
rect 398630 -21688 398716 -21632
rect 398772 -21688 398848 -21632
rect 398508 -21774 398848 -21688
rect 398508 -21830 398574 -21774
rect 398630 -21830 398716 -21774
rect 398772 -21830 398848 -21774
rect 398508 -21916 398848 -21830
rect 398508 -21972 398574 -21916
rect 398630 -21972 398716 -21916
rect 398772 -21972 398848 -21916
rect 398508 -22058 398848 -21972
rect 398508 -22114 398574 -22058
rect 398630 -22114 398716 -22058
rect 398772 -22114 398848 -22058
rect 398508 -22200 398848 -22114
rect 398508 -22256 398574 -22200
rect 398630 -22256 398716 -22200
rect 398772 -22256 398848 -22200
rect 398508 -22342 398848 -22256
rect 398508 -22398 398574 -22342
rect 398630 -22398 398716 -22342
rect 398772 -22398 398848 -22342
rect 398508 -22484 398848 -22398
rect 398508 -22540 398574 -22484
rect 398630 -22540 398716 -22484
rect 398772 -22540 398848 -22484
rect 398508 -22626 398848 -22540
rect 398508 -22682 398574 -22626
rect 398630 -22682 398716 -22626
rect 398772 -22682 398848 -22626
rect 398508 -22768 398848 -22682
rect 398508 -22824 398574 -22768
rect 398630 -22824 398716 -22768
rect 398772 -22824 398848 -22768
rect 398508 -22910 398848 -22824
rect 398508 -22966 398574 -22910
rect 398630 -22966 398716 -22910
rect 398772 -22966 398848 -22910
rect 398508 -23052 398848 -22966
rect 398508 -23108 398574 -23052
rect 398630 -23108 398716 -23052
rect 398772 -23108 398848 -23052
rect 398508 -23194 398848 -23108
rect 398508 -23250 398574 -23194
rect 398630 -23250 398716 -23194
rect 398772 -23250 398848 -23194
rect 398508 -23336 398848 -23250
rect 398508 -23392 398574 -23336
rect 398630 -23392 398716 -23336
rect 398772 -23392 398848 -23336
rect 398508 -23478 398848 -23392
rect 398508 -23534 398574 -23478
rect 398630 -23534 398716 -23478
rect 398772 -23534 398848 -23478
rect 398508 -23620 398848 -23534
rect 398508 -23676 398574 -23620
rect 398630 -23676 398716 -23620
rect 398772 -23676 398848 -23620
rect 398508 -23762 398848 -23676
rect 398508 -23818 398574 -23762
rect 398630 -23818 398716 -23762
rect 398772 -23818 398848 -23762
rect 398508 -23904 398848 -23818
rect 398508 -23960 398574 -23904
rect 398630 -23960 398716 -23904
rect 398772 -23960 398848 -23904
rect 398508 -24046 398848 -23960
rect 398508 -24102 398574 -24046
rect 398630 -24102 398716 -24046
rect 398772 -24102 398848 -24046
rect 398508 -24188 398848 -24102
rect 398508 -24244 398574 -24188
rect 398630 -24244 398716 -24188
rect 398772 -24244 398848 -24188
rect 398508 -24330 398848 -24244
rect 398508 -24386 398574 -24330
rect 398630 -24386 398716 -24330
rect 398772 -24386 398848 -24330
rect 398508 -24472 398848 -24386
rect 398508 -24528 398574 -24472
rect 398630 -24528 398716 -24472
rect 398772 -24528 398848 -24472
rect 398508 -24614 398848 -24528
rect 398508 -24670 398574 -24614
rect 398630 -24670 398716 -24614
rect 398772 -24670 398848 -24614
rect 398508 -24756 398848 -24670
rect 398508 -24812 398574 -24756
rect 398630 -24812 398716 -24756
rect 398772 -24812 398848 -24756
rect 398508 -24898 398848 -24812
rect 398508 -24954 398574 -24898
rect 398630 -24954 398716 -24898
rect 398772 -24954 398848 -24898
rect 398508 -25040 398848 -24954
rect 398508 -25096 398574 -25040
rect 398630 -25096 398716 -25040
rect 398772 -25096 398848 -25040
rect 398508 -25182 398848 -25096
rect 398508 -25238 398574 -25182
rect 398630 -25238 398716 -25182
rect 398772 -25238 398848 -25182
rect 398508 -25324 398848 -25238
rect 398508 -25380 398574 -25324
rect 398630 -25380 398716 -25324
rect 398772 -25380 398848 -25324
rect 398508 -25466 398848 -25380
rect 398508 -25522 398574 -25466
rect 398630 -25522 398716 -25466
rect 398772 -25522 398848 -25466
rect 398508 -25590 398848 -25522
rect 398908 -13680 399248 -13590
rect 398908 -13736 398971 -13680
rect 399027 -13736 399113 -13680
rect 399169 -13736 399248 -13680
rect 398908 -13822 399248 -13736
rect 398908 -13878 398971 -13822
rect 399027 -13878 399113 -13822
rect 399169 -13878 399248 -13822
rect 398908 -13964 399248 -13878
rect 398908 -14020 398971 -13964
rect 399027 -14020 399113 -13964
rect 399169 -14020 399248 -13964
rect 398908 -14106 399248 -14020
rect 398908 -14162 398971 -14106
rect 399027 -14162 399113 -14106
rect 399169 -14162 399248 -14106
rect 398908 -14248 399248 -14162
rect 398908 -14304 398971 -14248
rect 399027 -14304 399113 -14248
rect 399169 -14304 399248 -14248
rect 398908 -14390 399248 -14304
rect 398908 -14446 398971 -14390
rect 399027 -14446 399113 -14390
rect 399169 -14446 399248 -14390
rect 398908 -14532 399248 -14446
rect 398908 -14588 398971 -14532
rect 399027 -14588 399113 -14532
rect 399169 -14588 399248 -14532
rect 398908 -14674 399248 -14588
rect 398908 -14730 398971 -14674
rect 399027 -14730 399113 -14674
rect 399169 -14730 399248 -14674
rect 398908 -14816 399248 -14730
rect 398908 -14872 398971 -14816
rect 399027 -14872 399113 -14816
rect 399169 -14872 399248 -14816
rect 398908 -14958 399248 -14872
rect 398908 -15014 398971 -14958
rect 399027 -15014 399113 -14958
rect 399169 -15014 399248 -14958
rect 398908 -15100 399248 -15014
rect 398908 -15156 398971 -15100
rect 399027 -15156 399113 -15100
rect 399169 -15156 399248 -15100
rect 398908 -15242 399248 -15156
rect 398908 -15298 398971 -15242
rect 399027 -15298 399113 -15242
rect 399169 -15298 399248 -15242
rect 398908 -15384 399248 -15298
rect 398908 -15440 398971 -15384
rect 399027 -15440 399113 -15384
rect 399169 -15440 399248 -15384
rect 398908 -15526 399248 -15440
rect 398908 -15582 398971 -15526
rect 399027 -15582 399113 -15526
rect 399169 -15582 399248 -15526
rect 398908 -15668 399248 -15582
rect 398908 -15724 398971 -15668
rect 399027 -15724 399113 -15668
rect 399169 -15724 399248 -15668
rect 398908 -15810 399248 -15724
rect 398908 -15866 398971 -15810
rect 399027 -15866 399113 -15810
rect 399169 -15866 399248 -15810
rect 398908 -15952 399248 -15866
rect 398908 -16008 398971 -15952
rect 399027 -16008 399113 -15952
rect 399169 -16008 399248 -15952
rect 398908 -16094 399248 -16008
rect 398908 -16150 398971 -16094
rect 399027 -16150 399113 -16094
rect 399169 -16150 399248 -16094
rect 398908 -16236 399248 -16150
rect 398908 -16292 398971 -16236
rect 399027 -16292 399113 -16236
rect 399169 -16292 399248 -16236
rect 398908 -16378 399248 -16292
rect 398908 -16434 398971 -16378
rect 399027 -16434 399113 -16378
rect 399169 -16434 399248 -16378
rect 398908 -16520 399248 -16434
rect 398908 -16576 398971 -16520
rect 399027 -16576 399113 -16520
rect 399169 -16576 399248 -16520
rect 398908 -16662 399248 -16576
rect 398908 -16718 398971 -16662
rect 399027 -16718 399113 -16662
rect 399169 -16718 399248 -16662
rect 398908 -16804 399248 -16718
rect 398908 -16860 398971 -16804
rect 399027 -16860 399113 -16804
rect 399169 -16860 399248 -16804
rect 398908 -16946 399248 -16860
rect 398908 -17002 398971 -16946
rect 399027 -17002 399113 -16946
rect 399169 -17002 399248 -16946
rect 398908 -17088 399248 -17002
rect 398908 -17144 398971 -17088
rect 399027 -17144 399113 -17088
rect 399169 -17144 399248 -17088
rect 398908 -17230 399248 -17144
rect 398908 -17286 398971 -17230
rect 399027 -17286 399113 -17230
rect 399169 -17286 399248 -17230
rect 398908 -17372 399248 -17286
rect 398908 -17428 398971 -17372
rect 399027 -17428 399113 -17372
rect 399169 -17428 399248 -17372
rect 398908 -17514 399248 -17428
rect 398908 -17570 398971 -17514
rect 399027 -17570 399113 -17514
rect 399169 -17570 399248 -17514
rect 398908 -17656 399248 -17570
rect 398908 -17712 398971 -17656
rect 399027 -17712 399113 -17656
rect 399169 -17712 399248 -17656
rect 398908 -17798 399248 -17712
rect 398908 -17854 398971 -17798
rect 399027 -17854 399113 -17798
rect 399169 -17854 399248 -17798
rect 398908 -17940 399248 -17854
rect 398908 -17996 398971 -17940
rect 399027 -17996 399113 -17940
rect 399169 -17996 399248 -17940
rect 398908 -18082 399248 -17996
rect 398908 -18138 398971 -18082
rect 399027 -18138 399113 -18082
rect 399169 -18138 399248 -18082
rect 398908 -18224 399248 -18138
rect 398908 -18280 398971 -18224
rect 399027 -18280 399113 -18224
rect 399169 -18280 399248 -18224
rect 398908 -18366 399248 -18280
rect 398908 -18422 398971 -18366
rect 399027 -18422 399113 -18366
rect 399169 -18422 399248 -18366
rect 398908 -18508 399248 -18422
rect 398908 -18564 398971 -18508
rect 399027 -18564 399113 -18508
rect 399169 -18564 399248 -18508
rect 398908 -18650 399248 -18564
rect 398908 -18706 398971 -18650
rect 399027 -18706 399113 -18650
rect 399169 -18706 399248 -18650
rect 398908 -18792 399248 -18706
rect 398908 -18848 398971 -18792
rect 399027 -18848 399113 -18792
rect 399169 -18848 399248 -18792
rect 398908 -18934 399248 -18848
rect 398908 -18990 398971 -18934
rect 399027 -18990 399113 -18934
rect 399169 -18990 399248 -18934
rect 398908 -19076 399248 -18990
rect 398908 -19132 398971 -19076
rect 399027 -19132 399113 -19076
rect 399169 -19132 399248 -19076
rect 398908 -19218 399248 -19132
rect 398908 -19274 398971 -19218
rect 399027 -19274 399113 -19218
rect 399169 -19274 399248 -19218
rect 398908 -19360 399248 -19274
rect 398908 -19416 398971 -19360
rect 399027 -19416 399113 -19360
rect 399169 -19416 399248 -19360
rect 398908 -19502 399248 -19416
rect 398908 -19558 398971 -19502
rect 399027 -19558 399113 -19502
rect 399169 -19558 399248 -19502
rect 398908 -19644 399248 -19558
rect 398908 -19700 398971 -19644
rect 399027 -19700 399113 -19644
rect 399169 -19700 399248 -19644
rect 398908 -19786 399248 -19700
rect 398908 -19842 398971 -19786
rect 399027 -19842 399113 -19786
rect 399169 -19842 399248 -19786
rect 398908 -19928 399248 -19842
rect 398908 -19984 398971 -19928
rect 399027 -19984 399113 -19928
rect 399169 -19984 399248 -19928
rect 398908 -20070 399248 -19984
rect 398908 -20126 398971 -20070
rect 399027 -20126 399113 -20070
rect 399169 -20126 399248 -20070
rect 398908 -20212 399248 -20126
rect 398908 -20268 398971 -20212
rect 399027 -20268 399113 -20212
rect 399169 -20268 399248 -20212
rect 398908 -20354 399248 -20268
rect 398908 -20410 398971 -20354
rect 399027 -20410 399113 -20354
rect 399169 -20410 399248 -20354
rect 398908 -20496 399248 -20410
rect 398908 -20552 398971 -20496
rect 399027 -20552 399113 -20496
rect 399169 -20552 399248 -20496
rect 398908 -20638 399248 -20552
rect 398908 -20694 398971 -20638
rect 399027 -20694 399113 -20638
rect 399169 -20694 399248 -20638
rect 398908 -20780 399248 -20694
rect 398908 -20836 398971 -20780
rect 399027 -20836 399113 -20780
rect 399169 -20836 399248 -20780
rect 398908 -20922 399248 -20836
rect 398908 -20978 398971 -20922
rect 399027 -20978 399113 -20922
rect 399169 -20978 399248 -20922
rect 398908 -21064 399248 -20978
rect 398908 -21120 398971 -21064
rect 399027 -21120 399113 -21064
rect 399169 -21120 399248 -21064
rect 398908 -21206 399248 -21120
rect 398908 -21262 398971 -21206
rect 399027 -21262 399113 -21206
rect 399169 -21262 399248 -21206
rect 398908 -21348 399248 -21262
rect 398908 -21404 398971 -21348
rect 399027 -21404 399113 -21348
rect 399169 -21404 399248 -21348
rect 398908 -21490 399248 -21404
rect 398908 -21546 398971 -21490
rect 399027 -21546 399113 -21490
rect 399169 -21546 399248 -21490
rect 398908 -21632 399248 -21546
rect 398908 -21688 398971 -21632
rect 399027 -21688 399113 -21632
rect 399169 -21688 399248 -21632
rect 398908 -21774 399248 -21688
rect 398908 -21830 398971 -21774
rect 399027 -21830 399113 -21774
rect 399169 -21830 399248 -21774
rect 398908 -21916 399248 -21830
rect 398908 -21972 398971 -21916
rect 399027 -21972 399113 -21916
rect 399169 -21972 399248 -21916
rect 398908 -22058 399248 -21972
rect 398908 -22114 398971 -22058
rect 399027 -22114 399113 -22058
rect 399169 -22114 399248 -22058
rect 398908 -22200 399248 -22114
rect 398908 -22256 398971 -22200
rect 399027 -22256 399113 -22200
rect 399169 -22256 399248 -22200
rect 398908 -22342 399248 -22256
rect 398908 -22398 398971 -22342
rect 399027 -22398 399113 -22342
rect 399169 -22398 399248 -22342
rect 398908 -22484 399248 -22398
rect 398908 -22540 398971 -22484
rect 399027 -22540 399113 -22484
rect 399169 -22540 399248 -22484
rect 398908 -22626 399248 -22540
rect 398908 -22682 398971 -22626
rect 399027 -22682 399113 -22626
rect 399169 -22682 399248 -22626
rect 398908 -22768 399248 -22682
rect 398908 -22824 398971 -22768
rect 399027 -22824 399113 -22768
rect 399169 -22824 399248 -22768
rect 398908 -22910 399248 -22824
rect 398908 -22966 398971 -22910
rect 399027 -22966 399113 -22910
rect 399169 -22966 399248 -22910
rect 398908 -23052 399248 -22966
rect 398908 -23108 398971 -23052
rect 399027 -23108 399113 -23052
rect 399169 -23108 399248 -23052
rect 398908 -23194 399248 -23108
rect 398908 -23250 398971 -23194
rect 399027 -23250 399113 -23194
rect 399169 -23250 399248 -23194
rect 398908 -23336 399248 -23250
rect 398908 -23392 398971 -23336
rect 399027 -23392 399113 -23336
rect 399169 -23392 399248 -23336
rect 398908 -23478 399248 -23392
rect 398908 -23534 398971 -23478
rect 399027 -23534 399113 -23478
rect 399169 -23534 399248 -23478
rect 398908 -23620 399248 -23534
rect 398908 -23676 398971 -23620
rect 399027 -23676 399113 -23620
rect 399169 -23676 399248 -23620
rect 398908 -23762 399248 -23676
rect 398908 -23818 398971 -23762
rect 399027 -23818 399113 -23762
rect 399169 -23818 399248 -23762
rect 398908 -23904 399248 -23818
rect 398908 -23960 398971 -23904
rect 399027 -23960 399113 -23904
rect 399169 -23960 399248 -23904
rect 398908 -24046 399248 -23960
rect 398908 -24102 398971 -24046
rect 399027 -24102 399113 -24046
rect 399169 -24102 399248 -24046
rect 398908 -24188 399248 -24102
rect 398908 -24244 398971 -24188
rect 399027 -24244 399113 -24188
rect 399169 -24244 399248 -24188
rect 398908 -24330 399248 -24244
rect 398908 -24386 398971 -24330
rect 399027 -24386 399113 -24330
rect 399169 -24386 399248 -24330
rect 398908 -24472 399248 -24386
rect 398908 -24528 398971 -24472
rect 399027 -24528 399113 -24472
rect 399169 -24528 399248 -24472
rect 398908 -24614 399248 -24528
rect 398908 -24670 398971 -24614
rect 399027 -24670 399113 -24614
rect 399169 -24670 399248 -24614
rect 398908 -24756 399248 -24670
rect 398908 -24812 398971 -24756
rect 399027 -24812 399113 -24756
rect 399169 -24812 399248 -24756
rect 398908 -24898 399248 -24812
rect 398908 -24954 398971 -24898
rect 399027 -24954 399113 -24898
rect 399169 -24954 399248 -24898
rect 398908 -25040 399248 -24954
rect 398908 -25096 398971 -25040
rect 399027 -25096 399113 -25040
rect 399169 -25096 399248 -25040
rect 398908 -25182 399248 -25096
rect 398908 -25238 398971 -25182
rect 399027 -25238 399113 -25182
rect 399169 -25238 399248 -25182
rect 398908 -25324 399248 -25238
rect 398908 -25380 398971 -25324
rect 399027 -25380 399113 -25324
rect 399169 -25380 399248 -25324
rect 398908 -25466 399248 -25380
rect 398908 -25522 398971 -25466
rect 399027 -25522 399113 -25466
rect 399169 -25522 399248 -25466
rect 398908 -25590 399248 -25522
rect 399308 -13680 399648 -13590
rect 399308 -13736 399376 -13680
rect 399432 -13736 399518 -13680
rect 399574 -13736 399648 -13680
rect 399308 -13822 399648 -13736
rect 399308 -13878 399376 -13822
rect 399432 -13878 399518 -13822
rect 399574 -13878 399648 -13822
rect 399308 -13964 399648 -13878
rect 399308 -14020 399376 -13964
rect 399432 -14020 399518 -13964
rect 399574 -14020 399648 -13964
rect 399308 -14106 399648 -14020
rect 399308 -14162 399376 -14106
rect 399432 -14162 399518 -14106
rect 399574 -14162 399648 -14106
rect 399308 -14248 399648 -14162
rect 399308 -14304 399376 -14248
rect 399432 -14304 399518 -14248
rect 399574 -14304 399648 -14248
rect 399308 -14390 399648 -14304
rect 399308 -14446 399376 -14390
rect 399432 -14446 399518 -14390
rect 399574 -14446 399648 -14390
rect 399308 -14532 399648 -14446
rect 399308 -14588 399376 -14532
rect 399432 -14588 399518 -14532
rect 399574 -14588 399648 -14532
rect 399308 -14674 399648 -14588
rect 399308 -14730 399376 -14674
rect 399432 -14730 399518 -14674
rect 399574 -14730 399648 -14674
rect 399308 -14816 399648 -14730
rect 399308 -14872 399376 -14816
rect 399432 -14872 399518 -14816
rect 399574 -14872 399648 -14816
rect 399308 -14958 399648 -14872
rect 399308 -15014 399376 -14958
rect 399432 -15014 399518 -14958
rect 399574 -15014 399648 -14958
rect 399308 -15100 399648 -15014
rect 399308 -15156 399376 -15100
rect 399432 -15156 399518 -15100
rect 399574 -15156 399648 -15100
rect 399308 -15242 399648 -15156
rect 399308 -15298 399376 -15242
rect 399432 -15298 399518 -15242
rect 399574 -15298 399648 -15242
rect 399308 -15384 399648 -15298
rect 399308 -15440 399376 -15384
rect 399432 -15440 399518 -15384
rect 399574 -15440 399648 -15384
rect 399308 -15526 399648 -15440
rect 399308 -15582 399376 -15526
rect 399432 -15582 399518 -15526
rect 399574 -15582 399648 -15526
rect 399308 -15668 399648 -15582
rect 399308 -15724 399376 -15668
rect 399432 -15724 399518 -15668
rect 399574 -15724 399648 -15668
rect 399308 -15810 399648 -15724
rect 399308 -15866 399376 -15810
rect 399432 -15866 399518 -15810
rect 399574 -15866 399648 -15810
rect 399308 -15952 399648 -15866
rect 399308 -16008 399376 -15952
rect 399432 -16008 399518 -15952
rect 399574 -16008 399648 -15952
rect 399308 -16094 399648 -16008
rect 399308 -16150 399376 -16094
rect 399432 -16150 399518 -16094
rect 399574 -16150 399648 -16094
rect 399308 -16236 399648 -16150
rect 399308 -16292 399376 -16236
rect 399432 -16292 399518 -16236
rect 399574 -16292 399648 -16236
rect 399308 -16378 399648 -16292
rect 399308 -16434 399376 -16378
rect 399432 -16434 399518 -16378
rect 399574 -16434 399648 -16378
rect 399308 -16520 399648 -16434
rect 399308 -16576 399376 -16520
rect 399432 -16576 399518 -16520
rect 399574 -16576 399648 -16520
rect 399308 -16662 399648 -16576
rect 399308 -16718 399376 -16662
rect 399432 -16718 399518 -16662
rect 399574 -16718 399648 -16662
rect 399308 -16804 399648 -16718
rect 399308 -16860 399376 -16804
rect 399432 -16860 399518 -16804
rect 399574 -16860 399648 -16804
rect 399308 -16946 399648 -16860
rect 399308 -17002 399376 -16946
rect 399432 -17002 399518 -16946
rect 399574 -17002 399648 -16946
rect 399308 -17088 399648 -17002
rect 399308 -17144 399376 -17088
rect 399432 -17144 399518 -17088
rect 399574 -17144 399648 -17088
rect 399308 -17230 399648 -17144
rect 399308 -17286 399376 -17230
rect 399432 -17286 399518 -17230
rect 399574 -17286 399648 -17230
rect 399308 -17372 399648 -17286
rect 399308 -17428 399376 -17372
rect 399432 -17428 399518 -17372
rect 399574 -17428 399648 -17372
rect 399308 -17514 399648 -17428
rect 399308 -17570 399376 -17514
rect 399432 -17570 399518 -17514
rect 399574 -17570 399648 -17514
rect 399308 -17656 399648 -17570
rect 399308 -17712 399376 -17656
rect 399432 -17712 399518 -17656
rect 399574 -17712 399648 -17656
rect 399308 -17798 399648 -17712
rect 399308 -17854 399376 -17798
rect 399432 -17854 399518 -17798
rect 399574 -17854 399648 -17798
rect 399308 -17940 399648 -17854
rect 399308 -17996 399376 -17940
rect 399432 -17996 399518 -17940
rect 399574 -17996 399648 -17940
rect 399308 -18082 399648 -17996
rect 399308 -18138 399376 -18082
rect 399432 -18138 399518 -18082
rect 399574 -18138 399648 -18082
rect 399308 -18224 399648 -18138
rect 399308 -18280 399376 -18224
rect 399432 -18280 399518 -18224
rect 399574 -18280 399648 -18224
rect 399308 -18366 399648 -18280
rect 399308 -18422 399376 -18366
rect 399432 -18422 399518 -18366
rect 399574 -18422 399648 -18366
rect 399308 -18508 399648 -18422
rect 399308 -18564 399376 -18508
rect 399432 -18564 399518 -18508
rect 399574 -18564 399648 -18508
rect 399308 -18650 399648 -18564
rect 399308 -18706 399376 -18650
rect 399432 -18706 399518 -18650
rect 399574 -18706 399648 -18650
rect 399308 -18792 399648 -18706
rect 399308 -18848 399376 -18792
rect 399432 -18848 399518 -18792
rect 399574 -18848 399648 -18792
rect 399308 -18934 399648 -18848
rect 399308 -18990 399376 -18934
rect 399432 -18990 399518 -18934
rect 399574 -18990 399648 -18934
rect 399308 -19076 399648 -18990
rect 399308 -19132 399376 -19076
rect 399432 -19132 399518 -19076
rect 399574 -19132 399648 -19076
rect 399308 -19218 399648 -19132
rect 399308 -19274 399376 -19218
rect 399432 -19274 399518 -19218
rect 399574 -19274 399648 -19218
rect 399308 -19360 399648 -19274
rect 399308 -19416 399376 -19360
rect 399432 -19416 399518 -19360
rect 399574 -19416 399648 -19360
rect 399308 -19502 399648 -19416
rect 399308 -19558 399376 -19502
rect 399432 -19558 399518 -19502
rect 399574 -19558 399648 -19502
rect 399308 -19644 399648 -19558
rect 399308 -19700 399376 -19644
rect 399432 -19700 399518 -19644
rect 399574 -19700 399648 -19644
rect 399308 -19786 399648 -19700
rect 399308 -19842 399376 -19786
rect 399432 -19842 399518 -19786
rect 399574 -19842 399648 -19786
rect 399308 -19928 399648 -19842
rect 399308 -19984 399376 -19928
rect 399432 -19984 399518 -19928
rect 399574 -19984 399648 -19928
rect 399308 -20070 399648 -19984
rect 399308 -20126 399376 -20070
rect 399432 -20126 399518 -20070
rect 399574 -20126 399648 -20070
rect 399308 -20212 399648 -20126
rect 399308 -20268 399376 -20212
rect 399432 -20268 399518 -20212
rect 399574 -20268 399648 -20212
rect 399308 -20354 399648 -20268
rect 399308 -20410 399376 -20354
rect 399432 -20410 399518 -20354
rect 399574 -20410 399648 -20354
rect 399308 -20496 399648 -20410
rect 399308 -20552 399376 -20496
rect 399432 -20552 399518 -20496
rect 399574 -20552 399648 -20496
rect 399308 -20638 399648 -20552
rect 399308 -20694 399376 -20638
rect 399432 -20694 399518 -20638
rect 399574 -20694 399648 -20638
rect 399308 -20780 399648 -20694
rect 399308 -20836 399376 -20780
rect 399432 -20836 399518 -20780
rect 399574 -20836 399648 -20780
rect 399308 -20922 399648 -20836
rect 399308 -20978 399376 -20922
rect 399432 -20978 399518 -20922
rect 399574 -20978 399648 -20922
rect 399308 -21064 399648 -20978
rect 399308 -21120 399376 -21064
rect 399432 -21120 399518 -21064
rect 399574 -21120 399648 -21064
rect 399308 -21206 399648 -21120
rect 399308 -21262 399376 -21206
rect 399432 -21262 399518 -21206
rect 399574 -21262 399648 -21206
rect 399308 -21348 399648 -21262
rect 399308 -21404 399376 -21348
rect 399432 -21404 399518 -21348
rect 399574 -21404 399648 -21348
rect 399308 -21490 399648 -21404
rect 399308 -21546 399376 -21490
rect 399432 -21546 399518 -21490
rect 399574 -21546 399648 -21490
rect 399308 -21632 399648 -21546
rect 399308 -21688 399376 -21632
rect 399432 -21688 399518 -21632
rect 399574 -21688 399648 -21632
rect 399308 -21774 399648 -21688
rect 399308 -21830 399376 -21774
rect 399432 -21830 399518 -21774
rect 399574 -21830 399648 -21774
rect 399308 -21916 399648 -21830
rect 399308 -21972 399376 -21916
rect 399432 -21972 399518 -21916
rect 399574 -21972 399648 -21916
rect 399308 -22058 399648 -21972
rect 399308 -22114 399376 -22058
rect 399432 -22114 399518 -22058
rect 399574 -22114 399648 -22058
rect 399308 -22200 399648 -22114
rect 399308 -22256 399376 -22200
rect 399432 -22256 399518 -22200
rect 399574 -22256 399648 -22200
rect 399308 -22342 399648 -22256
rect 399308 -22398 399376 -22342
rect 399432 -22398 399518 -22342
rect 399574 -22398 399648 -22342
rect 399308 -22484 399648 -22398
rect 399308 -22540 399376 -22484
rect 399432 -22540 399518 -22484
rect 399574 -22540 399648 -22484
rect 399308 -22626 399648 -22540
rect 399308 -22682 399376 -22626
rect 399432 -22682 399518 -22626
rect 399574 -22682 399648 -22626
rect 399308 -22768 399648 -22682
rect 399308 -22824 399376 -22768
rect 399432 -22824 399518 -22768
rect 399574 -22824 399648 -22768
rect 399308 -22910 399648 -22824
rect 399308 -22966 399376 -22910
rect 399432 -22966 399518 -22910
rect 399574 -22966 399648 -22910
rect 399308 -23052 399648 -22966
rect 399308 -23108 399376 -23052
rect 399432 -23108 399518 -23052
rect 399574 -23108 399648 -23052
rect 399308 -23194 399648 -23108
rect 399308 -23250 399376 -23194
rect 399432 -23250 399518 -23194
rect 399574 -23250 399648 -23194
rect 399308 -23336 399648 -23250
rect 399308 -23392 399376 -23336
rect 399432 -23392 399518 -23336
rect 399574 -23392 399648 -23336
rect 399308 -23478 399648 -23392
rect 399308 -23534 399376 -23478
rect 399432 -23534 399518 -23478
rect 399574 -23534 399648 -23478
rect 399308 -23620 399648 -23534
rect 399308 -23676 399376 -23620
rect 399432 -23676 399518 -23620
rect 399574 -23676 399648 -23620
rect 399308 -23762 399648 -23676
rect 399308 -23818 399376 -23762
rect 399432 -23818 399518 -23762
rect 399574 -23818 399648 -23762
rect 399308 -23904 399648 -23818
rect 399308 -23960 399376 -23904
rect 399432 -23960 399518 -23904
rect 399574 -23960 399648 -23904
rect 399308 -24046 399648 -23960
rect 399308 -24102 399376 -24046
rect 399432 -24102 399518 -24046
rect 399574 -24102 399648 -24046
rect 399308 -24188 399648 -24102
rect 399308 -24244 399376 -24188
rect 399432 -24244 399518 -24188
rect 399574 -24244 399648 -24188
rect 399308 -24330 399648 -24244
rect 399308 -24386 399376 -24330
rect 399432 -24386 399518 -24330
rect 399574 -24386 399648 -24330
rect 399308 -24472 399648 -24386
rect 399308 -24528 399376 -24472
rect 399432 -24528 399518 -24472
rect 399574 -24528 399648 -24472
rect 399308 -24614 399648 -24528
rect 399308 -24670 399376 -24614
rect 399432 -24670 399518 -24614
rect 399574 -24670 399648 -24614
rect 399308 -24756 399648 -24670
rect 399308 -24812 399376 -24756
rect 399432 -24812 399518 -24756
rect 399574 -24812 399648 -24756
rect 399308 -24898 399648 -24812
rect 399308 -24954 399376 -24898
rect 399432 -24954 399518 -24898
rect 399574 -24954 399648 -24898
rect 399308 -25040 399648 -24954
rect 399308 -25096 399376 -25040
rect 399432 -25096 399518 -25040
rect 399574 -25096 399648 -25040
rect 399308 -25182 399648 -25096
rect 399308 -25238 399376 -25182
rect 399432 -25238 399518 -25182
rect 399574 -25238 399648 -25182
rect 399308 -25324 399648 -25238
rect 399308 -25380 399376 -25324
rect 399432 -25380 399518 -25324
rect 399574 -25380 399648 -25324
rect 399308 -25466 399648 -25380
rect 399308 -25522 399376 -25466
rect 399432 -25522 399518 -25466
rect 399574 -25522 399648 -25466
rect 399308 -25590 399648 -25522
rect 399708 -13680 400048 -13590
rect 399708 -13736 399776 -13680
rect 399832 -13736 399918 -13680
rect 399974 -13736 400048 -13680
rect 399708 -13822 400048 -13736
rect 399708 -13878 399776 -13822
rect 399832 -13878 399918 -13822
rect 399974 -13878 400048 -13822
rect 399708 -13964 400048 -13878
rect 399708 -14020 399776 -13964
rect 399832 -14020 399918 -13964
rect 399974 -14020 400048 -13964
rect 399708 -14106 400048 -14020
rect 399708 -14162 399776 -14106
rect 399832 -14162 399918 -14106
rect 399974 -14162 400048 -14106
rect 399708 -14248 400048 -14162
rect 399708 -14304 399776 -14248
rect 399832 -14304 399918 -14248
rect 399974 -14304 400048 -14248
rect 399708 -14390 400048 -14304
rect 399708 -14446 399776 -14390
rect 399832 -14446 399918 -14390
rect 399974 -14446 400048 -14390
rect 399708 -14532 400048 -14446
rect 399708 -14588 399776 -14532
rect 399832 -14588 399918 -14532
rect 399974 -14588 400048 -14532
rect 399708 -14674 400048 -14588
rect 399708 -14730 399776 -14674
rect 399832 -14730 399918 -14674
rect 399974 -14730 400048 -14674
rect 399708 -14816 400048 -14730
rect 399708 -14872 399776 -14816
rect 399832 -14872 399918 -14816
rect 399974 -14872 400048 -14816
rect 399708 -14958 400048 -14872
rect 399708 -15014 399776 -14958
rect 399832 -15014 399918 -14958
rect 399974 -15014 400048 -14958
rect 399708 -15100 400048 -15014
rect 399708 -15156 399776 -15100
rect 399832 -15156 399918 -15100
rect 399974 -15156 400048 -15100
rect 399708 -15242 400048 -15156
rect 399708 -15298 399776 -15242
rect 399832 -15298 399918 -15242
rect 399974 -15298 400048 -15242
rect 399708 -15384 400048 -15298
rect 399708 -15440 399776 -15384
rect 399832 -15440 399918 -15384
rect 399974 -15440 400048 -15384
rect 399708 -15526 400048 -15440
rect 399708 -15582 399776 -15526
rect 399832 -15582 399918 -15526
rect 399974 -15582 400048 -15526
rect 399708 -15668 400048 -15582
rect 399708 -15724 399776 -15668
rect 399832 -15724 399918 -15668
rect 399974 -15724 400048 -15668
rect 399708 -15810 400048 -15724
rect 399708 -15866 399776 -15810
rect 399832 -15866 399918 -15810
rect 399974 -15866 400048 -15810
rect 399708 -15952 400048 -15866
rect 399708 -16008 399776 -15952
rect 399832 -16008 399918 -15952
rect 399974 -16008 400048 -15952
rect 399708 -16094 400048 -16008
rect 399708 -16150 399776 -16094
rect 399832 -16150 399918 -16094
rect 399974 -16150 400048 -16094
rect 399708 -16236 400048 -16150
rect 399708 -16292 399776 -16236
rect 399832 -16292 399918 -16236
rect 399974 -16292 400048 -16236
rect 399708 -16378 400048 -16292
rect 399708 -16434 399776 -16378
rect 399832 -16434 399918 -16378
rect 399974 -16434 400048 -16378
rect 399708 -16520 400048 -16434
rect 399708 -16576 399776 -16520
rect 399832 -16576 399918 -16520
rect 399974 -16576 400048 -16520
rect 399708 -16662 400048 -16576
rect 399708 -16718 399776 -16662
rect 399832 -16718 399918 -16662
rect 399974 -16718 400048 -16662
rect 399708 -16804 400048 -16718
rect 399708 -16860 399776 -16804
rect 399832 -16860 399918 -16804
rect 399974 -16860 400048 -16804
rect 399708 -16946 400048 -16860
rect 399708 -17002 399776 -16946
rect 399832 -17002 399918 -16946
rect 399974 -17002 400048 -16946
rect 399708 -17088 400048 -17002
rect 399708 -17144 399776 -17088
rect 399832 -17144 399918 -17088
rect 399974 -17144 400048 -17088
rect 399708 -17230 400048 -17144
rect 399708 -17286 399776 -17230
rect 399832 -17286 399918 -17230
rect 399974 -17286 400048 -17230
rect 399708 -17372 400048 -17286
rect 399708 -17428 399776 -17372
rect 399832 -17428 399918 -17372
rect 399974 -17428 400048 -17372
rect 399708 -17514 400048 -17428
rect 399708 -17570 399776 -17514
rect 399832 -17570 399918 -17514
rect 399974 -17570 400048 -17514
rect 399708 -17656 400048 -17570
rect 399708 -17712 399776 -17656
rect 399832 -17712 399918 -17656
rect 399974 -17712 400048 -17656
rect 399708 -17798 400048 -17712
rect 399708 -17854 399776 -17798
rect 399832 -17854 399918 -17798
rect 399974 -17854 400048 -17798
rect 399708 -17940 400048 -17854
rect 399708 -17996 399776 -17940
rect 399832 -17996 399918 -17940
rect 399974 -17996 400048 -17940
rect 399708 -18082 400048 -17996
rect 399708 -18138 399776 -18082
rect 399832 -18138 399918 -18082
rect 399974 -18138 400048 -18082
rect 399708 -18224 400048 -18138
rect 399708 -18280 399776 -18224
rect 399832 -18280 399918 -18224
rect 399974 -18280 400048 -18224
rect 399708 -18366 400048 -18280
rect 399708 -18422 399776 -18366
rect 399832 -18422 399918 -18366
rect 399974 -18422 400048 -18366
rect 399708 -18508 400048 -18422
rect 399708 -18564 399776 -18508
rect 399832 -18564 399918 -18508
rect 399974 -18564 400048 -18508
rect 399708 -18650 400048 -18564
rect 399708 -18706 399776 -18650
rect 399832 -18706 399918 -18650
rect 399974 -18706 400048 -18650
rect 399708 -18792 400048 -18706
rect 399708 -18848 399776 -18792
rect 399832 -18848 399918 -18792
rect 399974 -18848 400048 -18792
rect 399708 -18934 400048 -18848
rect 399708 -18990 399776 -18934
rect 399832 -18990 399918 -18934
rect 399974 -18990 400048 -18934
rect 399708 -19076 400048 -18990
rect 399708 -19132 399776 -19076
rect 399832 -19132 399918 -19076
rect 399974 -19132 400048 -19076
rect 399708 -19218 400048 -19132
rect 399708 -19274 399776 -19218
rect 399832 -19274 399918 -19218
rect 399974 -19274 400048 -19218
rect 399708 -19360 400048 -19274
rect 399708 -19416 399776 -19360
rect 399832 -19416 399918 -19360
rect 399974 -19416 400048 -19360
rect 399708 -19502 400048 -19416
rect 399708 -19558 399776 -19502
rect 399832 -19558 399918 -19502
rect 399974 -19558 400048 -19502
rect 399708 -19644 400048 -19558
rect 399708 -19700 399776 -19644
rect 399832 -19700 399918 -19644
rect 399974 -19700 400048 -19644
rect 399708 -19786 400048 -19700
rect 399708 -19842 399776 -19786
rect 399832 -19842 399918 -19786
rect 399974 -19842 400048 -19786
rect 399708 -19928 400048 -19842
rect 399708 -19984 399776 -19928
rect 399832 -19984 399918 -19928
rect 399974 -19984 400048 -19928
rect 399708 -20070 400048 -19984
rect 399708 -20126 399776 -20070
rect 399832 -20126 399918 -20070
rect 399974 -20126 400048 -20070
rect 399708 -20212 400048 -20126
rect 399708 -20268 399776 -20212
rect 399832 -20268 399918 -20212
rect 399974 -20268 400048 -20212
rect 399708 -20354 400048 -20268
rect 399708 -20410 399776 -20354
rect 399832 -20410 399918 -20354
rect 399974 -20410 400048 -20354
rect 399708 -20496 400048 -20410
rect 399708 -20552 399776 -20496
rect 399832 -20552 399918 -20496
rect 399974 -20552 400048 -20496
rect 399708 -20638 400048 -20552
rect 399708 -20694 399776 -20638
rect 399832 -20694 399918 -20638
rect 399974 -20694 400048 -20638
rect 399708 -20780 400048 -20694
rect 399708 -20836 399776 -20780
rect 399832 -20836 399918 -20780
rect 399974 -20836 400048 -20780
rect 399708 -20922 400048 -20836
rect 399708 -20978 399776 -20922
rect 399832 -20978 399918 -20922
rect 399974 -20978 400048 -20922
rect 399708 -21064 400048 -20978
rect 399708 -21120 399776 -21064
rect 399832 -21120 399918 -21064
rect 399974 -21120 400048 -21064
rect 399708 -21206 400048 -21120
rect 399708 -21262 399776 -21206
rect 399832 -21262 399918 -21206
rect 399974 -21262 400048 -21206
rect 399708 -21348 400048 -21262
rect 399708 -21404 399776 -21348
rect 399832 -21404 399918 -21348
rect 399974 -21404 400048 -21348
rect 399708 -21490 400048 -21404
rect 399708 -21546 399776 -21490
rect 399832 -21546 399918 -21490
rect 399974 -21546 400048 -21490
rect 399708 -21632 400048 -21546
rect 399708 -21688 399776 -21632
rect 399832 -21688 399918 -21632
rect 399974 -21688 400048 -21632
rect 399708 -21774 400048 -21688
rect 399708 -21830 399776 -21774
rect 399832 -21830 399918 -21774
rect 399974 -21830 400048 -21774
rect 399708 -21916 400048 -21830
rect 399708 -21972 399776 -21916
rect 399832 -21972 399918 -21916
rect 399974 -21972 400048 -21916
rect 399708 -22058 400048 -21972
rect 399708 -22114 399776 -22058
rect 399832 -22114 399918 -22058
rect 399974 -22114 400048 -22058
rect 399708 -22200 400048 -22114
rect 399708 -22256 399776 -22200
rect 399832 -22256 399918 -22200
rect 399974 -22256 400048 -22200
rect 399708 -22342 400048 -22256
rect 399708 -22398 399776 -22342
rect 399832 -22398 399918 -22342
rect 399974 -22398 400048 -22342
rect 399708 -22484 400048 -22398
rect 399708 -22540 399776 -22484
rect 399832 -22540 399918 -22484
rect 399974 -22540 400048 -22484
rect 399708 -22626 400048 -22540
rect 399708 -22682 399776 -22626
rect 399832 -22682 399918 -22626
rect 399974 -22682 400048 -22626
rect 399708 -22768 400048 -22682
rect 399708 -22824 399776 -22768
rect 399832 -22824 399918 -22768
rect 399974 -22824 400048 -22768
rect 399708 -22910 400048 -22824
rect 399708 -22966 399776 -22910
rect 399832 -22966 399918 -22910
rect 399974 -22966 400048 -22910
rect 399708 -23052 400048 -22966
rect 399708 -23108 399776 -23052
rect 399832 -23108 399918 -23052
rect 399974 -23108 400048 -23052
rect 399708 -23194 400048 -23108
rect 399708 -23250 399776 -23194
rect 399832 -23250 399918 -23194
rect 399974 -23250 400048 -23194
rect 399708 -23336 400048 -23250
rect 399708 -23392 399776 -23336
rect 399832 -23392 399918 -23336
rect 399974 -23392 400048 -23336
rect 399708 -23478 400048 -23392
rect 399708 -23534 399776 -23478
rect 399832 -23534 399918 -23478
rect 399974 -23534 400048 -23478
rect 399708 -23620 400048 -23534
rect 399708 -23676 399776 -23620
rect 399832 -23676 399918 -23620
rect 399974 -23676 400048 -23620
rect 399708 -23762 400048 -23676
rect 399708 -23818 399776 -23762
rect 399832 -23818 399918 -23762
rect 399974 -23818 400048 -23762
rect 399708 -23904 400048 -23818
rect 399708 -23960 399776 -23904
rect 399832 -23960 399918 -23904
rect 399974 -23960 400048 -23904
rect 399708 -24046 400048 -23960
rect 399708 -24102 399776 -24046
rect 399832 -24102 399918 -24046
rect 399974 -24102 400048 -24046
rect 399708 -24188 400048 -24102
rect 399708 -24244 399776 -24188
rect 399832 -24244 399918 -24188
rect 399974 -24244 400048 -24188
rect 399708 -24330 400048 -24244
rect 399708 -24386 399776 -24330
rect 399832 -24386 399918 -24330
rect 399974 -24386 400048 -24330
rect 399708 -24472 400048 -24386
rect 399708 -24528 399776 -24472
rect 399832 -24528 399918 -24472
rect 399974 -24528 400048 -24472
rect 399708 -24614 400048 -24528
rect 399708 -24670 399776 -24614
rect 399832 -24670 399918 -24614
rect 399974 -24670 400048 -24614
rect 399708 -24756 400048 -24670
rect 399708 -24812 399776 -24756
rect 399832 -24812 399918 -24756
rect 399974 -24812 400048 -24756
rect 399708 -24898 400048 -24812
rect 399708 -24954 399776 -24898
rect 399832 -24954 399918 -24898
rect 399974 -24954 400048 -24898
rect 399708 -25040 400048 -24954
rect 399708 -25096 399776 -25040
rect 399832 -25096 399918 -25040
rect 399974 -25096 400048 -25040
rect 399708 -25182 400048 -25096
rect 399708 -25238 399776 -25182
rect 399832 -25238 399918 -25182
rect 399974 -25238 400048 -25182
rect 399708 -25324 400048 -25238
rect 399708 -25380 399776 -25324
rect 399832 -25380 399918 -25324
rect 399974 -25380 400048 -25324
rect 399708 -25466 400048 -25380
rect 399708 -25522 399776 -25466
rect 399832 -25522 399918 -25466
rect 399974 -25522 400048 -25466
rect 399708 -25590 400048 -25522
rect 400108 -13680 400448 -13590
rect 400108 -13736 400181 -13680
rect 400237 -13736 400323 -13680
rect 400379 -13736 400448 -13680
rect 400108 -13822 400448 -13736
rect 400108 -13878 400181 -13822
rect 400237 -13878 400323 -13822
rect 400379 -13878 400448 -13822
rect 400108 -13964 400448 -13878
rect 400108 -14020 400181 -13964
rect 400237 -14020 400323 -13964
rect 400379 -14020 400448 -13964
rect 400108 -14106 400448 -14020
rect 400108 -14162 400181 -14106
rect 400237 -14162 400323 -14106
rect 400379 -14162 400448 -14106
rect 400108 -14248 400448 -14162
rect 400108 -14304 400181 -14248
rect 400237 -14304 400323 -14248
rect 400379 -14304 400448 -14248
rect 400108 -14390 400448 -14304
rect 400108 -14446 400181 -14390
rect 400237 -14446 400323 -14390
rect 400379 -14446 400448 -14390
rect 400108 -14532 400448 -14446
rect 400108 -14588 400181 -14532
rect 400237 -14588 400323 -14532
rect 400379 -14588 400448 -14532
rect 400108 -14674 400448 -14588
rect 400108 -14730 400181 -14674
rect 400237 -14730 400323 -14674
rect 400379 -14730 400448 -14674
rect 400108 -14816 400448 -14730
rect 400108 -14872 400181 -14816
rect 400237 -14872 400323 -14816
rect 400379 -14872 400448 -14816
rect 400108 -14958 400448 -14872
rect 400108 -15014 400181 -14958
rect 400237 -15014 400323 -14958
rect 400379 -15014 400448 -14958
rect 400108 -15100 400448 -15014
rect 400108 -15156 400181 -15100
rect 400237 -15156 400323 -15100
rect 400379 -15156 400448 -15100
rect 400108 -15242 400448 -15156
rect 400108 -15298 400181 -15242
rect 400237 -15298 400323 -15242
rect 400379 -15298 400448 -15242
rect 400108 -15384 400448 -15298
rect 400108 -15440 400181 -15384
rect 400237 -15440 400323 -15384
rect 400379 -15440 400448 -15384
rect 400108 -15526 400448 -15440
rect 400108 -15582 400181 -15526
rect 400237 -15582 400323 -15526
rect 400379 -15582 400448 -15526
rect 400108 -15668 400448 -15582
rect 400108 -15724 400181 -15668
rect 400237 -15724 400323 -15668
rect 400379 -15724 400448 -15668
rect 400108 -15810 400448 -15724
rect 400108 -15866 400181 -15810
rect 400237 -15866 400323 -15810
rect 400379 -15866 400448 -15810
rect 400108 -15952 400448 -15866
rect 400108 -16008 400181 -15952
rect 400237 -16008 400323 -15952
rect 400379 -16008 400448 -15952
rect 400108 -16094 400448 -16008
rect 400108 -16150 400181 -16094
rect 400237 -16150 400323 -16094
rect 400379 -16150 400448 -16094
rect 400108 -16236 400448 -16150
rect 400108 -16292 400181 -16236
rect 400237 -16292 400323 -16236
rect 400379 -16292 400448 -16236
rect 400108 -16378 400448 -16292
rect 400108 -16434 400181 -16378
rect 400237 -16434 400323 -16378
rect 400379 -16434 400448 -16378
rect 400108 -16520 400448 -16434
rect 400108 -16576 400181 -16520
rect 400237 -16576 400323 -16520
rect 400379 -16576 400448 -16520
rect 400108 -16662 400448 -16576
rect 400108 -16718 400181 -16662
rect 400237 -16718 400323 -16662
rect 400379 -16718 400448 -16662
rect 400108 -16804 400448 -16718
rect 400108 -16860 400181 -16804
rect 400237 -16860 400323 -16804
rect 400379 -16860 400448 -16804
rect 400108 -16946 400448 -16860
rect 400108 -17002 400181 -16946
rect 400237 -17002 400323 -16946
rect 400379 -17002 400448 -16946
rect 400108 -17088 400448 -17002
rect 400108 -17144 400181 -17088
rect 400237 -17144 400323 -17088
rect 400379 -17144 400448 -17088
rect 400108 -17230 400448 -17144
rect 400108 -17286 400181 -17230
rect 400237 -17286 400323 -17230
rect 400379 -17286 400448 -17230
rect 400108 -17372 400448 -17286
rect 400108 -17428 400181 -17372
rect 400237 -17428 400323 -17372
rect 400379 -17428 400448 -17372
rect 400108 -17514 400448 -17428
rect 400108 -17570 400181 -17514
rect 400237 -17570 400323 -17514
rect 400379 -17570 400448 -17514
rect 400108 -17656 400448 -17570
rect 400108 -17712 400181 -17656
rect 400237 -17712 400323 -17656
rect 400379 -17712 400448 -17656
rect 400108 -17798 400448 -17712
rect 400108 -17854 400181 -17798
rect 400237 -17854 400323 -17798
rect 400379 -17854 400448 -17798
rect 400108 -17940 400448 -17854
rect 400108 -17996 400181 -17940
rect 400237 -17996 400323 -17940
rect 400379 -17996 400448 -17940
rect 400108 -18082 400448 -17996
rect 400108 -18138 400181 -18082
rect 400237 -18138 400323 -18082
rect 400379 -18138 400448 -18082
rect 400108 -18224 400448 -18138
rect 400108 -18280 400181 -18224
rect 400237 -18280 400323 -18224
rect 400379 -18280 400448 -18224
rect 400108 -18366 400448 -18280
rect 400108 -18422 400181 -18366
rect 400237 -18422 400323 -18366
rect 400379 -18422 400448 -18366
rect 400108 -18508 400448 -18422
rect 400108 -18564 400181 -18508
rect 400237 -18564 400323 -18508
rect 400379 -18564 400448 -18508
rect 400108 -18650 400448 -18564
rect 400108 -18706 400181 -18650
rect 400237 -18706 400323 -18650
rect 400379 -18706 400448 -18650
rect 400108 -18792 400448 -18706
rect 400108 -18848 400181 -18792
rect 400237 -18848 400323 -18792
rect 400379 -18848 400448 -18792
rect 400108 -18934 400448 -18848
rect 400108 -18990 400181 -18934
rect 400237 -18990 400323 -18934
rect 400379 -18990 400448 -18934
rect 400108 -19076 400448 -18990
rect 400108 -19132 400181 -19076
rect 400237 -19132 400323 -19076
rect 400379 -19132 400448 -19076
rect 400108 -19218 400448 -19132
rect 400108 -19274 400181 -19218
rect 400237 -19274 400323 -19218
rect 400379 -19274 400448 -19218
rect 400108 -19360 400448 -19274
rect 400108 -19416 400181 -19360
rect 400237 -19416 400323 -19360
rect 400379 -19416 400448 -19360
rect 400108 -19502 400448 -19416
rect 400108 -19558 400181 -19502
rect 400237 -19558 400323 -19502
rect 400379 -19558 400448 -19502
rect 400108 -19644 400448 -19558
rect 400108 -19700 400181 -19644
rect 400237 -19700 400323 -19644
rect 400379 -19700 400448 -19644
rect 400108 -19786 400448 -19700
rect 400108 -19842 400181 -19786
rect 400237 -19842 400323 -19786
rect 400379 -19842 400448 -19786
rect 400108 -19928 400448 -19842
rect 400108 -19984 400181 -19928
rect 400237 -19984 400323 -19928
rect 400379 -19984 400448 -19928
rect 400108 -20070 400448 -19984
rect 400108 -20126 400181 -20070
rect 400237 -20126 400323 -20070
rect 400379 -20126 400448 -20070
rect 400108 -20212 400448 -20126
rect 400108 -20268 400181 -20212
rect 400237 -20268 400323 -20212
rect 400379 -20268 400448 -20212
rect 400108 -20354 400448 -20268
rect 400108 -20410 400181 -20354
rect 400237 -20410 400323 -20354
rect 400379 -20410 400448 -20354
rect 400108 -20496 400448 -20410
rect 400108 -20552 400181 -20496
rect 400237 -20552 400323 -20496
rect 400379 -20552 400448 -20496
rect 400108 -20638 400448 -20552
rect 400108 -20694 400181 -20638
rect 400237 -20694 400323 -20638
rect 400379 -20694 400448 -20638
rect 400108 -20780 400448 -20694
rect 400108 -20836 400181 -20780
rect 400237 -20836 400323 -20780
rect 400379 -20836 400448 -20780
rect 400108 -20922 400448 -20836
rect 400108 -20978 400181 -20922
rect 400237 -20978 400323 -20922
rect 400379 -20978 400448 -20922
rect 400108 -21064 400448 -20978
rect 400108 -21120 400181 -21064
rect 400237 -21120 400323 -21064
rect 400379 -21120 400448 -21064
rect 400108 -21206 400448 -21120
rect 400108 -21262 400181 -21206
rect 400237 -21262 400323 -21206
rect 400379 -21262 400448 -21206
rect 400108 -21348 400448 -21262
rect 400108 -21404 400181 -21348
rect 400237 -21404 400323 -21348
rect 400379 -21404 400448 -21348
rect 400108 -21490 400448 -21404
rect 400108 -21546 400181 -21490
rect 400237 -21546 400323 -21490
rect 400379 -21546 400448 -21490
rect 400108 -21632 400448 -21546
rect 400108 -21688 400181 -21632
rect 400237 -21688 400323 -21632
rect 400379 -21688 400448 -21632
rect 400108 -21774 400448 -21688
rect 400108 -21830 400181 -21774
rect 400237 -21830 400323 -21774
rect 400379 -21830 400448 -21774
rect 400108 -21916 400448 -21830
rect 400108 -21972 400181 -21916
rect 400237 -21972 400323 -21916
rect 400379 -21972 400448 -21916
rect 400108 -22058 400448 -21972
rect 400108 -22114 400181 -22058
rect 400237 -22114 400323 -22058
rect 400379 -22114 400448 -22058
rect 400108 -22200 400448 -22114
rect 400108 -22256 400181 -22200
rect 400237 -22256 400323 -22200
rect 400379 -22256 400448 -22200
rect 400108 -22342 400448 -22256
rect 400108 -22398 400181 -22342
rect 400237 -22398 400323 -22342
rect 400379 -22398 400448 -22342
rect 400108 -22484 400448 -22398
rect 400108 -22540 400181 -22484
rect 400237 -22540 400323 -22484
rect 400379 -22540 400448 -22484
rect 400108 -22626 400448 -22540
rect 400108 -22682 400181 -22626
rect 400237 -22682 400323 -22626
rect 400379 -22682 400448 -22626
rect 400108 -22768 400448 -22682
rect 400108 -22824 400181 -22768
rect 400237 -22824 400323 -22768
rect 400379 -22824 400448 -22768
rect 400108 -22910 400448 -22824
rect 400108 -22966 400181 -22910
rect 400237 -22966 400323 -22910
rect 400379 -22966 400448 -22910
rect 400108 -23052 400448 -22966
rect 400108 -23108 400181 -23052
rect 400237 -23108 400323 -23052
rect 400379 -23108 400448 -23052
rect 400108 -23194 400448 -23108
rect 400108 -23250 400181 -23194
rect 400237 -23250 400323 -23194
rect 400379 -23250 400448 -23194
rect 400108 -23336 400448 -23250
rect 400108 -23392 400181 -23336
rect 400237 -23392 400323 -23336
rect 400379 -23392 400448 -23336
rect 400108 -23478 400448 -23392
rect 400108 -23534 400181 -23478
rect 400237 -23534 400323 -23478
rect 400379 -23534 400448 -23478
rect 400108 -23620 400448 -23534
rect 400108 -23676 400181 -23620
rect 400237 -23676 400323 -23620
rect 400379 -23676 400448 -23620
rect 400108 -23762 400448 -23676
rect 400108 -23818 400181 -23762
rect 400237 -23818 400323 -23762
rect 400379 -23818 400448 -23762
rect 400108 -23904 400448 -23818
rect 400108 -23960 400181 -23904
rect 400237 -23960 400323 -23904
rect 400379 -23960 400448 -23904
rect 400108 -24046 400448 -23960
rect 400108 -24102 400181 -24046
rect 400237 -24102 400323 -24046
rect 400379 -24102 400448 -24046
rect 400108 -24188 400448 -24102
rect 400108 -24244 400181 -24188
rect 400237 -24244 400323 -24188
rect 400379 -24244 400448 -24188
rect 400108 -24330 400448 -24244
rect 400108 -24386 400181 -24330
rect 400237 -24386 400323 -24330
rect 400379 -24386 400448 -24330
rect 400108 -24472 400448 -24386
rect 400108 -24528 400181 -24472
rect 400237 -24528 400323 -24472
rect 400379 -24528 400448 -24472
rect 400108 -24614 400448 -24528
rect 400108 -24670 400181 -24614
rect 400237 -24670 400323 -24614
rect 400379 -24670 400448 -24614
rect 400108 -24756 400448 -24670
rect 400108 -24812 400181 -24756
rect 400237 -24812 400323 -24756
rect 400379 -24812 400448 -24756
rect 400108 -24898 400448 -24812
rect 400108 -24954 400181 -24898
rect 400237 -24954 400323 -24898
rect 400379 -24954 400448 -24898
rect 400108 -25040 400448 -24954
rect 400108 -25096 400181 -25040
rect 400237 -25096 400323 -25040
rect 400379 -25096 400448 -25040
rect 400108 -25182 400448 -25096
rect 400108 -25238 400181 -25182
rect 400237 -25238 400323 -25182
rect 400379 -25238 400448 -25182
rect 400108 -25324 400448 -25238
rect 400108 -25380 400181 -25324
rect 400237 -25380 400323 -25324
rect 400379 -25380 400448 -25324
rect 400108 -25466 400448 -25380
rect 400108 -25522 400181 -25466
rect 400237 -25522 400323 -25466
rect 400379 -25522 400448 -25466
rect 400108 -25590 400448 -25522
rect 400640 -13632 401440 -13590
rect 400640 -13688 400766 -13632
rect 400822 -13688 400890 -13632
rect 400946 -13688 401014 -13632
rect 401070 -13688 401138 -13632
rect 401194 -13688 401262 -13632
rect 401318 -13688 401440 -13632
rect 400640 -13756 401440 -13688
rect 400640 -13812 400766 -13756
rect 400822 -13812 400890 -13756
rect 400946 -13812 401014 -13756
rect 401070 -13812 401138 -13756
rect 401194 -13812 401262 -13756
rect 401318 -13812 401440 -13756
rect 400640 -13880 401440 -13812
rect 400640 -13936 400766 -13880
rect 400822 -13936 400890 -13880
rect 400946 -13936 401014 -13880
rect 401070 -13936 401138 -13880
rect 401194 -13936 401262 -13880
rect 401318 -13936 401440 -13880
rect 400640 -14004 401440 -13936
rect 400640 -14060 400766 -14004
rect 400822 -14060 400890 -14004
rect 400946 -14060 401014 -14004
rect 401070 -14060 401138 -14004
rect 401194 -14060 401262 -14004
rect 401318 -14060 401440 -14004
rect 400640 -14128 401440 -14060
rect 400640 -14184 400766 -14128
rect 400822 -14184 400890 -14128
rect 400946 -14184 401014 -14128
rect 401070 -14184 401138 -14128
rect 401194 -14184 401262 -14128
rect 401318 -14184 401440 -14128
rect 400640 -14252 401440 -14184
rect 400640 -14308 400766 -14252
rect 400822 -14308 400890 -14252
rect 400946 -14308 401014 -14252
rect 401070 -14308 401138 -14252
rect 401194 -14308 401262 -14252
rect 401318 -14308 401440 -14252
rect 400640 -14376 401440 -14308
rect 400640 -14432 400766 -14376
rect 400822 -14432 400890 -14376
rect 400946 -14432 401014 -14376
rect 401070 -14432 401138 -14376
rect 401194 -14432 401262 -14376
rect 401318 -14432 401440 -14376
rect 400640 -14500 401440 -14432
rect 400640 -14556 400766 -14500
rect 400822 -14556 400890 -14500
rect 400946 -14556 401014 -14500
rect 401070 -14556 401138 -14500
rect 401194 -14556 401262 -14500
rect 401318 -14556 401440 -14500
rect 400640 -14624 401440 -14556
rect 400640 -14680 400766 -14624
rect 400822 -14680 400890 -14624
rect 400946 -14680 401014 -14624
rect 401070 -14680 401138 -14624
rect 401194 -14680 401262 -14624
rect 401318 -14680 401440 -14624
rect 400640 -14748 401440 -14680
rect 400640 -14804 400766 -14748
rect 400822 -14804 400890 -14748
rect 400946 -14804 401014 -14748
rect 401070 -14804 401138 -14748
rect 401194 -14804 401262 -14748
rect 401318 -14804 401440 -14748
rect 400640 -14872 401440 -14804
rect 400640 -14928 400766 -14872
rect 400822 -14928 400890 -14872
rect 400946 -14928 401014 -14872
rect 401070 -14928 401138 -14872
rect 401194 -14928 401262 -14872
rect 401318 -14928 401440 -14872
rect 400640 -14996 401440 -14928
rect 400640 -15052 400766 -14996
rect 400822 -15052 400890 -14996
rect 400946 -15052 401014 -14996
rect 401070 -15052 401138 -14996
rect 401194 -15052 401262 -14996
rect 401318 -15052 401440 -14996
rect 400640 -15120 401440 -15052
rect 400640 -15176 400766 -15120
rect 400822 -15176 400890 -15120
rect 400946 -15176 401014 -15120
rect 401070 -15176 401138 -15120
rect 401194 -15176 401262 -15120
rect 401318 -15176 401440 -15120
rect 400640 -15244 401440 -15176
rect 400640 -15300 400766 -15244
rect 400822 -15300 400890 -15244
rect 400946 -15300 401014 -15244
rect 401070 -15300 401138 -15244
rect 401194 -15300 401262 -15244
rect 401318 -15300 401440 -15244
rect 400640 -15368 401440 -15300
rect 400640 -15424 400766 -15368
rect 400822 -15424 400890 -15368
rect 400946 -15424 401014 -15368
rect 401070 -15424 401138 -15368
rect 401194 -15424 401262 -15368
rect 401318 -15424 401440 -15368
rect 400640 -15492 401440 -15424
rect 400640 -15548 400766 -15492
rect 400822 -15548 400890 -15492
rect 400946 -15548 401014 -15492
rect 401070 -15548 401138 -15492
rect 401194 -15548 401262 -15492
rect 401318 -15548 401440 -15492
rect 400640 -15616 401440 -15548
rect 400640 -15672 400766 -15616
rect 400822 -15672 400890 -15616
rect 400946 -15672 401014 -15616
rect 401070 -15672 401138 -15616
rect 401194 -15672 401262 -15616
rect 401318 -15672 401440 -15616
rect 400640 -15740 401440 -15672
rect 400640 -15796 400766 -15740
rect 400822 -15796 400890 -15740
rect 400946 -15796 401014 -15740
rect 401070 -15796 401138 -15740
rect 401194 -15796 401262 -15740
rect 401318 -15796 401440 -15740
rect 400640 -15864 401440 -15796
rect 400640 -15920 400766 -15864
rect 400822 -15920 400890 -15864
rect 400946 -15920 401014 -15864
rect 401070 -15920 401138 -15864
rect 401194 -15920 401262 -15864
rect 401318 -15920 401440 -15864
rect 400640 -15988 401440 -15920
rect 400640 -16044 400766 -15988
rect 400822 -16044 400890 -15988
rect 400946 -16044 401014 -15988
rect 401070 -16044 401138 -15988
rect 401194 -16044 401262 -15988
rect 401318 -16044 401440 -15988
rect 400640 -16112 401440 -16044
rect 400640 -16168 400766 -16112
rect 400822 -16168 400890 -16112
rect 400946 -16168 401014 -16112
rect 401070 -16168 401138 -16112
rect 401194 -16168 401262 -16112
rect 401318 -16168 401440 -16112
rect 400640 -16236 401440 -16168
rect 400640 -16292 400766 -16236
rect 400822 -16292 400890 -16236
rect 400946 -16292 401014 -16236
rect 401070 -16292 401138 -16236
rect 401194 -16292 401262 -16236
rect 401318 -16292 401440 -16236
rect 400640 -16360 401440 -16292
rect 400640 -16416 400766 -16360
rect 400822 -16416 400890 -16360
rect 400946 -16416 401014 -16360
rect 401070 -16416 401138 -16360
rect 401194 -16416 401262 -16360
rect 401318 -16416 401440 -16360
rect 400640 -16484 401440 -16416
rect 400640 -16540 400766 -16484
rect 400822 -16540 400890 -16484
rect 400946 -16540 401014 -16484
rect 401070 -16540 401138 -16484
rect 401194 -16540 401262 -16484
rect 401318 -16540 401440 -16484
rect 400640 -16608 401440 -16540
rect 400640 -16664 400766 -16608
rect 400822 -16664 400890 -16608
rect 400946 -16664 401014 -16608
rect 401070 -16664 401138 -16608
rect 401194 -16664 401262 -16608
rect 401318 -16664 401440 -16608
rect 400640 -16732 401440 -16664
rect 400640 -16788 400766 -16732
rect 400822 -16788 400890 -16732
rect 400946 -16788 401014 -16732
rect 401070 -16788 401138 -16732
rect 401194 -16788 401262 -16732
rect 401318 -16788 401440 -16732
rect 400640 -16856 401440 -16788
rect 400640 -16912 400766 -16856
rect 400822 -16912 400890 -16856
rect 400946 -16912 401014 -16856
rect 401070 -16912 401138 -16856
rect 401194 -16912 401262 -16856
rect 401318 -16912 401440 -16856
rect 400640 -16980 401440 -16912
rect 400640 -17036 400766 -16980
rect 400822 -17036 400890 -16980
rect 400946 -17036 401014 -16980
rect 401070 -17036 401138 -16980
rect 401194 -17036 401262 -16980
rect 401318 -17036 401440 -16980
rect 400640 -17104 401440 -17036
rect 400640 -17160 400766 -17104
rect 400822 -17160 400890 -17104
rect 400946 -17160 401014 -17104
rect 401070 -17160 401138 -17104
rect 401194 -17160 401262 -17104
rect 401318 -17160 401440 -17104
rect 400640 -17228 401440 -17160
rect 400640 -17284 400766 -17228
rect 400822 -17284 400890 -17228
rect 400946 -17284 401014 -17228
rect 401070 -17284 401138 -17228
rect 401194 -17284 401262 -17228
rect 401318 -17284 401440 -17228
rect 400640 -17352 401440 -17284
rect 400640 -17408 400766 -17352
rect 400822 -17408 400890 -17352
rect 400946 -17408 401014 -17352
rect 401070 -17408 401138 -17352
rect 401194 -17408 401262 -17352
rect 401318 -17408 401440 -17352
rect 400640 -17476 401440 -17408
rect 400640 -17532 400766 -17476
rect 400822 -17532 400890 -17476
rect 400946 -17532 401014 -17476
rect 401070 -17532 401138 -17476
rect 401194 -17532 401262 -17476
rect 401318 -17532 401440 -17476
rect 400640 -17600 401440 -17532
rect 400640 -17656 400766 -17600
rect 400822 -17656 400890 -17600
rect 400946 -17656 401014 -17600
rect 401070 -17656 401138 -17600
rect 401194 -17656 401262 -17600
rect 401318 -17656 401440 -17600
rect 400640 -17724 401440 -17656
rect 400640 -17780 400766 -17724
rect 400822 -17780 400890 -17724
rect 400946 -17780 401014 -17724
rect 401070 -17780 401138 -17724
rect 401194 -17780 401262 -17724
rect 401318 -17780 401440 -17724
rect 400640 -17848 401440 -17780
rect 400640 -17904 400766 -17848
rect 400822 -17904 400890 -17848
rect 400946 -17904 401014 -17848
rect 401070 -17904 401138 -17848
rect 401194 -17904 401262 -17848
rect 401318 -17904 401440 -17848
rect 400640 -17972 401440 -17904
rect 400640 -18028 400766 -17972
rect 400822 -18028 400890 -17972
rect 400946 -18028 401014 -17972
rect 401070 -18028 401138 -17972
rect 401194 -18028 401262 -17972
rect 401318 -18028 401440 -17972
rect 400640 -18096 401440 -18028
rect 400640 -18152 400766 -18096
rect 400822 -18152 400890 -18096
rect 400946 -18152 401014 -18096
rect 401070 -18152 401138 -18096
rect 401194 -18152 401262 -18096
rect 401318 -18152 401440 -18096
rect 400640 -18220 401440 -18152
rect 400640 -18276 400766 -18220
rect 400822 -18276 400890 -18220
rect 400946 -18276 401014 -18220
rect 401070 -18276 401138 -18220
rect 401194 -18276 401262 -18220
rect 401318 -18276 401440 -18220
rect 400640 -18344 401440 -18276
rect 400640 -18400 400766 -18344
rect 400822 -18400 400890 -18344
rect 400946 -18400 401014 -18344
rect 401070 -18400 401138 -18344
rect 401194 -18400 401262 -18344
rect 401318 -18400 401440 -18344
rect 400640 -18468 401440 -18400
rect 400640 -18524 400766 -18468
rect 400822 -18524 400890 -18468
rect 400946 -18524 401014 -18468
rect 401070 -18524 401138 -18468
rect 401194 -18524 401262 -18468
rect 401318 -18524 401440 -18468
rect 400640 -18592 401440 -18524
rect 400640 -18648 400766 -18592
rect 400822 -18648 400890 -18592
rect 400946 -18648 401014 -18592
rect 401070 -18648 401138 -18592
rect 401194 -18648 401262 -18592
rect 401318 -18648 401440 -18592
rect 400640 -18716 401440 -18648
rect 400640 -18772 400766 -18716
rect 400822 -18772 400890 -18716
rect 400946 -18772 401014 -18716
rect 401070 -18772 401138 -18716
rect 401194 -18772 401262 -18716
rect 401318 -18772 401440 -18716
rect 400640 -18840 401440 -18772
rect 400640 -18896 400766 -18840
rect 400822 -18896 400890 -18840
rect 400946 -18896 401014 -18840
rect 401070 -18896 401138 -18840
rect 401194 -18896 401262 -18840
rect 401318 -18896 401440 -18840
rect 400640 -18964 401440 -18896
rect 400640 -19020 400766 -18964
rect 400822 -19020 400890 -18964
rect 400946 -19020 401014 -18964
rect 401070 -19020 401138 -18964
rect 401194 -19020 401262 -18964
rect 401318 -19020 401440 -18964
rect 400640 -19088 401440 -19020
rect 400640 -19144 400766 -19088
rect 400822 -19144 400890 -19088
rect 400946 -19144 401014 -19088
rect 401070 -19144 401138 -19088
rect 401194 -19144 401262 -19088
rect 401318 -19144 401440 -19088
rect 400640 -19212 401440 -19144
rect 400640 -19268 400766 -19212
rect 400822 -19268 400890 -19212
rect 400946 -19268 401014 -19212
rect 401070 -19268 401138 -19212
rect 401194 -19268 401262 -19212
rect 401318 -19268 401440 -19212
rect 400640 -19336 401440 -19268
rect 400640 -19392 400766 -19336
rect 400822 -19392 400890 -19336
rect 400946 -19392 401014 -19336
rect 401070 -19392 401138 -19336
rect 401194 -19392 401262 -19336
rect 401318 -19392 401440 -19336
rect 400640 -19460 401440 -19392
rect 400640 -19516 400766 -19460
rect 400822 -19516 400890 -19460
rect 400946 -19516 401014 -19460
rect 401070 -19516 401138 -19460
rect 401194 -19516 401262 -19460
rect 401318 -19516 401440 -19460
rect 400640 -19584 401440 -19516
rect 400640 -19640 400766 -19584
rect 400822 -19640 400890 -19584
rect 400946 -19640 401014 -19584
rect 401070 -19640 401138 -19584
rect 401194 -19640 401262 -19584
rect 401318 -19640 401440 -19584
rect 400640 -19708 401440 -19640
rect 400640 -19764 400766 -19708
rect 400822 -19764 400890 -19708
rect 400946 -19764 401014 -19708
rect 401070 -19764 401138 -19708
rect 401194 -19764 401262 -19708
rect 401318 -19764 401440 -19708
rect 400640 -19832 401440 -19764
rect 400640 -19888 400766 -19832
rect 400822 -19888 400890 -19832
rect 400946 -19888 401014 -19832
rect 401070 -19888 401138 -19832
rect 401194 -19888 401262 -19832
rect 401318 -19888 401440 -19832
rect 400640 -19956 401440 -19888
rect 400640 -20012 400766 -19956
rect 400822 -20012 400890 -19956
rect 400946 -20012 401014 -19956
rect 401070 -20012 401138 -19956
rect 401194 -20012 401262 -19956
rect 401318 -20012 401440 -19956
rect 400640 -20080 401440 -20012
rect 400640 -20136 400766 -20080
rect 400822 -20136 400890 -20080
rect 400946 -20136 401014 -20080
rect 401070 -20136 401138 -20080
rect 401194 -20136 401262 -20080
rect 401318 -20136 401440 -20080
rect 400640 -20204 401440 -20136
rect 400640 -20260 400766 -20204
rect 400822 -20260 400890 -20204
rect 400946 -20260 401014 -20204
rect 401070 -20260 401138 -20204
rect 401194 -20260 401262 -20204
rect 401318 -20260 401440 -20204
rect 400640 -20328 401440 -20260
rect 400640 -20384 400766 -20328
rect 400822 -20384 400890 -20328
rect 400946 -20384 401014 -20328
rect 401070 -20384 401138 -20328
rect 401194 -20384 401262 -20328
rect 401318 -20384 401440 -20328
rect 400640 -20452 401440 -20384
rect 400640 -20508 400766 -20452
rect 400822 -20508 400890 -20452
rect 400946 -20508 401014 -20452
rect 401070 -20508 401138 -20452
rect 401194 -20508 401262 -20452
rect 401318 -20508 401440 -20452
rect 400640 -20576 401440 -20508
rect 400640 -20632 400766 -20576
rect 400822 -20632 400890 -20576
rect 400946 -20632 401014 -20576
rect 401070 -20632 401138 -20576
rect 401194 -20632 401262 -20576
rect 401318 -20632 401440 -20576
rect 400640 -20700 401440 -20632
rect 400640 -20756 400766 -20700
rect 400822 -20756 400890 -20700
rect 400946 -20756 401014 -20700
rect 401070 -20756 401138 -20700
rect 401194 -20756 401262 -20700
rect 401318 -20756 401440 -20700
rect 400640 -20824 401440 -20756
rect 400640 -20880 400766 -20824
rect 400822 -20880 400890 -20824
rect 400946 -20880 401014 -20824
rect 401070 -20880 401138 -20824
rect 401194 -20880 401262 -20824
rect 401318 -20880 401440 -20824
rect 400640 -20948 401440 -20880
rect 400640 -21004 400766 -20948
rect 400822 -21004 400890 -20948
rect 400946 -21004 401014 -20948
rect 401070 -21004 401138 -20948
rect 401194 -21004 401262 -20948
rect 401318 -21004 401440 -20948
rect 400640 -21072 401440 -21004
rect 400640 -21128 400766 -21072
rect 400822 -21128 400890 -21072
rect 400946 -21128 401014 -21072
rect 401070 -21128 401138 -21072
rect 401194 -21128 401262 -21072
rect 401318 -21128 401440 -21072
rect 400640 -21196 401440 -21128
rect 400640 -21252 400766 -21196
rect 400822 -21252 400890 -21196
rect 400946 -21252 401014 -21196
rect 401070 -21252 401138 -21196
rect 401194 -21252 401262 -21196
rect 401318 -21252 401440 -21196
rect 400640 -21320 401440 -21252
rect 400640 -21376 400766 -21320
rect 400822 -21376 400890 -21320
rect 400946 -21376 401014 -21320
rect 401070 -21376 401138 -21320
rect 401194 -21376 401262 -21320
rect 401318 -21376 401440 -21320
rect 400640 -21444 401440 -21376
rect 400640 -21500 400766 -21444
rect 400822 -21500 400890 -21444
rect 400946 -21500 401014 -21444
rect 401070 -21500 401138 -21444
rect 401194 -21500 401262 -21444
rect 401318 -21500 401440 -21444
rect 400640 -21568 401440 -21500
rect 400640 -21624 400766 -21568
rect 400822 -21624 400890 -21568
rect 400946 -21624 401014 -21568
rect 401070 -21624 401138 -21568
rect 401194 -21624 401262 -21568
rect 401318 -21624 401440 -21568
rect 400640 -21692 401440 -21624
rect 400640 -21748 400766 -21692
rect 400822 -21748 400890 -21692
rect 400946 -21748 401014 -21692
rect 401070 -21748 401138 -21692
rect 401194 -21748 401262 -21692
rect 401318 -21748 401440 -21692
rect 400640 -21816 401440 -21748
rect 400640 -21872 400766 -21816
rect 400822 -21872 400890 -21816
rect 400946 -21872 401014 -21816
rect 401070 -21872 401138 -21816
rect 401194 -21872 401262 -21816
rect 401318 -21872 401440 -21816
rect 400640 -21940 401440 -21872
rect 400640 -21996 400766 -21940
rect 400822 -21996 400890 -21940
rect 400946 -21996 401014 -21940
rect 401070 -21996 401138 -21940
rect 401194 -21996 401262 -21940
rect 401318 -21996 401440 -21940
rect 400640 -22064 401440 -21996
rect 400640 -22120 400766 -22064
rect 400822 -22120 400890 -22064
rect 400946 -22120 401014 -22064
rect 401070 -22120 401138 -22064
rect 401194 -22120 401262 -22064
rect 401318 -22120 401440 -22064
rect 400640 -22188 401440 -22120
rect 400640 -22244 400766 -22188
rect 400822 -22244 400890 -22188
rect 400946 -22244 401014 -22188
rect 401070 -22244 401138 -22188
rect 401194 -22244 401262 -22188
rect 401318 -22244 401440 -22188
rect 400640 -22312 401440 -22244
rect 400640 -22368 400766 -22312
rect 400822 -22368 400890 -22312
rect 400946 -22368 401014 -22312
rect 401070 -22368 401138 -22312
rect 401194 -22368 401262 -22312
rect 401318 -22368 401440 -22312
rect 400640 -22436 401440 -22368
rect 400640 -22492 400766 -22436
rect 400822 -22492 400890 -22436
rect 400946 -22492 401014 -22436
rect 401070 -22492 401138 -22436
rect 401194 -22492 401262 -22436
rect 401318 -22492 401440 -22436
rect 400640 -22560 401440 -22492
rect 400640 -22616 400766 -22560
rect 400822 -22616 400890 -22560
rect 400946 -22616 401014 -22560
rect 401070 -22616 401138 -22560
rect 401194 -22616 401262 -22560
rect 401318 -22616 401440 -22560
rect 400640 -22684 401440 -22616
rect 400640 -22740 400766 -22684
rect 400822 -22740 400890 -22684
rect 400946 -22740 401014 -22684
rect 401070 -22740 401138 -22684
rect 401194 -22740 401262 -22684
rect 401318 -22740 401440 -22684
rect 400640 -22808 401440 -22740
rect 400640 -22864 400766 -22808
rect 400822 -22864 400890 -22808
rect 400946 -22864 401014 -22808
rect 401070 -22864 401138 -22808
rect 401194 -22864 401262 -22808
rect 401318 -22864 401440 -22808
rect 400640 -22932 401440 -22864
rect 400640 -22988 400766 -22932
rect 400822 -22988 400890 -22932
rect 400946 -22988 401014 -22932
rect 401070 -22988 401138 -22932
rect 401194 -22988 401262 -22932
rect 401318 -22988 401440 -22932
rect 400640 -23056 401440 -22988
rect 400640 -23112 400766 -23056
rect 400822 -23112 400890 -23056
rect 400946 -23112 401014 -23056
rect 401070 -23112 401138 -23056
rect 401194 -23112 401262 -23056
rect 401318 -23112 401440 -23056
rect 400640 -23180 401440 -23112
rect 400640 -23236 400766 -23180
rect 400822 -23236 400890 -23180
rect 400946 -23236 401014 -23180
rect 401070 -23236 401138 -23180
rect 401194 -23236 401262 -23180
rect 401318 -23236 401440 -23180
rect 400640 -23304 401440 -23236
rect 400640 -23360 400766 -23304
rect 400822 -23360 400890 -23304
rect 400946 -23360 401014 -23304
rect 401070 -23360 401138 -23304
rect 401194 -23360 401262 -23304
rect 401318 -23360 401440 -23304
rect 400640 -23428 401440 -23360
rect 400640 -23484 400766 -23428
rect 400822 -23484 400890 -23428
rect 400946 -23484 401014 -23428
rect 401070 -23484 401138 -23428
rect 401194 -23484 401262 -23428
rect 401318 -23484 401440 -23428
rect 400640 -23552 401440 -23484
rect 400640 -23608 400766 -23552
rect 400822 -23608 400890 -23552
rect 400946 -23608 401014 -23552
rect 401070 -23608 401138 -23552
rect 401194 -23608 401262 -23552
rect 401318 -23608 401440 -23552
rect 400640 -23676 401440 -23608
rect 400640 -23732 400766 -23676
rect 400822 -23732 400890 -23676
rect 400946 -23732 401014 -23676
rect 401070 -23732 401138 -23676
rect 401194 -23732 401262 -23676
rect 401318 -23732 401440 -23676
rect 400640 -23800 401440 -23732
rect 400640 -23856 400766 -23800
rect 400822 -23856 400890 -23800
rect 400946 -23856 401014 -23800
rect 401070 -23856 401138 -23800
rect 401194 -23856 401262 -23800
rect 401318 -23856 401440 -23800
rect 400640 -23924 401440 -23856
rect 400640 -23980 400766 -23924
rect 400822 -23980 400890 -23924
rect 400946 -23980 401014 -23924
rect 401070 -23980 401138 -23924
rect 401194 -23980 401262 -23924
rect 401318 -23980 401440 -23924
rect 400640 -24048 401440 -23980
rect 400640 -24104 400766 -24048
rect 400822 -24104 400890 -24048
rect 400946 -24104 401014 -24048
rect 401070 -24104 401138 -24048
rect 401194 -24104 401262 -24048
rect 401318 -24104 401440 -24048
rect 400640 -24172 401440 -24104
rect 400640 -24228 400766 -24172
rect 400822 -24228 400890 -24172
rect 400946 -24228 401014 -24172
rect 401070 -24228 401138 -24172
rect 401194 -24228 401262 -24172
rect 401318 -24228 401440 -24172
rect 400640 -24296 401440 -24228
rect 400640 -24352 400766 -24296
rect 400822 -24352 400890 -24296
rect 400946 -24352 401014 -24296
rect 401070 -24352 401138 -24296
rect 401194 -24352 401262 -24296
rect 401318 -24352 401440 -24296
rect 400640 -24420 401440 -24352
rect 400640 -24476 400766 -24420
rect 400822 -24476 400890 -24420
rect 400946 -24476 401014 -24420
rect 401070 -24476 401138 -24420
rect 401194 -24476 401262 -24420
rect 401318 -24476 401440 -24420
rect 400640 -24544 401440 -24476
rect 400640 -24600 400766 -24544
rect 400822 -24600 400890 -24544
rect 400946 -24600 401014 -24544
rect 401070 -24600 401138 -24544
rect 401194 -24600 401262 -24544
rect 401318 -24600 401440 -24544
rect 400640 -24668 401440 -24600
rect 400640 -24724 400766 -24668
rect 400822 -24724 400890 -24668
rect 400946 -24724 401014 -24668
rect 401070 -24724 401138 -24668
rect 401194 -24724 401262 -24668
rect 401318 -24724 401440 -24668
rect 400640 -24792 401440 -24724
rect 400640 -24848 400766 -24792
rect 400822 -24848 400890 -24792
rect 400946 -24848 401014 -24792
rect 401070 -24848 401138 -24792
rect 401194 -24848 401262 -24792
rect 401318 -24848 401440 -24792
rect 400640 -24916 401440 -24848
rect 400640 -24972 400766 -24916
rect 400822 -24972 400890 -24916
rect 400946 -24972 401014 -24916
rect 401070 -24972 401138 -24916
rect 401194 -24972 401262 -24916
rect 401318 -24972 401440 -24916
rect 400640 -25040 401440 -24972
rect 400640 -25096 400766 -25040
rect 400822 -25096 400890 -25040
rect 400946 -25096 401014 -25040
rect 401070 -25096 401138 -25040
rect 401194 -25096 401262 -25040
rect 401318 -25096 401440 -25040
rect 400640 -25164 401440 -25096
rect 400640 -25220 400766 -25164
rect 400822 -25220 400890 -25164
rect 400946 -25220 401014 -25164
rect 401070 -25220 401138 -25164
rect 401194 -25220 401262 -25164
rect 401318 -25220 401440 -25164
rect 400640 -25288 401440 -25220
rect 400640 -25344 400766 -25288
rect 400822 -25344 400890 -25288
rect 400946 -25344 401014 -25288
rect 401070 -25344 401138 -25288
rect 401194 -25344 401262 -25288
rect 401318 -25344 401440 -25288
rect 400640 -25412 401440 -25344
rect 400640 -25468 400766 -25412
rect 400822 -25468 400890 -25412
rect 400946 -25468 401014 -25412
rect 401070 -25468 401138 -25412
rect 401194 -25468 401262 -25412
rect 401318 -25468 401440 -25412
rect 400640 -25536 401440 -25468
rect 400640 -25590 400766 -25536
rect 388506 -25592 400766 -25590
rect 400822 -25592 400890 -25536
rect 400946 -25592 401014 -25536
rect 401070 -25592 401138 -25536
rect 401194 -25592 401262 -25536
rect 401318 -25592 401440 -25536
rect 387840 -25660 401440 -25592
rect 387840 -25716 387954 -25660
rect 388010 -25716 388078 -25660
rect 388134 -25716 388202 -25660
rect 388258 -25716 388326 -25660
rect 388382 -25716 388450 -25660
rect 388506 -25688 400766 -25660
rect 388506 -25716 388655 -25688
rect 387840 -25744 388655 -25716
rect 388711 -25744 388797 -25688
rect 388853 -25744 388939 -25688
rect 388995 -25744 389081 -25688
rect 389137 -25744 389223 -25688
rect 389279 -25744 389365 -25688
rect 389421 -25744 389507 -25688
rect 389563 -25744 389649 -25688
rect 389705 -25744 389791 -25688
rect 389847 -25744 389933 -25688
rect 389989 -25744 390075 -25688
rect 390131 -25744 390217 -25688
rect 390273 -25744 390359 -25688
rect 390415 -25744 390501 -25688
rect 390557 -25744 390643 -25688
rect 390699 -25744 390785 -25688
rect 390841 -25744 390927 -25688
rect 390983 -25744 391069 -25688
rect 391125 -25744 391211 -25688
rect 391267 -25744 391353 -25688
rect 391409 -25744 391495 -25688
rect 391551 -25744 391637 -25688
rect 391693 -25744 391779 -25688
rect 391835 -25744 391921 -25688
rect 391977 -25744 392063 -25688
rect 392119 -25744 392205 -25688
rect 392261 -25744 392347 -25688
rect 392403 -25744 392489 -25688
rect 392545 -25744 392631 -25688
rect 392687 -25744 392773 -25688
rect 392829 -25744 392915 -25688
rect 392971 -25744 393057 -25688
rect 393113 -25744 393199 -25688
rect 393255 -25744 393341 -25688
rect 393397 -25744 393483 -25688
rect 393539 -25744 393625 -25688
rect 393681 -25744 393767 -25688
rect 393823 -25744 393909 -25688
rect 393965 -25744 394051 -25688
rect 394107 -25744 394193 -25688
rect 394249 -25744 394335 -25688
rect 394391 -25744 394477 -25688
rect 394533 -25744 394619 -25688
rect 394675 -25744 394761 -25688
rect 394817 -25744 394903 -25688
rect 394959 -25744 395045 -25688
rect 395101 -25744 395187 -25688
rect 395243 -25744 395329 -25688
rect 395385 -25744 395471 -25688
rect 395527 -25744 395613 -25688
rect 395669 -25744 395755 -25688
rect 395811 -25744 395897 -25688
rect 395953 -25744 396039 -25688
rect 396095 -25744 396181 -25688
rect 396237 -25744 396323 -25688
rect 396379 -25744 396465 -25688
rect 396521 -25744 396607 -25688
rect 396663 -25744 396749 -25688
rect 396805 -25744 396891 -25688
rect 396947 -25744 397033 -25688
rect 397089 -25744 397175 -25688
rect 397231 -25744 397317 -25688
rect 397373 -25744 397459 -25688
rect 397515 -25744 397601 -25688
rect 397657 -25744 397743 -25688
rect 397799 -25744 397885 -25688
rect 397941 -25744 398027 -25688
rect 398083 -25744 398169 -25688
rect 398225 -25744 398311 -25688
rect 398367 -25744 398453 -25688
rect 398509 -25744 398595 -25688
rect 398651 -25744 398737 -25688
rect 398793 -25744 398879 -25688
rect 398935 -25744 399021 -25688
rect 399077 -25744 399163 -25688
rect 399219 -25744 399305 -25688
rect 399361 -25744 399447 -25688
rect 399503 -25744 399589 -25688
rect 399645 -25744 399731 -25688
rect 399787 -25744 399873 -25688
rect 399929 -25744 400015 -25688
rect 400071 -25744 400157 -25688
rect 400213 -25744 400299 -25688
rect 400355 -25744 400441 -25688
rect 400497 -25744 400583 -25688
rect 400639 -25716 400766 -25688
rect 400822 -25716 400890 -25660
rect 400946 -25716 401014 -25660
rect 401070 -25716 401138 -25660
rect 401194 -25716 401262 -25660
rect 401318 -25716 401440 -25660
rect 400639 -25744 401440 -25716
rect 387840 -25784 401440 -25744
rect 387840 -25840 387954 -25784
rect 388010 -25840 388078 -25784
rect 388134 -25840 388202 -25784
rect 388258 -25840 388326 -25784
rect 388382 -25840 388450 -25784
rect 388506 -25830 400766 -25784
rect 388506 -25840 388655 -25830
rect 387840 -25886 388655 -25840
rect 388711 -25886 388797 -25830
rect 388853 -25886 388939 -25830
rect 388995 -25886 389081 -25830
rect 389137 -25886 389223 -25830
rect 389279 -25886 389365 -25830
rect 389421 -25886 389507 -25830
rect 389563 -25886 389649 -25830
rect 389705 -25886 389791 -25830
rect 389847 -25886 389933 -25830
rect 389989 -25886 390075 -25830
rect 390131 -25886 390217 -25830
rect 390273 -25886 390359 -25830
rect 390415 -25886 390501 -25830
rect 390557 -25886 390643 -25830
rect 390699 -25886 390785 -25830
rect 390841 -25886 390927 -25830
rect 390983 -25886 391069 -25830
rect 391125 -25886 391211 -25830
rect 391267 -25886 391353 -25830
rect 391409 -25886 391495 -25830
rect 391551 -25886 391637 -25830
rect 391693 -25886 391779 -25830
rect 391835 -25886 391921 -25830
rect 391977 -25886 392063 -25830
rect 392119 -25886 392205 -25830
rect 392261 -25886 392347 -25830
rect 392403 -25886 392489 -25830
rect 392545 -25886 392631 -25830
rect 392687 -25886 392773 -25830
rect 392829 -25886 392915 -25830
rect 392971 -25886 393057 -25830
rect 393113 -25886 393199 -25830
rect 393255 -25886 393341 -25830
rect 393397 -25886 393483 -25830
rect 393539 -25886 393625 -25830
rect 393681 -25886 393767 -25830
rect 393823 -25886 393909 -25830
rect 393965 -25886 394051 -25830
rect 394107 -25886 394193 -25830
rect 394249 -25886 394335 -25830
rect 394391 -25886 394477 -25830
rect 394533 -25886 394619 -25830
rect 394675 -25886 394761 -25830
rect 394817 -25886 394903 -25830
rect 394959 -25886 395045 -25830
rect 395101 -25886 395187 -25830
rect 395243 -25886 395329 -25830
rect 395385 -25886 395471 -25830
rect 395527 -25886 395613 -25830
rect 395669 -25886 395755 -25830
rect 395811 -25886 395897 -25830
rect 395953 -25886 396039 -25830
rect 396095 -25886 396181 -25830
rect 396237 -25886 396323 -25830
rect 396379 -25886 396465 -25830
rect 396521 -25886 396607 -25830
rect 396663 -25886 396749 -25830
rect 396805 -25886 396891 -25830
rect 396947 -25886 397033 -25830
rect 397089 -25886 397175 -25830
rect 397231 -25886 397317 -25830
rect 397373 -25886 397459 -25830
rect 397515 -25886 397601 -25830
rect 397657 -25886 397743 -25830
rect 397799 -25886 397885 -25830
rect 397941 -25886 398027 -25830
rect 398083 -25886 398169 -25830
rect 398225 -25886 398311 -25830
rect 398367 -25886 398453 -25830
rect 398509 -25886 398595 -25830
rect 398651 -25886 398737 -25830
rect 398793 -25886 398879 -25830
rect 398935 -25886 399021 -25830
rect 399077 -25886 399163 -25830
rect 399219 -25886 399305 -25830
rect 399361 -25886 399447 -25830
rect 399503 -25886 399589 -25830
rect 399645 -25886 399731 -25830
rect 399787 -25886 399873 -25830
rect 399929 -25886 400015 -25830
rect 400071 -25886 400157 -25830
rect 400213 -25886 400299 -25830
rect 400355 -25886 400441 -25830
rect 400497 -25886 400583 -25830
rect 400639 -25840 400766 -25830
rect 400822 -25840 400890 -25784
rect 400946 -25840 401014 -25784
rect 401070 -25840 401138 -25784
rect 401194 -25840 401262 -25784
rect 401318 -25840 401440 -25784
rect 400639 -25886 401440 -25840
rect 387840 -25990 401440 -25886
<< via2 >>
rect 387986 -13097 388042 -13041
rect 388110 -13097 388166 -13041
rect 388234 -13097 388290 -13041
rect 388358 -13097 388414 -13041
rect 388482 -13097 388538 -13041
rect 388606 -13097 388662 -13041
rect 388730 -13097 388786 -13041
rect 388854 -13097 388910 -13041
rect 388978 -13097 389034 -13041
rect 389102 -13097 389158 -13041
rect 389226 -13097 389282 -13041
rect 389350 -13097 389406 -13041
rect 389474 -13097 389530 -13041
rect 389598 -13097 389654 -13041
rect 389722 -13097 389778 -13041
rect 389846 -13097 389902 -13041
rect 389970 -13097 390026 -13041
rect 390094 -13097 390150 -13041
rect 390218 -13097 390274 -13041
rect 390342 -13097 390398 -13041
rect 390466 -13097 390522 -13041
rect 390590 -13097 390646 -13041
rect 390714 -13097 390770 -13041
rect 390838 -13097 390894 -13041
rect 390962 -13097 391018 -13041
rect 391086 -13097 391142 -13041
rect 391210 -13097 391266 -13041
rect 391334 -13097 391390 -13041
rect 391458 -13097 391514 -13041
rect 391582 -13097 391638 -13041
rect 391706 -13097 391762 -13041
rect 391830 -13097 391886 -13041
rect 391954 -13097 392010 -13041
rect 392078 -13097 392134 -13041
rect 392202 -13097 392258 -13041
rect 392326 -13097 392382 -13041
rect 392450 -13097 392506 -13041
rect 392574 -13097 392630 -13041
rect 392698 -13097 392754 -13041
rect 392822 -13097 392878 -13041
rect 392946 -13097 393002 -13041
rect 393070 -13097 393126 -13041
rect 393194 -13097 393250 -13041
rect 393318 -13097 393374 -13041
rect 393442 -13097 393498 -13041
rect 393566 -13097 393622 -13041
rect 393690 -13097 393746 -13041
rect 393814 -13097 393870 -13041
rect 393938 -13097 393994 -13041
rect 394062 -13097 394118 -13041
rect 394186 -13097 394242 -13041
rect 394310 -13097 394366 -13041
rect 394434 -13097 394490 -13041
rect 394558 -13097 394614 -13041
rect 394682 -13097 394738 -13041
rect 394806 -13097 394862 -13041
rect 394930 -13097 394986 -13041
rect 395054 -13097 395110 -13041
rect 395178 -13097 395234 -13041
rect 395302 -13097 395358 -13041
rect 395426 -13097 395482 -13041
rect 395550 -13097 395606 -13041
rect 395674 -13097 395730 -13041
rect 395798 -13097 395854 -13041
rect 395922 -13097 395978 -13041
rect 396046 -13097 396102 -13041
rect 396170 -13097 396226 -13041
rect 396294 -13097 396350 -13041
rect 396418 -13097 396474 -13041
rect 396542 -13097 396598 -13041
rect 396666 -13097 396722 -13041
rect 396790 -13097 396846 -13041
rect 396914 -13097 396970 -13041
rect 397038 -13097 397094 -13041
rect 397162 -13097 397218 -13041
rect 397286 -13097 397342 -13041
rect 397410 -13097 397466 -13041
rect 397534 -13097 397590 -13041
rect 397658 -13097 397714 -13041
rect 397782 -13097 397838 -13041
rect 397906 -13097 397962 -13041
rect 398030 -13097 398086 -13041
rect 398154 -13097 398210 -13041
rect 398278 -13097 398334 -13041
rect 398402 -13097 398458 -13041
rect 398526 -13097 398582 -13041
rect 398650 -13097 398706 -13041
rect 398774 -13097 398830 -13041
rect 398898 -13097 398954 -13041
rect 399022 -13097 399078 -13041
rect 399146 -13097 399202 -13041
rect 399270 -13097 399326 -13041
rect 399394 -13097 399450 -13041
rect 399518 -13097 399574 -13041
rect 399642 -13097 399698 -13041
rect 399766 -13097 399822 -13041
rect 399890 -13097 399946 -13041
rect 400014 -13097 400070 -13041
rect 400138 -13097 400194 -13041
rect 400262 -13097 400318 -13041
rect 400386 -13097 400442 -13041
rect 400510 -13097 400566 -13041
rect 400634 -13097 400690 -13041
rect 400758 -13097 400814 -13041
rect 400882 -13097 400938 -13041
rect 401006 -13097 401062 -13041
rect 401130 -13097 401186 -13041
rect 401254 -13097 401310 -13041
rect 387986 -13221 388042 -13165
rect 388110 -13221 388166 -13165
rect 388234 -13221 388290 -13165
rect 388358 -13221 388414 -13165
rect 388482 -13221 388538 -13165
rect 388606 -13221 388662 -13165
rect 388730 -13221 388786 -13165
rect 388854 -13221 388910 -13165
rect 388978 -13221 389034 -13165
rect 389102 -13221 389158 -13165
rect 389226 -13221 389282 -13165
rect 389350 -13221 389406 -13165
rect 389474 -13221 389530 -13165
rect 389598 -13221 389654 -13165
rect 389722 -13221 389778 -13165
rect 389846 -13221 389902 -13165
rect 389970 -13221 390026 -13165
rect 390094 -13221 390150 -13165
rect 390218 -13221 390274 -13165
rect 390342 -13221 390398 -13165
rect 390466 -13221 390522 -13165
rect 390590 -13221 390646 -13165
rect 390714 -13221 390770 -13165
rect 390838 -13221 390894 -13165
rect 390962 -13221 391018 -13165
rect 391086 -13221 391142 -13165
rect 391210 -13221 391266 -13165
rect 391334 -13221 391390 -13165
rect 391458 -13221 391514 -13165
rect 391582 -13221 391638 -13165
rect 391706 -13221 391762 -13165
rect 391830 -13221 391886 -13165
rect 391954 -13221 392010 -13165
rect 392078 -13221 392134 -13165
rect 392202 -13221 392258 -13165
rect 392326 -13221 392382 -13165
rect 392450 -13221 392506 -13165
rect 392574 -13221 392630 -13165
rect 392698 -13221 392754 -13165
rect 392822 -13221 392878 -13165
rect 392946 -13221 393002 -13165
rect 393070 -13221 393126 -13165
rect 393194 -13221 393250 -13165
rect 393318 -13221 393374 -13165
rect 393442 -13221 393498 -13165
rect 393566 -13221 393622 -13165
rect 393690 -13221 393746 -13165
rect 393814 -13221 393870 -13165
rect 393938 -13221 393994 -13165
rect 394062 -13221 394118 -13165
rect 394186 -13221 394242 -13165
rect 394310 -13221 394366 -13165
rect 394434 -13221 394490 -13165
rect 394558 -13221 394614 -13165
rect 394682 -13221 394738 -13165
rect 394806 -13221 394862 -13165
rect 394930 -13221 394986 -13165
rect 395054 -13221 395110 -13165
rect 395178 -13221 395234 -13165
rect 395302 -13221 395358 -13165
rect 395426 -13221 395482 -13165
rect 395550 -13221 395606 -13165
rect 395674 -13221 395730 -13165
rect 395798 -13221 395854 -13165
rect 395922 -13221 395978 -13165
rect 396046 -13221 396102 -13165
rect 396170 -13221 396226 -13165
rect 396294 -13221 396350 -13165
rect 396418 -13221 396474 -13165
rect 396542 -13221 396598 -13165
rect 396666 -13221 396722 -13165
rect 396790 -13221 396846 -13165
rect 396914 -13221 396970 -13165
rect 397038 -13221 397094 -13165
rect 397162 -13221 397218 -13165
rect 397286 -13221 397342 -13165
rect 397410 -13221 397466 -13165
rect 397534 -13221 397590 -13165
rect 397658 -13221 397714 -13165
rect 397782 -13221 397838 -13165
rect 397906 -13221 397962 -13165
rect 398030 -13221 398086 -13165
rect 398154 -13221 398210 -13165
rect 398278 -13221 398334 -13165
rect 398402 -13221 398458 -13165
rect 398526 -13221 398582 -13165
rect 398650 -13221 398706 -13165
rect 398774 -13221 398830 -13165
rect 398898 -13221 398954 -13165
rect 399022 -13221 399078 -13165
rect 399146 -13221 399202 -13165
rect 399270 -13221 399326 -13165
rect 399394 -13221 399450 -13165
rect 399518 -13221 399574 -13165
rect 399642 -13221 399698 -13165
rect 399766 -13221 399822 -13165
rect 399890 -13221 399946 -13165
rect 400014 -13221 400070 -13165
rect 400138 -13221 400194 -13165
rect 400262 -13221 400318 -13165
rect 400386 -13221 400442 -13165
rect 400510 -13221 400566 -13165
rect 400634 -13221 400690 -13165
rect 400758 -13221 400814 -13165
rect 400882 -13221 400938 -13165
rect 401006 -13221 401062 -13165
rect 401130 -13221 401186 -13165
rect 401254 -13221 401310 -13165
rect 387986 -13345 388042 -13289
rect 388110 -13345 388166 -13289
rect 388234 -13345 388290 -13289
rect 388358 -13345 388414 -13289
rect 388482 -13345 388538 -13289
rect 388606 -13345 388662 -13289
rect 388730 -13345 388786 -13289
rect 388854 -13345 388910 -13289
rect 388978 -13345 389034 -13289
rect 389102 -13345 389158 -13289
rect 389226 -13345 389282 -13289
rect 389350 -13345 389406 -13289
rect 389474 -13345 389530 -13289
rect 389598 -13345 389654 -13289
rect 389722 -13345 389778 -13289
rect 389846 -13345 389902 -13289
rect 389970 -13345 390026 -13289
rect 390094 -13345 390150 -13289
rect 390218 -13345 390274 -13289
rect 390342 -13345 390398 -13289
rect 390466 -13345 390522 -13289
rect 390590 -13345 390646 -13289
rect 390714 -13345 390770 -13289
rect 390838 -13345 390894 -13289
rect 390962 -13345 391018 -13289
rect 391086 -13345 391142 -13289
rect 391210 -13345 391266 -13289
rect 391334 -13345 391390 -13289
rect 391458 -13345 391514 -13289
rect 391582 -13345 391638 -13289
rect 391706 -13345 391762 -13289
rect 391830 -13345 391886 -13289
rect 391954 -13345 392010 -13289
rect 392078 -13345 392134 -13289
rect 392202 -13345 392258 -13289
rect 392326 -13345 392382 -13289
rect 392450 -13345 392506 -13289
rect 392574 -13345 392630 -13289
rect 392698 -13345 392754 -13289
rect 392822 -13345 392878 -13289
rect 392946 -13345 393002 -13289
rect 393070 -13345 393126 -13289
rect 393194 -13345 393250 -13289
rect 393318 -13345 393374 -13289
rect 393442 -13345 393498 -13289
rect 393566 -13345 393622 -13289
rect 393690 -13345 393746 -13289
rect 393814 -13345 393870 -13289
rect 393938 -13345 393994 -13289
rect 394062 -13345 394118 -13289
rect 394186 -13345 394242 -13289
rect 394310 -13345 394366 -13289
rect 394434 -13345 394490 -13289
rect 394558 -13345 394614 -13289
rect 394682 -13345 394738 -13289
rect 394806 -13345 394862 -13289
rect 394930 -13345 394986 -13289
rect 395054 -13345 395110 -13289
rect 395178 -13345 395234 -13289
rect 395302 -13345 395358 -13289
rect 395426 -13345 395482 -13289
rect 395550 -13345 395606 -13289
rect 395674 -13345 395730 -13289
rect 395798 -13345 395854 -13289
rect 395922 -13345 395978 -13289
rect 396046 -13345 396102 -13289
rect 396170 -13345 396226 -13289
rect 396294 -13345 396350 -13289
rect 396418 -13345 396474 -13289
rect 396542 -13345 396598 -13289
rect 396666 -13345 396722 -13289
rect 396790 -13345 396846 -13289
rect 396914 -13345 396970 -13289
rect 397038 -13345 397094 -13289
rect 397162 -13345 397218 -13289
rect 397286 -13345 397342 -13289
rect 397410 -13345 397466 -13289
rect 397534 -13345 397590 -13289
rect 397658 -13345 397714 -13289
rect 397782 -13345 397838 -13289
rect 397906 -13345 397962 -13289
rect 398030 -13345 398086 -13289
rect 398154 -13345 398210 -13289
rect 398278 -13345 398334 -13289
rect 398402 -13345 398458 -13289
rect 398526 -13345 398582 -13289
rect 398650 -13345 398706 -13289
rect 398774 -13345 398830 -13289
rect 398898 -13345 398954 -13289
rect 399022 -13345 399078 -13289
rect 399146 -13345 399202 -13289
rect 399270 -13345 399326 -13289
rect 399394 -13345 399450 -13289
rect 399518 -13345 399574 -13289
rect 399642 -13345 399698 -13289
rect 399766 -13345 399822 -13289
rect 399890 -13345 399946 -13289
rect 400014 -13345 400070 -13289
rect 400138 -13345 400194 -13289
rect 400262 -13345 400318 -13289
rect 400386 -13345 400442 -13289
rect 400510 -13345 400566 -13289
rect 400634 -13345 400690 -13289
rect 400758 -13345 400814 -13289
rect 400882 -13345 400938 -13289
rect 401006 -13345 401062 -13289
rect 401130 -13345 401186 -13289
rect 401254 -13345 401310 -13289
rect 387986 -13469 388042 -13413
rect 388110 -13469 388166 -13413
rect 388234 -13469 388290 -13413
rect 388358 -13469 388414 -13413
rect 388482 -13469 388538 -13413
rect 388606 -13469 388662 -13413
rect 388730 -13469 388786 -13413
rect 388854 -13469 388910 -13413
rect 388978 -13469 389034 -13413
rect 389102 -13469 389158 -13413
rect 389226 -13469 389282 -13413
rect 389350 -13469 389406 -13413
rect 389474 -13469 389530 -13413
rect 389598 -13469 389654 -13413
rect 389722 -13469 389778 -13413
rect 389846 -13469 389902 -13413
rect 389970 -13469 390026 -13413
rect 390094 -13469 390150 -13413
rect 390218 -13469 390274 -13413
rect 390342 -13469 390398 -13413
rect 390466 -13469 390522 -13413
rect 390590 -13469 390646 -13413
rect 390714 -13469 390770 -13413
rect 390838 -13469 390894 -13413
rect 390962 -13469 391018 -13413
rect 391086 -13469 391142 -13413
rect 391210 -13469 391266 -13413
rect 391334 -13469 391390 -13413
rect 391458 -13469 391514 -13413
rect 391582 -13469 391638 -13413
rect 391706 -13469 391762 -13413
rect 391830 -13469 391886 -13413
rect 391954 -13469 392010 -13413
rect 392078 -13469 392134 -13413
rect 392202 -13469 392258 -13413
rect 392326 -13469 392382 -13413
rect 392450 -13469 392506 -13413
rect 392574 -13469 392630 -13413
rect 392698 -13469 392754 -13413
rect 392822 -13469 392878 -13413
rect 392946 -13469 393002 -13413
rect 393070 -13469 393126 -13413
rect 393194 -13469 393250 -13413
rect 393318 -13469 393374 -13413
rect 393442 -13469 393498 -13413
rect 393566 -13469 393622 -13413
rect 393690 -13469 393746 -13413
rect 393814 -13469 393870 -13413
rect 393938 -13469 393994 -13413
rect 394062 -13469 394118 -13413
rect 394186 -13469 394242 -13413
rect 394310 -13469 394366 -13413
rect 394434 -13469 394490 -13413
rect 394558 -13469 394614 -13413
rect 394682 -13469 394738 -13413
rect 394806 -13469 394862 -13413
rect 394930 -13469 394986 -13413
rect 395054 -13469 395110 -13413
rect 395178 -13469 395234 -13413
rect 395302 -13469 395358 -13413
rect 395426 -13469 395482 -13413
rect 395550 -13469 395606 -13413
rect 395674 -13469 395730 -13413
rect 395798 -13469 395854 -13413
rect 395922 -13469 395978 -13413
rect 396046 -13469 396102 -13413
rect 396170 -13469 396226 -13413
rect 396294 -13469 396350 -13413
rect 396418 -13469 396474 -13413
rect 396542 -13469 396598 -13413
rect 396666 -13469 396722 -13413
rect 396790 -13469 396846 -13413
rect 396914 -13469 396970 -13413
rect 397038 -13469 397094 -13413
rect 397162 -13469 397218 -13413
rect 397286 -13469 397342 -13413
rect 397410 -13469 397466 -13413
rect 397534 -13469 397590 -13413
rect 397658 -13469 397714 -13413
rect 397782 -13469 397838 -13413
rect 397906 -13469 397962 -13413
rect 398030 -13469 398086 -13413
rect 398154 -13469 398210 -13413
rect 398278 -13469 398334 -13413
rect 398402 -13469 398458 -13413
rect 398526 -13469 398582 -13413
rect 398650 -13469 398706 -13413
rect 398774 -13469 398830 -13413
rect 398898 -13469 398954 -13413
rect 399022 -13469 399078 -13413
rect 399146 -13469 399202 -13413
rect 399270 -13469 399326 -13413
rect 399394 -13469 399450 -13413
rect 399518 -13469 399574 -13413
rect 399642 -13469 399698 -13413
rect 399766 -13469 399822 -13413
rect 399890 -13469 399946 -13413
rect 400014 -13469 400070 -13413
rect 400138 -13469 400194 -13413
rect 400262 -13469 400318 -13413
rect 400386 -13469 400442 -13413
rect 400510 -13469 400566 -13413
rect 400634 -13469 400690 -13413
rect 400758 -13469 400814 -13413
rect 400882 -13469 400938 -13413
rect 401006 -13469 401062 -13413
rect 401130 -13469 401186 -13413
rect 401254 -13469 401310 -13413
rect 387954 -13688 388010 -13632
rect 388078 -13688 388134 -13632
rect 388202 -13688 388258 -13632
rect 388326 -13688 388382 -13632
rect 388450 -13688 388506 -13632
rect 387954 -13812 388010 -13756
rect 388078 -13812 388134 -13756
rect 388202 -13812 388258 -13756
rect 388326 -13812 388382 -13756
rect 388450 -13812 388506 -13756
rect 387954 -13936 388010 -13880
rect 388078 -13936 388134 -13880
rect 388202 -13936 388258 -13880
rect 388326 -13936 388382 -13880
rect 388450 -13936 388506 -13880
rect 387954 -14060 388010 -14004
rect 388078 -14060 388134 -14004
rect 388202 -14060 388258 -14004
rect 388326 -14060 388382 -14004
rect 388450 -14060 388506 -14004
rect 387954 -14184 388010 -14128
rect 388078 -14184 388134 -14128
rect 388202 -14184 388258 -14128
rect 388326 -14184 388382 -14128
rect 388450 -14184 388506 -14128
rect 387954 -14308 388010 -14252
rect 388078 -14308 388134 -14252
rect 388202 -14308 388258 -14252
rect 388326 -14308 388382 -14252
rect 388450 -14308 388506 -14252
rect 387954 -14432 388010 -14376
rect 388078 -14432 388134 -14376
rect 388202 -14432 388258 -14376
rect 388326 -14432 388382 -14376
rect 388450 -14432 388506 -14376
rect 387954 -14556 388010 -14500
rect 388078 -14556 388134 -14500
rect 388202 -14556 388258 -14500
rect 388326 -14556 388382 -14500
rect 388450 -14556 388506 -14500
rect 387954 -14680 388010 -14624
rect 388078 -14680 388134 -14624
rect 388202 -14680 388258 -14624
rect 388326 -14680 388382 -14624
rect 388450 -14680 388506 -14624
rect 387954 -14804 388010 -14748
rect 388078 -14804 388134 -14748
rect 388202 -14804 388258 -14748
rect 388326 -14804 388382 -14748
rect 388450 -14804 388506 -14748
rect 387954 -14928 388010 -14872
rect 388078 -14928 388134 -14872
rect 388202 -14928 388258 -14872
rect 388326 -14928 388382 -14872
rect 388450 -14928 388506 -14872
rect 387954 -15052 388010 -14996
rect 388078 -15052 388134 -14996
rect 388202 -15052 388258 -14996
rect 388326 -15052 388382 -14996
rect 388450 -15052 388506 -14996
rect 387954 -15176 388010 -15120
rect 388078 -15176 388134 -15120
rect 388202 -15176 388258 -15120
rect 388326 -15176 388382 -15120
rect 388450 -15176 388506 -15120
rect 387954 -15300 388010 -15244
rect 388078 -15300 388134 -15244
rect 388202 -15300 388258 -15244
rect 388326 -15300 388382 -15244
rect 388450 -15300 388506 -15244
rect 387954 -15424 388010 -15368
rect 388078 -15424 388134 -15368
rect 388202 -15424 388258 -15368
rect 388326 -15424 388382 -15368
rect 388450 -15424 388506 -15368
rect 387954 -15548 388010 -15492
rect 388078 -15548 388134 -15492
rect 388202 -15548 388258 -15492
rect 388326 -15548 388382 -15492
rect 388450 -15548 388506 -15492
rect 387954 -15672 388010 -15616
rect 388078 -15672 388134 -15616
rect 388202 -15672 388258 -15616
rect 388326 -15672 388382 -15616
rect 388450 -15672 388506 -15616
rect 387954 -15796 388010 -15740
rect 388078 -15796 388134 -15740
rect 388202 -15796 388258 -15740
rect 388326 -15796 388382 -15740
rect 388450 -15796 388506 -15740
rect 387954 -15920 388010 -15864
rect 388078 -15920 388134 -15864
rect 388202 -15920 388258 -15864
rect 388326 -15920 388382 -15864
rect 388450 -15920 388506 -15864
rect 387954 -16044 388010 -15988
rect 388078 -16044 388134 -15988
rect 388202 -16044 388258 -15988
rect 388326 -16044 388382 -15988
rect 388450 -16044 388506 -15988
rect 387954 -16168 388010 -16112
rect 388078 -16168 388134 -16112
rect 388202 -16168 388258 -16112
rect 388326 -16168 388382 -16112
rect 388450 -16168 388506 -16112
rect 387954 -16292 388010 -16236
rect 388078 -16292 388134 -16236
rect 388202 -16292 388258 -16236
rect 388326 -16292 388382 -16236
rect 388450 -16292 388506 -16236
rect 387954 -16416 388010 -16360
rect 388078 -16416 388134 -16360
rect 388202 -16416 388258 -16360
rect 388326 -16416 388382 -16360
rect 388450 -16416 388506 -16360
rect 387954 -16540 388010 -16484
rect 388078 -16540 388134 -16484
rect 388202 -16540 388258 -16484
rect 388326 -16540 388382 -16484
rect 388450 -16540 388506 -16484
rect 387954 -16664 388010 -16608
rect 388078 -16664 388134 -16608
rect 388202 -16664 388258 -16608
rect 388326 -16664 388382 -16608
rect 388450 -16664 388506 -16608
rect 387954 -16788 388010 -16732
rect 388078 -16788 388134 -16732
rect 388202 -16788 388258 -16732
rect 388326 -16788 388382 -16732
rect 388450 -16788 388506 -16732
rect 387954 -16912 388010 -16856
rect 388078 -16912 388134 -16856
rect 388202 -16912 388258 -16856
rect 388326 -16912 388382 -16856
rect 388450 -16912 388506 -16856
rect 387954 -17036 388010 -16980
rect 388078 -17036 388134 -16980
rect 388202 -17036 388258 -16980
rect 388326 -17036 388382 -16980
rect 388450 -17036 388506 -16980
rect 387954 -17160 388010 -17104
rect 388078 -17160 388134 -17104
rect 388202 -17160 388258 -17104
rect 388326 -17160 388382 -17104
rect 388450 -17160 388506 -17104
rect 387954 -17284 388010 -17228
rect 388078 -17284 388134 -17228
rect 388202 -17284 388258 -17228
rect 388326 -17284 388382 -17228
rect 388450 -17284 388506 -17228
rect 387954 -17408 388010 -17352
rect 388078 -17408 388134 -17352
rect 388202 -17408 388258 -17352
rect 388326 -17408 388382 -17352
rect 388450 -17408 388506 -17352
rect 387954 -17532 388010 -17476
rect 388078 -17532 388134 -17476
rect 388202 -17532 388258 -17476
rect 388326 -17532 388382 -17476
rect 388450 -17532 388506 -17476
rect 387954 -17656 388010 -17600
rect 388078 -17656 388134 -17600
rect 388202 -17656 388258 -17600
rect 388326 -17656 388382 -17600
rect 388450 -17656 388506 -17600
rect 387954 -17780 388010 -17724
rect 388078 -17780 388134 -17724
rect 388202 -17780 388258 -17724
rect 388326 -17780 388382 -17724
rect 388450 -17780 388506 -17724
rect 387954 -17904 388010 -17848
rect 388078 -17904 388134 -17848
rect 388202 -17904 388258 -17848
rect 388326 -17904 388382 -17848
rect 388450 -17904 388506 -17848
rect 387954 -18028 388010 -17972
rect 388078 -18028 388134 -17972
rect 388202 -18028 388258 -17972
rect 388326 -18028 388382 -17972
rect 388450 -18028 388506 -17972
rect 387954 -18152 388010 -18096
rect 388078 -18152 388134 -18096
rect 388202 -18152 388258 -18096
rect 388326 -18152 388382 -18096
rect 388450 -18152 388506 -18096
rect 387954 -18276 388010 -18220
rect 388078 -18276 388134 -18220
rect 388202 -18276 388258 -18220
rect 388326 -18276 388382 -18220
rect 388450 -18276 388506 -18220
rect 387954 -18400 388010 -18344
rect 388078 -18400 388134 -18344
rect 388202 -18400 388258 -18344
rect 388326 -18400 388382 -18344
rect 388450 -18400 388506 -18344
rect 387954 -18524 388010 -18468
rect 388078 -18524 388134 -18468
rect 388202 -18524 388258 -18468
rect 388326 -18524 388382 -18468
rect 388450 -18524 388506 -18468
rect 387954 -18648 388010 -18592
rect 388078 -18648 388134 -18592
rect 388202 -18648 388258 -18592
rect 388326 -18648 388382 -18592
rect 388450 -18648 388506 -18592
rect 387954 -18772 388010 -18716
rect 388078 -18772 388134 -18716
rect 388202 -18772 388258 -18716
rect 388326 -18772 388382 -18716
rect 388450 -18772 388506 -18716
rect 387954 -18896 388010 -18840
rect 388078 -18896 388134 -18840
rect 388202 -18896 388258 -18840
rect 388326 -18896 388382 -18840
rect 388450 -18896 388506 -18840
rect 387954 -19020 388010 -18964
rect 388078 -19020 388134 -18964
rect 388202 -19020 388258 -18964
rect 388326 -19020 388382 -18964
rect 388450 -19020 388506 -18964
rect 387954 -19144 388010 -19088
rect 388078 -19144 388134 -19088
rect 388202 -19144 388258 -19088
rect 388326 -19144 388382 -19088
rect 388450 -19144 388506 -19088
rect 387954 -19268 388010 -19212
rect 388078 -19268 388134 -19212
rect 388202 -19268 388258 -19212
rect 388326 -19268 388382 -19212
rect 388450 -19268 388506 -19212
rect 387954 -19392 388010 -19336
rect 388078 -19392 388134 -19336
rect 388202 -19392 388258 -19336
rect 388326 -19392 388382 -19336
rect 388450 -19392 388506 -19336
rect 387954 -19516 388010 -19460
rect 388078 -19516 388134 -19460
rect 388202 -19516 388258 -19460
rect 388326 -19516 388382 -19460
rect 388450 -19516 388506 -19460
rect 387954 -19640 388010 -19584
rect 388078 -19640 388134 -19584
rect 388202 -19640 388258 -19584
rect 388326 -19640 388382 -19584
rect 388450 -19640 388506 -19584
rect 387954 -19764 388010 -19708
rect 388078 -19764 388134 -19708
rect 388202 -19764 388258 -19708
rect 388326 -19764 388382 -19708
rect 388450 -19764 388506 -19708
rect 387954 -19888 388010 -19832
rect 388078 -19888 388134 -19832
rect 388202 -19888 388258 -19832
rect 388326 -19888 388382 -19832
rect 388450 -19888 388506 -19832
rect 387954 -20012 388010 -19956
rect 388078 -20012 388134 -19956
rect 388202 -20012 388258 -19956
rect 388326 -20012 388382 -19956
rect 388450 -20012 388506 -19956
rect 387954 -20136 388010 -20080
rect 388078 -20136 388134 -20080
rect 388202 -20136 388258 -20080
rect 388326 -20136 388382 -20080
rect 388450 -20136 388506 -20080
rect 387954 -20260 388010 -20204
rect 388078 -20260 388134 -20204
rect 388202 -20260 388258 -20204
rect 388326 -20260 388382 -20204
rect 388450 -20260 388506 -20204
rect 387954 -20384 388010 -20328
rect 388078 -20384 388134 -20328
rect 388202 -20384 388258 -20328
rect 388326 -20384 388382 -20328
rect 388450 -20384 388506 -20328
rect 387954 -20508 388010 -20452
rect 388078 -20508 388134 -20452
rect 388202 -20508 388258 -20452
rect 388326 -20508 388382 -20452
rect 388450 -20508 388506 -20452
rect 387954 -20632 388010 -20576
rect 388078 -20632 388134 -20576
rect 388202 -20632 388258 -20576
rect 388326 -20632 388382 -20576
rect 388450 -20632 388506 -20576
rect 387954 -20756 388010 -20700
rect 388078 -20756 388134 -20700
rect 388202 -20756 388258 -20700
rect 388326 -20756 388382 -20700
rect 388450 -20756 388506 -20700
rect 387954 -20880 388010 -20824
rect 388078 -20880 388134 -20824
rect 388202 -20880 388258 -20824
rect 388326 -20880 388382 -20824
rect 388450 -20880 388506 -20824
rect 387954 -21004 388010 -20948
rect 388078 -21004 388134 -20948
rect 388202 -21004 388258 -20948
rect 388326 -21004 388382 -20948
rect 388450 -21004 388506 -20948
rect 387954 -21128 388010 -21072
rect 388078 -21128 388134 -21072
rect 388202 -21128 388258 -21072
rect 388326 -21128 388382 -21072
rect 388450 -21128 388506 -21072
rect 387954 -21252 388010 -21196
rect 388078 -21252 388134 -21196
rect 388202 -21252 388258 -21196
rect 388326 -21252 388382 -21196
rect 388450 -21252 388506 -21196
rect 387954 -21376 388010 -21320
rect 388078 -21376 388134 -21320
rect 388202 -21376 388258 -21320
rect 388326 -21376 388382 -21320
rect 388450 -21376 388506 -21320
rect 387954 -21500 388010 -21444
rect 388078 -21500 388134 -21444
rect 388202 -21500 388258 -21444
rect 388326 -21500 388382 -21444
rect 388450 -21500 388506 -21444
rect 387954 -21624 388010 -21568
rect 388078 -21624 388134 -21568
rect 388202 -21624 388258 -21568
rect 388326 -21624 388382 -21568
rect 388450 -21624 388506 -21568
rect 387954 -21748 388010 -21692
rect 388078 -21748 388134 -21692
rect 388202 -21748 388258 -21692
rect 388326 -21748 388382 -21692
rect 388450 -21748 388506 -21692
rect 387954 -21872 388010 -21816
rect 388078 -21872 388134 -21816
rect 388202 -21872 388258 -21816
rect 388326 -21872 388382 -21816
rect 388450 -21872 388506 -21816
rect 387954 -21996 388010 -21940
rect 388078 -21996 388134 -21940
rect 388202 -21996 388258 -21940
rect 388326 -21996 388382 -21940
rect 388450 -21996 388506 -21940
rect 387954 -22120 388010 -22064
rect 388078 -22120 388134 -22064
rect 388202 -22120 388258 -22064
rect 388326 -22120 388382 -22064
rect 388450 -22120 388506 -22064
rect 387954 -22244 388010 -22188
rect 388078 -22244 388134 -22188
rect 388202 -22244 388258 -22188
rect 388326 -22244 388382 -22188
rect 388450 -22244 388506 -22188
rect 387954 -22368 388010 -22312
rect 388078 -22368 388134 -22312
rect 388202 -22368 388258 -22312
rect 388326 -22368 388382 -22312
rect 388450 -22368 388506 -22312
rect 387954 -22492 388010 -22436
rect 388078 -22492 388134 -22436
rect 388202 -22492 388258 -22436
rect 388326 -22492 388382 -22436
rect 388450 -22492 388506 -22436
rect 387954 -22616 388010 -22560
rect 388078 -22616 388134 -22560
rect 388202 -22616 388258 -22560
rect 388326 -22616 388382 -22560
rect 388450 -22616 388506 -22560
rect 387954 -22740 388010 -22684
rect 388078 -22740 388134 -22684
rect 388202 -22740 388258 -22684
rect 388326 -22740 388382 -22684
rect 388450 -22740 388506 -22684
rect 387954 -22864 388010 -22808
rect 388078 -22864 388134 -22808
rect 388202 -22864 388258 -22808
rect 388326 -22864 388382 -22808
rect 388450 -22864 388506 -22808
rect 387954 -22988 388010 -22932
rect 388078 -22988 388134 -22932
rect 388202 -22988 388258 -22932
rect 388326 -22988 388382 -22932
rect 388450 -22988 388506 -22932
rect 387954 -23112 388010 -23056
rect 388078 -23112 388134 -23056
rect 388202 -23112 388258 -23056
rect 388326 -23112 388382 -23056
rect 388450 -23112 388506 -23056
rect 387954 -23236 388010 -23180
rect 388078 -23236 388134 -23180
rect 388202 -23236 388258 -23180
rect 388326 -23236 388382 -23180
rect 388450 -23236 388506 -23180
rect 387954 -23360 388010 -23304
rect 388078 -23360 388134 -23304
rect 388202 -23360 388258 -23304
rect 388326 -23360 388382 -23304
rect 388450 -23360 388506 -23304
rect 387954 -23484 388010 -23428
rect 388078 -23484 388134 -23428
rect 388202 -23484 388258 -23428
rect 388326 -23484 388382 -23428
rect 388450 -23484 388506 -23428
rect 387954 -23608 388010 -23552
rect 388078 -23608 388134 -23552
rect 388202 -23608 388258 -23552
rect 388326 -23608 388382 -23552
rect 388450 -23608 388506 -23552
rect 387954 -23732 388010 -23676
rect 388078 -23732 388134 -23676
rect 388202 -23732 388258 -23676
rect 388326 -23732 388382 -23676
rect 388450 -23732 388506 -23676
rect 387954 -23856 388010 -23800
rect 388078 -23856 388134 -23800
rect 388202 -23856 388258 -23800
rect 388326 -23856 388382 -23800
rect 388450 -23856 388506 -23800
rect 387954 -23980 388010 -23924
rect 388078 -23980 388134 -23924
rect 388202 -23980 388258 -23924
rect 388326 -23980 388382 -23924
rect 388450 -23980 388506 -23924
rect 387954 -24104 388010 -24048
rect 388078 -24104 388134 -24048
rect 388202 -24104 388258 -24048
rect 388326 -24104 388382 -24048
rect 388450 -24104 388506 -24048
rect 387954 -24228 388010 -24172
rect 388078 -24228 388134 -24172
rect 388202 -24228 388258 -24172
rect 388326 -24228 388382 -24172
rect 388450 -24228 388506 -24172
rect 387954 -24352 388010 -24296
rect 388078 -24352 388134 -24296
rect 388202 -24352 388258 -24296
rect 388326 -24352 388382 -24296
rect 388450 -24352 388506 -24296
rect 387954 -24476 388010 -24420
rect 388078 -24476 388134 -24420
rect 388202 -24476 388258 -24420
rect 388326 -24476 388382 -24420
rect 388450 -24476 388506 -24420
rect 387954 -24600 388010 -24544
rect 388078 -24600 388134 -24544
rect 388202 -24600 388258 -24544
rect 388326 -24600 388382 -24544
rect 388450 -24600 388506 -24544
rect 387954 -24724 388010 -24668
rect 388078 -24724 388134 -24668
rect 388202 -24724 388258 -24668
rect 388326 -24724 388382 -24668
rect 388450 -24724 388506 -24668
rect 387954 -24848 388010 -24792
rect 388078 -24848 388134 -24792
rect 388202 -24848 388258 -24792
rect 388326 -24848 388382 -24792
rect 388450 -24848 388506 -24792
rect 387954 -24972 388010 -24916
rect 388078 -24972 388134 -24916
rect 388202 -24972 388258 -24916
rect 388326 -24972 388382 -24916
rect 388450 -24972 388506 -24916
rect 387954 -25096 388010 -25040
rect 388078 -25096 388134 -25040
rect 388202 -25096 388258 -25040
rect 388326 -25096 388382 -25040
rect 388450 -25096 388506 -25040
rect 387954 -25220 388010 -25164
rect 388078 -25220 388134 -25164
rect 388202 -25220 388258 -25164
rect 388326 -25220 388382 -25164
rect 388450 -25220 388506 -25164
rect 387954 -25344 388010 -25288
rect 388078 -25344 388134 -25288
rect 388202 -25344 388258 -25288
rect 388326 -25344 388382 -25288
rect 388450 -25344 388506 -25288
rect 387954 -25468 388010 -25412
rect 388078 -25468 388134 -25412
rect 388202 -25468 388258 -25412
rect 388326 -25468 388382 -25412
rect 388450 -25468 388506 -25412
rect 387954 -25592 388010 -25536
rect 388078 -25592 388134 -25536
rect 388202 -25592 388258 -25536
rect 388326 -25592 388382 -25536
rect 388450 -25592 388506 -25536
rect 388981 -13736 389037 -13680
rect 389123 -13736 389179 -13680
rect 388981 -13878 389037 -13822
rect 389123 -13878 389179 -13822
rect 388981 -14020 389037 -13964
rect 389123 -14020 389179 -13964
rect 388981 -14162 389037 -14106
rect 389123 -14162 389179 -14106
rect 388981 -14304 389037 -14248
rect 389123 -14304 389179 -14248
rect 388981 -14446 389037 -14390
rect 389123 -14446 389179 -14390
rect 388981 -14588 389037 -14532
rect 389123 -14588 389179 -14532
rect 388981 -14730 389037 -14674
rect 389123 -14730 389179 -14674
rect 388981 -14872 389037 -14816
rect 389123 -14872 389179 -14816
rect 388981 -15014 389037 -14958
rect 389123 -15014 389179 -14958
rect 388981 -15156 389037 -15100
rect 389123 -15156 389179 -15100
rect 388981 -15298 389037 -15242
rect 389123 -15298 389179 -15242
rect 388981 -15440 389037 -15384
rect 389123 -15440 389179 -15384
rect 388981 -15582 389037 -15526
rect 389123 -15582 389179 -15526
rect 388981 -15724 389037 -15668
rect 389123 -15724 389179 -15668
rect 388981 -15866 389037 -15810
rect 389123 -15866 389179 -15810
rect 388981 -16008 389037 -15952
rect 389123 -16008 389179 -15952
rect 388981 -16150 389037 -16094
rect 389123 -16150 389179 -16094
rect 388981 -16292 389037 -16236
rect 389123 -16292 389179 -16236
rect 388981 -16434 389037 -16378
rect 389123 -16434 389179 -16378
rect 388981 -16576 389037 -16520
rect 389123 -16576 389179 -16520
rect 388981 -16718 389037 -16662
rect 389123 -16718 389179 -16662
rect 388981 -16860 389037 -16804
rect 389123 -16860 389179 -16804
rect 388981 -17002 389037 -16946
rect 389123 -17002 389179 -16946
rect 388981 -17144 389037 -17088
rect 389123 -17144 389179 -17088
rect 388981 -17286 389037 -17230
rect 389123 -17286 389179 -17230
rect 388981 -17428 389037 -17372
rect 389123 -17428 389179 -17372
rect 388981 -17570 389037 -17514
rect 389123 -17570 389179 -17514
rect 388981 -17712 389037 -17656
rect 389123 -17712 389179 -17656
rect 388981 -17854 389037 -17798
rect 389123 -17854 389179 -17798
rect 388981 -17996 389037 -17940
rect 389123 -17996 389179 -17940
rect 388981 -18138 389037 -18082
rect 389123 -18138 389179 -18082
rect 388981 -18280 389037 -18224
rect 389123 -18280 389179 -18224
rect 388981 -18422 389037 -18366
rect 389123 -18422 389179 -18366
rect 388981 -18564 389037 -18508
rect 389123 -18564 389179 -18508
rect 388981 -18706 389037 -18650
rect 389123 -18706 389179 -18650
rect 388981 -18848 389037 -18792
rect 389123 -18848 389179 -18792
rect 388981 -18990 389037 -18934
rect 389123 -18990 389179 -18934
rect 388981 -19132 389037 -19076
rect 389123 -19132 389179 -19076
rect 388981 -19274 389037 -19218
rect 389123 -19274 389179 -19218
rect 388981 -19416 389037 -19360
rect 389123 -19416 389179 -19360
rect 388981 -19558 389037 -19502
rect 389123 -19558 389179 -19502
rect 388981 -19700 389037 -19644
rect 389123 -19700 389179 -19644
rect 388981 -19842 389037 -19786
rect 389123 -19842 389179 -19786
rect 388981 -19984 389037 -19928
rect 389123 -19984 389179 -19928
rect 388981 -20126 389037 -20070
rect 389123 -20126 389179 -20070
rect 388981 -20268 389037 -20212
rect 389123 -20268 389179 -20212
rect 388981 -20410 389037 -20354
rect 389123 -20410 389179 -20354
rect 388981 -20552 389037 -20496
rect 389123 -20552 389179 -20496
rect 388981 -20694 389037 -20638
rect 389123 -20694 389179 -20638
rect 388981 -20836 389037 -20780
rect 389123 -20836 389179 -20780
rect 388981 -20978 389037 -20922
rect 389123 -20978 389179 -20922
rect 388981 -21120 389037 -21064
rect 389123 -21120 389179 -21064
rect 388981 -21262 389037 -21206
rect 389123 -21262 389179 -21206
rect 388981 -21404 389037 -21348
rect 389123 -21404 389179 -21348
rect 388981 -21546 389037 -21490
rect 389123 -21546 389179 -21490
rect 388981 -21688 389037 -21632
rect 389123 -21688 389179 -21632
rect 388981 -21830 389037 -21774
rect 389123 -21830 389179 -21774
rect 388981 -21972 389037 -21916
rect 389123 -21972 389179 -21916
rect 388981 -22114 389037 -22058
rect 389123 -22114 389179 -22058
rect 388981 -22256 389037 -22200
rect 389123 -22256 389179 -22200
rect 388981 -22398 389037 -22342
rect 389123 -22398 389179 -22342
rect 388981 -22540 389037 -22484
rect 389123 -22540 389179 -22484
rect 388981 -22682 389037 -22626
rect 389123 -22682 389179 -22626
rect 388981 -22824 389037 -22768
rect 389123 -22824 389179 -22768
rect 388981 -22966 389037 -22910
rect 389123 -22966 389179 -22910
rect 388981 -23108 389037 -23052
rect 389123 -23108 389179 -23052
rect 388981 -23250 389037 -23194
rect 389123 -23250 389179 -23194
rect 388981 -23392 389037 -23336
rect 389123 -23392 389179 -23336
rect 388981 -23534 389037 -23478
rect 389123 -23534 389179 -23478
rect 388981 -23676 389037 -23620
rect 389123 -23676 389179 -23620
rect 388981 -23818 389037 -23762
rect 389123 -23818 389179 -23762
rect 388981 -23960 389037 -23904
rect 389123 -23960 389179 -23904
rect 388981 -24102 389037 -24046
rect 389123 -24102 389179 -24046
rect 388981 -24244 389037 -24188
rect 389123 -24244 389179 -24188
rect 388981 -24386 389037 -24330
rect 389123 -24386 389179 -24330
rect 388981 -24528 389037 -24472
rect 389123 -24528 389179 -24472
rect 388981 -24670 389037 -24614
rect 389123 -24670 389179 -24614
rect 388981 -24812 389037 -24756
rect 389123 -24812 389179 -24756
rect 388981 -24954 389037 -24898
rect 389123 -24954 389179 -24898
rect 388981 -25096 389037 -25040
rect 389123 -25096 389179 -25040
rect 388981 -25238 389037 -25182
rect 389123 -25238 389179 -25182
rect 388981 -25380 389037 -25324
rect 389123 -25380 389179 -25324
rect 388981 -25522 389037 -25466
rect 389123 -25522 389179 -25466
rect 389382 -13736 389438 -13680
rect 389524 -13736 389580 -13680
rect 389382 -13878 389438 -13822
rect 389524 -13878 389580 -13822
rect 389382 -14020 389438 -13964
rect 389524 -14020 389580 -13964
rect 389382 -14162 389438 -14106
rect 389524 -14162 389580 -14106
rect 389382 -14304 389438 -14248
rect 389524 -14304 389580 -14248
rect 389382 -14446 389438 -14390
rect 389524 -14446 389580 -14390
rect 389382 -14588 389438 -14532
rect 389524 -14588 389580 -14532
rect 389382 -14730 389438 -14674
rect 389524 -14730 389580 -14674
rect 389382 -14872 389438 -14816
rect 389524 -14872 389580 -14816
rect 389382 -15014 389438 -14958
rect 389524 -15014 389580 -14958
rect 389382 -15156 389438 -15100
rect 389524 -15156 389580 -15100
rect 389382 -15298 389438 -15242
rect 389524 -15298 389580 -15242
rect 389382 -15440 389438 -15384
rect 389524 -15440 389580 -15384
rect 389382 -15582 389438 -15526
rect 389524 -15582 389580 -15526
rect 389382 -15724 389438 -15668
rect 389524 -15724 389580 -15668
rect 389382 -15866 389438 -15810
rect 389524 -15866 389580 -15810
rect 389382 -16008 389438 -15952
rect 389524 -16008 389580 -15952
rect 389382 -16150 389438 -16094
rect 389524 -16150 389580 -16094
rect 389382 -16292 389438 -16236
rect 389524 -16292 389580 -16236
rect 389382 -16434 389438 -16378
rect 389524 -16434 389580 -16378
rect 389382 -16576 389438 -16520
rect 389524 -16576 389580 -16520
rect 389382 -16718 389438 -16662
rect 389524 -16718 389580 -16662
rect 389382 -16860 389438 -16804
rect 389524 -16860 389580 -16804
rect 389382 -17002 389438 -16946
rect 389524 -17002 389580 -16946
rect 389382 -17144 389438 -17088
rect 389524 -17144 389580 -17088
rect 389382 -17286 389438 -17230
rect 389524 -17286 389580 -17230
rect 389382 -17428 389438 -17372
rect 389524 -17428 389580 -17372
rect 389382 -17570 389438 -17514
rect 389524 -17570 389580 -17514
rect 389382 -17712 389438 -17656
rect 389524 -17712 389580 -17656
rect 389382 -17854 389438 -17798
rect 389524 -17854 389580 -17798
rect 389382 -17996 389438 -17940
rect 389524 -17996 389580 -17940
rect 389382 -18138 389438 -18082
rect 389524 -18138 389580 -18082
rect 389382 -18280 389438 -18224
rect 389524 -18280 389580 -18224
rect 389382 -18422 389438 -18366
rect 389524 -18422 389580 -18366
rect 389382 -18564 389438 -18508
rect 389524 -18564 389580 -18508
rect 389382 -18706 389438 -18650
rect 389524 -18706 389580 -18650
rect 389382 -18848 389438 -18792
rect 389524 -18848 389580 -18792
rect 389382 -18990 389438 -18934
rect 389524 -18990 389580 -18934
rect 389382 -19132 389438 -19076
rect 389524 -19132 389580 -19076
rect 389382 -19274 389438 -19218
rect 389524 -19274 389580 -19218
rect 389382 -19416 389438 -19360
rect 389524 -19416 389580 -19360
rect 389382 -19558 389438 -19502
rect 389524 -19558 389580 -19502
rect 389382 -19700 389438 -19644
rect 389524 -19700 389580 -19644
rect 389382 -19842 389438 -19786
rect 389524 -19842 389580 -19786
rect 389382 -19984 389438 -19928
rect 389524 -19984 389580 -19928
rect 389382 -20126 389438 -20070
rect 389524 -20126 389580 -20070
rect 389382 -20268 389438 -20212
rect 389524 -20268 389580 -20212
rect 389382 -20410 389438 -20354
rect 389524 -20410 389580 -20354
rect 389382 -20552 389438 -20496
rect 389524 -20552 389580 -20496
rect 389382 -20694 389438 -20638
rect 389524 -20694 389580 -20638
rect 389382 -20836 389438 -20780
rect 389524 -20836 389580 -20780
rect 389382 -20978 389438 -20922
rect 389524 -20978 389580 -20922
rect 389382 -21120 389438 -21064
rect 389524 -21120 389580 -21064
rect 389382 -21262 389438 -21206
rect 389524 -21262 389580 -21206
rect 389382 -21404 389438 -21348
rect 389524 -21404 389580 -21348
rect 389382 -21546 389438 -21490
rect 389524 -21546 389580 -21490
rect 389382 -21688 389438 -21632
rect 389524 -21688 389580 -21632
rect 389382 -21830 389438 -21774
rect 389524 -21830 389580 -21774
rect 389382 -21972 389438 -21916
rect 389524 -21972 389580 -21916
rect 389382 -22114 389438 -22058
rect 389524 -22114 389580 -22058
rect 389382 -22256 389438 -22200
rect 389524 -22256 389580 -22200
rect 389382 -22398 389438 -22342
rect 389524 -22398 389580 -22342
rect 389382 -22540 389438 -22484
rect 389524 -22540 389580 -22484
rect 389382 -22682 389438 -22626
rect 389524 -22682 389580 -22626
rect 389382 -22824 389438 -22768
rect 389524 -22824 389580 -22768
rect 389382 -22966 389438 -22910
rect 389524 -22966 389580 -22910
rect 389382 -23108 389438 -23052
rect 389524 -23108 389580 -23052
rect 389382 -23250 389438 -23194
rect 389524 -23250 389580 -23194
rect 389382 -23392 389438 -23336
rect 389524 -23392 389580 -23336
rect 389382 -23534 389438 -23478
rect 389524 -23534 389580 -23478
rect 389382 -23676 389438 -23620
rect 389524 -23676 389580 -23620
rect 389382 -23818 389438 -23762
rect 389524 -23818 389580 -23762
rect 389382 -23960 389438 -23904
rect 389524 -23960 389580 -23904
rect 389382 -24102 389438 -24046
rect 389524 -24102 389580 -24046
rect 389382 -24244 389438 -24188
rect 389524 -24244 389580 -24188
rect 389382 -24386 389438 -24330
rect 389524 -24386 389580 -24330
rect 389382 -24528 389438 -24472
rect 389524 -24528 389580 -24472
rect 389382 -24670 389438 -24614
rect 389524 -24670 389580 -24614
rect 389382 -24812 389438 -24756
rect 389524 -24812 389580 -24756
rect 389382 -24954 389438 -24898
rect 389524 -24954 389580 -24898
rect 389382 -25096 389438 -25040
rect 389524 -25096 389580 -25040
rect 389382 -25238 389438 -25182
rect 389524 -25238 389580 -25182
rect 389382 -25380 389438 -25324
rect 389524 -25380 389580 -25324
rect 389382 -25522 389438 -25466
rect 389524 -25522 389580 -25466
rect 389782 -13736 389838 -13680
rect 389924 -13736 389980 -13680
rect 389782 -13878 389838 -13822
rect 389924 -13878 389980 -13822
rect 389782 -14020 389838 -13964
rect 389924 -14020 389980 -13964
rect 389782 -14162 389838 -14106
rect 389924 -14162 389980 -14106
rect 389782 -14304 389838 -14248
rect 389924 -14304 389980 -14248
rect 389782 -14446 389838 -14390
rect 389924 -14446 389980 -14390
rect 389782 -14588 389838 -14532
rect 389924 -14588 389980 -14532
rect 389782 -14730 389838 -14674
rect 389924 -14730 389980 -14674
rect 389782 -14872 389838 -14816
rect 389924 -14872 389980 -14816
rect 389782 -15014 389838 -14958
rect 389924 -15014 389980 -14958
rect 389782 -15156 389838 -15100
rect 389924 -15156 389980 -15100
rect 389782 -15298 389838 -15242
rect 389924 -15298 389980 -15242
rect 389782 -15440 389838 -15384
rect 389924 -15440 389980 -15384
rect 389782 -15582 389838 -15526
rect 389924 -15582 389980 -15526
rect 389782 -15724 389838 -15668
rect 389924 -15724 389980 -15668
rect 389782 -15866 389838 -15810
rect 389924 -15866 389980 -15810
rect 389782 -16008 389838 -15952
rect 389924 -16008 389980 -15952
rect 389782 -16150 389838 -16094
rect 389924 -16150 389980 -16094
rect 389782 -16292 389838 -16236
rect 389924 -16292 389980 -16236
rect 389782 -16434 389838 -16378
rect 389924 -16434 389980 -16378
rect 389782 -16576 389838 -16520
rect 389924 -16576 389980 -16520
rect 389782 -16718 389838 -16662
rect 389924 -16718 389980 -16662
rect 389782 -16860 389838 -16804
rect 389924 -16860 389980 -16804
rect 389782 -17002 389838 -16946
rect 389924 -17002 389980 -16946
rect 389782 -17144 389838 -17088
rect 389924 -17144 389980 -17088
rect 389782 -17286 389838 -17230
rect 389924 -17286 389980 -17230
rect 389782 -17428 389838 -17372
rect 389924 -17428 389980 -17372
rect 389782 -17570 389838 -17514
rect 389924 -17570 389980 -17514
rect 389782 -17712 389838 -17656
rect 389924 -17712 389980 -17656
rect 389782 -17854 389838 -17798
rect 389924 -17854 389980 -17798
rect 389782 -17996 389838 -17940
rect 389924 -17996 389980 -17940
rect 389782 -18138 389838 -18082
rect 389924 -18138 389980 -18082
rect 389782 -18280 389838 -18224
rect 389924 -18280 389980 -18224
rect 389782 -18422 389838 -18366
rect 389924 -18422 389980 -18366
rect 389782 -18564 389838 -18508
rect 389924 -18564 389980 -18508
rect 389782 -18706 389838 -18650
rect 389924 -18706 389980 -18650
rect 389782 -18848 389838 -18792
rect 389924 -18848 389980 -18792
rect 389782 -18990 389838 -18934
rect 389924 -18990 389980 -18934
rect 389782 -19132 389838 -19076
rect 389924 -19132 389980 -19076
rect 389782 -19274 389838 -19218
rect 389924 -19274 389980 -19218
rect 389782 -19416 389838 -19360
rect 389924 -19416 389980 -19360
rect 389782 -19558 389838 -19502
rect 389924 -19558 389980 -19502
rect 389782 -19700 389838 -19644
rect 389924 -19700 389980 -19644
rect 389782 -19842 389838 -19786
rect 389924 -19842 389980 -19786
rect 389782 -19984 389838 -19928
rect 389924 -19984 389980 -19928
rect 389782 -20126 389838 -20070
rect 389924 -20126 389980 -20070
rect 389782 -20268 389838 -20212
rect 389924 -20268 389980 -20212
rect 389782 -20410 389838 -20354
rect 389924 -20410 389980 -20354
rect 389782 -20552 389838 -20496
rect 389924 -20552 389980 -20496
rect 389782 -20694 389838 -20638
rect 389924 -20694 389980 -20638
rect 389782 -20836 389838 -20780
rect 389924 -20836 389980 -20780
rect 389782 -20978 389838 -20922
rect 389924 -20978 389980 -20922
rect 389782 -21120 389838 -21064
rect 389924 -21120 389980 -21064
rect 389782 -21262 389838 -21206
rect 389924 -21262 389980 -21206
rect 389782 -21404 389838 -21348
rect 389924 -21404 389980 -21348
rect 389782 -21546 389838 -21490
rect 389924 -21546 389980 -21490
rect 389782 -21688 389838 -21632
rect 389924 -21688 389980 -21632
rect 389782 -21830 389838 -21774
rect 389924 -21830 389980 -21774
rect 389782 -21972 389838 -21916
rect 389924 -21972 389980 -21916
rect 389782 -22114 389838 -22058
rect 389924 -22114 389980 -22058
rect 389782 -22256 389838 -22200
rect 389924 -22256 389980 -22200
rect 389782 -22398 389838 -22342
rect 389924 -22398 389980 -22342
rect 389782 -22540 389838 -22484
rect 389924 -22540 389980 -22484
rect 389782 -22682 389838 -22626
rect 389924 -22682 389980 -22626
rect 389782 -22824 389838 -22768
rect 389924 -22824 389980 -22768
rect 389782 -22966 389838 -22910
rect 389924 -22966 389980 -22910
rect 389782 -23108 389838 -23052
rect 389924 -23108 389980 -23052
rect 389782 -23250 389838 -23194
rect 389924 -23250 389980 -23194
rect 389782 -23392 389838 -23336
rect 389924 -23392 389980 -23336
rect 389782 -23534 389838 -23478
rect 389924 -23534 389980 -23478
rect 389782 -23676 389838 -23620
rect 389924 -23676 389980 -23620
rect 389782 -23818 389838 -23762
rect 389924 -23818 389980 -23762
rect 389782 -23960 389838 -23904
rect 389924 -23960 389980 -23904
rect 389782 -24102 389838 -24046
rect 389924 -24102 389980 -24046
rect 389782 -24244 389838 -24188
rect 389924 -24244 389980 -24188
rect 389782 -24386 389838 -24330
rect 389924 -24386 389980 -24330
rect 389782 -24528 389838 -24472
rect 389924 -24528 389980 -24472
rect 389782 -24670 389838 -24614
rect 389924 -24670 389980 -24614
rect 389782 -24812 389838 -24756
rect 389924 -24812 389980 -24756
rect 389782 -24954 389838 -24898
rect 389924 -24954 389980 -24898
rect 389782 -25096 389838 -25040
rect 389924 -25096 389980 -25040
rect 389782 -25238 389838 -25182
rect 389924 -25238 389980 -25182
rect 389782 -25380 389838 -25324
rect 389924 -25380 389980 -25324
rect 389782 -25522 389838 -25466
rect 389924 -25522 389980 -25466
rect 390179 -13736 390235 -13680
rect 390321 -13736 390377 -13680
rect 390179 -13878 390235 -13822
rect 390321 -13878 390377 -13822
rect 390179 -14020 390235 -13964
rect 390321 -14020 390377 -13964
rect 390179 -14162 390235 -14106
rect 390321 -14162 390377 -14106
rect 390179 -14304 390235 -14248
rect 390321 -14304 390377 -14248
rect 390179 -14446 390235 -14390
rect 390321 -14446 390377 -14390
rect 390179 -14588 390235 -14532
rect 390321 -14588 390377 -14532
rect 390179 -14730 390235 -14674
rect 390321 -14730 390377 -14674
rect 390179 -14872 390235 -14816
rect 390321 -14872 390377 -14816
rect 390179 -15014 390235 -14958
rect 390321 -15014 390377 -14958
rect 390179 -15156 390235 -15100
rect 390321 -15156 390377 -15100
rect 390179 -15298 390235 -15242
rect 390321 -15298 390377 -15242
rect 390179 -15440 390235 -15384
rect 390321 -15440 390377 -15384
rect 390179 -15582 390235 -15526
rect 390321 -15582 390377 -15526
rect 390179 -15724 390235 -15668
rect 390321 -15724 390377 -15668
rect 390179 -15866 390235 -15810
rect 390321 -15866 390377 -15810
rect 390179 -16008 390235 -15952
rect 390321 -16008 390377 -15952
rect 390179 -16150 390235 -16094
rect 390321 -16150 390377 -16094
rect 390179 -16292 390235 -16236
rect 390321 -16292 390377 -16236
rect 390179 -16434 390235 -16378
rect 390321 -16434 390377 -16378
rect 390179 -16576 390235 -16520
rect 390321 -16576 390377 -16520
rect 390179 -16718 390235 -16662
rect 390321 -16718 390377 -16662
rect 390179 -16860 390235 -16804
rect 390321 -16860 390377 -16804
rect 390179 -17002 390235 -16946
rect 390321 -17002 390377 -16946
rect 390179 -17144 390235 -17088
rect 390321 -17144 390377 -17088
rect 390179 -17286 390235 -17230
rect 390321 -17286 390377 -17230
rect 390179 -17428 390235 -17372
rect 390321 -17428 390377 -17372
rect 390179 -17570 390235 -17514
rect 390321 -17570 390377 -17514
rect 390179 -17712 390235 -17656
rect 390321 -17712 390377 -17656
rect 390179 -17854 390235 -17798
rect 390321 -17854 390377 -17798
rect 390179 -17996 390235 -17940
rect 390321 -17996 390377 -17940
rect 390179 -18138 390235 -18082
rect 390321 -18138 390377 -18082
rect 390179 -18280 390235 -18224
rect 390321 -18280 390377 -18224
rect 390179 -18422 390235 -18366
rect 390321 -18422 390377 -18366
rect 390179 -18564 390235 -18508
rect 390321 -18564 390377 -18508
rect 390179 -18706 390235 -18650
rect 390321 -18706 390377 -18650
rect 390179 -18848 390235 -18792
rect 390321 -18848 390377 -18792
rect 390179 -18990 390235 -18934
rect 390321 -18990 390377 -18934
rect 390179 -19132 390235 -19076
rect 390321 -19132 390377 -19076
rect 390179 -19274 390235 -19218
rect 390321 -19274 390377 -19218
rect 390179 -19416 390235 -19360
rect 390321 -19416 390377 -19360
rect 390179 -19558 390235 -19502
rect 390321 -19558 390377 -19502
rect 390179 -19700 390235 -19644
rect 390321 -19700 390377 -19644
rect 390179 -19842 390235 -19786
rect 390321 -19842 390377 -19786
rect 390179 -19984 390235 -19928
rect 390321 -19984 390377 -19928
rect 390179 -20126 390235 -20070
rect 390321 -20126 390377 -20070
rect 390179 -20268 390235 -20212
rect 390321 -20268 390377 -20212
rect 390179 -20410 390235 -20354
rect 390321 -20410 390377 -20354
rect 390179 -20552 390235 -20496
rect 390321 -20552 390377 -20496
rect 390179 -20694 390235 -20638
rect 390321 -20694 390377 -20638
rect 390179 -20836 390235 -20780
rect 390321 -20836 390377 -20780
rect 390179 -20978 390235 -20922
rect 390321 -20978 390377 -20922
rect 390179 -21120 390235 -21064
rect 390321 -21120 390377 -21064
rect 390179 -21262 390235 -21206
rect 390321 -21262 390377 -21206
rect 390179 -21404 390235 -21348
rect 390321 -21404 390377 -21348
rect 390179 -21546 390235 -21490
rect 390321 -21546 390377 -21490
rect 390179 -21688 390235 -21632
rect 390321 -21688 390377 -21632
rect 390179 -21830 390235 -21774
rect 390321 -21830 390377 -21774
rect 390179 -21972 390235 -21916
rect 390321 -21972 390377 -21916
rect 390179 -22114 390235 -22058
rect 390321 -22114 390377 -22058
rect 390179 -22256 390235 -22200
rect 390321 -22256 390377 -22200
rect 390179 -22398 390235 -22342
rect 390321 -22398 390377 -22342
rect 390179 -22540 390235 -22484
rect 390321 -22540 390377 -22484
rect 390179 -22682 390235 -22626
rect 390321 -22682 390377 -22626
rect 390179 -22824 390235 -22768
rect 390321 -22824 390377 -22768
rect 390179 -22966 390235 -22910
rect 390321 -22966 390377 -22910
rect 390179 -23108 390235 -23052
rect 390321 -23108 390377 -23052
rect 390179 -23250 390235 -23194
rect 390321 -23250 390377 -23194
rect 390179 -23392 390235 -23336
rect 390321 -23392 390377 -23336
rect 390179 -23534 390235 -23478
rect 390321 -23534 390377 -23478
rect 390179 -23676 390235 -23620
rect 390321 -23676 390377 -23620
rect 390179 -23818 390235 -23762
rect 390321 -23818 390377 -23762
rect 390179 -23960 390235 -23904
rect 390321 -23960 390377 -23904
rect 390179 -24102 390235 -24046
rect 390321 -24102 390377 -24046
rect 390179 -24244 390235 -24188
rect 390321 -24244 390377 -24188
rect 390179 -24386 390235 -24330
rect 390321 -24386 390377 -24330
rect 390179 -24528 390235 -24472
rect 390321 -24528 390377 -24472
rect 390179 -24670 390235 -24614
rect 390321 -24670 390377 -24614
rect 390179 -24812 390235 -24756
rect 390321 -24812 390377 -24756
rect 390179 -24954 390235 -24898
rect 390321 -24954 390377 -24898
rect 390179 -25096 390235 -25040
rect 390321 -25096 390377 -25040
rect 390179 -25238 390235 -25182
rect 390321 -25238 390377 -25182
rect 390179 -25380 390235 -25324
rect 390321 -25380 390377 -25324
rect 390179 -25522 390235 -25466
rect 390321 -25522 390377 -25466
rect 390576 -13736 390632 -13680
rect 390718 -13736 390774 -13680
rect 390576 -13878 390632 -13822
rect 390718 -13878 390774 -13822
rect 390576 -14020 390632 -13964
rect 390718 -14020 390774 -13964
rect 390576 -14162 390632 -14106
rect 390718 -14162 390774 -14106
rect 390576 -14304 390632 -14248
rect 390718 -14304 390774 -14248
rect 390576 -14446 390632 -14390
rect 390718 -14446 390774 -14390
rect 390576 -14588 390632 -14532
rect 390718 -14588 390774 -14532
rect 390576 -14730 390632 -14674
rect 390718 -14730 390774 -14674
rect 390576 -14872 390632 -14816
rect 390718 -14872 390774 -14816
rect 390576 -15014 390632 -14958
rect 390718 -15014 390774 -14958
rect 390576 -15156 390632 -15100
rect 390718 -15156 390774 -15100
rect 390576 -15298 390632 -15242
rect 390718 -15298 390774 -15242
rect 390576 -15440 390632 -15384
rect 390718 -15440 390774 -15384
rect 390576 -15582 390632 -15526
rect 390718 -15582 390774 -15526
rect 390576 -15724 390632 -15668
rect 390718 -15724 390774 -15668
rect 390576 -15866 390632 -15810
rect 390718 -15866 390774 -15810
rect 390576 -16008 390632 -15952
rect 390718 -16008 390774 -15952
rect 390576 -16150 390632 -16094
rect 390718 -16150 390774 -16094
rect 390576 -16292 390632 -16236
rect 390718 -16292 390774 -16236
rect 390576 -16434 390632 -16378
rect 390718 -16434 390774 -16378
rect 390576 -16576 390632 -16520
rect 390718 -16576 390774 -16520
rect 390576 -16718 390632 -16662
rect 390718 -16718 390774 -16662
rect 390576 -16860 390632 -16804
rect 390718 -16860 390774 -16804
rect 390576 -17002 390632 -16946
rect 390718 -17002 390774 -16946
rect 390576 -17144 390632 -17088
rect 390718 -17144 390774 -17088
rect 390576 -17286 390632 -17230
rect 390718 -17286 390774 -17230
rect 390576 -17428 390632 -17372
rect 390718 -17428 390774 -17372
rect 390576 -17570 390632 -17514
rect 390718 -17570 390774 -17514
rect 390576 -17712 390632 -17656
rect 390718 -17712 390774 -17656
rect 390576 -17854 390632 -17798
rect 390718 -17854 390774 -17798
rect 390576 -17996 390632 -17940
rect 390718 -17996 390774 -17940
rect 390576 -18138 390632 -18082
rect 390718 -18138 390774 -18082
rect 390576 -18280 390632 -18224
rect 390718 -18280 390774 -18224
rect 390576 -18422 390632 -18366
rect 390718 -18422 390774 -18366
rect 390576 -18564 390632 -18508
rect 390718 -18564 390774 -18508
rect 390576 -18706 390632 -18650
rect 390718 -18706 390774 -18650
rect 390576 -18848 390632 -18792
rect 390718 -18848 390774 -18792
rect 390576 -18990 390632 -18934
rect 390718 -18990 390774 -18934
rect 390576 -19132 390632 -19076
rect 390718 -19132 390774 -19076
rect 390576 -19274 390632 -19218
rect 390718 -19274 390774 -19218
rect 390576 -19416 390632 -19360
rect 390718 -19416 390774 -19360
rect 390576 -19558 390632 -19502
rect 390718 -19558 390774 -19502
rect 390576 -19700 390632 -19644
rect 390718 -19700 390774 -19644
rect 390576 -19842 390632 -19786
rect 390718 -19842 390774 -19786
rect 390576 -19984 390632 -19928
rect 390718 -19984 390774 -19928
rect 390576 -20126 390632 -20070
rect 390718 -20126 390774 -20070
rect 390576 -20268 390632 -20212
rect 390718 -20268 390774 -20212
rect 390576 -20410 390632 -20354
rect 390718 -20410 390774 -20354
rect 390576 -20552 390632 -20496
rect 390718 -20552 390774 -20496
rect 390576 -20694 390632 -20638
rect 390718 -20694 390774 -20638
rect 390576 -20836 390632 -20780
rect 390718 -20836 390774 -20780
rect 390576 -20978 390632 -20922
rect 390718 -20978 390774 -20922
rect 390576 -21120 390632 -21064
rect 390718 -21120 390774 -21064
rect 390576 -21262 390632 -21206
rect 390718 -21262 390774 -21206
rect 390576 -21404 390632 -21348
rect 390718 -21404 390774 -21348
rect 390576 -21546 390632 -21490
rect 390718 -21546 390774 -21490
rect 390576 -21688 390632 -21632
rect 390718 -21688 390774 -21632
rect 390576 -21830 390632 -21774
rect 390718 -21830 390774 -21774
rect 390576 -21972 390632 -21916
rect 390718 -21972 390774 -21916
rect 390576 -22114 390632 -22058
rect 390718 -22114 390774 -22058
rect 390576 -22256 390632 -22200
rect 390718 -22256 390774 -22200
rect 390576 -22398 390632 -22342
rect 390718 -22398 390774 -22342
rect 390576 -22540 390632 -22484
rect 390718 -22540 390774 -22484
rect 390576 -22682 390632 -22626
rect 390718 -22682 390774 -22626
rect 390576 -22824 390632 -22768
rect 390718 -22824 390774 -22768
rect 390576 -22966 390632 -22910
rect 390718 -22966 390774 -22910
rect 390576 -23108 390632 -23052
rect 390718 -23108 390774 -23052
rect 390576 -23250 390632 -23194
rect 390718 -23250 390774 -23194
rect 390576 -23392 390632 -23336
rect 390718 -23392 390774 -23336
rect 390576 -23534 390632 -23478
rect 390718 -23534 390774 -23478
rect 390576 -23676 390632 -23620
rect 390718 -23676 390774 -23620
rect 390576 -23818 390632 -23762
rect 390718 -23818 390774 -23762
rect 390576 -23960 390632 -23904
rect 390718 -23960 390774 -23904
rect 390576 -24102 390632 -24046
rect 390718 -24102 390774 -24046
rect 390576 -24244 390632 -24188
rect 390718 -24244 390774 -24188
rect 390576 -24386 390632 -24330
rect 390718 -24386 390774 -24330
rect 390576 -24528 390632 -24472
rect 390718 -24528 390774 -24472
rect 390576 -24670 390632 -24614
rect 390718 -24670 390774 -24614
rect 390576 -24812 390632 -24756
rect 390718 -24812 390774 -24756
rect 390576 -24954 390632 -24898
rect 390718 -24954 390774 -24898
rect 390576 -25096 390632 -25040
rect 390718 -25096 390774 -25040
rect 390576 -25238 390632 -25182
rect 390718 -25238 390774 -25182
rect 390576 -25380 390632 -25324
rect 390718 -25380 390774 -25324
rect 390576 -25522 390632 -25466
rect 390718 -25522 390774 -25466
rect 390980 -13736 391036 -13680
rect 391122 -13736 391178 -13680
rect 390980 -13878 391036 -13822
rect 391122 -13878 391178 -13822
rect 390980 -14020 391036 -13964
rect 391122 -14020 391178 -13964
rect 390980 -14162 391036 -14106
rect 391122 -14162 391178 -14106
rect 390980 -14304 391036 -14248
rect 391122 -14304 391178 -14248
rect 390980 -14446 391036 -14390
rect 391122 -14446 391178 -14390
rect 390980 -14588 391036 -14532
rect 391122 -14588 391178 -14532
rect 390980 -14730 391036 -14674
rect 391122 -14730 391178 -14674
rect 390980 -14872 391036 -14816
rect 391122 -14872 391178 -14816
rect 390980 -15014 391036 -14958
rect 391122 -15014 391178 -14958
rect 390980 -15156 391036 -15100
rect 391122 -15156 391178 -15100
rect 390980 -15298 391036 -15242
rect 391122 -15298 391178 -15242
rect 390980 -15440 391036 -15384
rect 391122 -15440 391178 -15384
rect 390980 -15582 391036 -15526
rect 391122 -15582 391178 -15526
rect 390980 -15724 391036 -15668
rect 391122 -15724 391178 -15668
rect 390980 -15866 391036 -15810
rect 391122 -15866 391178 -15810
rect 390980 -16008 391036 -15952
rect 391122 -16008 391178 -15952
rect 390980 -16150 391036 -16094
rect 391122 -16150 391178 -16094
rect 390980 -16292 391036 -16236
rect 391122 -16292 391178 -16236
rect 390980 -16434 391036 -16378
rect 391122 -16434 391178 -16378
rect 390980 -16576 391036 -16520
rect 391122 -16576 391178 -16520
rect 390980 -16718 391036 -16662
rect 391122 -16718 391178 -16662
rect 390980 -16860 391036 -16804
rect 391122 -16860 391178 -16804
rect 390980 -17002 391036 -16946
rect 391122 -17002 391178 -16946
rect 390980 -17144 391036 -17088
rect 391122 -17144 391178 -17088
rect 390980 -17286 391036 -17230
rect 391122 -17286 391178 -17230
rect 390980 -17428 391036 -17372
rect 391122 -17428 391178 -17372
rect 390980 -17570 391036 -17514
rect 391122 -17570 391178 -17514
rect 390980 -17712 391036 -17656
rect 391122 -17712 391178 -17656
rect 390980 -17854 391036 -17798
rect 391122 -17854 391178 -17798
rect 390980 -17996 391036 -17940
rect 391122 -17996 391178 -17940
rect 390980 -18138 391036 -18082
rect 391122 -18138 391178 -18082
rect 390980 -18280 391036 -18224
rect 391122 -18280 391178 -18224
rect 390980 -18422 391036 -18366
rect 391122 -18422 391178 -18366
rect 390980 -18564 391036 -18508
rect 391122 -18564 391178 -18508
rect 390980 -18706 391036 -18650
rect 391122 -18706 391178 -18650
rect 390980 -18848 391036 -18792
rect 391122 -18848 391178 -18792
rect 390980 -18990 391036 -18934
rect 391122 -18990 391178 -18934
rect 390980 -19132 391036 -19076
rect 391122 -19132 391178 -19076
rect 390980 -19274 391036 -19218
rect 391122 -19274 391178 -19218
rect 390980 -19416 391036 -19360
rect 391122 -19416 391178 -19360
rect 390980 -19558 391036 -19502
rect 391122 -19558 391178 -19502
rect 390980 -19700 391036 -19644
rect 391122 -19700 391178 -19644
rect 390980 -19842 391036 -19786
rect 391122 -19842 391178 -19786
rect 390980 -19984 391036 -19928
rect 391122 -19984 391178 -19928
rect 390980 -20126 391036 -20070
rect 391122 -20126 391178 -20070
rect 390980 -20268 391036 -20212
rect 391122 -20268 391178 -20212
rect 390980 -20410 391036 -20354
rect 391122 -20410 391178 -20354
rect 390980 -20552 391036 -20496
rect 391122 -20552 391178 -20496
rect 390980 -20694 391036 -20638
rect 391122 -20694 391178 -20638
rect 390980 -20836 391036 -20780
rect 391122 -20836 391178 -20780
rect 390980 -20978 391036 -20922
rect 391122 -20978 391178 -20922
rect 390980 -21120 391036 -21064
rect 391122 -21120 391178 -21064
rect 390980 -21262 391036 -21206
rect 391122 -21262 391178 -21206
rect 390980 -21404 391036 -21348
rect 391122 -21404 391178 -21348
rect 390980 -21546 391036 -21490
rect 391122 -21546 391178 -21490
rect 390980 -21688 391036 -21632
rect 391122 -21688 391178 -21632
rect 390980 -21830 391036 -21774
rect 391122 -21830 391178 -21774
rect 390980 -21972 391036 -21916
rect 391122 -21972 391178 -21916
rect 390980 -22114 391036 -22058
rect 391122 -22114 391178 -22058
rect 390980 -22256 391036 -22200
rect 391122 -22256 391178 -22200
rect 390980 -22398 391036 -22342
rect 391122 -22398 391178 -22342
rect 390980 -22540 391036 -22484
rect 391122 -22540 391178 -22484
rect 390980 -22682 391036 -22626
rect 391122 -22682 391178 -22626
rect 390980 -22824 391036 -22768
rect 391122 -22824 391178 -22768
rect 390980 -22966 391036 -22910
rect 391122 -22966 391178 -22910
rect 390980 -23108 391036 -23052
rect 391122 -23108 391178 -23052
rect 390980 -23250 391036 -23194
rect 391122 -23250 391178 -23194
rect 390980 -23392 391036 -23336
rect 391122 -23392 391178 -23336
rect 390980 -23534 391036 -23478
rect 391122 -23534 391178 -23478
rect 390980 -23676 391036 -23620
rect 391122 -23676 391178 -23620
rect 390980 -23818 391036 -23762
rect 391122 -23818 391178 -23762
rect 390980 -23960 391036 -23904
rect 391122 -23960 391178 -23904
rect 390980 -24102 391036 -24046
rect 391122 -24102 391178 -24046
rect 390980 -24244 391036 -24188
rect 391122 -24244 391178 -24188
rect 390980 -24386 391036 -24330
rect 391122 -24386 391178 -24330
rect 390980 -24528 391036 -24472
rect 391122 -24528 391178 -24472
rect 390980 -24670 391036 -24614
rect 391122 -24670 391178 -24614
rect 390980 -24812 391036 -24756
rect 391122 -24812 391178 -24756
rect 390980 -24954 391036 -24898
rect 391122 -24954 391178 -24898
rect 390980 -25096 391036 -25040
rect 391122 -25096 391178 -25040
rect 390980 -25238 391036 -25182
rect 391122 -25238 391178 -25182
rect 390980 -25380 391036 -25324
rect 391122 -25380 391178 -25324
rect 390980 -25522 391036 -25466
rect 391122 -25522 391178 -25466
rect 391376 -13736 391432 -13680
rect 391518 -13736 391574 -13680
rect 391376 -13878 391432 -13822
rect 391518 -13878 391574 -13822
rect 391376 -14020 391432 -13964
rect 391518 -14020 391574 -13964
rect 391376 -14162 391432 -14106
rect 391518 -14162 391574 -14106
rect 391376 -14304 391432 -14248
rect 391518 -14304 391574 -14248
rect 391376 -14446 391432 -14390
rect 391518 -14446 391574 -14390
rect 391376 -14588 391432 -14532
rect 391518 -14588 391574 -14532
rect 391376 -14730 391432 -14674
rect 391518 -14730 391574 -14674
rect 391376 -14872 391432 -14816
rect 391518 -14872 391574 -14816
rect 391376 -15014 391432 -14958
rect 391518 -15014 391574 -14958
rect 391376 -15156 391432 -15100
rect 391518 -15156 391574 -15100
rect 391376 -15298 391432 -15242
rect 391518 -15298 391574 -15242
rect 391376 -15440 391432 -15384
rect 391518 -15440 391574 -15384
rect 391376 -15582 391432 -15526
rect 391518 -15582 391574 -15526
rect 391376 -15724 391432 -15668
rect 391518 -15724 391574 -15668
rect 391376 -15866 391432 -15810
rect 391518 -15866 391574 -15810
rect 391376 -16008 391432 -15952
rect 391518 -16008 391574 -15952
rect 391376 -16150 391432 -16094
rect 391518 -16150 391574 -16094
rect 391376 -16292 391432 -16236
rect 391518 -16292 391574 -16236
rect 391376 -16434 391432 -16378
rect 391518 -16434 391574 -16378
rect 391376 -16576 391432 -16520
rect 391518 -16576 391574 -16520
rect 391376 -16718 391432 -16662
rect 391518 -16718 391574 -16662
rect 391376 -16860 391432 -16804
rect 391518 -16860 391574 -16804
rect 391376 -17002 391432 -16946
rect 391518 -17002 391574 -16946
rect 391376 -17144 391432 -17088
rect 391518 -17144 391574 -17088
rect 391376 -17286 391432 -17230
rect 391518 -17286 391574 -17230
rect 391376 -17428 391432 -17372
rect 391518 -17428 391574 -17372
rect 391376 -17570 391432 -17514
rect 391518 -17570 391574 -17514
rect 391376 -17712 391432 -17656
rect 391518 -17712 391574 -17656
rect 391376 -17854 391432 -17798
rect 391518 -17854 391574 -17798
rect 391376 -17996 391432 -17940
rect 391518 -17996 391574 -17940
rect 391376 -18138 391432 -18082
rect 391518 -18138 391574 -18082
rect 391376 -18280 391432 -18224
rect 391518 -18280 391574 -18224
rect 391376 -18422 391432 -18366
rect 391518 -18422 391574 -18366
rect 391376 -18564 391432 -18508
rect 391518 -18564 391574 -18508
rect 391376 -18706 391432 -18650
rect 391518 -18706 391574 -18650
rect 391376 -18848 391432 -18792
rect 391518 -18848 391574 -18792
rect 391376 -18990 391432 -18934
rect 391518 -18990 391574 -18934
rect 391376 -19132 391432 -19076
rect 391518 -19132 391574 -19076
rect 391376 -19274 391432 -19218
rect 391518 -19274 391574 -19218
rect 391376 -19416 391432 -19360
rect 391518 -19416 391574 -19360
rect 391376 -19558 391432 -19502
rect 391518 -19558 391574 -19502
rect 391376 -19700 391432 -19644
rect 391518 -19700 391574 -19644
rect 391376 -19842 391432 -19786
rect 391518 -19842 391574 -19786
rect 391376 -19984 391432 -19928
rect 391518 -19984 391574 -19928
rect 391376 -20126 391432 -20070
rect 391518 -20126 391574 -20070
rect 391376 -20268 391432 -20212
rect 391518 -20268 391574 -20212
rect 391376 -20410 391432 -20354
rect 391518 -20410 391574 -20354
rect 391376 -20552 391432 -20496
rect 391518 -20552 391574 -20496
rect 391376 -20694 391432 -20638
rect 391518 -20694 391574 -20638
rect 391376 -20836 391432 -20780
rect 391518 -20836 391574 -20780
rect 391376 -20978 391432 -20922
rect 391518 -20978 391574 -20922
rect 391376 -21120 391432 -21064
rect 391518 -21120 391574 -21064
rect 391376 -21262 391432 -21206
rect 391518 -21262 391574 -21206
rect 391376 -21404 391432 -21348
rect 391518 -21404 391574 -21348
rect 391376 -21546 391432 -21490
rect 391518 -21546 391574 -21490
rect 391376 -21688 391432 -21632
rect 391518 -21688 391574 -21632
rect 391376 -21830 391432 -21774
rect 391518 -21830 391574 -21774
rect 391376 -21972 391432 -21916
rect 391518 -21972 391574 -21916
rect 391376 -22114 391432 -22058
rect 391518 -22114 391574 -22058
rect 391376 -22256 391432 -22200
rect 391518 -22256 391574 -22200
rect 391376 -22398 391432 -22342
rect 391518 -22398 391574 -22342
rect 391376 -22540 391432 -22484
rect 391518 -22540 391574 -22484
rect 391376 -22682 391432 -22626
rect 391518 -22682 391574 -22626
rect 391376 -22824 391432 -22768
rect 391518 -22824 391574 -22768
rect 391376 -22966 391432 -22910
rect 391518 -22966 391574 -22910
rect 391376 -23108 391432 -23052
rect 391518 -23108 391574 -23052
rect 391376 -23250 391432 -23194
rect 391518 -23250 391574 -23194
rect 391376 -23392 391432 -23336
rect 391518 -23392 391574 -23336
rect 391376 -23534 391432 -23478
rect 391518 -23534 391574 -23478
rect 391376 -23676 391432 -23620
rect 391518 -23676 391574 -23620
rect 391376 -23818 391432 -23762
rect 391518 -23818 391574 -23762
rect 391376 -23960 391432 -23904
rect 391518 -23960 391574 -23904
rect 391376 -24102 391432 -24046
rect 391518 -24102 391574 -24046
rect 391376 -24244 391432 -24188
rect 391518 -24244 391574 -24188
rect 391376 -24386 391432 -24330
rect 391518 -24386 391574 -24330
rect 391376 -24528 391432 -24472
rect 391518 -24528 391574 -24472
rect 391376 -24670 391432 -24614
rect 391518 -24670 391574 -24614
rect 391376 -24812 391432 -24756
rect 391518 -24812 391574 -24756
rect 391376 -24954 391432 -24898
rect 391518 -24954 391574 -24898
rect 391376 -25096 391432 -25040
rect 391518 -25096 391574 -25040
rect 391376 -25238 391432 -25182
rect 391518 -25238 391574 -25182
rect 391376 -25380 391432 -25324
rect 391518 -25380 391574 -25324
rect 391376 -25522 391432 -25466
rect 391518 -25522 391574 -25466
rect 391776 -13736 391832 -13680
rect 391918 -13736 391974 -13680
rect 391776 -13878 391832 -13822
rect 391918 -13878 391974 -13822
rect 391776 -14020 391832 -13964
rect 391918 -14020 391974 -13964
rect 391776 -14162 391832 -14106
rect 391918 -14162 391974 -14106
rect 391776 -14304 391832 -14248
rect 391918 -14304 391974 -14248
rect 391776 -14446 391832 -14390
rect 391918 -14446 391974 -14390
rect 391776 -14588 391832 -14532
rect 391918 -14588 391974 -14532
rect 391776 -14730 391832 -14674
rect 391918 -14730 391974 -14674
rect 391776 -14872 391832 -14816
rect 391918 -14872 391974 -14816
rect 391776 -15014 391832 -14958
rect 391918 -15014 391974 -14958
rect 391776 -15156 391832 -15100
rect 391918 -15156 391974 -15100
rect 391776 -15298 391832 -15242
rect 391918 -15298 391974 -15242
rect 391776 -15440 391832 -15384
rect 391918 -15440 391974 -15384
rect 391776 -15582 391832 -15526
rect 391918 -15582 391974 -15526
rect 391776 -15724 391832 -15668
rect 391918 -15724 391974 -15668
rect 391776 -15866 391832 -15810
rect 391918 -15866 391974 -15810
rect 391776 -16008 391832 -15952
rect 391918 -16008 391974 -15952
rect 391776 -16150 391832 -16094
rect 391918 -16150 391974 -16094
rect 391776 -16292 391832 -16236
rect 391918 -16292 391974 -16236
rect 391776 -16434 391832 -16378
rect 391918 -16434 391974 -16378
rect 391776 -16576 391832 -16520
rect 391918 -16576 391974 -16520
rect 391776 -16718 391832 -16662
rect 391918 -16718 391974 -16662
rect 391776 -16860 391832 -16804
rect 391918 -16860 391974 -16804
rect 391776 -17002 391832 -16946
rect 391918 -17002 391974 -16946
rect 391776 -17144 391832 -17088
rect 391918 -17144 391974 -17088
rect 391776 -17286 391832 -17230
rect 391918 -17286 391974 -17230
rect 391776 -17428 391832 -17372
rect 391918 -17428 391974 -17372
rect 391776 -17570 391832 -17514
rect 391918 -17570 391974 -17514
rect 391776 -17712 391832 -17656
rect 391918 -17712 391974 -17656
rect 391776 -17854 391832 -17798
rect 391918 -17854 391974 -17798
rect 391776 -17996 391832 -17940
rect 391918 -17996 391974 -17940
rect 391776 -18138 391832 -18082
rect 391918 -18138 391974 -18082
rect 391776 -18280 391832 -18224
rect 391918 -18280 391974 -18224
rect 391776 -18422 391832 -18366
rect 391918 -18422 391974 -18366
rect 391776 -18564 391832 -18508
rect 391918 -18564 391974 -18508
rect 391776 -18706 391832 -18650
rect 391918 -18706 391974 -18650
rect 391776 -18848 391832 -18792
rect 391918 -18848 391974 -18792
rect 391776 -18990 391832 -18934
rect 391918 -18990 391974 -18934
rect 391776 -19132 391832 -19076
rect 391918 -19132 391974 -19076
rect 391776 -19274 391832 -19218
rect 391918 -19274 391974 -19218
rect 391776 -19416 391832 -19360
rect 391918 -19416 391974 -19360
rect 391776 -19558 391832 -19502
rect 391918 -19558 391974 -19502
rect 391776 -19700 391832 -19644
rect 391918 -19700 391974 -19644
rect 391776 -19842 391832 -19786
rect 391918 -19842 391974 -19786
rect 391776 -19984 391832 -19928
rect 391918 -19984 391974 -19928
rect 391776 -20126 391832 -20070
rect 391918 -20126 391974 -20070
rect 391776 -20268 391832 -20212
rect 391918 -20268 391974 -20212
rect 391776 -20410 391832 -20354
rect 391918 -20410 391974 -20354
rect 391776 -20552 391832 -20496
rect 391918 -20552 391974 -20496
rect 391776 -20694 391832 -20638
rect 391918 -20694 391974 -20638
rect 391776 -20836 391832 -20780
rect 391918 -20836 391974 -20780
rect 391776 -20978 391832 -20922
rect 391918 -20978 391974 -20922
rect 391776 -21120 391832 -21064
rect 391918 -21120 391974 -21064
rect 391776 -21262 391832 -21206
rect 391918 -21262 391974 -21206
rect 391776 -21404 391832 -21348
rect 391918 -21404 391974 -21348
rect 391776 -21546 391832 -21490
rect 391918 -21546 391974 -21490
rect 391776 -21688 391832 -21632
rect 391918 -21688 391974 -21632
rect 391776 -21830 391832 -21774
rect 391918 -21830 391974 -21774
rect 391776 -21972 391832 -21916
rect 391918 -21972 391974 -21916
rect 391776 -22114 391832 -22058
rect 391918 -22114 391974 -22058
rect 391776 -22256 391832 -22200
rect 391918 -22256 391974 -22200
rect 391776 -22398 391832 -22342
rect 391918 -22398 391974 -22342
rect 391776 -22540 391832 -22484
rect 391918 -22540 391974 -22484
rect 391776 -22682 391832 -22626
rect 391918 -22682 391974 -22626
rect 391776 -22824 391832 -22768
rect 391918 -22824 391974 -22768
rect 391776 -22966 391832 -22910
rect 391918 -22966 391974 -22910
rect 391776 -23108 391832 -23052
rect 391918 -23108 391974 -23052
rect 391776 -23250 391832 -23194
rect 391918 -23250 391974 -23194
rect 391776 -23392 391832 -23336
rect 391918 -23392 391974 -23336
rect 391776 -23534 391832 -23478
rect 391918 -23534 391974 -23478
rect 391776 -23676 391832 -23620
rect 391918 -23676 391974 -23620
rect 391776 -23818 391832 -23762
rect 391918 -23818 391974 -23762
rect 391776 -23960 391832 -23904
rect 391918 -23960 391974 -23904
rect 391776 -24102 391832 -24046
rect 391918 -24102 391974 -24046
rect 391776 -24244 391832 -24188
rect 391918 -24244 391974 -24188
rect 391776 -24386 391832 -24330
rect 391918 -24386 391974 -24330
rect 391776 -24528 391832 -24472
rect 391918 -24528 391974 -24472
rect 391776 -24670 391832 -24614
rect 391918 -24670 391974 -24614
rect 391776 -24812 391832 -24756
rect 391918 -24812 391974 -24756
rect 391776 -24954 391832 -24898
rect 391918 -24954 391974 -24898
rect 391776 -25096 391832 -25040
rect 391918 -25096 391974 -25040
rect 391776 -25238 391832 -25182
rect 391918 -25238 391974 -25182
rect 391776 -25380 391832 -25324
rect 391918 -25380 391974 -25324
rect 391776 -25522 391832 -25466
rect 391918 -25522 391974 -25466
rect 392173 -13736 392229 -13680
rect 392315 -13736 392371 -13680
rect 392173 -13878 392229 -13822
rect 392315 -13878 392371 -13822
rect 392173 -14020 392229 -13964
rect 392315 -14020 392371 -13964
rect 392173 -14162 392229 -14106
rect 392315 -14162 392371 -14106
rect 392173 -14304 392229 -14248
rect 392315 -14304 392371 -14248
rect 392173 -14446 392229 -14390
rect 392315 -14446 392371 -14390
rect 392173 -14588 392229 -14532
rect 392315 -14588 392371 -14532
rect 392173 -14730 392229 -14674
rect 392315 -14730 392371 -14674
rect 392173 -14872 392229 -14816
rect 392315 -14872 392371 -14816
rect 392173 -15014 392229 -14958
rect 392315 -15014 392371 -14958
rect 392173 -15156 392229 -15100
rect 392315 -15156 392371 -15100
rect 392173 -15298 392229 -15242
rect 392315 -15298 392371 -15242
rect 392173 -15440 392229 -15384
rect 392315 -15440 392371 -15384
rect 392173 -15582 392229 -15526
rect 392315 -15582 392371 -15526
rect 392173 -15724 392229 -15668
rect 392315 -15724 392371 -15668
rect 392173 -15866 392229 -15810
rect 392315 -15866 392371 -15810
rect 392173 -16008 392229 -15952
rect 392315 -16008 392371 -15952
rect 392173 -16150 392229 -16094
rect 392315 -16150 392371 -16094
rect 392173 -16292 392229 -16236
rect 392315 -16292 392371 -16236
rect 392173 -16434 392229 -16378
rect 392315 -16434 392371 -16378
rect 392173 -16576 392229 -16520
rect 392315 -16576 392371 -16520
rect 392173 -16718 392229 -16662
rect 392315 -16718 392371 -16662
rect 392173 -16860 392229 -16804
rect 392315 -16860 392371 -16804
rect 392173 -17002 392229 -16946
rect 392315 -17002 392371 -16946
rect 392173 -17144 392229 -17088
rect 392315 -17144 392371 -17088
rect 392173 -17286 392229 -17230
rect 392315 -17286 392371 -17230
rect 392173 -17428 392229 -17372
rect 392315 -17428 392371 -17372
rect 392173 -17570 392229 -17514
rect 392315 -17570 392371 -17514
rect 392173 -17712 392229 -17656
rect 392315 -17712 392371 -17656
rect 392173 -17854 392229 -17798
rect 392315 -17854 392371 -17798
rect 392173 -17996 392229 -17940
rect 392315 -17996 392371 -17940
rect 392173 -18138 392229 -18082
rect 392315 -18138 392371 -18082
rect 392173 -18280 392229 -18224
rect 392315 -18280 392371 -18224
rect 392173 -18422 392229 -18366
rect 392315 -18422 392371 -18366
rect 392173 -18564 392229 -18508
rect 392315 -18564 392371 -18508
rect 392173 -18706 392229 -18650
rect 392315 -18706 392371 -18650
rect 392173 -18848 392229 -18792
rect 392315 -18848 392371 -18792
rect 392173 -18990 392229 -18934
rect 392315 -18990 392371 -18934
rect 392173 -19132 392229 -19076
rect 392315 -19132 392371 -19076
rect 392173 -19274 392229 -19218
rect 392315 -19274 392371 -19218
rect 392173 -19416 392229 -19360
rect 392315 -19416 392371 -19360
rect 392173 -19558 392229 -19502
rect 392315 -19558 392371 -19502
rect 392173 -19700 392229 -19644
rect 392315 -19700 392371 -19644
rect 392173 -19842 392229 -19786
rect 392315 -19842 392371 -19786
rect 392173 -19984 392229 -19928
rect 392315 -19984 392371 -19928
rect 392173 -20126 392229 -20070
rect 392315 -20126 392371 -20070
rect 392173 -20268 392229 -20212
rect 392315 -20268 392371 -20212
rect 392173 -20410 392229 -20354
rect 392315 -20410 392371 -20354
rect 392173 -20552 392229 -20496
rect 392315 -20552 392371 -20496
rect 392173 -20694 392229 -20638
rect 392315 -20694 392371 -20638
rect 392173 -20836 392229 -20780
rect 392315 -20836 392371 -20780
rect 392173 -20978 392229 -20922
rect 392315 -20978 392371 -20922
rect 392173 -21120 392229 -21064
rect 392315 -21120 392371 -21064
rect 392173 -21262 392229 -21206
rect 392315 -21262 392371 -21206
rect 392173 -21404 392229 -21348
rect 392315 -21404 392371 -21348
rect 392173 -21546 392229 -21490
rect 392315 -21546 392371 -21490
rect 392173 -21688 392229 -21632
rect 392315 -21688 392371 -21632
rect 392173 -21830 392229 -21774
rect 392315 -21830 392371 -21774
rect 392173 -21972 392229 -21916
rect 392315 -21972 392371 -21916
rect 392173 -22114 392229 -22058
rect 392315 -22114 392371 -22058
rect 392173 -22256 392229 -22200
rect 392315 -22256 392371 -22200
rect 392173 -22398 392229 -22342
rect 392315 -22398 392371 -22342
rect 392173 -22540 392229 -22484
rect 392315 -22540 392371 -22484
rect 392173 -22682 392229 -22626
rect 392315 -22682 392371 -22626
rect 392173 -22824 392229 -22768
rect 392315 -22824 392371 -22768
rect 392173 -22966 392229 -22910
rect 392315 -22966 392371 -22910
rect 392173 -23108 392229 -23052
rect 392315 -23108 392371 -23052
rect 392173 -23250 392229 -23194
rect 392315 -23250 392371 -23194
rect 392173 -23392 392229 -23336
rect 392315 -23392 392371 -23336
rect 392173 -23534 392229 -23478
rect 392315 -23534 392371 -23478
rect 392173 -23676 392229 -23620
rect 392315 -23676 392371 -23620
rect 392173 -23818 392229 -23762
rect 392315 -23818 392371 -23762
rect 392173 -23960 392229 -23904
rect 392315 -23960 392371 -23904
rect 392173 -24102 392229 -24046
rect 392315 -24102 392371 -24046
rect 392173 -24244 392229 -24188
rect 392315 -24244 392371 -24188
rect 392173 -24386 392229 -24330
rect 392315 -24386 392371 -24330
rect 392173 -24528 392229 -24472
rect 392315 -24528 392371 -24472
rect 392173 -24670 392229 -24614
rect 392315 -24670 392371 -24614
rect 392173 -24812 392229 -24756
rect 392315 -24812 392371 -24756
rect 392173 -24954 392229 -24898
rect 392315 -24954 392371 -24898
rect 392173 -25096 392229 -25040
rect 392315 -25096 392371 -25040
rect 392173 -25238 392229 -25182
rect 392315 -25238 392371 -25182
rect 392173 -25380 392229 -25324
rect 392315 -25380 392371 -25324
rect 392173 -25522 392229 -25466
rect 392315 -25522 392371 -25466
rect 392578 -13736 392634 -13680
rect 392720 -13736 392776 -13680
rect 392578 -13878 392634 -13822
rect 392720 -13878 392776 -13822
rect 392578 -14020 392634 -13964
rect 392720 -14020 392776 -13964
rect 392578 -14162 392634 -14106
rect 392720 -14162 392776 -14106
rect 392578 -14304 392634 -14248
rect 392720 -14304 392776 -14248
rect 392578 -14446 392634 -14390
rect 392720 -14446 392776 -14390
rect 392578 -14588 392634 -14532
rect 392720 -14588 392776 -14532
rect 392578 -14730 392634 -14674
rect 392720 -14730 392776 -14674
rect 392578 -14872 392634 -14816
rect 392720 -14872 392776 -14816
rect 392578 -15014 392634 -14958
rect 392720 -15014 392776 -14958
rect 392578 -15156 392634 -15100
rect 392720 -15156 392776 -15100
rect 392578 -15298 392634 -15242
rect 392720 -15298 392776 -15242
rect 392578 -15440 392634 -15384
rect 392720 -15440 392776 -15384
rect 392578 -15582 392634 -15526
rect 392720 -15582 392776 -15526
rect 392578 -15724 392634 -15668
rect 392720 -15724 392776 -15668
rect 392578 -15866 392634 -15810
rect 392720 -15866 392776 -15810
rect 392578 -16008 392634 -15952
rect 392720 -16008 392776 -15952
rect 392578 -16150 392634 -16094
rect 392720 -16150 392776 -16094
rect 392578 -16292 392634 -16236
rect 392720 -16292 392776 -16236
rect 392578 -16434 392634 -16378
rect 392720 -16434 392776 -16378
rect 392578 -16576 392634 -16520
rect 392720 -16576 392776 -16520
rect 392578 -16718 392634 -16662
rect 392720 -16718 392776 -16662
rect 392578 -16860 392634 -16804
rect 392720 -16860 392776 -16804
rect 392578 -17002 392634 -16946
rect 392720 -17002 392776 -16946
rect 392578 -17144 392634 -17088
rect 392720 -17144 392776 -17088
rect 392578 -17286 392634 -17230
rect 392720 -17286 392776 -17230
rect 392578 -17428 392634 -17372
rect 392720 -17428 392776 -17372
rect 392578 -17570 392634 -17514
rect 392720 -17570 392776 -17514
rect 392578 -17712 392634 -17656
rect 392720 -17712 392776 -17656
rect 392578 -17854 392634 -17798
rect 392720 -17854 392776 -17798
rect 392578 -17996 392634 -17940
rect 392720 -17996 392776 -17940
rect 392578 -18138 392634 -18082
rect 392720 -18138 392776 -18082
rect 392578 -18280 392634 -18224
rect 392720 -18280 392776 -18224
rect 392578 -18422 392634 -18366
rect 392720 -18422 392776 -18366
rect 392578 -18564 392634 -18508
rect 392720 -18564 392776 -18508
rect 392578 -18706 392634 -18650
rect 392720 -18706 392776 -18650
rect 392578 -18848 392634 -18792
rect 392720 -18848 392776 -18792
rect 392578 -18990 392634 -18934
rect 392720 -18990 392776 -18934
rect 392578 -19132 392634 -19076
rect 392720 -19132 392776 -19076
rect 392578 -19274 392634 -19218
rect 392720 -19274 392776 -19218
rect 392578 -19416 392634 -19360
rect 392720 -19416 392776 -19360
rect 392578 -19558 392634 -19502
rect 392720 -19558 392776 -19502
rect 392578 -19700 392634 -19644
rect 392720 -19700 392776 -19644
rect 392578 -19842 392634 -19786
rect 392720 -19842 392776 -19786
rect 392578 -19984 392634 -19928
rect 392720 -19984 392776 -19928
rect 392578 -20126 392634 -20070
rect 392720 -20126 392776 -20070
rect 392578 -20268 392634 -20212
rect 392720 -20268 392776 -20212
rect 392578 -20410 392634 -20354
rect 392720 -20410 392776 -20354
rect 392578 -20552 392634 -20496
rect 392720 -20552 392776 -20496
rect 392578 -20694 392634 -20638
rect 392720 -20694 392776 -20638
rect 392578 -20836 392634 -20780
rect 392720 -20836 392776 -20780
rect 392578 -20978 392634 -20922
rect 392720 -20978 392776 -20922
rect 392578 -21120 392634 -21064
rect 392720 -21120 392776 -21064
rect 392578 -21262 392634 -21206
rect 392720 -21262 392776 -21206
rect 392578 -21404 392634 -21348
rect 392720 -21404 392776 -21348
rect 392578 -21546 392634 -21490
rect 392720 -21546 392776 -21490
rect 392578 -21688 392634 -21632
rect 392720 -21688 392776 -21632
rect 392578 -21830 392634 -21774
rect 392720 -21830 392776 -21774
rect 392578 -21972 392634 -21916
rect 392720 -21972 392776 -21916
rect 392578 -22114 392634 -22058
rect 392720 -22114 392776 -22058
rect 392578 -22256 392634 -22200
rect 392720 -22256 392776 -22200
rect 392578 -22398 392634 -22342
rect 392720 -22398 392776 -22342
rect 392578 -22540 392634 -22484
rect 392720 -22540 392776 -22484
rect 392578 -22682 392634 -22626
rect 392720 -22682 392776 -22626
rect 392578 -22824 392634 -22768
rect 392720 -22824 392776 -22768
rect 392578 -22966 392634 -22910
rect 392720 -22966 392776 -22910
rect 392578 -23108 392634 -23052
rect 392720 -23108 392776 -23052
rect 392578 -23250 392634 -23194
rect 392720 -23250 392776 -23194
rect 392578 -23392 392634 -23336
rect 392720 -23392 392776 -23336
rect 392578 -23534 392634 -23478
rect 392720 -23534 392776 -23478
rect 392578 -23676 392634 -23620
rect 392720 -23676 392776 -23620
rect 392578 -23818 392634 -23762
rect 392720 -23818 392776 -23762
rect 392578 -23960 392634 -23904
rect 392720 -23960 392776 -23904
rect 392578 -24102 392634 -24046
rect 392720 -24102 392776 -24046
rect 392578 -24244 392634 -24188
rect 392720 -24244 392776 -24188
rect 392578 -24386 392634 -24330
rect 392720 -24386 392776 -24330
rect 392578 -24528 392634 -24472
rect 392720 -24528 392776 -24472
rect 392578 -24670 392634 -24614
rect 392720 -24670 392776 -24614
rect 392578 -24812 392634 -24756
rect 392720 -24812 392776 -24756
rect 392578 -24954 392634 -24898
rect 392720 -24954 392776 -24898
rect 392578 -25096 392634 -25040
rect 392720 -25096 392776 -25040
rect 392578 -25238 392634 -25182
rect 392720 -25238 392776 -25182
rect 392578 -25380 392634 -25324
rect 392720 -25380 392776 -25324
rect 392578 -25522 392634 -25466
rect 392720 -25522 392776 -25466
rect 392978 -13736 393034 -13680
rect 393120 -13736 393176 -13680
rect 392978 -13878 393034 -13822
rect 393120 -13878 393176 -13822
rect 392978 -14020 393034 -13964
rect 393120 -14020 393176 -13964
rect 392978 -14162 393034 -14106
rect 393120 -14162 393176 -14106
rect 392978 -14304 393034 -14248
rect 393120 -14304 393176 -14248
rect 392978 -14446 393034 -14390
rect 393120 -14446 393176 -14390
rect 392978 -14588 393034 -14532
rect 393120 -14588 393176 -14532
rect 392978 -14730 393034 -14674
rect 393120 -14730 393176 -14674
rect 392978 -14872 393034 -14816
rect 393120 -14872 393176 -14816
rect 392978 -15014 393034 -14958
rect 393120 -15014 393176 -14958
rect 392978 -15156 393034 -15100
rect 393120 -15156 393176 -15100
rect 392978 -15298 393034 -15242
rect 393120 -15298 393176 -15242
rect 392978 -15440 393034 -15384
rect 393120 -15440 393176 -15384
rect 392978 -15582 393034 -15526
rect 393120 -15582 393176 -15526
rect 392978 -15724 393034 -15668
rect 393120 -15724 393176 -15668
rect 392978 -15866 393034 -15810
rect 393120 -15866 393176 -15810
rect 392978 -16008 393034 -15952
rect 393120 -16008 393176 -15952
rect 392978 -16150 393034 -16094
rect 393120 -16150 393176 -16094
rect 392978 -16292 393034 -16236
rect 393120 -16292 393176 -16236
rect 392978 -16434 393034 -16378
rect 393120 -16434 393176 -16378
rect 392978 -16576 393034 -16520
rect 393120 -16576 393176 -16520
rect 392978 -16718 393034 -16662
rect 393120 -16718 393176 -16662
rect 392978 -16860 393034 -16804
rect 393120 -16860 393176 -16804
rect 392978 -17002 393034 -16946
rect 393120 -17002 393176 -16946
rect 392978 -17144 393034 -17088
rect 393120 -17144 393176 -17088
rect 392978 -17286 393034 -17230
rect 393120 -17286 393176 -17230
rect 392978 -17428 393034 -17372
rect 393120 -17428 393176 -17372
rect 392978 -17570 393034 -17514
rect 393120 -17570 393176 -17514
rect 392978 -17712 393034 -17656
rect 393120 -17712 393176 -17656
rect 392978 -17854 393034 -17798
rect 393120 -17854 393176 -17798
rect 392978 -17996 393034 -17940
rect 393120 -17996 393176 -17940
rect 392978 -18138 393034 -18082
rect 393120 -18138 393176 -18082
rect 392978 -18280 393034 -18224
rect 393120 -18280 393176 -18224
rect 392978 -18422 393034 -18366
rect 393120 -18422 393176 -18366
rect 392978 -18564 393034 -18508
rect 393120 -18564 393176 -18508
rect 392978 -18706 393034 -18650
rect 393120 -18706 393176 -18650
rect 392978 -18848 393034 -18792
rect 393120 -18848 393176 -18792
rect 392978 -18990 393034 -18934
rect 393120 -18990 393176 -18934
rect 392978 -19132 393034 -19076
rect 393120 -19132 393176 -19076
rect 392978 -19274 393034 -19218
rect 393120 -19274 393176 -19218
rect 392978 -19416 393034 -19360
rect 393120 -19416 393176 -19360
rect 392978 -19558 393034 -19502
rect 393120 -19558 393176 -19502
rect 392978 -19700 393034 -19644
rect 393120 -19700 393176 -19644
rect 392978 -19842 393034 -19786
rect 393120 -19842 393176 -19786
rect 392978 -19984 393034 -19928
rect 393120 -19984 393176 -19928
rect 392978 -20126 393034 -20070
rect 393120 -20126 393176 -20070
rect 392978 -20268 393034 -20212
rect 393120 -20268 393176 -20212
rect 392978 -20410 393034 -20354
rect 393120 -20410 393176 -20354
rect 392978 -20552 393034 -20496
rect 393120 -20552 393176 -20496
rect 392978 -20694 393034 -20638
rect 393120 -20694 393176 -20638
rect 392978 -20836 393034 -20780
rect 393120 -20836 393176 -20780
rect 392978 -20978 393034 -20922
rect 393120 -20978 393176 -20922
rect 392978 -21120 393034 -21064
rect 393120 -21120 393176 -21064
rect 392978 -21262 393034 -21206
rect 393120 -21262 393176 -21206
rect 392978 -21404 393034 -21348
rect 393120 -21404 393176 -21348
rect 392978 -21546 393034 -21490
rect 393120 -21546 393176 -21490
rect 392978 -21688 393034 -21632
rect 393120 -21688 393176 -21632
rect 392978 -21830 393034 -21774
rect 393120 -21830 393176 -21774
rect 392978 -21972 393034 -21916
rect 393120 -21972 393176 -21916
rect 392978 -22114 393034 -22058
rect 393120 -22114 393176 -22058
rect 392978 -22256 393034 -22200
rect 393120 -22256 393176 -22200
rect 392978 -22398 393034 -22342
rect 393120 -22398 393176 -22342
rect 392978 -22540 393034 -22484
rect 393120 -22540 393176 -22484
rect 392978 -22682 393034 -22626
rect 393120 -22682 393176 -22626
rect 392978 -22824 393034 -22768
rect 393120 -22824 393176 -22768
rect 392978 -22966 393034 -22910
rect 393120 -22966 393176 -22910
rect 392978 -23108 393034 -23052
rect 393120 -23108 393176 -23052
rect 392978 -23250 393034 -23194
rect 393120 -23250 393176 -23194
rect 392978 -23392 393034 -23336
rect 393120 -23392 393176 -23336
rect 392978 -23534 393034 -23478
rect 393120 -23534 393176 -23478
rect 392978 -23676 393034 -23620
rect 393120 -23676 393176 -23620
rect 392978 -23818 393034 -23762
rect 393120 -23818 393176 -23762
rect 392978 -23960 393034 -23904
rect 393120 -23960 393176 -23904
rect 392978 -24102 393034 -24046
rect 393120 -24102 393176 -24046
rect 392978 -24244 393034 -24188
rect 393120 -24244 393176 -24188
rect 392978 -24386 393034 -24330
rect 393120 -24386 393176 -24330
rect 392978 -24528 393034 -24472
rect 393120 -24528 393176 -24472
rect 392978 -24670 393034 -24614
rect 393120 -24670 393176 -24614
rect 392978 -24812 393034 -24756
rect 393120 -24812 393176 -24756
rect 392978 -24954 393034 -24898
rect 393120 -24954 393176 -24898
rect 392978 -25096 393034 -25040
rect 393120 -25096 393176 -25040
rect 392978 -25238 393034 -25182
rect 393120 -25238 393176 -25182
rect 392978 -25380 393034 -25324
rect 393120 -25380 393176 -25324
rect 392978 -25522 393034 -25466
rect 393120 -25522 393176 -25466
rect 393383 -13736 393439 -13680
rect 393525 -13736 393581 -13680
rect 393383 -13878 393439 -13822
rect 393525 -13878 393581 -13822
rect 393383 -14020 393439 -13964
rect 393525 -14020 393581 -13964
rect 393383 -14162 393439 -14106
rect 393525 -14162 393581 -14106
rect 393383 -14304 393439 -14248
rect 393525 -14304 393581 -14248
rect 393383 -14446 393439 -14390
rect 393525 -14446 393581 -14390
rect 393383 -14588 393439 -14532
rect 393525 -14588 393581 -14532
rect 393383 -14730 393439 -14674
rect 393525 -14730 393581 -14674
rect 393383 -14872 393439 -14816
rect 393525 -14872 393581 -14816
rect 393383 -15014 393439 -14958
rect 393525 -15014 393581 -14958
rect 393383 -15156 393439 -15100
rect 393525 -15156 393581 -15100
rect 393383 -15298 393439 -15242
rect 393525 -15298 393581 -15242
rect 393383 -15440 393439 -15384
rect 393525 -15440 393581 -15384
rect 393383 -15582 393439 -15526
rect 393525 -15582 393581 -15526
rect 393383 -15724 393439 -15668
rect 393525 -15724 393581 -15668
rect 393383 -15866 393439 -15810
rect 393525 -15866 393581 -15810
rect 393383 -16008 393439 -15952
rect 393525 -16008 393581 -15952
rect 393383 -16150 393439 -16094
rect 393525 -16150 393581 -16094
rect 393383 -16292 393439 -16236
rect 393525 -16292 393581 -16236
rect 393383 -16434 393439 -16378
rect 393525 -16434 393581 -16378
rect 393383 -16576 393439 -16520
rect 393525 -16576 393581 -16520
rect 393383 -16718 393439 -16662
rect 393525 -16718 393581 -16662
rect 393383 -16860 393439 -16804
rect 393525 -16860 393581 -16804
rect 393383 -17002 393439 -16946
rect 393525 -17002 393581 -16946
rect 393383 -17144 393439 -17088
rect 393525 -17144 393581 -17088
rect 393383 -17286 393439 -17230
rect 393525 -17286 393581 -17230
rect 393383 -17428 393439 -17372
rect 393525 -17428 393581 -17372
rect 393383 -17570 393439 -17514
rect 393525 -17570 393581 -17514
rect 393383 -17712 393439 -17656
rect 393525 -17712 393581 -17656
rect 393383 -17854 393439 -17798
rect 393525 -17854 393581 -17798
rect 393383 -17996 393439 -17940
rect 393525 -17996 393581 -17940
rect 393383 -18138 393439 -18082
rect 393525 -18138 393581 -18082
rect 393383 -18280 393439 -18224
rect 393525 -18280 393581 -18224
rect 393383 -18422 393439 -18366
rect 393525 -18422 393581 -18366
rect 393383 -18564 393439 -18508
rect 393525 -18564 393581 -18508
rect 393383 -18706 393439 -18650
rect 393525 -18706 393581 -18650
rect 393383 -18848 393439 -18792
rect 393525 -18848 393581 -18792
rect 393383 -18990 393439 -18934
rect 393525 -18990 393581 -18934
rect 393383 -19132 393439 -19076
rect 393525 -19132 393581 -19076
rect 393383 -19274 393439 -19218
rect 393525 -19274 393581 -19218
rect 393383 -19416 393439 -19360
rect 393525 -19416 393581 -19360
rect 393383 -19558 393439 -19502
rect 393525 -19558 393581 -19502
rect 393383 -19700 393439 -19644
rect 393525 -19700 393581 -19644
rect 393383 -19842 393439 -19786
rect 393525 -19842 393581 -19786
rect 393383 -19984 393439 -19928
rect 393525 -19984 393581 -19928
rect 393383 -20126 393439 -20070
rect 393525 -20126 393581 -20070
rect 393383 -20268 393439 -20212
rect 393525 -20268 393581 -20212
rect 393383 -20410 393439 -20354
rect 393525 -20410 393581 -20354
rect 393383 -20552 393439 -20496
rect 393525 -20552 393581 -20496
rect 393383 -20694 393439 -20638
rect 393525 -20694 393581 -20638
rect 393383 -20836 393439 -20780
rect 393525 -20836 393581 -20780
rect 393383 -20978 393439 -20922
rect 393525 -20978 393581 -20922
rect 393383 -21120 393439 -21064
rect 393525 -21120 393581 -21064
rect 393383 -21262 393439 -21206
rect 393525 -21262 393581 -21206
rect 393383 -21404 393439 -21348
rect 393525 -21404 393581 -21348
rect 393383 -21546 393439 -21490
rect 393525 -21546 393581 -21490
rect 393383 -21688 393439 -21632
rect 393525 -21688 393581 -21632
rect 393383 -21830 393439 -21774
rect 393525 -21830 393581 -21774
rect 393383 -21972 393439 -21916
rect 393525 -21972 393581 -21916
rect 393383 -22114 393439 -22058
rect 393525 -22114 393581 -22058
rect 393383 -22256 393439 -22200
rect 393525 -22256 393581 -22200
rect 393383 -22398 393439 -22342
rect 393525 -22398 393581 -22342
rect 393383 -22540 393439 -22484
rect 393525 -22540 393581 -22484
rect 393383 -22682 393439 -22626
rect 393525 -22682 393581 -22626
rect 393383 -22824 393439 -22768
rect 393525 -22824 393581 -22768
rect 393383 -22966 393439 -22910
rect 393525 -22966 393581 -22910
rect 393383 -23108 393439 -23052
rect 393525 -23108 393581 -23052
rect 393383 -23250 393439 -23194
rect 393525 -23250 393581 -23194
rect 393383 -23392 393439 -23336
rect 393525 -23392 393581 -23336
rect 393383 -23534 393439 -23478
rect 393525 -23534 393581 -23478
rect 393383 -23676 393439 -23620
rect 393525 -23676 393581 -23620
rect 393383 -23818 393439 -23762
rect 393525 -23818 393581 -23762
rect 393383 -23960 393439 -23904
rect 393525 -23960 393581 -23904
rect 393383 -24102 393439 -24046
rect 393525 -24102 393581 -24046
rect 393383 -24244 393439 -24188
rect 393525 -24244 393581 -24188
rect 393383 -24386 393439 -24330
rect 393525 -24386 393581 -24330
rect 393383 -24528 393439 -24472
rect 393525 -24528 393581 -24472
rect 393383 -24670 393439 -24614
rect 393525 -24670 393581 -24614
rect 393383 -24812 393439 -24756
rect 393525 -24812 393581 -24756
rect 393383 -24954 393439 -24898
rect 393525 -24954 393581 -24898
rect 393383 -25096 393439 -25040
rect 393525 -25096 393581 -25040
rect 393383 -25238 393439 -25182
rect 393525 -25238 393581 -25182
rect 393383 -25380 393439 -25324
rect 393525 -25380 393581 -25324
rect 393383 -25522 393439 -25466
rect 393525 -25522 393581 -25466
rect 393780 -13736 393836 -13680
rect 393922 -13736 393978 -13680
rect 393780 -13878 393836 -13822
rect 393922 -13878 393978 -13822
rect 393780 -14020 393836 -13964
rect 393922 -14020 393978 -13964
rect 393780 -14162 393836 -14106
rect 393922 -14162 393978 -14106
rect 393780 -14304 393836 -14248
rect 393922 -14304 393978 -14248
rect 393780 -14446 393836 -14390
rect 393922 -14446 393978 -14390
rect 393780 -14588 393836 -14532
rect 393922 -14588 393978 -14532
rect 393780 -14730 393836 -14674
rect 393922 -14730 393978 -14674
rect 393780 -14872 393836 -14816
rect 393922 -14872 393978 -14816
rect 393780 -15014 393836 -14958
rect 393922 -15014 393978 -14958
rect 393780 -15156 393836 -15100
rect 393922 -15156 393978 -15100
rect 393780 -15298 393836 -15242
rect 393922 -15298 393978 -15242
rect 393780 -15440 393836 -15384
rect 393922 -15440 393978 -15384
rect 393780 -15582 393836 -15526
rect 393922 -15582 393978 -15526
rect 393780 -15724 393836 -15668
rect 393922 -15724 393978 -15668
rect 393780 -15866 393836 -15810
rect 393922 -15866 393978 -15810
rect 393780 -16008 393836 -15952
rect 393922 -16008 393978 -15952
rect 393780 -16150 393836 -16094
rect 393922 -16150 393978 -16094
rect 393780 -16292 393836 -16236
rect 393922 -16292 393978 -16236
rect 393780 -16434 393836 -16378
rect 393922 -16434 393978 -16378
rect 393780 -16576 393836 -16520
rect 393922 -16576 393978 -16520
rect 393780 -16718 393836 -16662
rect 393922 -16718 393978 -16662
rect 393780 -16860 393836 -16804
rect 393922 -16860 393978 -16804
rect 393780 -17002 393836 -16946
rect 393922 -17002 393978 -16946
rect 393780 -17144 393836 -17088
rect 393922 -17144 393978 -17088
rect 393780 -17286 393836 -17230
rect 393922 -17286 393978 -17230
rect 393780 -17428 393836 -17372
rect 393922 -17428 393978 -17372
rect 393780 -17570 393836 -17514
rect 393922 -17570 393978 -17514
rect 393780 -17712 393836 -17656
rect 393922 -17712 393978 -17656
rect 393780 -17854 393836 -17798
rect 393922 -17854 393978 -17798
rect 393780 -17996 393836 -17940
rect 393922 -17996 393978 -17940
rect 393780 -18138 393836 -18082
rect 393922 -18138 393978 -18082
rect 393780 -18280 393836 -18224
rect 393922 -18280 393978 -18224
rect 393780 -18422 393836 -18366
rect 393922 -18422 393978 -18366
rect 393780 -18564 393836 -18508
rect 393922 -18564 393978 -18508
rect 393780 -18706 393836 -18650
rect 393922 -18706 393978 -18650
rect 393780 -18848 393836 -18792
rect 393922 -18848 393978 -18792
rect 393780 -18990 393836 -18934
rect 393922 -18990 393978 -18934
rect 393780 -19132 393836 -19076
rect 393922 -19132 393978 -19076
rect 393780 -19274 393836 -19218
rect 393922 -19274 393978 -19218
rect 393780 -19416 393836 -19360
rect 393922 -19416 393978 -19360
rect 393780 -19558 393836 -19502
rect 393922 -19558 393978 -19502
rect 393780 -19700 393836 -19644
rect 393922 -19700 393978 -19644
rect 393780 -19842 393836 -19786
rect 393922 -19842 393978 -19786
rect 393780 -19984 393836 -19928
rect 393922 -19984 393978 -19928
rect 393780 -20126 393836 -20070
rect 393922 -20126 393978 -20070
rect 393780 -20268 393836 -20212
rect 393922 -20268 393978 -20212
rect 393780 -20410 393836 -20354
rect 393922 -20410 393978 -20354
rect 393780 -20552 393836 -20496
rect 393922 -20552 393978 -20496
rect 393780 -20694 393836 -20638
rect 393922 -20694 393978 -20638
rect 393780 -20836 393836 -20780
rect 393922 -20836 393978 -20780
rect 393780 -20978 393836 -20922
rect 393922 -20978 393978 -20922
rect 393780 -21120 393836 -21064
rect 393922 -21120 393978 -21064
rect 393780 -21262 393836 -21206
rect 393922 -21262 393978 -21206
rect 393780 -21404 393836 -21348
rect 393922 -21404 393978 -21348
rect 393780 -21546 393836 -21490
rect 393922 -21546 393978 -21490
rect 393780 -21688 393836 -21632
rect 393922 -21688 393978 -21632
rect 393780 -21830 393836 -21774
rect 393922 -21830 393978 -21774
rect 393780 -21972 393836 -21916
rect 393922 -21972 393978 -21916
rect 393780 -22114 393836 -22058
rect 393922 -22114 393978 -22058
rect 393780 -22256 393836 -22200
rect 393922 -22256 393978 -22200
rect 393780 -22398 393836 -22342
rect 393922 -22398 393978 -22342
rect 393780 -22540 393836 -22484
rect 393922 -22540 393978 -22484
rect 393780 -22682 393836 -22626
rect 393922 -22682 393978 -22626
rect 393780 -22824 393836 -22768
rect 393922 -22824 393978 -22768
rect 393780 -22966 393836 -22910
rect 393922 -22966 393978 -22910
rect 393780 -23108 393836 -23052
rect 393922 -23108 393978 -23052
rect 393780 -23250 393836 -23194
rect 393922 -23250 393978 -23194
rect 393780 -23392 393836 -23336
rect 393922 -23392 393978 -23336
rect 393780 -23534 393836 -23478
rect 393922 -23534 393978 -23478
rect 393780 -23676 393836 -23620
rect 393922 -23676 393978 -23620
rect 393780 -23818 393836 -23762
rect 393922 -23818 393978 -23762
rect 393780 -23960 393836 -23904
rect 393922 -23960 393978 -23904
rect 393780 -24102 393836 -24046
rect 393922 -24102 393978 -24046
rect 393780 -24244 393836 -24188
rect 393922 -24244 393978 -24188
rect 393780 -24386 393836 -24330
rect 393922 -24386 393978 -24330
rect 393780 -24528 393836 -24472
rect 393922 -24528 393978 -24472
rect 393780 -24670 393836 -24614
rect 393922 -24670 393978 -24614
rect 393780 -24812 393836 -24756
rect 393922 -24812 393978 -24756
rect 393780 -24954 393836 -24898
rect 393922 -24954 393978 -24898
rect 393780 -25096 393836 -25040
rect 393922 -25096 393978 -25040
rect 393780 -25238 393836 -25182
rect 393922 -25238 393978 -25182
rect 393780 -25380 393836 -25324
rect 393922 -25380 393978 -25324
rect 393780 -25522 393836 -25466
rect 393922 -25522 393978 -25466
rect 394177 -13736 394233 -13680
rect 394319 -13736 394375 -13680
rect 394177 -13878 394233 -13822
rect 394319 -13878 394375 -13822
rect 394177 -14020 394233 -13964
rect 394319 -14020 394375 -13964
rect 394177 -14162 394233 -14106
rect 394319 -14162 394375 -14106
rect 394177 -14304 394233 -14248
rect 394319 -14304 394375 -14248
rect 394177 -14446 394233 -14390
rect 394319 -14446 394375 -14390
rect 394177 -14588 394233 -14532
rect 394319 -14588 394375 -14532
rect 394177 -14730 394233 -14674
rect 394319 -14730 394375 -14674
rect 394177 -14872 394233 -14816
rect 394319 -14872 394375 -14816
rect 394177 -15014 394233 -14958
rect 394319 -15014 394375 -14958
rect 394177 -15156 394233 -15100
rect 394319 -15156 394375 -15100
rect 394177 -15298 394233 -15242
rect 394319 -15298 394375 -15242
rect 394177 -15440 394233 -15384
rect 394319 -15440 394375 -15384
rect 394177 -15582 394233 -15526
rect 394319 -15582 394375 -15526
rect 394177 -15724 394233 -15668
rect 394319 -15724 394375 -15668
rect 394177 -15866 394233 -15810
rect 394319 -15866 394375 -15810
rect 394177 -16008 394233 -15952
rect 394319 -16008 394375 -15952
rect 394177 -16150 394233 -16094
rect 394319 -16150 394375 -16094
rect 394177 -16292 394233 -16236
rect 394319 -16292 394375 -16236
rect 394177 -16434 394233 -16378
rect 394319 -16434 394375 -16378
rect 394177 -16576 394233 -16520
rect 394319 -16576 394375 -16520
rect 394177 -16718 394233 -16662
rect 394319 -16718 394375 -16662
rect 394177 -16860 394233 -16804
rect 394319 -16860 394375 -16804
rect 394177 -17002 394233 -16946
rect 394319 -17002 394375 -16946
rect 394177 -17144 394233 -17088
rect 394319 -17144 394375 -17088
rect 394177 -17286 394233 -17230
rect 394319 -17286 394375 -17230
rect 394177 -17428 394233 -17372
rect 394319 -17428 394375 -17372
rect 394177 -17570 394233 -17514
rect 394319 -17570 394375 -17514
rect 394177 -17712 394233 -17656
rect 394319 -17712 394375 -17656
rect 394177 -17854 394233 -17798
rect 394319 -17854 394375 -17798
rect 394177 -17996 394233 -17940
rect 394319 -17996 394375 -17940
rect 394177 -18138 394233 -18082
rect 394319 -18138 394375 -18082
rect 394177 -18280 394233 -18224
rect 394319 -18280 394375 -18224
rect 394177 -18422 394233 -18366
rect 394319 -18422 394375 -18366
rect 394177 -18564 394233 -18508
rect 394319 -18564 394375 -18508
rect 394177 -18706 394233 -18650
rect 394319 -18706 394375 -18650
rect 394177 -18848 394233 -18792
rect 394319 -18848 394375 -18792
rect 394177 -18990 394233 -18934
rect 394319 -18990 394375 -18934
rect 394177 -19132 394233 -19076
rect 394319 -19132 394375 -19076
rect 394177 -19274 394233 -19218
rect 394319 -19274 394375 -19218
rect 394177 -19416 394233 -19360
rect 394319 -19416 394375 -19360
rect 394177 -19558 394233 -19502
rect 394319 -19558 394375 -19502
rect 394177 -19700 394233 -19644
rect 394319 -19700 394375 -19644
rect 394177 -19842 394233 -19786
rect 394319 -19842 394375 -19786
rect 394177 -19984 394233 -19928
rect 394319 -19984 394375 -19928
rect 394177 -20126 394233 -20070
rect 394319 -20126 394375 -20070
rect 394177 -20268 394233 -20212
rect 394319 -20268 394375 -20212
rect 394177 -20410 394233 -20354
rect 394319 -20410 394375 -20354
rect 394177 -20552 394233 -20496
rect 394319 -20552 394375 -20496
rect 394177 -20694 394233 -20638
rect 394319 -20694 394375 -20638
rect 394177 -20836 394233 -20780
rect 394319 -20836 394375 -20780
rect 394177 -20978 394233 -20922
rect 394319 -20978 394375 -20922
rect 394177 -21120 394233 -21064
rect 394319 -21120 394375 -21064
rect 394177 -21262 394233 -21206
rect 394319 -21262 394375 -21206
rect 394177 -21404 394233 -21348
rect 394319 -21404 394375 -21348
rect 394177 -21546 394233 -21490
rect 394319 -21546 394375 -21490
rect 394177 -21688 394233 -21632
rect 394319 -21688 394375 -21632
rect 394177 -21830 394233 -21774
rect 394319 -21830 394375 -21774
rect 394177 -21972 394233 -21916
rect 394319 -21972 394375 -21916
rect 394177 -22114 394233 -22058
rect 394319 -22114 394375 -22058
rect 394177 -22256 394233 -22200
rect 394319 -22256 394375 -22200
rect 394177 -22398 394233 -22342
rect 394319 -22398 394375 -22342
rect 394177 -22540 394233 -22484
rect 394319 -22540 394375 -22484
rect 394177 -22682 394233 -22626
rect 394319 -22682 394375 -22626
rect 394177 -22824 394233 -22768
rect 394319 -22824 394375 -22768
rect 394177 -22966 394233 -22910
rect 394319 -22966 394375 -22910
rect 394177 -23108 394233 -23052
rect 394319 -23108 394375 -23052
rect 394177 -23250 394233 -23194
rect 394319 -23250 394375 -23194
rect 394177 -23392 394233 -23336
rect 394319 -23392 394375 -23336
rect 394177 -23534 394233 -23478
rect 394319 -23534 394375 -23478
rect 394177 -23676 394233 -23620
rect 394319 -23676 394375 -23620
rect 394177 -23818 394233 -23762
rect 394319 -23818 394375 -23762
rect 394177 -23960 394233 -23904
rect 394319 -23960 394375 -23904
rect 394177 -24102 394233 -24046
rect 394319 -24102 394375 -24046
rect 394177 -24244 394233 -24188
rect 394319 -24244 394375 -24188
rect 394177 -24386 394233 -24330
rect 394319 -24386 394375 -24330
rect 394177 -24528 394233 -24472
rect 394319 -24528 394375 -24472
rect 394177 -24670 394233 -24614
rect 394319 -24670 394375 -24614
rect 394177 -24812 394233 -24756
rect 394319 -24812 394375 -24756
rect 394177 -24954 394233 -24898
rect 394319 -24954 394375 -24898
rect 394177 -25096 394233 -25040
rect 394319 -25096 394375 -25040
rect 394177 -25238 394233 -25182
rect 394319 -25238 394375 -25182
rect 394177 -25380 394233 -25324
rect 394319 -25380 394375 -25324
rect 394177 -25522 394233 -25466
rect 394319 -25522 394375 -25466
rect 394580 -13736 394636 -13680
rect 394722 -13736 394778 -13680
rect 394580 -13878 394636 -13822
rect 394722 -13878 394778 -13822
rect 394580 -14020 394636 -13964
rect 394722 -14020 394778 -13964
rect 394580 -14162 394636 -14106
rect 394722 -14162 394778 -14106
rect 394580 -14304 394636 -14248
rect 394722 -14304 394778 -14248
rect 394580 -14446 394636 -14390
rect 394722 -14446 394778 -14390
rect 394580 -14588 394636 -14532
rect 394722 -14588 394778 -14532
rect 394580 -14730 394636 -14674
rect 394722 -14730 394778 -14674
rect 394580 -14872 394636 -14816
rect 394722 -14872 394778 -14816
rect 394580 -15014 394636 -14958
rect 394722 -15014 394778 -14958
rect 394580 -15156 394636 -15100
rect 394722 -15156 394778 -15100
rect 394580 -15298 394636 -15242
rect 394722 -15298 394778 -15242
rect 394580 -15440 394636 -15384
rect 394722 -15440 394778 -15384
rect 394580 -15582 394636 -15526
rect 394722 -15582 394778 -15526
rect 394580 -15724 394636 -15668
rect 394722 -15724 394778 -15668
rect 394580 -15866 394636 -15810
rect 394722 -15866 394778 -15810
rect 394580 -16008 394636 -15952
rect 394722 -16008 394778 -15952
rect 394580 -16150 394636 -16094
rect 394722 -16150 394778 -16094
rect 394580 -16292 394636 -16236
rect 394722 -16292 394778 -16236
rect 394580 -16434 394636 -16378
rect 394722 -16434 394778 -16378
rect 394580 -16576 394636 -16520
rect 394722 -16576 394778 -16520
rect 394580 -16718 394636 -16662
rect 394722 -16718 394778 -16662
rect 394580 -16860 394636 -16804
rect 394722 -16860 394778 -16804
rect 394580 -17002 394636 -16946
rect 394722 -17002 394778 -16946
rect 394580 -17144 394636 -17088
rect 394722 -17144 394778 -17088
rect 394580 -17286 394636 -17230
rect 394722 -17286 394778 -17230
rect 394580 -17428 394636 -17372
rect 394722 -17428 394778 -17372
rect 394580 -17570 394636 -17514
rect 394722 -17570 394778 -17514
rect 394580 -17712 394636 -17656
rect 394722 -17712 394778 -17656
rect 394580 -17854 394636 -17798
rect 394722 -17854 394778 -17798
rect 394580 -17996 394636 -17940
rect 394722 -17996 394778 -17940
rect 394580 -18138 394636 -18082
rect 394722 -18138 394778 -18082
rect 394580 -18280 394636 -18224
rect 394722 -18280 394778 -18224
rect 394580 -18422 394636 -18366
rect 394722 -18422 394778 -18366
rect 394580 -18564 394636 -18508
rect 394722 -18564 394778 -18508
rect 394580 -18706 394636 -18650
rect 394722 -18706 394778 -18650
rect 394580 -18848 394636 -18792
rect 394722 -18848 394778 -18792
rect 394580 -18990 394636 -18934
rect 394722 -18990 394778 -18934
rect 394580 -19132 394636 -19076
rect 394722 -19132 394778 -19076
rect 394580 -19274 394636 -19218
rect 394722 -19274 394778 -19218
rect 394580 -19416 394636 -19360
rect 394722 -19416 394778 -19360
rect 394580 -19558 394636 -19502
rect 394722 -19558 394778 -19502
rect 394580 -19700 394636 -19644
rect 394722 -19700 394778 -19644
rect 394580 -19842 394636 -19786
rect 394722 -19842 394778 -19786
rect 394580 -19984 394636 -19928
rect 394722 -19984 394778 -19928
rect 394580 -20126 394636 -20070
rect 394722 -20126 394778 -20070
rect 394580 -20268 394636 -20212
rect 394722 -20268 394778 -20212
rect 394580 -20410 394636 -20354
rect 394722 -20410 394778 -20354
rect 394580 -20552 394636 -20496
rect 394722 -20552 394778 -20496
rect 394580 -20694 394636 -20638
rect 394722 -20694 394778 -20638
rect 394580 -20836 394636 -20780
rect 394722 -20836 394778 -20780
rect 394580 -20978 394636 -20922
rect 394722 -20978 394778 -20922
rect 394580 -21120 394636 -21064
rect 394722 -21120 394778 -21064
rect 394580 -21262 394636 -21206
rect 394722 -21262 394778 -21206
rect 394580 -21404 394636 -21348
rect 394722 -21404 394778 -21348
rect 394580 -21546 394636 -21490
rect 394722 -21546 394778 -21490
rect 394580 -21688 394636 -21632
rect 394722 -21688 394778 -21632
rect 394580 -21830 394636 -21774
rect 394722 -21830 394778 -21774
rect 394580 -21972 394636 -21916
rect 394722 -21972 394778 -21916
rect 394580 -22114 394636 -22058
rect 394722 -22114 394778 -22058
rect 394580 -22256 394636 -22200
rect 394722 -22256 394778 -22200
rect 394580 -22398 394636 -22342
rect 394722 -22398 394778 -22342
rect 394580 -22540 394636 -22484
rect 394722 -22540 394778 -22484
rect 394580 -22682 394636 -22626
rect 394722 -22682 394778 -22626
rect 394580 -22824 394636 -22768
rect 394722 -22824 394778 -22768
rect 394580 -22966 394636 -22910
rect 394722 -22966 394778 -22910
rect 394580 -23108 394636 -23052
rect 394722 -23108 394778 -23052
rect 394580 -23250 394636 -23194
rect 394722 -23250 394778 -23194
rect 394580 -23392 394636 -23336
rect 394722 -23392 394778 -23336
rect 394580 -23534 394636 -23478
rect 394722 -23534 394778 -23478
rect 394580 -23676 394636 -23620
rect 394722 -23676 394778 -23620
rect 394580 -23818 394636 -23762
rect 394722 -23818 394778 -23762
rect 394580 -23960 394636 -23904
rect 394722 -23960 394778 -23904
rect 394580 -24102 394636 -24046
rect 394722 -24102 394778 -24046
rect 394580 -24244 394636 -24188
rect 394722 -24244 394778 -24188
rect 394580 -24386 394636 -24330
rect 394722 -24386 394778 -24330
rect 394580 -24528 394636 -24472
rect 394722 -24528 394778 -24472
rect 394580 -24670 394636 -24614
rect 394722 -24670 394778 -24614
rect 394580 -24812 394636 -24756
rect 394722 -24812 394778 -24756
rect 394580 -24954 394636 -24898
rect 394722 -24954 394778 -24898
rect 394580 -25096 394636 -25040
rect 394722 -25096 394778 -25040
rect 394580 -25238 394636 -25182
rect 394722 -25238 394778 -25182
rect 394580 -25380 394636 -25324
rect 394722 -25380 394778 -25324
rect 394580 -25522 394636 -25466
rect 394722 -25522 394778 -25466
rect 394982 -13736 395038 -13680
rect 395124 -13736 395180 -13680
rect 394982 -13878 395038 -13822
rect 395124 -13878 395180 -13822
rect 394982 -14020 395038 -13964
rect 395124 -14020 395180 -13964
rect 394982 -14162 395038 -14106
rect 395124 -14162 395180 -14106
rect 394982 -14304 395038 -14248
rect 395124 -14304 395180 -14248
rect 394982 -14446 395038 -14390
rect 395124 -14446 395180 -14390
rect 394982 -14588 395038 -14532
rect 395124 -14588 395180 -14532
rect 394982 -14730 395038 -14674
rect 395124 -14730 395180 -14674
rect 394982 -14872 395038 -14816
rect 395124 -14872 395180 -14816
rect 394982 -15014 395038 -14958
rect 395124 -15014 395180 -14958
rect 394982 -15156 395038 -15100
rect 395124 -15156 395180 -15100
rect 394982 -15298 395038 -15242
rect 395124 -15298 395180 -15242
rect 394982 -15440 395038 -15384
rect 395124 -15440 395180 -15384
rect 394982 -15582 395038 -15526
rect 395124 -15582 395180 -15526
rect 394982 -15724 395038 -15668
rect 395124 -15724 395180 -15668
rect 394982 -15866 395038 -15810
rect 395124 -15866 395180 -15810
rect 394982 -16008 395038 -15952
rect 395124 -16008 395180 -15952
rect 394982 -16150 395038 -16094
rect 395124 -16150 395180 -16094
rect 394982 -16292 395038 -16236
rect 395124 -16292 395180 -16236
rect 394982 -16434 395038 -16378
rect 395124 -16434 395180 -16378
rect 394982 -16576 395038 -16520
rect 395124 -16576 395180 -16520
rect 394982 -16718 395038 -16662
rect 395124 -16718 395180 -16662
rect 394982 -16860 395038 -16804
rect 395124 -16860 395180 -16804
rect 394982 -17002 395038 -16946
rect 395124 -17002 395180 -16946
rect 394982 -17144 395038 -17088
rect 395124 -17144 395180 -17088
rect 394982 -17286 395038 -17230
rect 395124 -17286 395180 -17230
rect 394982 -17428 395038 -17372
rect 395124 -17428 395180 -17372
rect 394982 -17570 395038 -17514
rect 395124 -17570 395180 -17514
rect 394982 -17712 395038 -17656
rect 395124 -17712 395180 -17656
rect 394982 -17854 395038 -17798
rect 395124 -17854 395180 -17798
rect 394982 -17996 395038 -17940
rect 395124 -17996 395180 -17940
rect 394982 -18138 395038 -18082
rect 395124 -18138 395180 -18082
rect 394982 -18280 395038 -18224
rect 395124 -18280 395180 -18224
rect 394982 -18422 395038 -18366
rect 395124 -18422 395180 -18366
rect 394982 -18564 395038 -18508
rect 395124 -18564 395180 -18508
rect 394982 -18706 395038 -18650
rect 395124 -18706 395180 -18650
rect 394982 -18848 395038 -18792
rect 395124 -18848 395180 -18792
rect 394982 -18990 395038 -18934
rect 395124 -18990 395180 -18934
rect 394982 -19132 395038 -19076
rect 395124 -19132 395180 -19076
rect 394982 -19274 395038 -19218
rect 395124 -19274 395180 -19218
rect 394982 -19416 395038 -19360
rect 395124 -19416 395180 -19360
rect 394982 -19558 395038 -19502
rect 395124 -19558 395180 -19502
rect 394982 -19700 395038 -19644
rect 395124 -19700 395180 -19644
rect 394982 -19842 395038 -19786
rect 395124 -19842 395180 -19786
rect 394982 -19984 395038 -19928
rect 395124 -19984 395180 -19928
rect 394982 -20126 395038 -20070
rect 395124 -20126 395180 -20070
rect 394982 -20268 395038 -20212
rect 395124 -20268 395180 -20212
rect 394982 -20410 395038 -20354
rect 395124 -20410 395180 -20354
rect 394982 -20552 395038 -20496
rect 395124 -20552 395180 -20496
rect 394982 -20694 395038 -20638
rect 395124 -20694 395180 -20638
rect 394982 -20836 395038 -20780
rect 395124 -20836 395180 -20780
rect 394982 -20978 395038 -20922
rect 395124 -20978 395180 -20922
rect 394982 -21120 395038 -21064
rect 395124 -21120 395180 -21064
rect 394982 -21262 395038 -21206
rect 395124 -21262 395180 -21206
rect 394982 -21404 395038 -21348
rect 395124 -21404 395180 -21348
rect 394982 -21546 395038 -21490
rect 395124 -21546 395180 -21490
rect 394982 -21688 395038 -21632
rect 395124 -21688 395180 -21632
rect 394982 -21830 395038 -21774
rect 395124 -21830 395180 -21774
rect 394982 -21972 395038 -21916
rect 395124 -21972 395180 -21916
rect 394982 -22114 395038 -22058
rect 395124 -22114 395180 -22058
rect 394982 -22256 395038 -22200
rect 395124 -22256 395180 -22200
rect 394982 -22398 395038 -22342
rect 395124 -22398 395180 -22342
rect 394982 -22540 395038 -22484
rect 395124 -22540 395180 -22484
rect 394982 -22682 395038 -22626
rect 395124 -22682 395180 -22626
rect 394982 -22824 395038 -22768
rect 395124 -22824 395180 -22768
rect 394982 -22966 395038 -22910
rect 395124 -22966 395180 -22910
rect 394982 -23108 395038 -23052
rect 395124 -23108 395180 -23052
rect 394982 -23250 395038 -23194
rect 395124 -23250 395180 -23194
rect 394982 -23392 395038 -23336
rect 395124 -23392 395180 -23336
rect 394982 -23534 395038 -23478
rect 395124 -23534 395180 -23478
rect 394982 -23676 395038 -23620
rect 395124 -23676 395180 -23620
rect 394982 -23818 395038 -23762
rect 395124 -23818 395180 -23762
rect 394982 -23960 395038 -23904
rect 395124 -23960 395180 -23904
rect 394982 -24102 395038 -24046
rect 395124 -24102 395180 -24046
rect 394982 -24244 395038 -24188
rect 395124 -24244 395180 -24188
rect 394982 -24386 395038 -24330
rect 395124 -24386 395180 -24330
rect 394982 -24528 395038 -24472
rect 395124 -24528 395180 -24472
rect 394982 -24670 395038 -24614
rect 395124 -24670 395180 -24614
rect 394982 -24812 395038 -24756
rect 395124 -24812 395180 -24756
rect 394982 -24954 395038 -24898
rect 395124 -24954 395180 -24898
rect 394982 -25096 395038 -25040
rect 395124 -25096 395180 -25040
rect 394982 -25238 395038 -25182
rect 395124 -25238 395180 -25182
rect 394982 -25380 395038 -25324
rect 395124 -25380 395180 -25324
rect 394982 -25522 395038 -25466
rect 395124 -25522 395180 -25466
rect 395385 -13736 395441 -13680
rect 395527 -13736 395583 -13680
rect 395385 -13878 395441 -13822
rect 395527 -13878 395583 -13822
rect 395385 -14020 395441 -13964
rect 395527 -14020 395583 -13964
rect 395385 -14162 395441 -14106
rect 395527 -14162 395583 -14106
rect 395385 -14304 395441 -14248
rect 395527 -14304 395583 -14248
rect 395385 -14446 395441 -14390
rect 395527 -14446 395583 -14390
rect 395385 -14588 395441 -14532
rect 395527 -14588 395583 -14532
rect 395385 -14730 395441 -14674
rect 395527 -14730 395583 -14674
rect 395385 -14872 395441 -14816
rect 395527 -14872 395583 -14816
rect 395385 -15014 395441 -14958
rect 395527 -15014 395583 -14958
rect 395385 -15156 395441 -15100
rect 395527 -15156 395583 -15100
rect 395385 -15298 395441 -15242
rect 395527 -15298 395583 -15242
rect 395385 -15440 395441 -15384
rect 395527 -15440 395583 -15384
rect 395385 -15582 395441 -15526
rect 395527 -15582 395583 -15526
rect 395385 -15724 395441 -15668
rect 395527 -15724 395583 -15668
rect 395385 -15866 395441 -15810
rect 395527 -15866 395583 -15810
rect 395385 -16008 395441 -15952
rect 395527 -16008 395583 -15952
rect 395385 -16150 395441 -16094
rect 395527 -16150 395583 -16094
rect 395385 -16292 395441 -16236
rect 395527 -16292 395583 -16236
rect 395385 -16434 395441 -16378
rect 395527 -16434 395583 -16378
rect 395385 -16576 395441 -16520
rect 395527 -16576 395583 -16520
rect 395385 -16718 395441 -16662
rect 395527 -16718 395583 -16662
rect 395385 -16860 395441 -16804
rect 395527 -16860 395583 -16804
rect 395385 -17002 395441 -16946
rect 395527 -17002 395583 -16946
rect 395385 -17144 395441 -17088
rect 395527 -17144 395583 -17088
rect 395385 -17286 395441 -17230
rect 395527 -17286 395583 -17230
rect 395385 -17428 395441 -17372
rect 395527 -17428 395583 -17372
rect 395385 -17570 395441 -17514
rect 395527 -17570 395583 -17514
rect 395385 -17712 395441 -17656
rect 395527 -17712 395583 -17656
rect 395385 -17854 395441 -17798
rect 395527 -17854 395583 -17798
rect 395385 -17996 395441 -17940
rect 395527 -17996 395583 -17940
rect 395385 -18138 395441 -18082
rect 395527 -18138 395583 -18082
rect 395385 -18280 395441 -18224
rect 395527 -18280 395583 -18224
rect 395385 -18422 395441 -18366
rect 395527 -18422 395583 -18366
rect 395385 -18564 395441 -18508
rect 395527 -18564 395583 -18508
rect 395385 -18706 395441 -18650
rect 395527 -18706 395583 -18650
rect 395385 -18848 395441 -18792
rect 395527 -18848 395583 -18792
rect 395385 -18990 395441 -18934
rect 395527 -18990 395583 -18934
rect 395385 -19132 395441 -19076
rect 395527 -19132 395583 -19076
rect 395385 -19274 395441 -19218
rect 395527 -19274 395583 -19218
rect 395385 -19416 395441 -19360
rect 395527 -19416 395583 -19360
rect 395385 -19558 395441 -19502
rect 395527 -19558 395583 -19502
rect 395385 -19700 395441 -19644
rect 395527 -19700 395583 -19644
rect 395385 -19842 395441 -19786
rect 395527 -19842 395583 -19786
rect 395385 -19984 395441 -19928
rect 395527 -19984 395583 -19928
rect 395385 -20126 395441 -20070
rect 395527 -20126 395583 -20070
rect 395385 -20268 395441 -20212
rect 395527 -20268 395583 -20212
rect 395385 -20410 395441 -20354
rect 395527 -20410 395583 -20354
rect 395385 -20552 395441 -20496
rect 395527 -20552 395583 -20496
rect 395385 -20694 395441 -20638
rect 395527 -20694 395583 -20638
rect 395385 -20836 395441 -20780
rect 395527 -20836 395583 -20780
rect 395385 -20978 395441 -20922
rect 395527 -20978 395583 -20922
rect 395385 -21120 395441 -21064
rect 395527 -21120 395583 -21064
rect 395385 -21262 395441 -21206
rect 395527 -21262 395583 -21206
rect 395385 -21404 395441 -21348
rect 395527 -21404 395583 -21348
rect 395385 -21546 395441 -21490
rect 395527 -21546 395583 -21490
rect 395385 -21688 395441 -21632
rect 395527 -21688 395583 -21632
rect 395385 -21830 395441 -21774
rect 395527 -21830 395583 -21774
rect 395385 -21972 395441 -21916
rect 395527 -21972 395583 -21916
rect 395385 -22114 395441 -22058
rect 395527 -22114 395583 -22058
rect 395385 -22256 395441 -22200
rect 395527 -22256 395583 -22200
rect 395385 -22398 395441 -22342
rect 395527 -22398 395583 -22342
rect 395385 -22540 395441 -22484
rect 395527 -22540 395583 -22484
rect 395385 -22682 395441 -22626
rect 395527 -22682 395583 -22626
rect 395385 -22824 395441 -22768
rect 395527 -22824 395583 -22768
rect 395385 -22966 395441 -22910
rect 395527 -22966 395583 -22910
rect 395385 -23108 395441 -23052
rect 395527 -23108 395583 -23052
rect 395385 -23250 395441 -23194
rect 395527 -23250 395583 -23194
rect 395385 -23392 395441 -23336
rect 395527 -23392 395583 -23336
rect 395385 -23534 395441 -23478
rect 395527 -23534 395583 -23478
rect 395385 -23676 395441 -23620
rect 395527 -23676 395583 -23620
rect 395385 -23818 395441 -23762
rect 395527 -23818 395583 -23762
rect 395385 -23960 395441 -23904
rect 395527 -23960 395583 -23904
rect 395385 -24102 395441 -24046
rect 395527 -24102 395583 -24046
rect 395385 -24244 395441 -24188
rect 395527 -24244 395583 -24188
rect 395385 -24386 395441 -24330
rect 395527 -24386 395583 -24330
rect 395385 -24528 395441 -24472
rect 395527 -24528 395583 -24472
rect 395385 -24670 395441 -24614
rect 395527 -24670 395583 -24614
rect 395385 -24812 395441 -24756
rect 395527 -24812 395583 -24756
rect 395385 -24954 395441 -24898
rect 395527 -24954 395583 -24898
rect 395385 -25096 395441 -25040
rect 395527 -25096 395583 -25040
rect 395385 -25238 395441 -25182
rect 395527 -25238 395583 -25182
rect 395385 -25380 395441 -25324
rect 395527 -25380 395583 -25324
rect 395385 -25522 395441 -25466
rect 395527 -25522 395583 -25466
rect 395779 -13736 395835 -13680
rect 395921 -13736 395977 -13680
rect 395779 -13878 395835 -13822
rect 395921 -13878 395977 -13822
rect 395779 -14020 395835 -13964
rect 395921 -14020 395977 -13964
rect 395779 -14162 395835 -14106
rect 395921 -14162 395977 -14106
rect 395779 -14304 395835 -14248
rect 395921 -14304 395977 -14248
rect 395779 -14446 395835 -14390
rect 395921 -14446 395977 -14390
rect 395779 -14588 395835 -14532
rect 395921 -14588 395977 -14532
rect 395779 -14730 395835 -14674
rect 395921 -14730 395977 -14674
rect 395779 -14872 395835 -14816
rect 395921 -14872 395977 -14816
rect 395779 -15014 395835 -14958
rect 395921 -15014 395977 -14958
rect 395779 -15156 395835 -15100
rect 395921 -15156 395977 -15100
rect 395779 -15298 395835 -15242
rect 395921 -15298 395977 -15242
rect 395779 -15440 395835 -15384
rect 395921 -15440 395977 -15384
rect 395779 -15582 395835 -15526
rect 395921 -15582 395977 -15526
rect 395779 -15724 395835 -15668
rect 395921 -15724 395977 -15668
rect 395779 -15866 395835 -15810
rect 395921 -15866 395977 -15810
rect 395779 -16008 395835 -15952
rect 395921 -16008 395977 -15952
rect 395779 -16150 395835 -16094
rect 395921 -16150 395977 -16094
rect 395779 -16292 395835 -16236
rect 395921 -16292 395977 -16236
rect 395779 -16434 395835 -16378
rect 395921 -16434 395977 -16378
rect 395779 -16576 395835 -16520
rect 395921 -16576 395977 -16520
rect 395779 -16718 395835 -16662
rect 395921 -16718 395977 -16662
rect 395779 -16860 395835 -16804
rect 395921 -16860 395977 -16804
rect 395779 -17002 395835 -16946
rect 395921 -17002 395977 -16946
rect 395779 -17144 395835 -17088
rect 395921 -17144 395977 -17088
rect 395779 -17286 395835 -17230
rect 395921 -17286 395977 -17230
rect 395779 -17428 395835 -17372
rect 395921 -17428 395977 -17372
rect 395779 -17570 395835 -17514
rect 395921 -17570 395977 -17514
rect 395779 -17712 395835 -17656
rect 395921 -17712 395977 -17656
rect 395779 -17854 395835 -17798
rect 395921 -17854 395977 -17798
rect 395779 -17996 395835 -17940
rect 395921 -17996 395977 -17940
rect 395779 -18138 395835 -18082
rect 395921 -18138 395977 -18082
rect 395779 -18280 395835 -18224
rect 395921 -18280 395977 -18224
rect 395779 -18422 395835 -18366
rect 395921 -18422 395977 -18366
rect 395779 -18564 395835 -18508
rect 395921 -18564 395977 -18508
rect 395779 -18706 395835 -18650
rect 395921 -18706 395977 -18650
rect 395779 -18848 395835 -18792
rect 395921 -18848 395977 -18792
rect 395779 -18990 395835 -18934
rect 395921 -18990 395977 -18934
rect 395779 -19132 395835 -19076
rect 395921 -19132 395977 -19076
rect 395779 -19274 395835 -19218
rect 395921 -19274 395977 -19218
rect 395779 -19416 395835 -19360
rect 395921 -19416 395977 -19360
rect 395779 -19558 395835 -19502
rect 395921 -19558 395977 -19502
rect 395779 -19700 395835 -19644
rect 395921 -19700 395977 -19644
rect 395779 -19842 395835 -19786
rect 395921 -19842 395977 -19786
rect 395779 -19984 395835 -19928
rect 395921 -19984 395977 -19928
rect 395779 -20126 395835 -20070
rect 395921 -20126 395977 -20070
rect 395779 -20268 395835 -20212
rect 395921 -20268 395977 -20212
rect 395779 -20410 395835 -20354
rect 395921 -20410 395977 -20354
rect 395779 -20552 395835 -20496
rect 395921 -20552 395977 -20496
rect 395779 -20694 395835 -20638
rect 395921 -20694 395977 -20638
rect 395779 -20836 395835 -20780
rect 395921 -20836 395977 -20780
rect 395779 -20978 395835 -20922
rect 395921 -20978 395977 -20922
rect 395779 -21120 395835 -21064
rect 395921 -21120 395977 -21064
rect 395779 -21262 395835 -21206
rect 395921 -21262 395977 -21206
rect 395779 -21404 395835 -21348
rect 395921 -21404 395977 -21348
rect 395779 -21546 395835 -21490
rect 395921 -21546 395977 -21490
rect 395779 -21688 395835 -21632
rect 395921 -21688 395977 -21632
rect 395779 -21830 395835 -21774
rect 395921 -21830 395977 -21774
rect 395779 -21972 395835 -21916
rect 395921 -21972 395977 -21916
rect 395779 -22114 395835 -22058
rect 395921 -22114 395977 -22058
rect 395779 -22256 395835 -22200
rect 395921 -22256 395977 -22200
rect 395779 -22398 395835 -22342
rect 395921 -22398 395977 -22342
rect 395779 -22540 395835 -22484
rect 395921 -22540 395977 -22484
rect 395779 -22682 395835 -22626
rect 395921 -22682 395977 -22626
rect 395779 -22824 395835 -22768
rect 395921 -22824 395977 -22768
rect 395779 -22966 395835 -22910
rect 395921 -22966 395977 -22910
rect 395779 -23108 395835 -23052
rect 395921 -23108 395977 -23052
rect 395779 -23250 395835 -23194
rect 395921 -23250 395977 -23194
rect 395779 -23392 395835 -23336
rect 395921 -23392 395977 -23336
rect 395779 -23534 395835 -23478
rect 395921 -23534 395977 -23478
rect 395779 -23676 395835 -23620
rect 395921 -23676 395977 -23620
rect 395779 -23818 395835 -23762
rect 395921 -23818 395977 -23762
rect 395779 -23960 395835 -23904
rect 395921 -23960 395977 -23904
rect 395779 -24102 395835 -24046
rect 395921 -24102 395977 -24046
rect 395779 -24244 395835 -24188
rect 395921 -24244 395977 -24188
rect 395779 -24386 395835 -24330
rect 395921 -24386 395977 -24330
rect 395779 -24528 395835 -24472
rect 395921 -24528 395977 -24472
rect 395779 -24670 395835 -24614
rect 395921 -24670 395977 -24614
rect 395779 -24812 395835 -24756
rect 395921 -24812 395977 -24756
rect 395779 -24954 395835 -24898
rect 395921 -24954 395977 -24898
rect 395779 -25096 395835 -25040
rect 395921 -25096 395977 -25040
rect 395779 -25238 395835 -25182
rect 395921 -25238 395977 -25182
rect 395779 -25380 395835 -25324
rect 395921 -25380 395977 -25324
rect 395779 -25522 395835 -25466
rect 395921 -25522 395977 -25466
rect 396180 -13736 396236 -13680
rect 396322 -13736 396378 -13680
rect 396180 -13878 396236 -13822
rect 396322 -13878 396378 -13822
rect 396180 -14020 396236 -13964
rect 396322 -14020 396378 -13964
rect 396180 -14162 396236 -14106
rect 396322 -14162 396378 -14106
rect 396180 -14304 396236 -14248
rect 396322 -14304 396378 -14248
rect 396180 -14446 396236 -14390
rect 396322 -14446 396378 -14390
rect 396180 -14588 396236 -14532
rect 396322 -14588 396378 -14532
rect 396180 -14730 396236 -14674
rect 396322 -14730 396378 -14674
rect 396180 -14872 396236 -14816
rect 396322 -14872 396378 -14816
rect 396180 -15014 396236 -14958
rect 396322 -15014 396378 -14958
rect 396180 -15156 396236 -15100
rect 396322 -15156 396378 -15100
rect 396180 -15298 396236 -15242
rect 396322 -15298 396378 -15242
rect 396180 -15440 396236 -15384
rect 396322 -15440 396378 -15384
rect 396180 -15582 396236 -15526
rect 396322 -15582 396378 -15526
rect 396180 -15724 396236 -15668
rect 396322 -15724 396378 -15668
rect 396180 -15866 396236 -15810
rect 396322 -15866 396378 -15810
rect 396180 -16008 396236 -15952
rect 396322 -16008 396378 -15952
rect 396180 -16150 396236 -16094
rect 396322 -16150 396378 -16094
rect 396180 -16292 396236 -16236
rect 396322 -16292 396378 -16236
rect 396180 -16434 396236 -16378
rect 396322 -16434 396378 -16378
rect 396180 -16576 396236 -16520
rect 396322 -16576 396378 -16520
rect 396180 -16718 396236 -16662
rect 396322 -16718 396378 -16662
rect 396180 -16860 396236 -16804
rect 396322 -16860 396378 -16804
rect 396180 -17002 396236 -16946
rect 396322 -17002 396378 -16946
rect 396180 -17144 396236 -17088
rect 396322 -17144 396378 -17088
rect 396180 -17286 396236 -17230
rect 396322 -17286 396378 -17230
rect 396180 -17428 396236 -17372
rect 396322 -17428 396378 -17372
rect 396180 -17570 396236 -17514
rect 396322 -17570 396378 -17514
rect 396180 -17712 396236 -17656
rect 396322 -17712 396378 -17656
rect 396180 -17854 396236 -17798
rect 396322 -17854 396378 -17798
rect 396180 -17996 396236 -17940
rect 396322 -17996 396378 -17940
rect 396180 -18138 396236 -18082
rect 396322 -18138 396378 -18082
rect 396180 -18280 396236 -18224
rect 396322 -18280 396378 -18224
rect 396180 -18422 396236 -18366
rect 396322 -18422 396378 -18366
rect 396180 -18564 396236 -18508
rect 396322 -18564 396378 -18508
rect 396180 -18706 396236 -18650
rect 396322 -18706 396378 -18650
rect 396180 -18848 396236 -18792
rect 396322 -18848 396378 -18792
rect 396180 -18990 396236 -18934
rect 396322 -18990 396378 -18934
rect 396180 -19132 396236 -19076
rect 396322 -19132 396378 -19076
rect 396180 -19274 396236 -19218
rect 396322 -19274 396378 -19218
rect 396180 -19416 396236 -19360
rect 396322 -19416 396378 -19360
rect 396180 -19558 396236 -19502
rect 396322 -19558 396378 -19502
rect 396180 -19700 396236 -19644
rect 396322 -19700 396378 -19644
rect 396180 -19842 396236 -19786
rect 396322 -19842 396378 -19786
rect 396180 -19984 396236 -19928
rect 396322 -19984 396378 -19928
rect 396180 -20126 396236 -20070
rect 396322 -20126 396378 -20070
rect 396180 -20268 396236 -20212
rect 396322 -20268 396378 -20212
rect 396180 -20410 396236 -20354
rect 396322 -20410 396378 -20354
rect 396180 -20552 396236 -20496
rect 396322 -20552 396378 -20496
rect 396180 -20694 396236 -20638
rect 396322 -20694 396378 -20638
rect 396180 -20836 396236 -20780
rect 396322 -20836 396378 -20780
rect 396180 -20978 396236 -20922
rect 396322 -20978 396378 -20922
rect 396180 -21120 396236 -21064
rect 396322 -21120 396378 -21064
rect 396180 -21262 396236 -21206
rect 396322 -21262 396378 -21206
rect 396180 -21404 396236 -21348
rect 396322 -21404 396378 -21348
rect 396180 -21546 396236 -21490
rect 396322 -21546 396378 -21490
rect 396180 -21688 396236 -21632
rect 396322 -21688 396378 -21632
rect 396180 -21830 396236 -21774
rect 396322 -21830 396378 -21774
rect 396180 -21972 396236 -21916
rect 396322 -21972 396378 -21916
rect 396180 -22114 396236 -22058
rect 396322 -22114 396378 -22058
rect 396180 -22256 396236 -22200
rect 396322 -22256 396378 -22200
rect 396180 -22398 396236 -22342
rect 396322 -22398 396378 -22342
rect 396180 -22540 396236 -22484
rect 396322 -22540 396378 -22484
rect 396180 -22682 396236 -22626
rect 396322 -22682 396378 -22626
rect 396180 -22824 396236 -22768
rect 396322 -22824 396378 -22768
rect 396180 -22966 396236 -22910
rect 396322 -22966 396378 -22910
rect 396180 -23108 396236 -23052
rect 396322 -23108 396378 -23052
rect 396180 -23250 396236 -23194
rect 396322 -23250 396378 -23194
rect 396180 -23392 396236 -23336
rect 396322 -23392 396378 -23336
rect 396180 -23534 396236 -23478
rect 396322 -23534 396378 -23478
rect 396180 -23676 396236 -23620
rect 396322 -23676 396378 -23620
rect 396180 -23818 396236 -23762
rect 396322 -23818 396378 -23762
rect 396180 -23960 396236 -23904
rect 396322 -23960 396378 -23904
rect 396180 -24102 396236 -24046
rect 396322 -24102 396378 -24046
rect 396180 -24244 396236 -24188
rect 396322 -24244 396378 -24188
rect 396180 -24386 396236 -24330
rect 396322 -24386 396378 -24330
rect 396180 -24528 396236 -24472
rect 396322 -24528 396378 -24472
rect 396180 -24670 396236 -24614
rect 396322 -24670 396378 -24614
rect 396180 -24812 396236 -24756
rect 396322 -24812 396378 -24756
rect 396180 -24954 396236 -24898
rect 396322 -24954 396378 -24898
rect 396180 -25096 396236 -25040
rect 396322 -25096 396378 -25040
rect 396180 -25238 396236 -25182
rect 396322 -25238 396378 -25182
rect 396180 -25380 396236 -25324
rect 396322 -25380 396378 -25324
rect 396180 -25522 396236 -25466
rect 396322 -25522 396378 -25466
rect 396580 -13736 396636 -13680
rect 396722 -13736 396778 -13680
rect 396580 -13878 396636 -13822
rect 396722 -13878 396778 -13822
rect 396580 -14020 396636 -13964
rect 396722 -14020 396778 -13964
rect 396580 -14162 396636 -14106
rect 396722 -14162 396778 -14106
rect 396580 -14304 396636 -14248
rect 396722 -14304 396778 -14248
rect 396580 -14446 396636 -14390
rect 396722 -14446 396778 -14390
rect 396580 -14588 396636 -14532
rect 396722 -14588 396778 -14532
rect 396580 -14730 396636 -14674
rect 396722 -14730 396778 -14674
rect 396580 -14872 396636 -14816
rect 396722 -14872 396778 -14816
rect 396580 -15014 396636 -14958
rect 396722 -15014 396778 -14958
rect 396580 -15156 396636 -15100
rect 396722 -15156 396778 -15100
rect 396580 -15298 396636 -15242
rect 396722 -15298 396778 -15242
rect 396580 -15440 396636 -15384
rect 396722 -15440 396778 -15384
rect 396580 -15582 396636 -15526
rect 396722 -15582 396778 -15526
rect 396580 -15724 396636 -15668
rect 396722 -15724 396778 -15668
rect 396580 -15866 396636 -15810
rect 396722 -15866 396778 -15810
rect 396580 -16008 396636 -15952
rect 396722 -16008 396778 -15952
rect 396580 -16150 396636 -16094
rect 396722 -16150 396778 -16094
rect 396580 -16292 396636 -16236
rect 396722 -16292 396778 -16236
rect 396580 -16434 396636 -16378
rect 396722 -16434 396778 -16378
rect 396580 -16576 396636 -16520
rect 396722 -16576 396778 -16520
rect 396580 -16718 396636 -16662
rect 396722 -16718 396778 -16662
rect 396580 -16860 396636 -16804
rect 396722 -16860 396778 -16804
rect 396580 -17002 396636 -16946
rect 396722 -17002 396778 -16946
rect 396580 -17144 396636 -17088
rect 396722 -17144 396778 -17088
rect 396580 -17286 396636 -17230
rect 396722 -17286 396778 -17230
rect 396580 -17428 396636 -17372
rect 396722 -17428 396778 -17372
rect 396580 -17570 396636 -17514
rect 396722 -17570 396778 -17514
rect 396580 -17712 396636 -17656
rect 396722 -17712 396778 -17656
rect 396580 -17854 396636 -17798
rect 396722 -17854 396778 -17798
rect 396580 -17996 396636 -17940
rect 396722 -17996 396778 -17940
rect 396580 -18138 396636 -18082
rect 396722 -18138 396778 -18082
rect 396580 -18280 396636 -18224
rect 396722 -18280 396778 -18224
rect 396580 -18422 396636 -18366
rect 396722 -18422 396778 -18366
rect 396580 -18564 396636 -18508
rect 396722 -18564 396778 -18508
rect 396580 -18706 396636 -18650
rect 396722 -18706 396778 -18650
rect 396580 -18848 396636 -18792
rect 396722 -18848 396778 -18792
rect 396580 -18990 396636 -18934
rect 396722 -18990 396778 -18934
rect 396580 -19132 396636 -19076
rect 396722 -19132 396778 -19076
rect 396580 -19274 396636 -19218
rect 396722 -19274 396778 -19218
rect 396580 -19416 396636 -19360
rect 396722 -19416 396778 -19360
rect 396580 -19558 396636 -19502
rect 396722 -19558 396778 -19502
rect 396580 -19700 396636 -19644
rect 396722 -19700 396778 -19644
rect 396580 -19842 396636 -19786
rect 396722 -19842 396778 -19786
rect 396580 -19984 396636 -19928
rect 396722 -19984 396778 -19928
rect 396580 -20126 396636 -20070
rect 396722 -20126 396778 -20070
rect 396580 -20268 396636 -20212
rect 396722 -20268 396778 -20212
rect 396580 -20410 396636 -20354
rect 396722 -20410 396778 -20354
rect 396580 -20552 396636 -20496
rect 396722 -20552 396778 -20496
rect 396580 -20694 396636 -20638
rect 396722 -20694 396778 -20638
rect 396580 -20836 396636 -20780
rect 396722 -20836 396778 -20780
rect 396580 -20978 396636 -20922
rect 396722 -20978 396778 -20922
rect 396580 -21120 396636 -21064
rect 396722 -21120 396778 -21064
rect 396580 -21262 396636 -21206
rect 396722 -21262 396778 -21206
rect 396580 -21404 396636 -21348
rect 396722 -21404 396778 -21348
rect 396580 -21546 396636 -21490
rect 396722 -21546 396778 -21490
rect 396580 -21688 396636 -21632
rect 396722 -21688 396778 -21632
rect 396580 -21830 396636 -21774
rect 396722 -21830 396778 -21774
rect 396580 -21972 396636 -21916
rect 396722 -21972 396778 -21916
rect 396580 -22114 396636 -22058
rect 396722 -22114 396778 -22058
rect 396580 -22256 396636 -22200
rect 396722 -22256 396778 -22200
rect 396580 -22398 396636 -22342
rect 396722 -22398 396778 -22342
rect 396580 -22540 396636 -22484
rect 396722 -22540 396778 -22484
rect 396580 -22682 396636 -22626
rect 396722 -22682 396778 -22626
rect 396580 -22824 396636 -22768
rect 396722 -22824 396778 -22768
rect 396580 -22966 396636 -22910
rect 396722 -22966 396778 -22910
rect 396580 -23108 396636 -23052
rect 396722 -23108 396778 -23052
rect 396580 -23250 396636 -23194
rect 396722 -23250 396778 -23194
rect 396580 -23392 396636 -23336
rect 396722 -23392 396778 -23336
rect 396580 -23534 396636 -23478
rect 396722 -23534 396778 -23478
rect 396580 -23676 396636 -23620
rect 396722 -23676 396778 -23620
rect 396580 -23818 396636 -23762
rect 396722 -23818 396778 -23762
rect 396580 -23960 396636 -23904
rect 396722 -23960 396778 -23904
rect 396580 -24102 396636 -24046
rect 396722 -24102 396778 -24046
rect 396580 -24244 396636 -24188
rect 396722 -24244 396778 -24188
rect 396580 -24386 396636 -24330
rect 396722 -24386 396778 -24330
rect 396580 -24528 396636 -24472
rect 396722 -24528 396778 -24472
rect 396580 -24670 396636 -24614
rect 396722 -24670 396778 -24614
rect 396580 -24812 396636 -24756
rect 396722 -24812 396778 -24756
rect 396580 -24954 396636 -24898
rect 396722 -24954 396778 -24898
rect 396580 -25096 396636 -25040
rect 396722 -25096 396778 -25040
rect 396580 -25238 396636 -25182
rect 396722 -25238 396778 -25182
rect 396580 -25380 396636 -25324
rect 396722 -25380 396778 -25324
rect 396580 -25522 396636 -25466
rect 396722 -25522 396778 -25466
rect 396977 -13736 397033 -13680
rect 397119 -13736 397175 -13680
rect 396977 -13878 397033 -13822
rect 397119 -13878 397175 -13822
rect 396977 -14020 397033 -13964
rect 397119 -14020 397175 -13964
rect 396977 -14162 397033 -14106
rect 397119 -14162 397175 -14106
rect 396977 -14304 397033 -14248
rect 397119 -14304 397175 -14248
rect 396977 -14446 397033 -14390
rect 397119 -14446 397175 -14390
rect 396977 -14588 397033 -14532
rect 397119 -14588 397175 -14532
rect 396977 -14730 397033 -14674
rect 397119 -14730 397175 -14674
rect 396977 -14872 397033 -14816
rect 397119 -14872 397175 -14816
rect 396977 -15014 397033 -14958
rect 397119 -15014 397175 -14958
rect 396977 -15156 397033 -15100
rect 397119 -15156 397175 -15100
rect 396977 -15298 397033 -15242
rect 397119 -15298 397175 -15242
rect 396977 -15440 397033 -15384
rect 397119 -15440 397175 -15384
rect 396977 -15582 397033 -15526
rect 397119 -15582 397175 -15526
rect 396977 -15724 397033 -15668
rect 397119 -15724 397175 -15668
rect 396977 -15866 397033 -15810
rect 397119 -15866 397175 -15810
rect 396977 -16008 397033 -15952
rect 397119 -16008 397175 -15952
rect 396977 -16150 397033 -16094
rect 397119 -16150 397175 -16094
rect 396977 -16292 397033 -16236
rect 397119 -16292 397175 -16236
rect 396977 -16434 397033 -16378
rect 397119 -16434 397175 -16378
rect 396977 -16576 397033 -16520
rect 397119 -16576 397175 -16520
rect 396977 -16718 397033 -16662
rect 397119 -16718 397175 -16662
rect 396977 -16860 397033 -16804
rect 397119 -16860 397175 -16804
rect 396977 -17002 397033 -16946
rect 397119 -17002 397175 -16946
rect 396977 -17144 397033 -17088
rect 397119 -17144 397175 -17088
rect 396977 -17286 397033 -17230
rect 397119 -17286 397175 -17230
rect 396977 -17428 397033 -17372
rect 397119 -17428 397175 -17372
rect 396977 -17570 397033 -17514
rect 397119 -17570 397175 -17514
rect 396977 -17712 397033 -17656
rect 397119 -17712 397175 -17656
rect 396977 -17854 397033 -17798
rect 397119 -17854 397175 -17798
rect 396977 -17996 397033 -17940
rect 397119 -17996 397175 -17940
rect 396977 -18138 397033 -18082
rect 397119 -18138 397175 -18082
rect 396977 -18280 397033 -18224
rect 397119 -18280 397175 -18224
rect 396977 -18422 397033 -18366
rect 397119 -18422 397175 -18366
rect 396977 -18564 397033 -18508
rect 397119 -18564 397175 -18508
rect 396977 -18706 397033 -18650
rect 397119 -18706 397175 -18650
rect 396977 -18848 397033 -18792
rect 397119 -18848 397175 -18792
rect 396977 -18990 397033 -18934
rect 397119 -18990 397175 -18934
rect 396977 -19132 397033 -19076
rect 397119 -19132 397175 -19076
rect 396977 -19274 397033 -19218
rect 397119 -19274 397175 -19218
rect 396977 -19416 397033 -19360
rect 397119 -19416 397175 -19360
rect 396977 -19558 397033 -19502
rect 397119 -19558 397175 -19502
rect 396977 -19700 397033 -19644
rect 397119 -19700 397175 -19644
rect 396977 -19842 397033 -19786
rect 397119 -19842 397175 -19786
rect 396977 -19984 397033 -19928
rect 397119 -19984 397175 -19928
rect 396977 -20126 397033 -20070
rect 397119 -20126 397175 -20070
rect 396977 -20268 397033 -20212
rect 397119 -20268 397175 -20212
rect 396977 -20410 397033 -20354
rect 397119 -20410 397175 -20354
rect 396977 -20552 397033 -20496
rect 397119 -20552 397175 -20496
rect 396977 -20694 397033 -20638
rect 397119 -20694 397175 -20638
rect 396977 -20836 397033 -20780
rect 397119 -20836 397175 -20780
rect 396977 -20978 397033 -20922
rect 397119 -20978 397175 -20922
rect 396977 -21120 397033 -21064
rect 397119 -21120 397175 -21064
rect 396977 -21262 397033 -21206
rect 397119 -21262 397175 -21206
rect 396977 -21404 397033 -21348
rect 397119 -21404 397175 -21348
rect 396977 -21546 397033 -21490
rect 397119 -21546 397175 -21490
rect 396977 -21688 397033 -21632
rect 397119 -21688 397175 -21632
rect 396977 -21830 397033 -21774
rect 397119 -21830 397175 -21774
rect 396977 -21972 397033 -21916
rect 397119 -21972 397175 -21916
rect 396977 -22114 397033 -22058
rect 397119 -22114 397175 -22058
rect 396977 -22256 397033 -22200
rect 397119 -22256 397175 -22200
rect 396977 -22398 397033 -22342
rect 397119 -22398 397175 -22342
rect 396977 -22540 397033 -22484
rect 397119 -22540 397175 -22484
rect 396977 -22682 397033 -22626
rect 397119 -22682 397175 -22626
rect 396977 -22824 397033 -22768
rect 397119 -22824 397175 -22768
rect 396977 -22966 397033 -22910
rect 397119 -22966 397175 -22910
rect 396977 -23108 397033 -23052
rect 397119 -23108 397175 -23052
rect 396977 -23250 397033 -23194
rect 397119 -23250 397175 -23194
rect 396977 -23392 397033 -23336
rect 397119 -23392 397175 -23336
rect 396977 -23534 397033 -23478
rect 397119 -23534 397175 -23478
rect 396977 -23676 397033 -23620
rect 397119 -23676 397175 -23620
rect 396977 -23818 397033 -23762
rect 397119 -23818 397175 -23762
rect 396977 -23960 397033 -23904
rect 397119 -23960 397175 -23904
rect 396977 -24102 397033 -24046
rect 397119 -24102 397175 -24046
rect 396977 -24244 397033 -24188
rect 397119 -24244 397175 -24188
rect 396977 -24386 397033 -24330
rect 397119 -24386 397175 -24330
rect 396977 -24528 397033 -24472
rect 397119 -24528 397175 -24472
rect 396977 -24670 397033 -24614
rect 397119 -24670 397175 -24614
rect 396977 -24812 397033 -24756
rect 397119 -24812 397175 -24756
rect 396977 -24954 397033 -24898
rect 397119 -24954 397175 -24898
rect 396977 -25096 397033 -25040
rect 397119 -25096 397175 -25040
rect 396977 -25238 397033 -25182
rect 397119 -25238 397175 -25182
rect 396977 -25380 397033 -25324
rect 397119 -25380 397175 -25324
rect 396977 -25522 397033 -25466
rect 397119 -25522 397175 -25466
rect 397374 -13736 397430 -13680
rect 397516 -13736 397572 -13680
rect 397374 -13878 397430 -13822
rect 397516 -13878 397572 -13822
rect 397374 -14020 397430 -13964
rect 397516 -14020 397572 -13964
rect 397374 -14162 397430 -14106
rect 397516 -14162 397572 -14106
rect 397374 -14304 397430 -14248
rect 397516 -14304 397572 -14248
rect 397374 -14446 397430 -14390
rect 397516 -14446 397572 -14390
rect 397374 -14588 397430 -14532
rect 397516 -14588 397572 -14532
rect 397374 -14730 397430 -14674
rect 397516 -14730 397572 -14674
rect 397374 -14872 397430 -14816
rect 397516 -14872 397572 -14816
rect 397374 -15014 397430 -14958
rect 397516 -15014 397572 -14958
rect 397374 -15156 397430 -15100
rect 397516 -15156 397572 -15100
rect 397374 -15298 397430 -15242
rect 397516 -15298 397572 -15242
rect 397374 -15440 397430 -15384
rect 397516 -15440 397572 -15384
rect 397374 -15582 397430 -15526
rect 397516 -15582 397572 -15526
rect 397374 -15724 397430 -15668
rect 397516 -15724 397572 -15668
rect 397374 -15866 397430 -15810
rect 397516 -15866 397572 -15810
rect 397374 -16008 397430 -15952
rect 397516 -16008 397572 -15952
rect 397374 -16150 397430 -16094
rect 397516 -16150 397572 -16094
rect 397374 -16292 397430 -16236
rect 397516 -16292 397572 -16236
rect 397374 -16434 397430 -16378
rect 397516 -16434 397572 -16378
rect 397374 -16576 397430 -16520
rect 397516 -16576 397572 -16520
rect 397374 -16718 397430 -16662
rect 397516 -16718 397572 -16662
rect 397374 -16860 397430 -16804
rect 397516 -16860 397572 -16804
rect 397374 -17002 397430 -16946
rect 397516 -17002 397572 -16946
rect 397374 -17144 397430 -17088
rect 397516 -17144 397572 -17088
rect 397374 -17286 397430 -17230
rect 397516 -17286 397572 -17230
rect 397374 -17428 397430 -17372
rect 397516 -17428 397572 -17372
rect 397374 -17570 397430 -17514
rect 397516 -17570 397572 -17514
rect 397374 -17712 397430 -17656
rect 397516 -17712 397572 -17656
rect 397374 -17854 397430 -17798
rect 397516 -17854 397572 -17798
rect 397374 -17996 397430 -17940
rect 397516 -17996 397572 -17940
rect 397374 -18138 397430 -18082
rect 397516 -18138 397572 -18082
rect 397374 -18280 397430 -18224
rect 397516 -18280 397572 -18224
rect 397374 -18422 397430 -18366
rect 397516 -18422 397572 -18366
rect 397374 -18564 397430 -18508
rect 397516 -18564 397572 -18508
rect 397374 -18706 397430 -18650
rect 397516 -18706 397572 -18650
rect 397374 -18848 397430 -18792
rect 397516 -18848 397572 -18792
rect 397374 -18990 397430 -18934
rect 397516 -18990 397572 -18934
rect 397374 -19132 397430 -19076
rect 397516 -19132 397572 -19076
rect 397374 -19274 397430 -19218
rect 397516 -19274 397572 -19218
rect 397374 -19416 397430 -19360
rect 397516 -19416 397572 -19360
rect 397374 -19558 397430 -19502
rect 397516 -19558 397572 -19502
rect 397374 -19700 397430 -19644
rect 397516 -19700 397572 -19644
rect 397374 -19842 397430 -19786
rect 397516 -19842 397572 -19786
rect 397374 -19984 397430 -19928
rect 397516 -19984 397572 -19928
rect 397374 -20126 397430 -20070
rect 397516 -20126 397572 -20070
rect 397374 -20268 397430 -20212
rect 397516 -20268 397572 -20212
rect 397374 -20410 397430 -20354
rect 397516 -20410 397572 -20354
rect 397374 -20552 397430 -20496
rect 397516 -20552 397572 -20496
rect 397374 -20694 397430 -20638
rect 397516 -20694 397572 -20638
rect 397374 -20836 397430 -20780
rect 397516 -20836 397572 -20780
rect 397374 -20978 397430 -20922
rect 397516 -20978 397572 -20922
rect 397374 -21120 397430 -21064
rect 397516 -21120 397572 -21064
rect 397374 -21262 397430 -21206
rect 397516 -21262 397572 -21206
rect 397374 -21404 397430 -21348
rect 397516 -21404 397572 -21348
rect 397374 -21546 397430 -21490
rect 397516 -21546 397572 -21490
rect 397374 -21688 397430 -21632
rect 397516 -21688 397572 -21632
rect 397374 -21830 397430 -21774
rect 397516 -21830 397572 -21774
rect 397374 -21972 397430 -21916
rect 397516 -21972 397572 -21916
rect 397374 -22114 397430 -22058
rect 397516 -22114 397572 -22058
rect 397374 -22256 397430 -22200
rect 397516 -22256 397572 -22200
rect 397374 -22398 397430 -22342
rect 397516 -22398 397572 -22342
rect 397374 -22540 397430 -22484
rect 397516 -22540 397572 -22484
rect 397374 -22682 397430 -22626
rect 397516 -22682 397572 -22626
rect 397374 -22824 397430 -22768
rect 397516 -22824 397572 -22768
rect 397374 -22966 397430 -22910
rect 397516 -22966 397572 -22910
rect 397374 -23108 397430 -23052
rect 397516 -23108 397572 -23052
rect 397374 -23250 397430 -23194
rect 397516 -23250 397572 -23194
rect 397374 -23392 397430 -23336
rect 397516 -23392 397572 -23336
rect 397374 -23534 397430 -23478
rect 397516 -23534 397572 -23478
rect 397374 -23676 397430 -23620
rect 397516 -23676 397572 -23620
rect 397374 -23818 397430 -23762
rect 397516 -23818 397572 -23762
rect 397374 -23960 397430 -23904
rect 397516 -23960 397572 -23904
rect 397374 -24102 397430 -24046
rect 397516 -24102 397572 -24046
rect 397374 -24244 397430 -24188
rect 397516 -24244 397572 -24188
rect 397374 -24386 397430 -24330
rect 397516 -24386 397572 -24330
rect 397374 -24528 397430 -24472
rect 397516 -24528 397572 -24472
rect 397374 -24670 397430 -24614
rect 397516 -24670 397572 -24614
rect 397374 -24812 397430 -24756
rect 397516 -24812 397572 -24756
rect 397374 -24954 397430 -24898
rect 397516 -24954 397572 -24898
rect 397374 -25096 397430 -25040
rect 397516 -25096 397572 -25040
rect 397374 -25238 397430 -25182
rect 397516 -25238 397572 -25182
rect 397374 -25380 397430 -25324
rect 397516 -25380 397572 -25324
rect 397374 -25522 397430 -25466
rect 397516 -25522 397572 -25466
rect 397778 -13736 397834 -13680
rect 397920 -13736 397976 -13680
rect 397778 -13878 397834 -13822
rect 397920 -13878 397976 -13822
rect 397778 -14020 397834 -13964
rect 397920 -14020 397976 -13964
rect 397778 -14162 397834 -14106
rect 397920 -14162 397976 -14106
rect 397778 -14304 397834 -14248
rect 397920 -14304 397976 -14248
rect 397778 -14446 397834 -14390
rect 397920 -14446 397976 -14390
rect 397778 -14588 397834 -14532
rect 397920 -14588 397976 -14532
rect 397778 -14730 397834 -14674
rect 397920 -14730 397976 -14674
rect 397778 -14872 397834 -14816
rect 397920 -14872 397976 -14816
rect 397778 -15014 397834 -14958
rect 397920 -15014 397976 -14958
rect 397778 -15156 397834 -15100
rect 397920 -15156 397976 -15100
rect 397778 -15298 397834 -15242
rect 397920 -15298 397976 -15242
rect 397778 -15440 397834 -15384
rect 397920 -15440 397976 -15384
rect 397778 -15582 397834 -15526
rect 397920 -15582 397976 -15526
rect 397778 -15724 397834 -15668
rect 397920 -15724 397976 -15668
rect 397778 -15866 397834 -15810
rect 397920 -15866 397976 -15810
rect 397778 -16008 397834 -15952
rect 397920 -16008 397976 -15952
rect 397778 -16150 397834 -16094
rect 397920 -16150 397976 -16094
rect 397778 -16292 397834 -16236
rect 397920 -16292 397976 -16236
rect 397778 -16434 397834 -16378
rect 397920 -16434 397976 -16378
rect 397778 -16576 397834 -16520
rect 397920 -16576 397976 -16520
rect 397778 -16718 397834 -16662
rect 397920 -16718 397976 -16662
rect 397778 -16860 397834 -16804
rect 397920 -16860 397976 -16804
rect 397778 -17002 397834 -16946
rect 397920 -17002 397976 -16946
rect 397778 -17144 397834 -17088
rect 397920 -17144 397976 -17088
rect 397778 -17286 397834 -17230
rect 397920 -17286 397976 -17230
rect 397778 -17428 397834 -17372
rect 397920 -17428 397976 -17372
rect 397778 -17570 397834 -17514
rect 397920 -17570 397976 -17514
rect 397778 -17712 397834 -17656
rect 397920 -17712 397976 -17656
rect 397778 -17854 397834 -17798
rect 397920 -17854 397976 -17798
rect 397778 -17996 397834 -17940
rect 397920 -17996 397976 -17940
rect 397778 -18138 397834 -18082
rect 397920 -18138 397976 -18082
rect 397778 -18280 397834 -18224
rect 397920 -18280 397976 -18224
rect 397778 -18422 397834 -18366
rect 397920 -18422 397976 -18366
rect 397778 -18564 397834 -18508
rect 397920 -18564 397976 -18508
rect 397778 -18706 397834 -18650
rect 397920 -18706 397976 -18650
rect 397778 -18848 397834 -18792
rect 397920 -18848 397976 -18792
rect 397778 -18990 397834 -18934
rect 397920 -18990 397976 -18934
rect 397778 -19132 397834 -19076
rect 397920 -19132 397976 -19076
rect 397778 -19274 397834 -19218
rect 397920 -19274 397976 -19218
rect 397778 -19416 397834 -19360
rect 397920 -19416 397976 -19360
rect 397778 -19558 397834 -19502
rect 397920 -19558 397976 -19502
rect 397778 -19700 397834 -19644
rect 397920 -19700 397976 -19644
rect 397778 -19842 397834 -19786
rect 397920 -19842 397976 -19786
rect 397778 -19984 397834 -19928
rect 397920 -19984 397976 -19928
rect 397778 -20126 397834 -20070
rect 397920 -20126 397976 -20070
rect 397778 -20268 397834 -20212
rect 397920 -20268 397976 -20212
rect 397778 -20410 397834 -20354
rect 397920 -20410 397976 -20354
rect 397778 -20552 397834 -20496
rect 397920 -20552 397976 -20496
rect 397778 -20694 397834 -20638
rect 397920 -20694 397976 -20638
rect 397778 -20836 397834 -20780
rect 397920 -20836 397976 -20780
rect 397778 -20978 397834 -20922
rect 397920 -20978 397976 -20922
rect 397778 -21120 397834 -21064
rect 397920 -21120 397976 -21064
rect 397778 -21262 397834 -21206
rect 397920 -21262 397976 -21206
rect 397778 -21404 397834 -21348
rect 397920 -21404 397976 -21348
rect 397778 -21546 397834 -21490
rect 397920 -21546 397976 -21490
rect 397778 -21688 397834 -21632
rect 397920 -21688 397976 -21632
rect 397778 -21830 397834 -21774
rect 397920 -21830 397976 -21774
rect 397778 -21972 397834 -21916
rect 397920 -21972 397976 -21916
rect 397778 -22114 397834 -22058
rect 397920 -22114 397976 -22058
rect 397778 -22256 397834 -22200
rect 397920 -22256 397976 -22200
rect 397778 -22398 397834 -22342
rect 397920 -22398 397976 -22342
rect 397778 -22540 397834 -22484
rect 397920 -22540 397976 -22484
rect 397778 -22682 397834 -22626
rect 397920 -22682 397976 -22626
rect 397778 -22824 397834 -22768
rect 397920 -22824 397976 -22768
rect 397778 -22966 397834 -22910
rect 397920 -22966 397976 -22910
rect 397778 -23108 397834 -23052
rect 397920 -23108 397976 -23052
rect 397778 -23250 397834 -23194
rect 397920 -23250 397976 -23194
rect 397778 -23392 397834 -23336
rect 397920 -23392 397976 -23336
rect 397778 -23534 397834 -23478
rect 397920 -23534 397976 -23478
rect 397778 -23676 397834 -23620
rect 397920 -23676 397976 -23620
rect 397778 -23818 397834 -23762
rect 397920 -23818 397976 -23762
rect 397778 -23960 397834 -23904
rect 397920 -23960 397976 -23904
rect 397778 -24102 397834 -24046
rect 397920 -24102 397976 -24046
rect 397778 -24244 397834 -24188
rect 397920 -24244 397976 -24188
rect 397778 -24386 397834 -24330
rect 397920 -24386 397976 -24330
rect 397778 -24528 397834 -24472
rect 397920 -24528 397976 -24472
rect 397778 -24670 397834 -24614
rect 397920 -24670 397976 -24614
rect 397778 -24812 397834 -24756
rect 397920 -24812 397976 -24756
rect 397778 -24954 397834 -24898
rect 397920 -24954 397976 -24898
rect 397778 -25096 397834 -25040
rect 397920 -25096 397976 -25040
rect 397778 -25238 397834 -25182
rect 397920 -25238 397976 -25182
rect 397778 -25380 397834 -25324
rect 397920 -25380 397976 -25324
rect 397778 -25522 397834 -25466
rect 397920 -25522 397976 -25466
rect 398174 -13736 398230 -13680
rect 398316 -13736 398372 -13680
rect 398174 -13878 398230 -13822
rect 398316 -13878 398372 -13822
rect 398174 -14020 398230 -13964
rect 398316 -14020 398372 -13964
rect 398174 -14162 398230 -14106
rect 398316 -14162 398372 -14106
rect 398174 -14304 398230 -14248
rect 398316 -14304 398372 -14248
rect 398174 -14446 398230 -14390
rect 398316 -14446 398372 -14390
rect 398174 -14588 398230 -14532
rect 398316 -14588 398372 -14532
rect 398174 -14730 398230 -14674
rect 398316 -14730 398372 -14674
rect 398174 -14872 398230 -14816
rect 398316 -14872 398372 -14816
rect 398174 -15014 398230 -14958
rect 398316 -15014 398372 -14958
rect 398174 -15156 398230 -15100
rect 398316 -15156 398372 -15100
rect 398174 -15298 398230 -15242
rect 398316 -15298 398372 -15242
rect 398174 -15440 398230 -15384
rect 398316 -15440 398372 -15384
rect 398174 -15582 398230 -15526
rect 398316 -15582 398372 -15526
rect 398174 -15724 398230 -15668
rect 398316 -15724 398372 -15668
rect 398174 -15866 398230 -15810
rect 398316 -15866 398372 -15810
rect 398174 -16008 398230 -15952
rect 398316 -16008 398372 -15952
rect 398174 -16150 398230 -16094
rect 398316 -16150 398372 -16094
rect 398174 -16292 398230 -16236
rect 398316 -16292 398372 -16236
rect 398174 -16434 398230 -16378
rect 398316 -16434 398372 -16378
rect 398174 -16576 398230 -16520
rect 398316 -16576 398372 -16520
rect 398174 -16718 398230 -16662
rect 398316 -16718 398372 -16662
rect 398174 -16860 398230 -16804
rect 398316 -16860 398372 -16804
rect 398174 -17002 398230 -16946
rect 398316 -17002 398372 -16946
rect 398174 -17144 398230 -17088
rect 398316 -17144 398372 -17088
rect 398174 -17286 398230 -17230
rect 398316 -17286 398372 -17230
rect 398174 -17428 398230 -17372
rect 398316 -17428 398372 -17372
rect 398174 -17570 398230 -17514
rect 398316 -17570 398372 -17514
rect 398174 -17712 398230 -17656
rect 398316 -17712 398372 -17656
rect 398174 -17854 398230 -17798
rect 398316 -17854 398372 -17798
rect 398174 -17996 398230 -17940
rect 398316 -17996 398372 -17940
rect 398174 -18138 398230 -18082
rect 398316 -18138 398372 -18082
rect 398174 -18280 398230 -18224
rect 398316 -18280 398372 -18224
rect 398174 -18422 398230 -18366
rect 398316 -18422 398372 -18366
rect 398174 -18564 398230 -18508
rect 398316 -18564 398372 -18508
rect 398174 -18706 398230 -18650
rect 398316 -18706 398372 -18650
rect 398174 -18848 398230 -18792
rect 398316 -18848 398372 -18792
rect 398174 -18990 398230 -18934
rect 398316 -18990 398372 -18934
rect 398174 -19132 398230 -19076
rect 398316 -19132 398372 -19076
rect 398174 -19274 398230 -19218
rect 398316 -19274 398372 -19218
rect 398174 -19416 398230 -19360
rect 398316 -19416 398372 -19360
rect 398174 -19558 398230 -19502
rect 398316 -19558 398372 -19502
rect 398174 -19700 398230 -19644
rect 398316 -19700 398372 -19644
rect 398174 -19842 398230 -19786
rect 398316 -19842 398372 -19786
rect 398174 -19984 398230 -19928
rect 398316 -19984 398372 -19928
rect 398174 -20126 398230 -20070
rect 398316 -20126 398372 -20070
rect 398174 -20268 398230 -20212
rect 398316 -20268 398372 -20212
rect 398174 -20410 398230 -20354
rect 398316 -20410 398372 -20354
rect 398174 -20552 398230 -20496
rect 398316 -20552 398372 -20496
rect 398174 -20694 398230 -20638
rect 398316 -20694 398372 -20638
rect 398174 -20836 398230 -20780
rect 398316 -20836 398372 -20780
rect 398174 -20978 398230 -20922
rect 398316 -20978 398372 -20922
rect 398174 -21120 398230 -21064
rect 398316 -21120 398372 -21064
rect 398174 -21262 398230 -21206
rect 398316 -21262 398372 -21206
rect 398174 -21404 398230 -21348
rect 398316 -21404 398372 -21348
rect 398174 -21546 398230 -21490
rect 398316 -21546 398372 -21490
rect 398174 -21688 398230 -21632
rect 398316 -21688 398372 -21632
rect 398174 -21830 398230 -21774
rect 398316 -21830 398372 -21774
rect 398174 -21972 398230 -21916
rect 398316 -21972 398372 -21916
rect 398174 -22114 398230 -22058
rect 398316 -22114 398372 -22058
rect 398174 -22256 398230 -22200
rect 398316 -22256 398372 -22200
rect 398174 -22398 398230 -22342
rect 398316 -22398 398372 -22342
rect 398174 -22540 398230 -22484
rect 398316 -22540 398372 -22484
rect 398174 -22682 398230 -22626
rect 398316 -22682 398372 -22626
rect 398174 -22824 398230 -22768
rect 398316 -22824 398372 -22768
rect 398174 -22966 398230 -22910
rect 398316 -22966 398372 -22910
rect 398174 -23108 398230 -23052
rect 398316 -23108 398372 -23052
rect 398174 -23250 398230 -23194
rect 398316 -23250 398372 -23194
rect 398174 -23392 398230 -23336
rect 398316 -23392 398372 -23336
rect 398174 -23534 398230 -23478
rect 398316 -23534 398372 -23478
rect 398174 -23676 398230 -23620
rect 398316 -23676 398372 -23620
rect 398174 -23818 398230 -23762
rect 398316 -23818 398372 -23762
rect 398174 -23960 398230 -23904
rect 398316 -23960 398372 -23904
rect 398174 -24102 398230 -24046
rect 398316 -24102 398372 -24046
rect 398174 -24244 398230 -24188
rect 398316 -24244 398372 -24188
rect 398174 -24386 398230 -24330
rect 398316 -24386 398372 -24330
rect 398174 -24528 398230 -24472
rect 398316 -24528 398372 -24472
rect 398174 -24670 398230 -24614
rect 398316 -24670 398372 -24614
rect 398174 -24812 398230 -24756
rect 398316 -24812 398372 -24756
rect 398174 -24954 398230 -24898
rect 398316 -24954 398372 -24898
rect 398174 -25096 398230 -25040
rect 398316 -25096 398372 -25040
rect 398174 -25238 398230 -25182
rect 398316 -25238 398372 -25182
rect 398174 -25380 398230 -25324
rect 398316 -25380 398372 -25324
rect 398174 -25522 398230 -25466
rect 398316 -25522 398372 -25466
rect 398574 -13736 398630 -13680
rect 398716 -13736 398772 -13680
rect 398574 -13878 398630 -13822
rect 398716 -13878 398772 -13822
rect 398574 -14020 398630 -13964
rect 398716 -14020 398772 -13964
rect 398574 -14162 398630 -14106
rect 398716 -14162 398772 -14106
rect 398574 -14304 398630 -14248
rect 398716 -14304 398772 -14248
rect 398574 -14446 398630 -14390
rect 398716 -14446 398772 -14390
rect 398574 -14588 398630 -14532
rect 398716 -14588 398772 -14532
rect 398574 -14730 398630 -14674
rect 398716 -14730 398772 -14674
rect 398574 -14872 398630 -14816
rect 398716 -14872 398772 -14816
rect 398574 -15014 398630 -14958
rect 398716 -15014 398772 -14958
rect 398574 -15156 398630 -15100
rect 398716 -15156 398772 -15100
rect 398574 -15298 398630 -15242
rect 398716 -15298 398772 -15242
rect 398574 -15440 398630 -15384
rect 398716 -15440 398772 -15384
rect 398574 -15582 398630 -15526
rect 398716 -15582 398772 -15526
rect 398574 -15724 398630 -15668
rect 398716 -15724 398772 -15668
rect 398574 -15866 398630 -15810
rect 398716 -15866 398772 -15810
rect 398574 -16008 398630 -15952
rect 398716 -16008 398772 -15952
rect 398574 -16150 398630 -16094
rect 398716 -16150 398772 -16094
rect 398574 -16292 398630 -16236
rect 398716 -16292 398772 -16236
rect 398574 -16434 398630 -16378
rect 398716 -16434 398772 -16378
rect 398574 -16576 398630 -16520
rect 398716 -16576 398772 -16520
rect 398574 -16718 398630 -16662
rect 398716 -16718 398772 -16662
rect 398574 -16860 398630 -16804
rect 398716 -16860 398772 -16804
rect 398574 -17002 398630 -16946
rect 398716 -17002 398772 -16946
rect 398574 -17144 398630 -17088
rect 398716 -17144 398772 -17088
rect 398574 -17286 398630 -17230
rect 398716 -17286 398772 -17230
rect 398574 -17428 398630 -17372
rect 398716 -17428 398772 -17372
rect 398574 -17570 398630 -17514
rect 398716 -17570 398772 -17514
rect 398574 -17712 398630 -17656
rect 398716 -17712 398772 -17656
rect 398574 -17854 398630 -17798
rect 398716 -17854 398772 -17798
rect 398574 -17996 398630 -17940
rect 398716 -17996 398772 -17940
rect 398574 -18138 398630 -18082
rect 398716 -18138 398772 -18082
rect 398574 -18280 398630 -18224
rect 398716 -18280 398772 -18224
rect 398574 -18422 398630 -18366
rect 398716 -18422 398772 -18366
rect 398574 -18564 398630 -18508
rect 398716 -18564 398772 -18508
rect 398574 -18706 398630 -18650
rect 398716 -18706 398772 -18650
rect 398574 -18848 398630 -18792
rect 398716 -18848 398772 -18792
rect 398574 -18990 398630 -18934
rect 398716 -18990 398772 -18934
rect 398574 -19132 398630 -19076
rect 398716 -19132 398772 -19076
rect 398574 -19274 398630 -19218
rect 398716 -19274 398772 -19218
rect 398574 -19416 398630 -19360
rect 398716 -19416 398772 -19360
rect 398574 -19558 398630 -19502
rect 398716 -19558 398772 -19502
rect 398574 -19700 398630 -19644
rect 398716 -19700 398772 -19644
rect 398574 -19842 398630 -19786
rect 398716 -19842 398772 -19786
rect 398574 -19984 398630 -19928
rect 398716 -19984 398772 -19928
rect 398574 -20126 398630 -20070
rect 398716 -20126 398772 -20070
rect 398574 -20268 398630 -20212
rect 398716 -20268 398772 -20212
rect 398574 -20410 398630 -20354
rect 398716 -20410 398772 -20354
rect 398574 -20552 398630 -20496
rect 398716 -20552 398772 -20496
rect 398574 -20694 398630 -20638
rect 398716 -20694 398772 -20638
rect 398574 -20836 398630 -20780
rect 398716 -20836 398772 -20780
rect 398574 -20978 398630 -20922
rect 398716 -20978 398772 -20922
rect 398574 -21120 398630 -21064
rect 398716 -21120 398772 -21064
rect 398574 -21262 398630 -21206
rect 398716 -21262 398772 -21206
rect 398574 -21404 398630 -21348
rect 398716 -21404 398772 -21348
rect 398574 -21546 398630 -21490
rect 398716 -21546 398772 -21490
rect 398574 -21688 398630 -21632
rect 398716 -21688 398772 -21632
rect 398574 -21830 398630 -21774
rect 398716 -21830 398772 -21774
rect 398574 -21972 398630 -21916
rect 398716 -21972 398772 -21916
rect 398574 -22114 398630 -22058
rect 398716 -22114 398772 -22058
rect 398574 -22256 398630 -22200
rect 398716 -22256 398772 -22200
rect 398574 -22398 398630 -22342
rect 398716 -22398 398772 -22342
rect 398574 -22540 398630 -22484
rect 398716 -22540 398772 -22484
rect 398574 -22682 398630 -22626
rect 398716 -22682 398772 -22626
rect 398574 -22824 398630 -22768
rect 398716 -22824 398772 -22768
rect 398574 -22966 398630 -22910
rect 398716 -22966 398772 -22910
rect 398574 -23108 398630 -23052
rect 398716 -23108 398772 -23052
rect 398574 -23250 398630 -23194
rect 398716 -23250 398772 -23194
rect 398574 -23392 398630 -23336
rect 398716 -23392 398772 -23336
rect 398574 -23534 398630 -23478
rect 398716 -23534 398772 -23478
rect 398574 -23676 398630 -23620
rect 398716 -23676 398772 -23620
rect 398574 -23818 398630 -23762
rect 398716 -23818 398772 -23762
rect 398574 -23960 398630 -23904
rect 398716 -23960 398772 -23904
rect 398574 -24102 398630 -24046
rect 398716 -24102 398772 -24046
rect 398574 -24244 398630 -24188
rect 398716 -24244 398772 -24188
rect 398574 -24386 398630 -24330
rect 398716 -24386 398772 -24330
rect 398574 -24528 398630 -24472
rect 398716 -24528 398772 -24472
rect 398574 -24670 398630 -24614
rect 398716 -24670 398772 -24614
rect 398574 -24812 398630 -24756
rect 398716 -24812 398772 -24756
rect 398574 -24954 398630 -24898
rect 398716 -24954 398772 -24898
rect 398574 -25096 398630 -25040
rect 398716 -25096 398772 -25040
rect 398574 -25238 398630 -25182
rect 398716 -25238 398772 -25182
rect 398574 -25380 398630 -25324
rect 398716 -25380 398772 -25324
rect 398574 -25522 398630 -25466
rect 398716 -25522 398772 -25466
rect 398971 -13736 399027 -13680
rect 399113 -13736 399169 -13680
rect 398971 -13878 399027 -13822
rect 399113 -13878 399169 -13822
rect 398971 -14020 399027 -13964
rect 399113 -14020 399169 -13964
rect 398971 -14162 399027 -14106
rect 399113 -14162 399169 -14106
rect 398971 -14304 399027 -14248
rect 399113 -14304 399169 -14248
rect 398971 -14446 399027 -14390
rect 399113 -14446 399169 -14390
rect 398971 -14588 399027 -14532
rect 399113 -14588 399169 -14532
rect 398971 -14730 399027 -14674
rect 399113 -14730 399169 -14674
rect 398971 -14872 399027 -14816
rect 399113 -14872 399169 -14816
rect 398971 -15014 399027 -14958
rect 399113 -15014 399169 -14958
rect 398971 -15156 399027 -15100
rect 399113 -15156 399169 -15100
rect 398971 -15298 399027 -15242
rect 399113 -15298 399169 -15242
rect 398971 -15440 399027 -15384
rect 399113 -15440 399169 -15384
rect 398971 -15582 399027 -15526
rect 399113 -15582 399169 -15526
rect 398971 -15724 399027 -15668
rect 399113 -15724 399169 -15668
rect 398971 -15866 399027 -15810
rect 399113 -15866 399169 -15810
rect 398971 -16008 399027 -15952
rect 399113 -16008 399169 -15952
rect 398971 -16150 399027 -16094
rect 399113 -16150 399169 -16094
rect 398971 -16292 399027 -16236
rect 399113 -16292 399169 -16236
rect 398971 -16434 399027 -16378
rect 399113 -16434 399169 -16378
rect 398971 -16576 399027 -16520
rect 399113 -16576 399169 -16520
rect 398971 -16718 399027 -16662
rect 399113 -16718 399169 -16662
rect 398971 -16860 399027 -16804
rect 399113 -16860 399169 -16804
rect 398971 -17002 399027 -16946
rect 399113 -17002 399169 -16946
rect 398971 -17144 399027 -17088
rect 399113 -17144 399169 -17088
rect 398971 -17286 399027 -17230
rect 399113 -17286 399169 -17230
rect 398971 -17428 399027 -17372
rect 399113 -17428 399169 -17372
rect 398971 -17570 399027 -17514
rect 399113 -17570 399169 -17514
rect 398971 -17712 399027 -17656
rect 399113 -17712 399169 -17656
rect 398971 -17854 399027 -17798
rect 399113 -17854 399169 -17798
rect 398971 -17996 399027 -17940
rect 399113 -17996 399169 -17940
rect 398971 -18138 399027 -18082
rect 399113 -18138 399169 -18082
rect 398971 -18280 399027 -18224
rect 399113 -18280 399169 -18224
rect 398971 -18422 399027 -18366
rect 399113 -18422 399169 -18366
rect 398971 -18564 399027 -18508
rect 399113 -18564 399169 -18508
rect 398971 -18706 399027 -18650
rect 399113 -18706 399169 -18650
rect 398971 -18848 399027 -18792
rect 399113 -18848 399169 -18792
rect 398971 -18990 399027 -18934
rect 399113 -18990 399169 -18934
rect 398971 -19132 399027 -19076
rect 399113 -19132 399169 -19076
rect 398971 -19274 399027 -19218
rect 399113 -19274 399169 -19218
rect 398971 -19416 399027 -19360
rect 399113 -19416 399169 -19360
rect 398971 -19558 399027 -19502
rect 399113 -19558 399169 -19502
rect 398971 -19700 399027 -19644
rect 399113 -19700 399169 -19644
rect 398971 -19842 399027 -19786
rect 399113 -19842 399169 -19786
rect 398971 -19984 399027 -19928
rect 399113 -19984 399169 -19928
rect 398971 -20126 399027 -20070
rect 399113 -20126 399169 -20070
rect 398971 -20268 399027 -20212
rect 399113 -20268 399169 -20212
rect 398971 -20410 399027 -20354
rect 399113 -20410 399169 -20354
rect 398971 -20552 399027 -20496
rect 399113 -20552 399169 -20496
rect 398971 -20694 399027 -20638
rect 399113 -20694 399169 -20638
rect 398971 -20836 399027 -20780
rect 399113 -20836 399169 -20780
rect 398971 -20978 399027 -20922
rect 399113 -20978 399169 -20922
rect 398971 -21120 399027 -21064
rect 399113 -21120 399169 -21064
rect 398971 -21262 399027 -21206
rect 399113 -21262 399169 -21206
rect 398971 -21404 399027 -21348
rect 399113 -21404 399169 -21348
rect 398971 -21546 399027 -21490
rect 399113 -21546 399169 -21490
rect 398971 -21688 399027 -21632
rect 399113 -21688 399169 -21632
rect 398971 -21830 399027 -21774
rect 399113 -21830 399169 -21774
rect 398971 -21972 399027 -21916
rect 399113 -21972 399169 -21916
rect 398971 -22114 399027 -22058
rect 399113 -22114 399169 -22058
rect 398971 -22256 399027 -22200
rect 399113 -22256 399169 -22200
rect 398971 -22398 399027 -22342
rect 399113 -22398 399169 -22342
rect 398971 -22540 399027 -22484
rect 399113 -22540 399169 -22484
rect 398971 -22682 399027 -22626
rect 399113 -22682 399169 -22626
rect 398971 -22824 399027 -22768
rect 399113 -22824 399169 -22768
rect 398971 -22966 399027 -22910
rect 399113 -22966 399169 -22910
rect 398971 -23108 399027 -23052
rect 399113 -23108 399169 -23052
rect 398971 -23250 399027 -23194
rect 399113 -23250 399169 -23194
rect 398971 -23392 399027 -23336
rect 399113 -23392 399169 -23336
rect 398971 -23534 399027 -23478
rect 399113 -23534 399169 -23478
rect 398971 -23676 399027 -23620
rect 399113 -23676 399169 -23620
rect 398971 -23818 399027 -23762
rect 399113 -23818 399169 -23762
rect 398971 -23960 399027 -23904
rect 399113 -23960 399169 -23904
rect 398971 -24102 399027 -24046
rect 399113 -24102 399169 -24046
rect 398971 -24244 399027 -24188
rect 399113 -24244 399169 -24188
rect 398971 -24386 399027 -24330
rect 399113 -24386 399169 -24330
rect 398971 -24528 399027 -24472
rect 399113 -24528 399169 -24472
rect 398971 -24670 399027 -24614
rect 399113 -24670 399169 -24614
rect 398971 -24812 399027 -24756
rect 399113 -24812 399169 -24756
rect 398971 -24954 399027 -24898
rect 399113 -24954 399169 -24898
rect 398971 -25096 399027 -25040
rect 399113 -25096 399169 -25040
rect 398971 -25238 399027 -25182
rect 399113 -25238 399169 -25182
rect 398971 -25380 399027 -25324
rect 399113 -25380 399169 -25324
rect 398971 -25522 399027 -25466
rect 399113 -25522 399169 -25466
rect 399376 -13736 399432 -13680
rect 399518 -13736 399574 -13680
rect 399376 -13878 399432 -13822
rect 399518 -13878 399574 -13822
rect 399376 -14020 399432 -13964
rect 399518 -14020 399574 -13964
rect 399376 -14162 399432 -14106
rect 399518 -14162 399574 -14106
rect 399376 -14304 399432 -14248
rect 399518 -14304 399574 -14248
rect 399376 -14446 399432 -14390
rect 399518 -14446 399574 -14390
rect 399376 -14588 399432 -14532
rect 399518 -14588 399574 -14532
rect 399376 -14730 399432 -14674
rect 399518 -14730 399574 -14674
rect 399376 -14872 399432 -14816
rect 399518 -14872 399574 -14816
rect 399376 -15014 399432 -14958
rect 399518 -15014 399574 -14958
rect 399376 -15156 399432 -15100
rect 399518 -15156 399574 -15100
rect 399376 -15298 399432 -15242
rect 399518 -15298 399574 -15242
rect 399376 -15440 399432 -15384
rect 399518 -15440 399574 -15384
rect 399376 -15582 399432 -15526
rect 399518 -15582 399574 -15526
rect 399376 -15724 399432 -15668
rect 399518 -15724 399574 -15668
rect 399376 -15866 399432 -15810
rect 399518 -15866 399574 -15810
rect 399376 -16008 399432 -15952
rect 399518 -16008 399574 -15952
rect 399376 -16150 399432 -16094
rect 399518 -16150 399574 -16094
rect 399376 -16292 399432 -16236
rect 399518 -16292 399574 -16236
rect 399376 -16434 399432 -16378
rect 399518 -16434 399574 -16378
rect 399376 -16576 399432 -16520
rect 399518 -16576 399574 -16520
rect 399376 -16718 399432 -16662
rect 399518 -16718 399574 -16662
rect 399376 -16860 399432 -16804
rect 399518 -16860 399574 -16804
rect 399376 -17002 399432 -16946
rect 399518 -17002 399574 -16946
rect 399376 -17144 399432 -17088
rect 399518 -17144 399574 -17088
rect 399376 -17286 399432 -17230
rect 399518 -17286 399574 -17230
rect 399376 -17428 399432 -17372
rect 399518 -17428 399574 -17372
rect 399376 -17570 399432 -17514
rect 399518 -17570 399574 -17514
rect 399376 -17712 399432 -17656
rect 399518 -17712 399574 -17656
rect 399376 -17854 399432 -17798
rect 399518 -17854 399574 -17798
rect 399376 -17996 399432 -17940
rect 399518 -17996 399574 -17940
rect 399376 -18138 399432 -18082
rect 399518 -18138 399574 -18082
rect 399376 -18280 399432 -18224
rect 399518 -18280 399574 -18224
rect 399376 -18422 399432 -18366
rect 399518 -18422 399574 -18366
rect 399376 -18564 399432 -18508
rect 399518 -18564 399574 -18508
rect 399376 -18706 399432 -18650
rect 399518 -18706 399574 -18650
rect 399376 -18848 399432 -18792
rect 399518 -18848 399574 -18792
rect 399376 -18990 399432 -18934
rect 399518 -18990 399574 -18934
rect 399376 -19132 399432 -19076
rect 399518 -19132 399574 -19076
rect 399376 -19274 399432 -19218
rect 399518 -19274 399574 -19218
rect 399376 -19416 399432 -19360
rect 399518 -19416 399574 -19360
rect 399376 -19558 399432 -19502
rect 399518 -19558 399574 -19502
rect 399376 -19700 399432 -19644
rect 399518 -19700 399574 -19644
rect 399376 -19842 399432 -19786
rect 399518 -19842 399574 -19786
rect 399376 -19984 399432 -19928
rect 399518 -19984 399574 -19928
rect 399376 -20126 399432 -20070
rect 399518 -20126 399574 -20070
rect 399376 -20268 399432 -20212
rect 399518 -20268 399574 -20212
rect 399376 -20410 399432 -20354
rect 399518 -20410 399574 -20354
rect 399376 -20552 399432 -20496
rect 399518 -20552 399574 -20496
rect 399376 -20694 399432 -20638
rect 399518 -20694 399574 -20638
rect 399376 -20836 399432 -20780
rect 399518 -20836 399574 -20780
rect 399376 -20978 399432 -20922
rect 399518 -20978 399574 -20922
rect 399376 -21120 399432 -21064
rect 399518 -21120 399574 -21064
rect 399376 -21262 399432 -21206
rect 399518 -21262 399574 -21206
rect 399376 -21404 399432 -21348
rect 399518 -21404 399574 -21348
rect 399376 -21546 399432 -21490
rect 399518 -21546 399574 -21490
rect 399376 -21688 399432 -21632
rect 399518 -21688 399574 -21632
rect 399376 -21830 399432 -21774
rect 399518 -21830 399574 -21774
rect 399376 -21972 399432 -21916
rect 399518 -21972 399574 -21916
rect 399376 -22114 399432 -22058
rect 399518 -22114 399574 -22058
rect 399376 -22256 399432 -22200
rect 399518 -22256 399574 -22200
rect 399376 -22398 399432 -22342
rect 399518 -22398 399574 -22342
rect 399376 -22540 399432 -22484
rect 399518 -22540 399574 -22484
rect 399376 -22682 399432 -22626
rect 399518 -22682 399574 -22626
rect 399376 -22824 399432 -22768
rect 399518 -22824 399574 -22768
rect 399376 -22966 399432 -22910
rect 399518 -22966 399574 -22910
rect 399376 -23108 399432 -23052
rect 399518 -23108 399574 -23052
rect 399376 -23250 399432 -23194
rect 399518 -23250 399574 -23194
rect 399376 -23392 399432 -23336
rect 399518 -23392 399574 -23336
rect 399376 -23534 399432 -23478
rect 399518 -23534 399574 -23478
rect 399376 -23676 399432 -23620
rect 399518 -23676 399574 -23620
rect 399376 -23818 399432 -23762
rect 399518 -23818 399574 -23762
rect 399376 -23960 399432 -23904
rect 399518 -23960 399574 -23904
rect 399376 -24102 399432 -24046
rect 399518 -24102 399574 -24046
rect 399376 -24244 399432 -24188
rect 399518 -24244 399574 -24188
rect 399376 -24386 399432 -24330
rect 399518 -24386 399574 -24330
rect 399376 -24528 399432 -24472
rect 399518 -24528 399574 -24472
rect 399376 -24670 399432 -24614
rect 399518 -24670 399574 -24614
rect 399376 -24812 399432 -24756
rect 399518 -24812 399574 -24756
rect 399376 -24954 399432 -24898
rect 399518 -24954 399574 -24898
rect 399376 -25096 399432 -25040
rect 399518 -25096 399574 -25040
rect 399376 -25238 399432 -25182
rect 399518 -25238 399574 -25182
rect 399376 -25380 399432 -25324
rect 399518 -25380 399574 -25324
rect 399376 -25522 399432 -25466
rect 399518 -25522 399574 -25466
rect 399776 -13736 399832 -13680
rect 399918 -13736 399974 -13680
rect 399776 -13878 399832 -13822
rect 399918 -13878 399974 -13822
rect 399776 -14020 399832 -13964
rect 399918 -14020 399974 -13964
rect 399776 -14162 399832 -14106
rect 399918 -14162 399974 -14106
rect 399776 -14304 399832 -14248
rect 399918 -14304 399974 -14248
rect 399776 -14446 399832 -14390
rect 399918 -14446 399974 -14390
rect 399776 -14588 399832 -14532
rect 399918 -14588 399974 -14532
rect 399776 -14730 399832 -14674
rect 399918 -14730 399974 -14674
rect 399776 -14872 399832 -14816
rect 399918 -14872 399974 -14816
rect 399776 -15014 399832 -14958
rect 399918 -15014 399974 -14958
rect 399776 -15156 399832 -15100
rect 399918 -15156 399974 -15100
rect 399776 -15298 399832 -15242
rect 399918 -15298 399974 -15242
rect 399776 -15440 399832 -15384
rect 399918 -15440 399974 -15384
rect 399776 -15582 399832 -15526
rect 399918 -15582 399974 -15526
rect 399776 -15724 399832 -15668
rect 399918 -15724 399974 -15668
rect 399776 -15866 399832 -15810
rect 399918 -15866 399974 -15810
rect 399776 -16008 399832 -15952
rect 399918 -16008 399974 -15952
rect 399776 -16150 399832 -16094
rect 399918 -16150 399974 -16094
rect 399776 -16292 399832 -16236
rect 399918 -16292 399974 -16236
rect 399776 -16434 399832 -16378
rect 399918 -16434 399974 -16378
rect 399776 -16576 399832 -16520
rect 399918 -16576 399974 -16520
rect 399776 -16718 399832 -16662
rect 399918 -16718 399974 -16662
rect 399776 -16860 399832 -16804
rect 399918 -16860 399974 -16804
rect 399776 -17002 399832 -16946
rect 399918 -17002 399974 -16946
rect 399776 -17144 399832 -17088
rect 399918 -17144 399974 -17088
rect 399776 -17286 399832 -17230
rect 399918 -17286 399974 -17230
rect 399776 -17428 399832 -17372
rect 399918 -17428 399974 -17372
rect 399776 -17570 399832 -17514
rect 399918 -17570 399974 -17514
rect 399776 -17712 399832 -17656
rect 399918 -17712 399974 -17656
rect 399776 -17854 399832 -17798
rect 399918 -17854 399974 -17798
rect 399776 -17996 399832 -17940
rect 399918 -17996 399974 -17940
rect 399776 -18138 399832 -18082
rect 399918 -18138 399974 -18082
rect 399776 -18280 399832 -18224
rect 399918 -18280 399974 -18224
rect 399776 -18422 399832 -18366
rect 399918 -18422 399974 -18366
rect 399776 -18564 399832 -18508
rect 399918 -18564 399974 -18508
rect 399776 -18706 399832 -18650
rect 399918 -18706 399974 -18650
rect 399776 -18848 399832 -18792
rect 399918 -18848 399974 -18792
rect 399776 -18990 399832 -18934
rect 399918 -18990 399974 -18934
rect 399776 -19132 399832 -19076
rect 399918 -19132 399974 -19076
rect 399776 -19274 399832 -19218
rect 399918 -19274 399974 -19218
rect 399776 -19416 399832 -19360
rect 399918 -19416 399974 -19360
rect 399776 -19558 399832 -19502
rect 399918 -19558 399974 -19502
rect 399776 -19700 399832 -19644
rect 399918 -19700 399974 -19644
rect 399776 -19842 399832 -19786
rect 399918 -19842 399974 -19786
rect 399776 -19984 399832 -19928
rect 399918 -19984 399974 -19928
rect 399776 -20126 399832 -20070
rect 399918 -20126 399974 -20070
rect 399776 -20268 399832 -20212
rect 399918 -20268 399974 -20212
rect 399776 -20410 399832 -20354
rect 399918 -20410 399974 -20354
rect 399776 -20552 399832 -20496
rect 399918 -20552 399974 -20496
rect 399776 -20694 399832 -20638
rect 399918 -20694 399974 -20638
rect 399776 -20836 399832 -20780
rect 399918 -20836 399974 -20780
rect 399776 -20978 399832 -20922
rect 399918 -20978 399974 -20922
rect 399776 -21120 399832 -21064
rect 399918 -21120 399974 -21064
rect 399776 -21262 399832 -21206
rect 399918 -21262 399974 -21206
rect 399776 -21404 399832 -21348
rect 399918 -21404 399974 -21348
rect 399776 -21546 399832 -21490
rect 399918 -21546 399974 -21490
rect 399776 -21688 399832 -21632
rect 399918 -21688 399974 -21632
rect 399776 -21830 399832 -21774
rect 399918 -21830 399974 -21774
rect 399776 -21972 399832 -21916
rect 399918 -21972 399974 -21916
rect 399776 -22114 399832 -22058
rect 399918 -22114 399974 -22058
rect 399776 -22256 399832 -22200
rect 399918 -22256 399974 -22200
rect 399776 -22398 399832 -22342
rect 399918 -22398 399974 -22342
rect 399776 -22540 399832 -22484
rect 399918 -22540 399974 -22484
rect 399776 -22682 399832 -22626
rect 399918 -22682 399974 -22626
rect 399776 -22824 399832 -22768
rect 399918 -22824 399974 -22768
rect 399776 -22966 399832 -22910
rect 399918 -22966 399974 -22910
rect 399776 -23108 399832 -23052
rect 399918 -23108 399974 -23052
rect 399776 -23250 399832 -23194
rect 399918 -23250 399974 -23194
rect 399776 -23392 399832 -23336
rect 399918 -23392 399974 -23336
rect 399776 -23534 399832 -23478
rect 399918 -23534 399974 -23478
rect 399776 -23676 399832 -23620
rect 399918 -23676 399974 -23620
rect 399776 -23818 399832 -23762
rect 399918 -23818 399974 -23762
rect 399776 -23960 399832 -23904
rect 399918 -23960 399974 -23904
rect 399776 -24102 399832 -24046
rect 399918 -24102 399974 -24046
rect 399776 -24244 399832 -24188
rect 399918 -24244 399974 -24188
rect 399776 -24386 399832 -24330
rect 399918 -24386 399974 -24330
rect 399776 -24528 399832 -24472
rect 399918 -24528 399974 -24472
rect 399776 -24670 399832 -24614
rect 399918 -24670 399974 -24614
rect 399776 -24812 399832 -24756
rect 399918 -24812 399974 -24756
rect 399776 -24954 399832 -24898
rect 399918 -24954 399974 -24898
rect 399776 -25096 399832 -25040
rect 399918 -25096 399974 -25040
rect 399776 -25238 399832 -25182
rect 399918 -25238 399974 -25182
rect 399776 -25380 399832 -25324
rect 399918 -25380 399974 -25324
rect 399776 -25522 399832 -25466
rect 399918 -25522 399974 -25466
rect 400181 -13736 400237 -13680
rect 400323 -13736 400379 -13680
rect 400181 -13878 400237 -13822
rect 400323 -13878 400379 -13822
rect 400181 -14020 400237 -13964
rect 400323 -14020 400379 -13964
rect 400181 -14162 400237 -14106
rect 400323 -14162 400379 -14106
rect 400181 -14304 400237 -14248
rect 400323 -14304 400379 -14248
rect 400181 -14446 400237 -14390
rect 400323 -14446 400379 -14390
rect 400181 -14588 400237 -14532
rect 400323 -14588 400379 -14532
rect 400181 -14730 400237 -14674
rect 400323 -14730 400379 -14674
rect 400181 -14872 400237 -14816
rect 400323 -14872 400379 -14816
rect 400181 -15014 400237 -14958
rect 400323 -15014 400379 -14958
rect 400181 -15156 400237 -15100
rect 400323 -15156 400379 -15100
rect 400181 -15298 400237 -15242
rect 400323 -15298 400379 -15242
rect 400181 -15440 400237 -15384
rect 400323 -15440 400379 -15384
rect 400181 -15582 400237 -15526
rect 400323 -15582 400379 -15526
rect 400181 -15724 400237 -15668
rect 400323 -15724 400379 -15668
rect 400181 -15866 400237 -15810
rect 400323 -15866 400379 -15810
rect 400181 -16008 400237 -15952
rect 400323 -16008 400379 -15952
rect 400181 -16150 400237 -16094
rect 400323 -16150 400379 -16094
rect 400181 -16292 400237 -16236
rect 400323 -16292 400379 -16236
rect 400181 -16434 400237 -16378
rect 400323 -16434 400379 -16378
rect 400181 -16576 400237 -16520
rect 400323 -16576 400379 -16520
rect 400181 -16718 400237 -16662
rect 400323 -16718 400379 -16662
rect 400181 -16860 400237 -16804
rect 400323 -16860 400379 -16804
rect 400181 -17002 400237 -16946
rect 400323 -17002 400379 -16946
rect 400181 -17144 400237 -17088
rect 400323 -17144 400379 -17088
rect 400181 -17286 400237 -17230
rect 400323 -17286 400379 -17230
rect 400181 -17428 400237 -17372
rect 400323 -17428 400379 -17372
rect 400181 -17570 400237 -17514
rect 400323 -17570 400379 -17514
rect 400181 -17712 400237 -17656
rect 400323 -17712 400379 -17656
rect 400181 -17854 400237 -17798
rect 400323 -17854 400379 -17798
rect 400181 -17996 400237 -17940
rect 400323 -17996 400379 -17940
rect 400181 -18138 400237 -18082
rect 400323 -18138 400379 -18082
rect 400181 -18280 400237 -18224
rect 400323 -18280 400379 -18224
rect 400181 -18422 400237 -18366
rect 400323 -18422 400379 -18366
rect 400181 -18564 400237 -18508
rect 400323 -18564 400379 -18508
rect 400181 -18706 400237 -18650
rect 400323 -18706 400379 -18650
rect 400181 -18848 400237 -18792
rect 400323 -18848 400379 -18792
rect 400181 -18990 400237 -18934
rect 400323 -18990 400379 -18934
rect 400181 -19132 400237 -19076
rect 400323 -19132 400379 -19076
rect 400181 -19274 400237 -19218
rect 400323 -19274 400379 -19218
rect 400181 -19416 400237 -19360
rect 400323 -19416 400379 -19360
rect 400181 -19558 400237 -19502
rect 400323 -19558 400379 -19502
rect 400181 -19700 400237 -19644
rect 400323 -19700 400379 -19644
rect 400181 -19842 400237 -19786
rect 400323 -19842 400379 -19786
rect 400181 -19984 400237 -19928
rect 400323 -19984 400379 -19928
rect 400181 -20126 400237 -20070
rect 400323 -20126 400379 -20070
rect 400181 -20268 400237 -20212
rect 400323 -20268 400379 -20212
rect 400181 -20410 400237 -20354
rect 400323 -20410 400379 -20354
rect 400181 -20552 400237 -20496
rect 400323 -20552 400379 -20496
rect 400181 -20694 400237 -20638
rect 400323 -20694 400379 -20638
rect 400181 -20836 400237 -20780
rect 400323 -20836 400379 -20780
rect 400181 -20978 400237 -20922
rect 400323 -20978 400379 -20922
rect 400181 -21120 400237 -21064
rect 400323 -21120 400379 -21064
rect 400181 -21262 400237 -21206
rect 400323 -21262 400379 -21206
rect 400181 -21404 400237 -21348
rect 400323 -21404 400379 -21348
rect 400181 -21546 400237 -21490
rect 400323 -21546 400379 -21490
rect 400181 -21688 400237 -21632
rect 400323 -21688 400379 -21632
rect 400181 -21830 400237 -21774
rect 400323 -21830 400379 -21774
rect 400181 -21972 400237 -21916
rect 400323 -21972 400379 -21916
rect 400181 -22114 400237 -22058
rect 400323 -22114 400379 -22058
rect 400181 -22256 400237 -22200
rect 400323 -22256 400379 -22200
rect 400181 -22398 400237 -22342
rect 400323 -22398 400379 -22342
rect 400181 -22540 400237 -22484
rect 400323 -22540 400379 -22484
rect 400181 -22682 400237 -22626
rect 400323 -22682 400379 -22626
rect 400181 -22824 400237 -22768
rect 400323 -22824 400379 -22768
rect 400181 -22966 400237 -22910
rect 400323 -22966 400379 -22910
rect 400181 -23108 400237 -23052
rect 400323 -23108 400379 -23052
rect 400181 -23250 400237 -23194
rect 400323 -23250 400379 -23194
rect 400181 -23392 400237 -23336
rect 400323 -23392 400379 -23336
rect 400181 -23534 400237 -23478
rect 400323 -23534 400379 -23478
rect 400181 -23676 400237 -23620
rect 400323 -23676 400379 -23620
rect 400181 -23818 400237 -23762
rect 400323 -23818 400379 -23762
rect 400181 -23960 400237 -23904
rect 400323 -23960 400379 -23904
rect 400181 -24102 400237 -24046
rect 400323 -24102 400379 -24046
rect 400181 -24244 400237 -24188
rect 400323 -24244 400379 -24188
rect 400181 -24386 400237 -24330
rect 400323 -24386 400379 -24330
rect 400181 -24528 400237 -24472
rect 400323 -24528 400379 -24472
rect 400181 -24670 400237 -24614
rect 400323 -24670 400379 -24614
rect 400181 -24812 400237 -24756
rect 400323 -24812 400379 -24756
rect 400181 -24954 400237 -24898
rect 400323 -24954 400379 -24898
rect 400181 -25096 400237 -25040
rect 400323 -25096 400379 -25040
rect 400181 -25238 400237 -25182
rect 400323 -25238 400379 -25182
rect 400181 -25380 400237 -25324
rect 400323 -25380 400379 -25324
rect 400181 -25522 400237 -25466
rect 400323 -25522 400379 -25466
rect 400766 -13688 400822 -13632
rect 400890 -13688 400946 -13632
rect 401014 -13688 401070 -13632
rect 401138 -13688 401194 -13632
rect 401262 -13688 401318 -13632
rect 400766 -13812 400822 -13756
rect 400890 -13812 400946 -13756
rect 401014 -13812 401070 -13756
rect 401138 -13812 401194 -13756
rect 401262 -13812 401318 -13756
rect 400766 -13936 400822 -13880
rect 400890 -13936 400946 -13880
rect 401014 -13936 401070 -13880
rect 401138 -13936 401194 -13880
rect 401262 -13936 401318 -13880
rect 400766 -14060 400822 -14004
rect 400890 -14060 400946 -14004
rect 401014 -14060 401070 -14004
rect 401138 -14060 401194 -14004
rect 401262 -14060 401318 -14004
rect 400766 -14184 400822 -14128
rect 400890 -14184 400946 -14128
rect 401014 -14184 401070 -14128
rect 401138 -14184 401194 -14128
rect 401262 -14184 401318 -14128
rect 400766 -14308 400822 -14252
rect 400890 -14308 400946 -14252
rect 401014 -14308 401070 -14252
rect 401138 -14308 401194 -14252
rect 401262 -14308 401318 -14252
rect 400766 -14432 400822 -14376
rect 400890 -14432 400946 -14376
rect 401014 -14432 401070 -14376
rect 401138 -14432 401194 -14376
rect 401262 -14432 401318 -14376
rect 400766 -14556 400822 -14500
rect 400890 -14556 400946 -14500
rect 401014 -14556 401070 -14500
rect 401138 -14556 401194 -14500
rect 401262 -14556 401318 -14500
rect 400766 -14680 400822 -14624
rect 400890 -14680 400946 -14624
rect 401014 -14680 401070 -14624
rect 401138 -14680 401194 -14624
rect 401262 -14680 401318 -14624
rect 400766 -14804 400822 -14748
rect 400890 -14804 400946 -14748
rect 401014 -14804 401070 -14748
rect 401138 -14804 401194 -14748
rect 401262 -14804 401318 -14748
rect 400766 -14928 400822 -14872
rect 400890 -14928 400946 -14872
rect 401014 -14928 401070 -14872
rect 401138 -14928 401194 -14872
rect 401262 -14928 401318 -14872
rect 400766 -15052 400822 -14996
rect 400890 -15052 400946 -14996
rect 401014 -15052 401070 -14996
rect 401138 -15052 401194 -14996
rect 401262 -15052 401318 -14996
rect 400766 -15176 400822 -15120
rect 400890 -15176 400946 -15120
rect 401014 -15176 401070 -15120
rect 401138 -15176 401194 -15120
rect 401262 -15176 401318 -15120
rect 400766 -15300 400822 -15244
rect 400890 -15300 400946 -15244
rect 401014 -15300 401070 -15244
rect 401138 -15300 401194 -15244
rect 401262 -15300 401318 -15244
rect 400766 -15424 400822 -15368
rect 400890 -15424 400946 -15368
rect 401014 -15424 401070 -15368
rect 401138 -15424 401194 -15368
rect 401262 -15424 401318 -15368
rect 400766 -15548 400822 -15492
rect 400890 -15548 400946 -15492
rect 401014 -15548 401070 -15492
rect 401138 -15548 401194 -15492
rect 401262 -15548 401318 -15492
rect 400766 -15672 400822 -15616
rect 400890 -15672 400946 -15616
rect 401014 -15672 401070 -15616
rect 401138 -15672 401194 -15616
rect 401262 -15672 401318 -15616
rect 400766 -15796 400822 -15740
rect 400890 -15796 400946 -15740
rect 401014 -15796 401070 -15740
rect 401138 -15796 401194 -15740
rect 401262 -15796 401318 -15740
rect 400766 -15920 400822 -15864
rect 400890 -15920 400946 -15864
rect 401014 -15920 401070 -15864
rect 401138 -15920 401194 -15864
rect 401262 -15920 401318 -15864
rect 400766 -16044 400822 -15988
rect 400890 -16044 400946 -15988
rect 401014 -16044 401070 -15988
rect 401138 -16044 401194 -15988
rect 401262 -16044 401318 -15988
rect 400766 -16168 400822 -16112
rect 400890 -16168 400946 -16112
rect 401014 -16168 401070 -16112
rect 401138 -16168 401194 -16112
rect 401262 -16168 401318 -16112
rect 400766 -16292 400822 -16236
rect 400890 -16292 400946 -16236
rect 401014 -16292 401070 -16236
rect 401138 -16292 401194 -16236
rect 401262 -16292 401318 -16236
rect 400766 -16416 400822 -16360
rect 400890 -16416 400946 -16360
rect 401014 -16416 401070 -16360
rect 401138 -16416 401194 -16360
rect 401262 -16416 401318 -16360
rect 400766 -16540 400822 -16484
rect 400890 -16540 400946 -16484
rect 401014 -16540 401070 -16484
rect 401138 -16540 401194 -16484
rect 401262 -16540 401318 -16484
rect 400766 -16664 400822 -16608
rect 400890 -16664 400946 -16608
rect 401014 -16664 401070 -16608
rect 401138 -16664 401194 -16608
rect 401262 -16664 401318 -16608
rect 400766 -16788 400822 -16732
rect 400890 -16788 400946 -16732
rect 401014 -16788 401070 -16732
rect 401138 -16788 401194 -16732
rect 401262 -16788 401318 -16732
rect 400766 -16912 400822 -16856
rect 400890 -16912 400946 -16856
rect 401014 -16912 401070 -16856
rect 401138 -16912 401194 -16856
rect 401262 -16912 401318 -16856
rect 400766 -17036 400822 -16980
rect 400890 -17036 400946 -16980
rect 401014 -17036 401070 -16980
rect 401138 -17036 401194 -16980
rect 401262 -17036 401318 -16980
rect 400766 -17160 400822 -17104
rect 400890 -17160 400946 -17104
rect 401014 -17160 401070 -17104
rect 401138 -17160 401194 -17104
rect 401262 -17160 401318 -17104
rect 400766 -17284 400822 -17228
rect 400890 -17284 400946 -17228
rect 401014 -17284 401070 -17228
rect 401138 -17284 401194 -17228
rect 401262 -17284 401318 -17228
rect 400766 -17408 400822 -17352
rect 400890 -17408 400946 -17352
rect 401014 -17408 401070 -17352
rect 401138 -17408 401194 -17352
rect 401262 -17408 401318 -17352
rect 400766 -17532 400822 -17476
rect 400890 -17532 400946 -17476
rect 401014 -17532 401070 -17476
rect 401138 -17532 401194 -17476
rect 401262 -17532 401318 -17476
rect 400766 -17656 400822 -17600
rect 400890 -17656 400946 -17600
rect 401014 -17656 401070 -17600
rect 401138 -17656 401194 -17600
rect 401262 -17656 401318 -17600
rect 400766 -17780 400822 -17724
rect 400890 -17780 400946 -17724
rect 401014 -17780 401070 -17724
rect 401138 -17780 401194 -17724
rect 401262 -17780 401318 -17724
rect 400766 -17904 400822 -17848
rect 400890 -17904 400946 -17848
rect 401014 -17904 401070 -17848
rect 401138 -17904 401194 -17848
rect 401262 -17904 401318 -17848
rect 400766 -18028 400822 -17972
rect 400890 -18028 400946 -17972
rect 401014 -18028 401070 -17972
rect 401138 -18028 401194 -17972
rect 401262 -18028 401318 -17972
rect 400766 -18152 400822 -18096
rect 400890 -18152 400946 -18096
rect 401014 -18152 401070 -18096
rect 401138 -18152 401194 -18096
rect 401262 -18152 401318 -18096
rect 400766 -18276 400822 -18220
rect 400890 -18276 400946 -18220
rect 401014 -18276 401070 -18220
rect 401138 -18276 401194 -18220
rect 401262 -18276 401318 -18220
rect 400766 -18400 400822 -18344
rect 400890 -18400 400946 -18344
rect 401014 -18400 401070 -18344
rect 401138 -18400 401194 -18344
rect 401262 -18400 401318 -18344
rect 400766 -18524 400822 -18468
rect 400890 -18524 400946 -18468
rect 401014 -18524 401070 -18468
rect 401138 -18524 401194 -18468
rect 401262 -18524 401318 -18468
rect 400766 -18648 400822 -18592
rect 400890 -18648 400946 -18592
rect 401014 -18648 401070 -18592
rect 401138 -18648 401194 -18592
rect 401262 -18648 401318 -18592
rect 400766 -18772 400822 -18716
rect 400890 -18772 400946 -18716
rect 401014 -18772 401070 -18716
rect 401138 -18772 401194 -18716
rect 401262 -18772 401318 -18716
rect 400766 -18896 400822 -18840
rect 400890 -18896 400946 -18840
rect 401014 -18896 401070 -18840
rect 401138 -18896 401194 -18840
rect 401262 -18896 401318 -18840
rect 400766 -19020 400822 -18964
rect 400890 -19020 400946 -18964
rect 401014 -19020 401070 -18964
rect 401138 -19020 401194 -18964
rect 401262 -19020 401318 -18964
rect 400766 -19144 400822 -19088
rect 400890 -19144 400946 -19088
rect 401014 -19144 401070 -19088
rect 401138 -19144 401194 -19088
rect 401262 -19144 401318 -19088
rect 400766 -19268 400822 -19212
rect 400890 -19268 400946 -19212
rect 401014 -19268 401070 -19212
rect 401138 -19268 401194 -19212
rect 401262 -19268 401318 -19212
rect 400766 -19392 400822 -19336
rect 400890 -19392 400946 -19336
rect 401014 -19392 401070 -19336
rect 401138 -19392 401194 -19336
rect 401262 -19392 401318 -19336
rect 400766 -19516 400822 -19460
rect 400890 -19516 400946 -19460
rect 401014 -19516 401070 -19460
rect 401138 -19516 401194 -19460
rect 401262 -19516 401318 -19460
rect 400766 -19640 400822 -19584
rect 400890 -19640 400946 -19584
rect 401014 -19640 401070 -19584
rect 401138 -19640 401194 -19584
rect 401262 -19640 401318 -19584
rect 400766 -19764 400822 -19708
rect 400890 -19764 400946 -19708
rect 401014 -19764 401070 -19708
rect 401138 -19764 401194 -19708
rect 401262 -19764 401318 -19708
rect 400766 -19888 400822 -19832
rect 400890 -19888 400946 -19832
rect 401014 -19888 401070 -19832
rect 401138 -19888 401194 -19832
rect 401262 -19888 401318 -19832
rect 400766 -20012 400822 -19956
rect 400890 -20012 400946 -19956
rect 401014 -20012 401070 -19956
rect 401138 -20012 401194 -19956
rect 401262 -20012 401318 -19956
rect 400766 -20136 400822 -20080
rect 400890 -20136 400946 -20080
rect 401014 -20136 401070 -20080
rect 401138 -20136 401194 -20080
rect 401262 -20136 401318 -20080
rect 400766 -20260 400822 -20204
rect 400890 -20260 400946 -20204
rect 401014 -20260 401070 -20204
rect 401138 -20260 401194 -20204
rect 401262 -20260 401318 -20204
rect 400766 -20384 400822 -20328
rect 400890 -20384 400946 -20328
rect 401014 -20384 401070 -20328
rect 401138 -20384 401194 -20328
rect 401262 -20384 401318 -20328
rect 400766 -20508 400822 -20452
rect 400890 -20508 400946 -20452
rect 401014 -20508 401070 -20452
rect 401138 -20508 401194 -20452
rect 401262 -20508 401318 -20452
rect 400766 -20632 400822 -20576
rect 400890 -20632 400946 -20576
rect 401014 -20632 401070 -20576
rect 401138 -20632 401194 -20576
rect 401262 -20632 401318 -20576
rect 400766 -20756 400822 -20700
rect 400890 -20756 400946 -20700
rect 401014 -20756 401070 -20700
rect 401138 -20756 401194 -20700
rect 401262 -20756 401318 -20700
rect 400766 -20880 400822 -20824
rect 400890 -20880 400946 -20824
rect 401014 -20880 401070 -20824
rect 401138 -20880 401194 -20824
rect 401262 -20880 401318 -20824
rect 400766 -21004 400822 -20948
rect 400890 -21004 400946 -20948
rect 401014 -21004 401070 -20948
rect 401138 -21004 401194 -20948
rect 401262 -21004 401318 -20948
rect 400766 -21128 400822 -21072
rect 400890 -21128 400946 -21072
rect 401014 -21128 401070 -21072
rect 401138 -21128 401194 -21072
rect 401262 -21128 401318 -21072
rect 400766 -21252 400822 -21196
rect 400890 -21252 400946 -21196
rect 401014 -21252 401070 -21196
rect 401138 -21252 401194 -21196
rect 401262 -21252 401318 -21196
rect 400766 -21376 400822 -21320
rect 400890 -21376 400946 -21320
rect 401014 -21376 401070 -21320
rect 401138 -21376 401194 -21320
rect 401262 -21376 401318 -21320
rect 400766 -21500 400822 -21444
rect 400890 -21500 400946 -21444
rect 401014 -21500 401070 -21444
rect 401138 -21500 401194 -21444
rect 401262 -21500 401318 -21444
rect 400766 -21624 400822 -21568
rect 400890 -21624 400946 -21568
rect 401014 -21624 401070 -21568
rect 401138 -21624 401194 -21568
rect 401262 -21624 401318 -21568
rect 400766 -21748 400822 -21692
rect 400890 -21748 400946 -21692
rect 401014 -21748 401070 -21692
rect 401138 -21748 401194 -21692
rect 401262 -21748 401318 -21692
rect 400766 -21872 400822 -21816
rect 400890 -21872 400946 -21816
rect 401014 -21872 401070 -21816
rect 401138 -21872 401194 -21816
rect 401262 -21872 401318 -21816
rect 400766 -21996 400822 -21940
rect 400890 -21996 400946 -21940
rect 401014 -21996 401070 -21940
rect 401138 -21996 401194 -21940
rect 401262 -21996 401318 -21940
rect 400766 -22120 400822 -22064
rect 400890 -22120 400946 -22064
rect 401014 -22120 401070 -22064
rect 401138 -22120 401194 -22064
rect 401262 -22120 401318 -22064
rect 400766 -22244 400822 -22188
rect 400890 -22244 400946 -22188
rect 401014 -22244 401070 -22188
rect 401138 -22244 401194 -22188
rect 401262 -22244 401318 -22188
rect 400766 -22368 400822 -22312
rect 400890 -22368 400946 -22312
rect 401014 -22368 401070 -22312
rect 401138 -22368 401194 -22312
rect 401262 -22368 401318 -22312
rect 400766 -22492 400822 -22436
rect 400890 -22492 400946 -22436
rect 401014 -22492 401070 -22436
rect 401138 -22492 401194 -22436
rect 401262 -22492 401318 -22436
rect 400766 -22616 400822 -22560
rect 400890 -22616 400946 -22560
rect 401014 -22616 401070 -22560
rect 401138 -22616 401194 -22560
rect 401262 -22616 401318 -22560
rect 400766 -22740 400822 -22684
rect 400890 -22740 400946 -22684
rect 401014 -22740 401070 -22684
rect 401138 -22740 401194 -22684
rect 401262 -22740 401318 -22684
rect 400766 -22864 400822 -22808
rect 400890 -22864 400946 -22808
rect 401014 -22864 401070 -22808
rect 401138 -22864 401194 -22808
rect 401262 -22864 401318 -22808
rect 400766 -22988 400822 -22932
rect 400890 -22988 400946 -22932
rect 401014 -22988 401070 -22932
rect 401138 -22988 401194 -22932
rect 401262 -22988 401318 -22932
rect 400766 -23112 400822 -23056
rect 400890 -23112 400946 -23056
rect 401014 -23112 401070 -23056
rect 401138 -23112 401194 -23056
rect 401262 -23112 401318 -23056
rect 400766 -23236 400822 -23180
rect 400890 -23236 400946 -23180
rect 401014 -23236 401070 -23180
rect 401138 -23236 401194 -23180
rect 401262 -23236 401318 -23180
rect 400766 -23360 400822 -23304
rect 400890 -23360 400946 -23304
rect 401014 -23360 401070 -23304
rect 401138 -23360 401194 -23304
rect 401262 -23360 401318 -23304
rect 400766 -23484 400822 -23428
rect 400890 -23484 400946 -23428
rect 401014 -23484 401070 -23428
rect 401138 -23484 401194 -23428
rect 401262 -23484 401318 -23428
rect 400766 -23608 400822 -23552
rect 400890 -23608 400946 -23552
rect 401014 -23608 401070 -23552
rect 401138 -23608 401194 -23552
rect 401262 -23608 401318 -23552
rect 400766 -23732 400822 -23676
rect 400890 -23732 400946 -23676
rect 401014 -23732 401070 -23676
rect 401138 -23732 401194 -23676
rect 401262 -23732 401318 -23676
rect 400766 -23856 400822 -23800
rect 400890 -23856 400946 -23800
rect 401014 -23856 401070 -23800
rect 401138 -23856 401194 -23800
rect 401262 -23856 401318 -23800
rect 400766 -23980 400822 -23924
rect 400890 -23980 400946 -23924
rect 401014 -23980 401070 -23924
rect 401138 -23980 401194 -23924
rect 401262 -23980 401318 -23924
rect 400766 -24104 400822 -24048
rect 400890 -24104 400946 -24048
rect 401014 -24104 401070 -24048
rect 401138 -24104 401194 -24048
rect 401262 -24104 401318 -24048
rect 400766 -24228 400822 -24172
rect 400890 -24228 400946 -24172
rect 401014 -24228 401070 -24172
rect 401138 -24228 401194 -24172
rect 401262 -24228 401318 -24172
rect 400766 -24352 400822 -24296
rect 400890 -24352 400946 -24296
rect 401014 -24352 401070 -24296
rect 401138 -24352 401194 -24296
rect 401262 -24352 401318 -24296
rect 400766 -24476 400822 -24420
rect 400890 -24476 400946 -24420
rect 401014 -24476 401070 -24420
rect 401138 -24476 401194 -24420
rect 401262 -24476 401318 -24420
rect 400766 -24600 400822 -24544
rect 400890 -24600 400946 -24544
rect 401014 -24600 401070 -24544
rect 401138 -24600 401194 -24544
rect 401262 -24600 401318 -24544
rect 400766 -24724 400822 -24668
rect 400890 -24724 400946 -24668
rect 401014 -24724 401070 -24668
rect 401138 -24724 401194 -24668
rect 401262 -24724 401318 -24668
rect 400766 -24848 400822 -24792
rect 400890 -24848 400946 -24792
rect 401014 -24848 401070 -24792
rect 401138 -24848 401194 -24792
rect 401262 -24848 401318 -24792
rect 400766 -24972 400822 -24916
rect 400890 -24972 400946 -24916
rect 401014 -24972 401070 -24916
rect 401138 -24972 401194 -24916
rect 401262 -24972 401318 -24916
rect 400766 -25096 400822 -25040
rect 400890 -25096 400946 -25040
rect 401014 -25096 401070 -25040
rect 401138 -25096 401194 -25040
rect 401262 -25096 401318 -25040
rect 400766 -25220 400822 -25164
rect 400890 -25220 400946 -25164
rect 401014 -25220 401070 -25164
rect 401138 -25220 401194 -25164
rect 401262 -25220 401318 -25164
rect 400766 -25344 400822 -25288
rect 400890 -25344 400946 -25288
rect 401014 -25344 401070 -25288
rect 401138 -25344 401194 -25288
rect 401262 -25344 401318 -25288
rect 400766 -25468 400822 -25412
rect 400890 -25468 400946 -25412
rect 401014 -25468 401070 -25412
rect 401138 -25468 401194 -25412
rect 401262 -25468 401318 -25412
rect 400766 -25592 400822 -25536
rect 400890 -25592 400946 -25536
rect 401014 -25592 401070 -25536
rect 401138 -25592 401194 -25536
rect 401262 -25592 401318 -25536
rect 387954 -25716 388010 -25660
rect 388078 -25716 388134 -25660
rect 388202 -25716 388258 -25660
rect 388326 -25716 388382 -25660
rect 388450 -25716 388506 -25660
rect 388655 -25744 388711 -25688
rect 388797 -25744 388853 -25688
rect 388939 -25744 388995 -25688
rect 389081 -25744 389137 -25688
rect 389223 -25744 389279 -25688
rect 389365 -25744 389421 -25688
rect 389507 -25744 389563 -25688
rect 389649 -25744 389705 -25688
rect 389791 -25744 389847 -25688
rect 389933 -25744 389989 -25688
rect 390075 -25744 390131 -25688
rect 390217 -25744 390273 -25688
rect 390359 -25744 390415 -25688
rect 390501 -25744 390557 -25688
rect 390643 -25744 390699 -25688
rect 390785 -25744 390841 -25688
rect 390927 -25744 390983 -25688
rect 391069 -25744 391125 -25688
rect 391211 -25744 391267 -25688
rect 391353 -25744 391409 -25688
rect 391495 -25744 391551 -25688
rect 391637 -25744 391693 -25688
rect 391779 -25744 391835 -25688
rect 391921 -25744 391977 -25688
rect 392063 -25744 392119 -25688
rect 392205 -25744 392261 -25688
rect 392347 -25744 392403 -25688
rect 392489 -25744 392545 -25688
rect 392631 -25744 392687 -25688
rect 392773 -25744 392829 -25688
rect 392915 -25744 392971 -25688
rect 393057 -25744 393113 -25688
rect 393199 -25744 393255 -25688
rect 393341 -25744 393397 -25688
rect 393483 -25744 393539 -25688
rect 393625 -25744 393681 -25688
rect 393767 -25744 393823 -25688
rect 393909 -25744 393965 -25688
rect 394051 -25744 394107 -25688
rect 394193 -25744 394249 -25688
rect 394335 -25744 394391 -25688
rect 394477 -25744 394533 -25688
rect 394619 -25744 394675 -25688
rect 394761 -25744 394817 -25688
rect 394903 -25744 394959 -25688
rect 395045 -25744 395101 -25688
rect 395187 -25744 395243 -25688
rect 395329 -25744 395385 -25688
rect 395471 -25744 395527 -25688
rect 395613 -25744 395669 -25688
rect 395755 -25744 395811 -25688
rect 395897 -25744 395953 -25688
rect 396039 -25744 396095 -25688
rect 396181 -25744 396237 -25688
rect 396323 -25744 396379 -25688
rect 396465 -25744 396521 -25688
rect 396607 -25744 396663 -25688
rect 396749 -25744 396805 -25688
rect 396891 -25744 396947 -25688
rect 397033 -25744 397089 -25688
rect 397175 -25744 397231 -25688
rect 397317 -25744 397373 -25688
rect 397459 -25744 397515 -25688
rect 397601 -25744 397657 -25688
rect 397743 -25744 397799 -25688
rect 397885 -25744 397941 -25688
rect 398027 -25744 398083 -25688
rect 398169 -25744 398225 -25688
rect 398311 -25744 398367 -25688
rect 398453 -25744 398509 -25688
rect 398595 -25744 398651 -25688
rect 398737 -25744 398793 -25688
rect 398879 -25744 398935 -25688
rect 399021 -25744 399077 -25688
rect 399163 -25744 399219 -25688
rect 399305 -25744 399361 -25688
rect 399447 -25744 399503 -25688
rect 399589 -25744 399645 -25688
rect 399731 -25744 399787 -25688
rect 399873 -25744 399929 -25688
rect 400015 -25744 400071 -25688
rect 400157 -25744 400213 -25688
rect 400299 -25744 400355 -25688
rect 400441 -25744 400497 -25688
rect 400583 -25744 400639 -25688
rect 400766 -25716 400822 -25660
rect 400890 -25716 400946 -25660
rect 401014 -25716 401070 -25660
rect 401138 -25716 401194 -25660
rect 401262 -25716 401318 -25660
rect 387954 -25840 388010 -25784
rect 388078 -25840 388134 -25784
rect 388202 -25840 388258 -25784
rect 388326 -25840 388382 -25784
rect 388450 -25840 388506 -25784
rect 388655 -25886 388711 -25830
rect 388797 -25886 388853 -25830
rect 388939 -25886 388995 -25830
rect 389081 -25886 389137 -25830
rect 389223 -25886 389279 -25830
rect 389365 -25886 389421 -25830
rect 389507 -25886 389563 -25830
rect 389649 -25886 389705 -25830
rect 389791 -25886 389847 -25830
rect 389933 -25886 389989 -25830
rect 390075 -25886 390131 -25830
rect 390217 -25886 390273 -25830
rect 390359 -25886 390415 -25830
rect 390501 -25886 390557 -25830
rect 390643 -25886 390699 -25830
rect 390785 -25886 390841 -25830
rect 390927 -25886 390983 -25830
rect 391069 -25886 391125 -25830
rect 391211 -25886 391267 -25830
rect 391353 -25886 391409 -25830
rect 391495 -25886 391551 -25830
rect 391637 -25886 391693 -25830
rect 391779 -25886 391835 -25830
rect 391921 -25886 391977 -25830
rect 392063 -25886 392119 -25830
rect 392205 -25886 392261 -25830
rect 392347 -25886 392403 -25830
rect 392489 -25886 392545 -25830
rect 392631 -25886 392687 -25830
rect 392773 -25886 392829 -25830
rect 392915 -25886 392971 -25830
rect 393057 -25886 393113 -25830
rect 393199 -25886 393255 -25830
rect 393341 -25886 393397 -25830
rect 393483 -25886 393539 -25830
rect 393625 -25886 393681 -25830
rect 393767 -25886 393823 -25830
rect 393909 -25886 393965 -25830
rect 394051 -25886 394107 -25830
rect 394193 -25886 394249 -25830
rect 394335 -25886 394391 -25830
rect 394477 -25886 394533 -25830
rect 394619 -25886 394675 -25830
rect 394761 -25886 394817 -25830
rect 394903 -25886 394959 -25830
rect 395045 -25886 395101 -25830
rect 395187 -25886 395243 -25830
rect 395329 -25886 395385 -25830
rect 395471 -25886 395527 -25830
rect 395613 -25886 395669 -25830
rect 395755 -25886 395811 -25830
rect 395897 -25886 395953 -25830
rect 396039 -25886 396095 -25830
rect 396181 -25886 396237 -25830
rect 396323 -25886 396379 -25830
rect 396465 -25886 396521 -25830
rect 396607 -25886 396663 -25830
rect 396749 -25886 396805 -25830
rect 396891 -25886 396947 -25830
rect 397033 -25886 397089 -25830
rect 397175 -25886 397231 -25830
rect 397317 -25886 397373 -25830
rect 397459 -25886 397515 -25830
rect 397601 -25886 397657 -25830
rect 397743 -25886 397799 -25830
rect 397885 -25886 397941 -25830
rect 398027 -25886 398083 -25830
rect 398169 -25886 398225 -25830
rect 398311 -25886 398367 -25830
rect 398453 -25886 398509 -25830
rect 398595 -25886 398651 -25830
rect 398737 -25886 398793 -25830
rect 398879 -25886 398935 -25830
rect 399021 -25886 399077 -25830
rect 399163 -25886 399219 -25830
rect 399305 -25886 399361 -25830
rect 399447 -25886 399503 -25830
rect 399589 -25886 399645 -25830
rect 399731 -25886 399787 -25830
rect 399873 -25886 399929 -25830
rect 400015 -25886 400071 -25830
rect 400157 -25886 400213 -25830
rect 400299 -25886 400355 -25830
rect 400441 -25886 400497 -25830
rect 400583 -25886 400639 -25830
rect 400766 -25840 400822 -25784
rect 400890 -25840 400946 -25784
rect 401014 -25840 401070 -25784
rect 401138 -25840 401194 -25784
rect 401262 -25840 401318 -25784
<< metal3 >>
rect 387840 -13041 401440 -12925
rect 387840 -13097 387986 -13041
rect 388042 -13097 388110 -13041
rect 388166 -13097 388234 -13041
rect 388290 -13097 388358 -13041
rect 388414 -13097 388482 -13041
rect 388538 -13097 388606 -13041
rect 388662 -13097 388730 -13041
rect 388786 -13097 388854 -13041
rect 388910 -13097 388978 -13041
rect 389034 -13097 389102 -13041
rect 389158 -13097 389226 -13041
rect 389282 -13097 389350 -13041
rect 389406 -13097 389474 -13041
rect 389530 -13097 389598 -13041
rect 389654 -13097 389722 -13041
rect 389778 -13097 389846 -13041
rect 389902 -13097 389970 -13041
rect 390026 -13097 390094 -13041
rect 390150 -13097 390218 -13041
rect 390274 -13097 390342 -13041
rect 390398 -13097 390466 -13041
rect 390522 -13097 390590 -13041
rect 390646 -13097 390714 -13041
rect 390770 -13097 390838 -13041
rect 390894 -13097 390962 -13041
rect 391018 -13097 391086 -13041
rect 391142 -13097 391210 -13041
rect 391266 -13097 391334 -13041
rect 391390 -13097 391458 -13041
rect 391514 -13097 391582 -13041
rect 391638 -13097 391706 -13041
rect 391762 -13097 391830 -13041
rect 391886 -13097 391954 -13041
rect 392010 -13097 392078 -13041
rect 392134 -13097 392202 -13041
rect 392258 -13097 392326 -13041
rect 392382 -13097 392450 -13041
rect 392506 -13097 392574 -13041
rect 392630 -13097 392698 -13041
rect 392754 -13097 392822 -13041
rect 392878 -13097 392946 -13041
rect 393002 -13097 393070 -13041
rect 393126 -13097 393194 -13041
rect 393250 -13097 393318 -13041
rect 393374 -13097 393442 -13041
rect 393498 -13097 393566 -13041
rect 393622 -13097 393690 -13041
rect 393746 -13097 393814 -13041
rect 393870 -13097 393938 -13041
rect 393994 -13097 394062 -13041
rect 394118 -13097 394186 -13041
rect 394242 -13097 394310 -13041
rect 394366 -13097 394434 -13041
rect 394490 -13097 394558 -13041
rect 394614 -13097 394682 -13041
rect 394738 -13097 394806 -13041
rect 394862 -13097 394930 -13041
rect 394986 -13097 395054 -13041
rect 395110 -13097 395178 -13041
rect 395234 -13097 395302 -13041
rect 395358 -13097 395426 -13041
rect 395482 -13097 395550 -13041
rect 395606 -13097 395674 -13041
rect 395730 -13097 395798 -13041
rect 395854 -13097 395922 -13041
rect 395978 -13097 396046 -13041
rect 396102 -13097 396170 -13041
rect 396226 -13097 396294 -13041
rect 396350 -13097 396418 -13041
rect 396474 -13097 396542 -13041
rect 396598 -13097 396666 -13041
rect 396722 -13097 396790 -13041
rect 396846 -13097 396914 -13041
rect 396970 -13097 397038 -13041
rect 397094 -13097 397162 -13041
rect 397218 -13097 397286 -13041
rect 397342 -13097 397410 -13041
rect 397466 -13097 397534 -13041
rect 397590 -13097 397658 -13041
rect 397714 -13097 397782 -13041
rect 397838 -13097 397906 -13041
rect 397962 -13097 398030 -13041
rect 398086 -13097 398154 -13041
rect 398210 -13097 398278 -13041
rect 398334 -13097 398402 -13041
rect 398458 -13097 398526 -13041
rect 398582 -13097 398650 -13041
rect 398706 -13097 398774 -13041
rect 398830 -13097 398898 -13041
rect 398954 -13097 399022 -13041
rect 399078 -13097 399146 -13041
rect 399202 -13097 399270 -13041
rect 399326 -13097 399394 -13041
rect 399450 -13097 399518 -13041
rect 399574 -13097 399642 -13041
rect 399698 -13097 399766 -13041
rect 399822 -13097 399890 -13041
rect 399946 -13097 400014 -13041
rect 400070 -13097 400138 -13041
rect 400194 -13097 400262 -13041
rect 400318 -13097 400386 -13041
rect 400442 -13097 400510 -13041
rect 400566 -13097 400634 -13041
rect 400690 -13097 400758 -13041
rect 400814 -13097 400882 -13041
rect 400938 -13097 401006 -13041
rect 401062 -13097 401130 -13041
rect 401186 -13097 401254 -13041
rect 401310 -13097 401440 -13041
rect 387840 -13165 401440 -13097
rect 387840 -13221 387986 -13165
rect 388042 -13221 388110 -13165
rect 388166 -13221 388234 -13165
rect 388290 -13221 388358 -13165
rect 388414 -13221 388482 -13165
rect 388538 -13221 388606 -13165
rect 388662 -13221 388730 -13165
rect 388786 -13221 388854 -13165
rect 388910 -13221 388978 -13165
rect 389034 -13221 389102 -13165
rect 389158 -13221 389226 -13165
rect 389282 -13221 389350 -13165
rect 389406 -13221 389474 -13165
rect 389530 -13221 389598 -13165
rect 389654 -13221 389722 -13165
rect 389778 -13221 389846 -13165
rect 389902 -13221 389970 -13165
rect 390026 -13221 390094 -13165
rect 390150 -13221 390218 -13165
rect 390274 -13221 390342 -13165
rect 390398 -13221 390466 -13165
rect 390522 -13221 390590 -13165
rect 390646 -13221 390714 -13165
rect 390770 -13221 390838 -13165
rect 390894 -13221 390962 -13165
rect 391018 -13221 391086 -13165
rect 391142 -13221 391210 -13165
rect 391266 -13221 391334 -13165
rect 391390 -13221 391458 -13165
rect 391514 -13221 391582 -13165
rect 391638 -13221 391706 -13165
rect 391762 -13221 391830 -13165
rect 391886 -13221 391954 -13165
rect 392010 -13221 392078 -13165
rect 392134 -13221 392202 -13165
rect 392258 -13221 392326 -13165
rect 392382 -13221 392450 -13165
rect 392506 -13221 392574 -13165
rect 392630 -13221 392698 -13165
rect 392754 -13221 392822 -13165
rect 392878 -13221 392946 -13165
rect 393002 -13221 393070 -13165
rect 393126 -13221 393194 -13165
rect 393250 -13221 393318 -13165
rect 393374 -13221 393442 -13165
rect 393498 -13221 393566 -13165
rect 393622 -13221 393690 -13165
rect 393746 -13221 393814 -13165
rect 393870 -13221 393938 -13165
rect 393994 -13221 394062 -13165
rect 394118 -13221 394186 -13165
rect 394242 -13221 394310 -13165
rect 394366 -13221 394434 -13165
rect 394490 -13221 394558 -13165
rect 394614 -13221 394682 -13165
rect 394738 -13221 394806 -13165
rect 394862 -13221 394930 -13165
rect 394986 -13221 395054 -13165
rect 395110 -13221 395178 -13165
rect 395234 -13221 395302 -13165
rect 395358 -13221 395426 -13165
rect 395482 -13221 395550 -13165
rect 395606 -13221 395674 -13165
rect 395730 -13221 395798 -13165
rect 395854 -13221 395922 -13165
rect 395978 -13221 396046 -13165
rect 396102 -13221 396170 -13165
rect 396226 -13221 396294 -13165
rect 396350 -13221 396418 -13165
rect 396474 -13221 396542 -13165
rect 396598 -13221 396666 -13165
rect 396722 -13221 396790 -13165
rect 396846 -13221 396914 -13165
rect 396970 -13221 397038 -13165
rect 397094 -13221 397162 -13165
rect 397218 -13221 397286 -13165
rect 397342 -13221 397410 -13165
rect 397466 -13221 397534 -13165
rect 397590 -13221 397658 -13165
rect 397714 -13221 397782 -13165
rect 397838 -13221 397906 -13165
rect 397962 -13221 398030 -13165
rect 398086 -13221 398154 -13165
rect 398210 -13221 398278 -13165
rect 398334 -13221 398402 -13165
rect 398458 -13221 398526 -13165
rect 398582 -13221 398650 -13165
rect 398706 -13221 398774 -13165
rect 398830 -13221 398898 -13165
rect 398954 -13221 399022 -13165
rect 399078 -13221 399146 -13165
rect 399202 -13221 399270 -13165
rect 399326 -13221 399394 -13165
rect 399450 -13221 399518 -13165
rect 399574 -13221 399642 -13165
rect 399698 -13221 399766 -13165
rect 399822 -13221 399890 -13165
rect 399946 -13221 400014 -13165
rect 400070 -13221 400138 -13165
rect 400194 -13221 400262 -13165
rect 400318 -13221 400386 -13165
rect 400442 -13221 400510 -13165
rect 400566 -13221 400634 -13165
rect 400690 -13221 400758 -13165
rect 400814 -13221 400882 -13165
rect 400938 -13221 401006 -13165
rect 401062 -13221 401130 -13165
rect 401186 -13221 401254 -13165
rect 401310 -13221 401440 -13165
rect 387840 -13289 401440 -13221
rect 387840 -13345 387986 -13289
rect 388042 -13345 388110 -13289
rect 388166 -13345 388234 -13289
rect 388290 -13345 388358 -13289
rect 388414 -13345 388482 -13289
rect 388538 -13345 388606 -13289
rect 388662 -13345 388730 -13289
rect 388786 -13345 388854 -13289
rect 388910 -13345 388978 -13289
rect 389034 -13345 389102 -13289
rect 389158 -13345 389226 -13289
rect 389282 -13345 389350 -13289
rect 389406 -13345 389474 -13289
rect 389530 -13345 389598 -13289
rect 389654 -13345 389722 -13289
rect 389778 -13345 389846 -13289
rect 389902 -13345 389970 -13289
rect 390026 -13345 390094 -13289
rect 390150 -13345 390218 -13289
rect 390274 -13345 390342 -13289
rect 390398 -13345 390466 -13289
rect 390522 -13345 390590 -13289
rect 390646 -13345 390714 -13289
rect 390770 -13345 390838 -13289
rect 390894 -13345 390962 -13289
rect 391018 -13345 391086 -13289
rect 391142 -13345 391210 -13289
rect 391266 -13345 391334 -13289
rect 391390 -13345 391458 -13289
rect 391514 -13345 391582 -13289
rect 391638 -13345 391706 -13289
rect 391762 -13345 391830 -13289
rect 391886 -13345 391954 -13289
rect 392010 -13345 392078 -13289
rect 392134 -13345 392202 -13289
rect 392258 -13345 392326 -13289
rect 392382 -13345 392450 -13289
rect 392506 -13345 392574 -13289
rect 392630 -13345 392698 -13289
rect 392754 -13345 392822 -13289
rect 392878 -13345 392946 -13289
rect 393002 -13345 393070 -13289
rect 393126 -13345 393194 -13289
rect 393250 -13345 393318 -13289
rect 393374 -13345 393442 -13289
rect 393498 -13345 393566 -13289
rect 393622 -13345 393690 -13289
rect 393746 -13345 393814 -13289
rect 393870 -13345 393938 -13289
rect 393994 -13345 394062 -13289
rect 394118 -13345 394186 -13289
rect 394242 -13345 394310 -13289
rect 394366 -13345 394434 -13289
rect 394490 -13345 394558 -13289
rect 394614 -13345 394682 -13289
rect 394738 -13345 394806 -13289
rect 394862 -13345 394930 -13289
rect 394986 -13345 395054 -13289
rect 395110 -13345 395178 -13289
rect 395234 -13345 395302 -13289
rect 395358 -13345 395426 -13289
rect 395482 -13345 395550 -13289
rect 395606 -13345 395674 -13289
rect 395730 -13345 395798 -13289
rect 395854 -13345 395922 -13289
rect 395978 -13345 396046 -13289
rect 396102 -13345 396170 -13289
rect 396226 -13345 396294 -13289
rect 396350 -13345 396418 -13289
rect 396474 -13345 396542 -13289
rect 396598 -13345 396666 -13289
rect 396722 -13345 396790 -13289
rect 396846 -13345 396914 -13289
rect 396970 -13345 397038 -13289
rect 397094 -13345 397162 -13289
rect 397218 -13345 397286 -13289
rect 397342 -13345 397410 -13289
rect 397466 -13345 397534 -13289
rect 397590 -13345 397658 -13289
rect 397714 -13345 397782 -13289
rect 397838 -13345 397906 -13289
rect 397962 -13345 398030 -13289
rect 398086 -13345 398154 -13289
rect 398210 -13345 398278 -13289
rect 398334 -13345 398402 -13289
rect 398458 -13345 398526 -13289
rect 398582 -13345 398650 -13289
rect 398706 -13345 398774 -13289
rect 398830 -13345 398898 -13289
rect 398954 -13345 399022 -13289
rect 399078 -13345 399146 -13289
rect 399202 -13345 399270 -13289
rect 399326 -13345 399394 -13289
rect 399450 -13345 399518 -13289
rect 399574 -13345 399642 -13289
rect 399698 -13345 399766 -13289
rect 399822 -13345 399890 -13289
rect 399946 -13345 400014 -13289
rect 400070 -13345 400138 -13289
rect 400194 -13345 400262 -13289
rect 400318 -13345 400386 -13289
rect 400442 -13345 400510 -13289
rect 400566 -13345 400634 -13289
rect 400690 -13345 400758 -13289
rect 400814 -13345 400882 -13289
rect 400938 -13345 401006 -13289
rect 401062 -13345 401130 -13289
rect 401186 -13345 401254 -13289
rect 401310 -13345 401440 -13289
rect 387840 -13413 401440 -13345
rect 387840 -13469 387986 -13413
rect 388042 -13469 388110 -13413
rect 388166 -13469 388234 -13413
rect 388290 -13469 388358 -13413
rect 388414 -13469 388482 -13413
rect 388538 -13469 388606 -13413
rect 388662 -13469 388730 -13413
rect 388786 -13469 388854 -13413
rect 388910 -13469 388978 -13413
rect 389034 -13469 389102 -13413
rect 389158 -13469 389226 -13413
rect 389282 -13469 389350 -13413
rect 389406 -13469 389474 -13413
rect 389530 -13469 389598 -13413
rect 389654 -13469 389722 -13413
rect 389778 -13469 389846 -13413
rect 389902 -13469 389970 -13413
rect 390026 -13469 390094 -13413
rect 390150 -13469 390218 -13413
rect 390274 -13469 390342 -13413
rect 390398 -13469 390466 -13413
rect 390522 -13469 390590 -13413
rect 390646 -13469 390714 -13413
rect 390770 -13469 390838 -13413
rect 390894 -13469 390962 -13413
rect 391018 -13469 391086 -13413
rect 391142 -13469 391210 -13413
rect 391266 -13469 391334 -13413
rect 391390 -13469 391458 -13413
rect 391514 -13469 391582 -13413
rect 391638 -13469 391706 -13413
rect 391762 -13469 391830 -13413
rect 391886 -13469 391954 -13413
rect 392010 -13469 392078 -13413
rect 392134 -13469 392202 -13413
rect 392258 -13469 392326 -13413
rect 392382 -13469 392450 -13413
rect 392506 -13469 392574 -13413
rect 392630 -13469 392698 -13413
rect 392754 -13469 392822 -13413
rect 392878 -13469 392946 -13413
rect 393002 -13469 393070 -13413
rect 393126 -13469 393194 -13413
rect 393250 -13469 393318 -13413
rect 393374 -13469 393442 -13413
rect 393498 -13469 393566 -13413
rect 393622 -13469 393690 -13413
rect 393746 -13469 393814 -13413
rect 393870 -13469 393938 -13413
rect 393994 -13469 394062 -13413
rect 394118 -13469 394186 -13413
rect 394242 -13469 394310 -13413
rect 394366 -13469 394434 -13413
rect 394490 -13469 394558 -13413
rect 394614 -13469 394682 -13413
rect 394738 -13469 394806 -13413
rect 394862 -13469 394930 -13413
rect 394986 -13469 395054 -13413
rect 395110 -13469 395178 -13413
rect 395234 -13469 395302 -13413
rect 395358 -13469 395426 -13413
rect 395482 -13469 395550 -13413
rect 395606 -13469 395674 -13413
rect 395730 -13469 395798 -13413
rect 395854 -13469 395922 -13413
rect 395978 -13469 396046 -13413
rect 396102 -13469 396170 -13413
rect 396226 -13469 396294 -13413
rect 396350 -13469 396418 -13413
rect 396474 -13469 396542 -13413
rect 396598 -13469 396666 -13413
rect 396722 -13469 396790 -13413
rect 396846 -13469 396914 -13413
rect 396970 -13469 397038 -13413
rect 397094 -13469 397162 -13413
rect 397218 -13469 397286 -13413
rect 397342 -13469 397410 -13413
rect 397466 -13469 397534 -13413
rect 397590 -13469 397658 -13413
rect 397714 -13469 397782 -13413
rect 397838 -13469 397906 -13413
rect 397962 -13469 398030 -13413
rect 398086 -13469 398154 -13413
rect 398210 -13469 398278 -13413
rect 398334 -13469 398402 -13413
rect 398458 -13469 398526 -13413
rect 398582 -13469 398650 -13413
rect 398706 -13469 398774 -13413
rect 398830 -13469 398898 -13413
rect 398954 -13469 399022 -13413
rect 399078 -13469 399146 -13413
rect 399202 -13469 399270 -13413
rect 399326 -13469 399394 -13413
rect 399450 -13469 399518 -13413
rect 399574 -13469 399642 -13413
rect 399698 -13469 399766 -13413
rect 399822 -13469 399890 -13413
rect 399946 -13469 400014 -13413
rect 400070 -13469 400138 -13413
rect 400194 -13469 400262 -13413
rect 400318 -13469 400386 -13413
rect 400442 -13469 400510 -13413
rect 400566 -13469 400634 -13413
rect 400690 -13469 400758 -13413
rect 400814 -13469 400882 -13413
rect 400938 -13469 401006 -13413
rect 401062 -13469 401130 -13413
rect 401186 -13469 401254 -13413
rect 401310 -13469 401440 -13413
rect 387840 -13632 401440 -13469
rect 387840 -13688 387954 -13632
rect 388010 -13688 388078 -13632
rect 388134 -13688 388202 -13632
rect 388258 -13688 388326 -13632
rect 388382 -13688 388450 -13632
rect 388506 -13670 400766 -13632
rect 388506 -13688 388640 -13670
rect 387840 -13756 388640 -13688
rect 387840 -13812 387954 -13756
rect 388010 -13812 388078 -13756
rect 388134 -13812 388202 -13756
rect 388258 -13812 388326 -13756
rect 388382 -13812 388450 -13756
rect 388506 -13812 388640 -13756
rect 387840 -13880 388640 -13812
rect 387840 -13936 387954 -13880
rect 388010 -13936 388078 -13880
rect 388134 -13936 388202 -13880
rect 388258 -13936 388326 -13880
rect 388382 -13936 388450 -13880
rect 388506 -13936 388640 -13880
rect 387840 -14004 388640 -13936
rect 387840 -14060 387954 -14004
rect 388010 -14060 388078 -14004
rect 388134 -14060 388202 -14004
rect 388258 -14060 388326 -14004
rect 388382 -14060 388450 -14004
rect 388506 -14060 388640 -14004
rect 387840 -14128 388640 -14060
rect 387840 -14184 387954 -14128
rect 388010 -14184 388078 -14128
rect 388134 -14184 388202 -14128
rect 388258 -14184 388326 -14128
rect 388382 -14184 388450 -14128
rect 388506 -14184 388640 -14128
rect 387840 -14252 388640 -14184
rect 387840 -14308 387954 -14252
rect 388010 -14308 388078 -14252
rect 388134 -14308 388202 -14252
rect 388258 -14308 388326 -14252
rect 388382 -14308 388450 -14252
rect 388506 -14308 388640 -14252
rect 387840 -14376 388640 -14308
rect 387840 -14432 387954 -14376
rect 388010 -14432 388078 -14376
rect 388134 -14432 388202 -14376
rect 388258 -14432 388326 -14376
rect 388382 -14432 388450 -14376
rect 388506 -14432 388640 -14376
rect 387840 -14500 388640 -14432
rect 387840 -14556 387954 -14500
rect 388010 -14556 388078 -14500
rect 388134 -14556 388202 -14500
rect 388258 -14556 388326 -14500
rect 388382 -14556 388450 -14500
rect 388506 -14556 388640 -14500
rect 387840 -14624 388640 -14556
rect 387840 -14680 387954 -14624
rect 388010 -14680 388078 -14624
rect 388134 -14680 388202 -14624
rect 388258 -14680 388326 -14624
rect 388382 -14680 388450 -14624
rect 388506 -14680 388640 -14624
rect 387840 -14748 388640 -14680
rect 387840 -14804 387954 -14748
rect 388010 -14804 388078 -14748
rect 388134 -14804 388202 -14748
rect 388258 -14804 388326 -14748
rect 388382 -14804 388450 -14748
rect 388506 -14804 388640 -14748
rect 387840 -14872 388640 -14804
rect 387840 -14928 387954 -14872
rect 388010 -14928 388078 -14872
rect 388134 -14928 388202 -14872
rect 388258 -14928 388326 -14872
rect 388382 -14928 388450 -14872
rect 388506 -14928 388640 -14872
rect 387840 -14996 388640 -14928
rect 387840 -15052 387954 -14996
rect 388010 -15052 388078 -14996
rect 388134 -15052 388202 -14996
rect 388258 -15052 388326 -14996
rect 388382 -15052 388450 -14996
rect 388506 -15052 388640 -14996
rect 387840 -15120 388640 -15052
rect 387840 -15176 387954 -15120
rect 388010 -15176 388078 -15120
rect 388134 -15176 388202 -15120
rect 388258 -15176 388326 -15120
rect 388382 -15176 388450 -15120
rect 388506 -15176 388640 -15120
rect 387840 -15244 388640 -15176
rect 387840 -15300 387954 -15244
rect 388010 -15300 388078 -15244
rect 388134 -15300 388202 -15244
rect 388258 -15300 388326 -15244
rect 388382 -15300 388450 -15244
rect 388506 -15300 388640 -15244
rect 387840 -15368 388640 -15300
rect 387840 -15424 387954 -15368
rect 388010 -15424 388078 -15368
rect 388134 -15424 388202 -15368
rect 388258 -15424 388326 -15368
rect 388382 -15424 388450 -15368
rect 388506 -15424 388640 -15368
rect 387840 -15492 388640 -15424
rect 387840 -15548 387954 -15492
rect 388010 -15548 388078 -15492
rect 388134 -15548 388202 -15492
rect 388258 -15548 388326 -15492
rect 388382 -15548 388450 -15492
rect 388506 -15548 388640 -15492
rect 387840 -15616 388640 -15548
rect 387840 -15672 387954 -15616
rect 388010 -15672 388078 -15616
rect 388134 -15672 388202 -15616
rect 388258 -15672 388326 -15616
rect 388382 -15672 388450 -15616
rect 388506 -15672 388640 -15616
rect 387840 -15740 388640 -15672
rect 387840 -15796 387954 -15740
rect 388010 -15796 388078 -15740
rect 388134 -15796 388202 -15740
rect 388258 -15796 388326 -15740
rect 388382 -15796 388450 -15740
rect 388506 -15796 388640 -15740
rect 387840 -15864 388640 -15796
rect 387840 -15920 387954 -15864
rect 388010 -15920 388078 -15864
rect 388134 -15920 388202 -15864
rect 388258 -15920 388326 -15864
rect 388382 -15920 388450 -15864
rect 388506 -15920 388640 -15864
rect 387840 -15988 388640 -15920
rect 387840 -16044 387954 -15988
rect 388010 -16044 388078 -15988
rect 388134 -16044 388202 -15988
rect 388258 -16044 388326 -15988
rect 388382 -16044 388450 -15988
rect 388506 -16044 388640 -15988
rect 387840 -16112 388640 -16044
rect 387840 -16168 387954 -16112
rect 388010 -16168 388078 -16112
rect 388134 -16168 388202 -16112
rect 388258 -16168 388326 -16112
rect 388382 -16168 388450 -16112
rect 388506 -16168 388640 -16112
rect 387840 -16236 388640 -16168
rect 387840 -16292 387954 -16236
rect 388010 -16292 388078 -16236
rect 388134 -16292 388202 -16236
rect 388258 -16292 388326 -16236
rect 388382 -16292 388450 -16236
rect 388506 -16292 388640 -16236
rect 387840 -16360 388640 -16292
rect 387840 -16416 387954 -16360
rect 388010 -16416 388078 -16360
rect 388134 -16416 388202 -16360
rect 388258 -16416 388326 -16360
rect 388382 -16416 388450 -16360
rect 388506 -16416 388640 -16360
rect 387840 -16484 388640 -16416
rect 387840 -16540 387954 -16484
rect 388010 -16540 388078 -16484
rect 388134 -16540 388202 -16484
rect 388258 -16540 388326 -16484
rect 388382 -16540 388450 -16484
rect 388506 -16540 388640 -16484
rect 387840 -16608 388640 -16540
rect 387840 -16664 387954 -16608
rect 388010 -16664 388078 -16608
rect 388134 -16664 388202 -16608
rect 388258 -16664 388326 -16608
rect 388382 -16664 388450 -16608
rect 388506 -16664 388640 -16608
rect 387840 -16732 388640 -16664
rect 387840 -16788 387954 -16732
rect 388010 -16788 388078 -16732
rect 388134 -16788 388202 -16732
rect 388258 -16788 388326 -16732
rect 388382 -16788 388450 -16732
rect 388506 -16788 388640 -16732
rect 387840 -16856 388640 -16788
rect 387840 -16912 387954 -16856
rect 388010 -16912 388078 -16856
rect 388134 -16912 388202 -16856
rect 388258 -16912 388326 -16856
rect 388382 -16912 388450 -16856
rect 388506 -16912 388640 -16856
rect 387840 -16980 388640 -16912
rect 387840 -17036 387954 -16980
rect 388010 -17036 388078 -16980
rect 388134 -17036 388202 -16980
rect 388258 -17036 388326 -16980
rect 388382 -17036 388450 -16980
rect 388506 -17036 388640 -16980
rect 387840 -17104 388640 -17036
rect 387840 -17160 387954 -17104
rect 388010 -17160 388078 -17104
rect 388134 -17160 388202 -17104
rect 388258 -17160 388326 -17104
rect 388382 -17160 388450 -17104
rect 388506 -17160 388640 -17104
rect 387840 -17228 388640 -17160
rect 387840 -17284 387954 -17228
rect 388010 -17284 388078 -17228
rect 388134 -17284 388202 -17228
rect 388258 -17284 388326 -17228
rect 388382 -17284 388450 -17228
rect 388506 -17284 388640 -17228
rect 387840 -17352 388640 -17284
rect 387840 -17408 387954 -17352
rect 388010 -17408 388078 -17352
rect 388134 -17408 388202 -17352
rect 388258 -17408 388326 -17352
rect 388382 -17408 388450 -17352
rect 388506 -17408 388640 -17352
rect 387840 -17476 388640 -17408
rect 387840 -17532 387954 -17476
rect 388010 -17532 388078 -17476
rect 388134 -17532 388202 -17476
rect 388258 -17532 388326 -17476
rect 388382 -17532 388450 -17476
rect 388506 -17532 388640 -17476
rect 387840 -17600 388640 -17532
rect 387840 -17656 387954 -17600
rect 388010 -17656 388078 -17600
rect 388134 -17656 388202 -17600
rect 388258 -17656 388326 -17600
rect 388382 -17656 388450 -17600
rect 388506 -17656 388640 -17600
rect 387840 -17724 388640 -17656
rect 387840 -17780 387954 -17724
rect 388010 -17780 388078 -17724
rect 388134 -17780 388202 -17724
rect 388258 -17780 388326 -17724
rect 388382 -17780 388450 -17724
rect 388506 -17780 388640 -17724
rect 387840 -17848 388640 -17780
rect 387840 -17904 387954 -17848
rect 388010 -17904 388078 -17848
rect 388134 -17904 388202 -17848
rect 388258 -17904 388326 -17848
rect 388382 -17904 388450 -17848
rect 388506 -17904 388640 -17848
rect 387840 -17972 388640 -17904
rect 387840 -18028 387954 -17972
rect 388010 -18028 388078 -17972
rect 388134 -18028 388202 -17972
rect 388258 -18028 388326 -17972
rect 388382 -18028 388450 -17972
rect 388506 -18028 388640 -17972
rect 387840 -18096 388640 -18028
rect 387840 -18152 387954 -18096
rect 388010 -18152 388078 -18096
rect 388134 -18152 388202 -18096
rect 388258 -18152 388326 -18096
rect 388382 -18152 388450 -18096
rect 388506 -18152 388640 -18096
rect 387840 -18220 388640 -18152
rect 387840 -18276 387954 -18220
rect 388010 -18276 388078 -18220
rect 388134 -18276 388202 -18220
rect 388258 -18276 388326 -18220
rect 388382 -18276 388450 -18220
rect 388506 -18276 388640 -18220
rect 387840 -18344 388640 -18276
rect 387840 -18400 387954 -18344
rect 388010 -18400 388078 -18344
rect 388134 -18400 388202 -18344
rect 388258 -18400 388326 -18344
rect 388382 -18400 388450 -18344
rect 388506 -18400 388640 -18344
rect 387840 -18468 388640 -18400
rect 387840 -18524 387954 -18468
rect 388010 -18524 388078 -18468
rect 388134 -18524 388202 -18468
rect 388258 -18524 388326 -18468
rect 388382 -18524 388450 -18468
rect 388506 -18524 388640 -18468
rect 387840 -18592 388640 -18524
rect 387840 -18648 387954 -18592
rect 388010 -18648 388078 -18592
rect 388134 -18648 388202 -18592
rect 388258 -18648 388326 -18592
rect 388382 -18648 388450 -18592
rect 388506 -18648 388640 -18592
rect 387840 -18716 388640 -18648
rect 387840 -18772 387954 -18716
rect 388010 -18772 388078 -18716
rect 388134 -18772 388202 -18716
rect 388258 -18772 388326 -18716
rect 388382 -18772 388450 -18716
rect 388506 -18772 388640 -18716
rect 387840 -18840 388640 -18772
rect 387840 -18896 387954 -18840
rect 388010 -18896 388078 -18840
rect 388134 -18896 388202 -18840
rect 388258 -18896 388326 -18840
rect 388382 -18896 388450 -18840
rect 388506 -18896 388640 -18840
rect 387840 -18964 388640 -18896
rect 387840 -19020 387954 -18964
rect 388010 -19020 388078 -18964
rect 388134 -19020 388202 -18964
rect 388258 -19020 388326 -18964
rect 388382 -19020 388450 -18964
rect 388506 -19020 388640 -18964
rect 387840 -19088 388640 -19020
rect 387840 -19144 387954 -19088
rect 388010 -19144 388078 -19088
rect 388134 -19144 388202 -19088
rect 388258 -19144 388326 -19088
rect 388382 -19144 388450 -19088
rect 388506 -19144 388640 -19088
rect 387840 -19212 388640 -19144
rect 387840 -19268 387954 -19212
rect 388010 -19268 388078 -19212
rect 388134 -19268 388202 -19212
rect 388258 -19268 388326 -19212
rect 388382 -19268 388450 -19212
rect 388506 -19268 388640 -19212
rect 387840 -19336 388640 -19268
rect 387840 -19392 387954 -19336
rect 388010 -19392 388078 -19336
rect 388134 -19392 388202 -19336
rect 388258 -19392 388326 -19336
rect 388382 -19392 388450 -19336
rect 388506 -19392 388640 -19336
rect 387840 -19460 388640 -19392
rect 387840 -19516 387954 -19460
rect 388010 -19516 388078 -19460
rect 388134 -19516 388202 -19460
rect 388258 -19516 388326 -19460
rect 388382 -19516 388450 -19460
rect 388506 -19516 388640 -19460
rect 387840 -19584 388640 -19516
rect 387840 -19640 387954 -19584
rect 388010 -19640 388078 -19584
rect 388134 -19640 388202 -19584
rect 388258 -19640 388326 -19584
rect 388382 -19640 388450 -19584
rect 388506 -19640 388640 -19584
rect 387840 -19708 388640 -19640
rect 387840 -19764 387954 -19708
rect 388010 -19764 388078 -19708
rect 388134 -19764 388202 -19708
rect 388258 -19764 388326 -19708
rect 388382 -19764 388450 -19708
rect 388506 -19764 388640 -19708
rect 387840 -19832 388640 -19764
rect 387840 -19888 387954 -19832
rect 388010 -19888 388078 -19832
rect 388134 -19888 388202 -19832
rect 388258 -19888 388326 -19832
rect 388382 -19888 388450 -19832
rect 388506 -19888 388640 -19832
rect 387840 -19956 388640 -19888
rect 387840 -20012 387954 -19956
rect 388010 -20012 388078 -19956
rect 388134 -20012 388202 -19956
rect 388258 -20012 388326 -19956
rect 388382 -20012 388450 -19956
rect 388506 -20012 388640 -19956
rect 387840 -20080 388640 -20012
rect 387840 -20136 387954 -20080
rect 388010 -20136 388078 -20080
rect 388134 -20136 388202 -20080
rect 388258 -20136 388326 -20080
rect 388382 -20136 388450 -20080
rect 388506 -20136 388640 -20080
rect 387840 -20204 388640 -20136
rect 387840 -20260 387954 -20204
rect 388010 -20260 388078 -20204
rect 388134 -20260 388202 -20204
rect 388258 -20260 388326 -20204
rect 388382 -20260 388450 -20204
rect 388506 -20260 388640 -20204
rect 387840 -20328 388640 -20260
rect 387840 -20384 387954 -20328
rect 388010 -20384 388078 -20328
rect 388134 -20384 388202 -20328
rect 388258 -20384 388326 -20328
rect 388382 -20384 388450 -20328
rect 388506 -20384 388640 -20328
rect 387840 -20452 388640 -20384
rect 387840 -20508 387954 -20452
rect 388010 -20508 388078 -20452
rect 388134 -20508 388202 -20452
rect 388258 -20508 388326 -20452
rect 388382 -20508 388450 -20452
rect 388506 -20508 388640 -20452
rect 387840 -20576 388640 -20508
rect 387840 -20632 387954 -20576
rect 388010 -20632 388078 -20576
rect 388134 -20632 388202 -20576
rect 388258 -20632 388326 -20576
rect 388382 -20632 388450 -20576
rect 388506 -20632 388640 -20576
rect 387840 -20700 388640 -20632
rect 387840 -20756 387954 -20700
rect 388010 -20756 388078 -20700
rect 388134 -20756 388202 -20700
rect 388258 -20756 388326 -20700
rect 388382 -20756 388450 -20700
rect 388506 -20756 388640 -20700
rect 387840 -20824 388640 -20756
rect 387840 -20880 387954 -20824
rect 388010 -20880 388078 -20824
rect 388134 -20880 388202 -20824
rect 388258 -20880 388326 -20824
rect 388382 -20880 388450 -20824
rect 388506 -20880 388640 -20824
rect 387840 -20948 388640 -20880
rect 387840 -21004 387954 -20948
rect 388010 -21004 388078 -20948
rect 388134 -21004 388202 -20948
rect 388258 -21004 388326 -20948
rect 388382 -21004 388450 -20948
rect 388506 -21004 388640 -20948
rect 387840 -21072 388640 -21004
rect 387840 -21128 387954 -21072
rect 388010 -21128 388078 -21072
rect 388134 -21128 388202 -21072
rect 388258 -21128 388326 -21072
rect 388382 -21128 388450 -21072
rect 388506 -21128 388640 -21072
rect 387840 -21196 388640 -21128
rect 387840 -21252 387954 -21196
rect 388010 -21252 388078 -21196
rect 388134 -21252 388202 -21196
rect 388258 -21252 388326 -21196
rect 388382 -21252 388450 -21196
rect 388506 -21252 388640 -21196
rect 387840 -21320 388640 -21252
rect 387840 -21376 387954 -21320
rect 388010 -21376 388078 -21320
rect 388134 -21376 388202 -21320
rect 388258 -21376 388326 -21320
rect 388382 -21376 388450 -21320
rect 388506 -21376 388640 -21320
rect 387840 -21444 388640 -21376
rect 387840 -21500 387954 -21444
rect 388010 -21500 388078 -21444
rect 388134 -21500 388202 -21444
rect 388258 -21500 388326 -21444
rect 388382 -21500 388450 -21444
rect 388506 -21500 388640 -21444
rect 387840 -21568 388640 -21500
rect 387840 -21624 387954 -21568
rect 388010 -21624 388078 -21568
rect 388134 -21624 388202 -21568
rect 388258 -21624 388326 -21568
rect 388382 -21624 388450 -21568
rect 388506 -21624 388640 -21568
rect 387840 -21692 388640 -21624
rect 387840 -21748 387954 -21692
rect 388010 -21748 388078 -21692
rect 388134 -21748 388202 -21692
rect 388258 -21748 388326 -21692
rect 388382 -21748 388450 -21692
rect 388506 -21748 388640 -21692
rect 387840 -21816 388640 -21748
rect 387840 -21872 387954 -21816
rect 388010 -21872 388078 -21816
rect 388134 -21872 388202 -21816
rect 388258 -21872 388326 -21816
rect 388382 -21872 388450 -21816
rect 388506 -21872 388640 -21816
rect 387840 -21940 388640 -21872
rect 387840 -21996 387954 -21940
rect 388010 -21996 388078 -21940
rect 388134 -21996 388202 -21940
rect 388258 -21996 388326 -21940
rect 388382 -21996 388450 -21940
rect 388506 -21996 388640 -21940
rect 387840 -22064 388640 -21996
rect 387840 -22120 387954 -22064
rect 388010 -22120 388078 -22064
rect 388134 -22120 388202 -22064
rect 388258 -22120 388326 -22064
rect 388382 -22120 388450 -22064
rect 388506 -22120 388640 -22064
rect 387840 -22188 388640 -22120
rect 387840 -22244 387954 -22188
rect 388010 -22244 388078 -22188
rect 388134 -22244 388202 -22188
rect 388258 -22244 388326 -22188
rect 388382 -22244 388450 -22188
rect 388506 -22244 388640 -22188
rect 387840 -22312 388640 -22244
rect 387840 -22368 387954 -22312
rect 388010 -22368 388078 -22312
rect 388134 -22368 388202 -22312
rect 388258 -22368 388326 -22312
rect 388382 -22368 388450 -22312
rect 388506 -22368 388640 -22312
rect 387840 -22436 388640 -22368
rect 387840 -22492 387954 -22436
rect 388010 -22492 388078 -22436
rect 388134 -22492 388202 -22436
rect 388258 -22492 388326 -22436
rect 388382 -22492 388450 -22436
rect 388506 -22492 388640 -22436
rect 387840 -22560 388640 -22492
rect 387840 -22616 387954 -22560
rect 388010 -22616 388078 -22560
rect 388134 -22616 388202 -22560
rect 388258 -22616 388326 -22560
rect 388382 -22616 388450 -22560
rect 388506 -22616 388640 -22560
rect 387840 -22684 388640 -22616
rect 387840 -22740 387954 -22684
rect 388010 -22740 388078 -22684
rect 388134 -22740 388202 -22684
rect 388258 -22740 388326 -22684
rect 388382 -22740 388450 -22684
rect 388506 -22740 388640 -22684
rect 387840 -22808 388640 -22740
rect 387840 -22864 387954 -22808
rect 388010 -22864 388078 -22808
rect 388134 -22864 388202 -22808
rect 388258 -22864 388326 -22808
rect 388382 -22864 388450 -22808
rect 388506 -22864 388640 -22808
rect 387840 -22932 388640 -22864
rect 387840 -22988 387954 -22932
rect 388010 -22988 388078 -22932
rect 388134 -22988 388202 -22932
rect 388258 -22988 388326 -22932
rect 388382 -22988 388450 -22932
rect 388506 -22988 388640 -22932
rect 387840 -23056 388640 -22988
rect 387840 -23112 387954 -23056
rect 388010 -23112 388078 -23056
rect 388134 -23112 388202 -23056
rect 388258 -23112 388326 -23056
rect 388382 -23112 388450 -23056
rect 388506 -23112 388640 -23056
rect 387840 -23180 388640 -23112
rect 387840 -23236 387954 -23180
rect 388010 -23236 388078 -23180
rect 388134 -23236 388202 -23180
rect 388258 -23236 388326 -23180
rect 388382 -23236 388450 -23180
rect 388506 -23236 388640 -23180
rect 387840 -23304 388640 -23236
rect 387840 -23360 387954 -23304
rect 388010 -23360 388078 -23304
rect 388134 -23360 388202 -23304
rect 388258 -23360 388326 -23304
rect 388382 -23360 388450 -23304
rect 388506 -23360 388640 -23304
rect 387840 -23428 388640 -23360
rect 387840 -23484 387954 -23428
rect 388010 -23484 388078 -23428
rect 388134 -23484 388202 -23428
rect 388258 -23484 388326 -23428
rect 388382 -23484 388450 -23428
rect 388506 -23484 388640 -23428
rect 387840 -23552 388640 -23484
rect 387840 -23608 387954 -23552
rect 388010 -23608 388078 -23552
rect 388134 -23608 388202 -23552
rect 388258 -23608 388326 -23552
rect 388382 -23608 388450 -23552
rect 388506 -23608 388640 -23552
rect 387840 -23676 388640 -23608
rect 387840 -23732 387954 -23676
rect 388010 -23732 388078 -23676
rect 388134 -23732 388202 -23676
rect 388258 -23732 388326 -23676
rect 388382 -23732 388450 -23676
rect 388506 -23732 388640 -23676
rect 387840 -23800 388640 -23732
rect 387840 -23856 387954 -23800
rect 388010 -23856 388078 -23800
rect 388134 -23856 388202 -23800
rect 388258 -23856 388326 -23800
rect 388382 -23856 388450 -23800
rect 388506 -23856 388640 -23800
rect 387840 -23924 388640 -23856
rect 387840 -23980 387954 -23924
rect 388010 -23980 388078 -23924
rect 388134 -23980 388202 -23924
rect 388258 -23980 388326 -23924
rect 388382 -23980 388450 -23924
rect 388506 -23980 388640 -23924
rect 387840 -24048 388640 -23980
rect 387840 -24104 387954 -24048
rect 388010 -24104 388078 -24048
rect 388134 -24104 388202 -24048
rect 388258 -24104 388326 -24048
rect 388382 -24104 388450 -24048
rect 388506 -24104 388640 -24048
rect 387840 -24172 388640 -24104
rect 387840 -24228 387954 -24172
rect 388010 -24228 388078 -24172
rect 388134 -24228 388202 -24172
rect 388258 -24228 388326 -24172
rect 388382 -24228 388450 -24172
rect 388506 -24228 388640 -24172
rect 387840 -24296 388640 -24228
rect 387840 -24352 387954 -24296
rect 388010 -24352 388078 -24296
rect 388134 -24352 388202 -24296
rect 388258 -24352 388326 -24296
rect 388382 -24352 388450 -24296
rect 388506 -24352 388640 -24296
rect 387840 -24420 388640 -24352
rect 387840 -24476 387954 -24420
rect 388010 -24476 388078 -24420
rect 388134 -24476 388202 -24420
rect 388258 -24476 388326 -24420
rect 388382 -24476 388450 -24420
rect 388506 -24476 388640 -24420
rect 387840 -24544 388640 -24476
rect 387840 -24600 387954 -24544
rect 388010 -24600 388078 -24544
rect 388134 -24600 388202 -24544
rect 388258 -24600 388326 -24544
rect 388382 -24600 388450 -24544
rect 388506 -24600 388640 -24544
rect 387840 -24668 388640 -24600
rect 387840 -24724 387954 -24668
rect 388010 -24724 388078 -24668
rect 388134 -24724 388202 -24668
rect 388258 -24724 388326 -24668
rect 388382 -24724 388450 -24668
rect 388506 -24724 388640 -24668
rect 387840 -24792 388640 -24724
rect 387840 -24848 387954 -24792
rect 388010 -24848 388078 -24792
rect 388134 -24848 388202 -24792
rect 388258 -24848 388326 -24792
rect 388382 -24848 388450 -24792
rect 388506 -24848 388640 -24792
rect 387840 -24916 388640 -24848
rect 387840 -24972 387954 -24916
rect 388010 -24972 388078 -24916
rect 388134 -24972 388202 -24916
rect 388258 -24972 388326 -24916
rect 388382 -24972 388450 -24916
rect 388506 -24972 388640 -24916
rect 387840 -25040 388640 -24972
rect 387840 -25096 387954 -25040
rect 388010 -25096 388078 -25040
rect 388134 -25096 388202 -25040
rect 388258 -25096 388326 -25040
rect 388382 -25096 388450 -25040
rect 388506 -25096 388640 -25040
rect 387840 -25164 388640 -25096
rect 387840 -25220 387954 -25164
rect 388010 -25220 388078 -25164
rect 388134 -25220 388202 -25164
rect 388258 -25220 388326 -25164
rect 388382 -25220 388450 -25164
rect 388506 -25220 388640 -25164
rect 387840 -25288 388640 -25220
rect 387840 -25344 387954 -25288
rect 388010 -25344 388078 -25288
rect 388134 -25344 388202 -25288
rect 388258 -25344 388326 -25288
rect 388382 -25344 388450 -25288
rect 388506 -25344 388640 -25288
rect 387840 -25412 388640 -25344
rect 387840 -25468 387954 -25412
rect 388010 -25468 388078 -25412
rect 388134 -25468 388202 -25412
rect 388258 -25468 388326 -25412
rect 388382 -25468 388450 -25412
rect 388506 -25468 388640 -25412
rect 387840 -25532 388640 -25468
rect 388908 -13680 389248 -13670
rect 388908 -13736 388981 -13680
rect 389037 -13736 389123 -13680
rect 389179 -13736 389248 -13680
rect 388908 -13822 389248 -13736
rect 388908 -13878 388981 -13822
rect 389037 -13878 389123 -13822
rect 389179 -13878 389248 -13822
rect 388908 -13964 389248 -13878
rect 388908 -14020 388981 -13964
rect 389037 -14020 389123 -13964
rect 389179 -14020 389248 -13964
rect 388908 -14106 389248 -14020
rect 388908 -14162 388981 -14106
rect 389037 -14162 389123 -14106
rect 389179 -14162 389248 -14106
rect 388908 -14248 389248 -14162
rect 388908 -14304 388981 -14248
rect 389037 -14304 389123 -14248
rect 389179 -14304 389248 -14248
rect 388908 -14390 389248 -14304
rect 388908 -14446 388981 -14390
rect 389037 -14446 389123 -14390
rect 389179 -14446 389248 -14390
rect 388908 -14532 389248 -14446
rect 388908 -14588 388981 -14532
rect 389037 -14588 389123 -14532
rect 389179 -14588 389248 -14532
rect 388908 -14674 389248 -14588
rect 388908 -14730 388981 -14674
rect 389037 -14730 389123 -14674
rect 389179 -14730 389248 -14674
rect 388908 -14816 389248 -14730
rect 388908 -14872 388981 -14816
rect 389037 -14872 389123 -14816
rect 389179 -14872 389248 -14816
rect 388908 -14958 389248 -14872
rect 388908 -15014 388981 -14958
rect 389037 -15014 389123 -14958
rect 389179 -15014 389248 -14958
rect 388908 -15100 389248 -15014
rect 388908 -15156 388981 -15100
rect 389037 -15156 389123 -15100
rect 389179 -15156 389248 -15100
rect 388908 -15242 389248 -15156
rect 388908 -15298 388981 -15242
rect 389037 -15298 389123 -15242
rect 389179 -15298 389248 -15242
rect 388908 -15384 389248 -15298
rect 388908 -15440 388981 -15384
rect 389037 -15440 389123 -15384
rect 389179 -15440 389248 -15384
rect 388908 -15526 389248 -15440
rect 388908 -15582 388981 -15526
rect 389037 -15582 389123 -15526
rect 389179 -15582 389248 -15526
rect 388908 -15668 389248 -15582
rect 388908 -15724 388981 -15668
rect 389037 -15724 389123 -15668
rect 389179 -15724 389248 -15668
rect 388908 -15810 389248 -15724
rect 388908 -15866 388981 -15810
rect 389037 -15866 389123 -15810
rect 389179 -15866 389248 -15810
rect 388908 -15952 389248 -15866
rect 388908 -16008 388981 -15952
rect 389037 -16008 389123 -15952
rect 389179 -16008 389248 -15952
rect 388908 -16094 389248 -16008
rect 388908 -16150 388981 -16094
rect 389037 -16150 389123 -16094
rect 389179 -16150 389248 -16094
rect 388908 -16236 389248 -16150
rect 388908 -16292 388981 -16236
rect 389037 -16292 389123 -16236
rect 389179 -16292 389248 -16236
rect 388908 -16378 389248 -16292
rect 388908 -16434 388981 -16378
rect 389037 -16434 389123 -16378
rect 389179 -16434 389248 -16378
rect 388908 -16520 389248 -16434
rect 388908 -16576 388981 -16520
rect 389037 -16576 389123 -16520
rect 389179 -16576 389248 -16520
rect 388908 -16662 389248 -16576
rect 388908 -16718 388981 -16662
rect 389037 -16718 389123 -16662
rect 389179 -16718 389248 -16662
rect 388908 -16804 389248 -16718
rect 388908 -16860 388981 -16804
rect 389037 -16860 389123 -16804
rect 389179 -16860 389248 -16804
rect 388908 -16946 389248 -16860
rect 388908 -17002 388981 -16946
rect 389037 -17002 389123 -16946
rect 389179 -17002 389248 -16946
rect 388908 -17088 389248 -17002
rect 388908 -17144 388981 -17088
rect 389037 -17144 389123 -17088
rect 389179 -17144 389248 -17088
rect 388908 -17230 389248 -17144
rect 388908 -17286 388981 -17230
rect 389037 -17286 389123 -17230
rect 389179 -17286 389248 -17230
rect 388908 -17372 389248 -17286
rect 388908 -17428 388981 -17372
rect 389037 -17428 389123 -17372
rect 389179 -17428 389248 -17372
rect 388908 -17514 389248 -17428
rect 388908 -17570 388981 -17514
rect 389037 -17570 389123 -17514
rect 389179 -17570 389248 -17514
rect 388908 -17656 389248 -17570
rect 388908 -17712 388981 -17656
rect 389037 -17712 389123 -17656
rect 389179 -17712 389248 -17656
rect 388908 -17798 389248 -17712
rect 388908 -17854 388981 -17798
rect 389037 -17854 389123 -17798
rect 389179 -17854 389248 -17798
rect 388908 -17940 389248 -17854
rect 388908 -17996 388981 -17940
rect 389037 -17996 389123 -17940
rect 389179 -17996 389248 -17940
rect 388908 -18082 389248 -17996
rect 388908 -18138 388981 -18082
rect 389037 -18138 389123 -18082
rect 389179 -18138 389248 -18082
rect 388908 -18224 389248 -18138
rect 388908 -18280 388981 -18224
rect 389037 -18280 389123 -18224
rect 389179 -18280 389248 -18224
rect 388908 -18366 389248 -18280
rect 388908 -18422 388981 -18366
rect 389037 -18422 389123 -18366
rect 389179 -18422 389248 -18366
rect 388908 -18508 389248 -18422
rect 388908 -18564 388981 -18508
rect 389037 -18564 389123 -18508
rect 389179 -18564 389248 -18508
rect 388908 -18650 389248 -18564
rect 388908 -18706 388981 -18650
rect 389037 -18706 389123 -18650
rect 389179 -18706 389248 -18650
rect 388908 -18792 389248 -18706
rect 388908 -18848 388981 -18792
rect 389037 -18848 389123 -18792
rect 389179 -18848 389248 -18792
rect 388908 -18934 389248 -18848
rect 388908 -18990 388981 -18934
rect 389037 -18990 389123 -18934
rect 389179 -18990 389248 -18934
rect 388908 -19076 389248 -18990
rect 388908 -19132 388981 -19076
rect 389037 -19132 389123 -19076
rect 389179 -19132 389248 -19076
rect 388908 -19218 389248 -19132
rect 388908 -19274 388981 -19218
rect 389037 -19274 389123 -19218
rect 389179 -19274 389248 -19218
rect 388908 -19360 389248 -19274
rect 388908 -19416 388981 -19360
rect 389037 -19416 389123 -19360
rect 389179 -19416 389248 -19360
rect 388908 -19502 389248 -19416
rect 388908 -19558 388981 -19502
rect 389037 -19558 389123 -19502
rect 389179 -19558 389248 -19502
rect 388908 -19644 389248 -19558
rect 388908 -19700 388981 -19644
rect 389037 -19700 389123 -19644
rect 389179 -19700 389248 -19644
rect 388908 -19786 389248 -19700
rect 388908 -19842 388981 -19786
rect 389037 -19842 389123 -19786
rect 389179 -19842 389248 -19786
rect 388908 -19928 389248 -19842
rect 388908 -19984 388981 -19928
rect 389037 -19984 389123 -19928
rect 389179 -19984 389248 -19928
rect 388908 -20070 389248 -19984
rect 388908 -20126 388981 -20070
rect 389037 -20126 389123 -20070
rect 389179 -20126 389248 -20070
rect 388908 -20212 389248 -20126
rect 388908 -20268 388981 -20212
rect 389037 -20268 389123 -20212
rect 389179 -20268 389248 -20212
rect 388908 -20354 389248 -20268
rect 388908 -20410 388981 -20354
rect 389037 -20410 389123 -20354
rect 389179 -20410 389248 -20354
rect 388908 -20496 389248 -20410
rect 388908 -20552 388981 -20496
rect 389037 -20552 389123 -20496
rect 389179 -20552 389248 -20496
rect 388908 -20638 389248 -20552
rect 388908 -20694 388981 -20638
rect 389037 -20694 389123 -20638
rect 389179 -20694 389248 -20638
rect 388908 -20780 389248 -20694
rect 388908 -20836 388981 -20780
rect 389037 -20836 389123 -20780
rect 389179 -20836 389248 -20780
rect 388908 -20922 389248 -20836
rect 388908 -20978 388981 -20922
rect 389037 -20978 389123 -20922
rect 389179 -20978 389248 -20922
rect 388908 -21064 389248 -20978
rect 388908 -21120 388981 -21064
rect 389037 -21120 389123 -21064
rect 389179 -21120 389248 -21064
rect 388908 -21206 389248 -21120
rect 388908 -21262 388981 -21206
rect 389037 -21262 389123 -21206
rect 389179 -21262 389248 -21206
rect 388908 -21348 389248 -21262
rect 388908 -21404 388981 -21348
rect 389037 -21404 389123 -21348
rect 389179 -21404 389248 -21348
rect 388908 -21490 389248 -21404
rect 388908 -21546 388981 -21490
rect 389037 -21546 389123 -21490
rect 389179 -21546 389248 -21490
rect 388908 -21632 389248 -21546
rect 388908 -21688 388981 -21632
rect 389037 -21688 389123 -21632
rect 389179 -21688 389248 -21632
rect 388908 -21774 389248 -21688
rect 388908 -21830 388981 -21774
rect 389037 -21830 389123 -21774
rect 389179 -21830 389248 -21774
rect 388908 -21916 389248 -21830
rect 388908 -21972 388981 -21916
rect 389037 -21972 389123 -21916
rect 389179 -21972 389248 -21916
rect 388908 -22058 389248 -21972
rect 388908 -22114 388981 -22058
rect 389037 -22114 389123 -22058
rect 389179 -22114 389248 -22058
rect 388908 -22200 389248 -22114
rect 388908 -22256 388981 -22200
rect 389037 -22256 389123 -22200
rect 389179 -22256 389248 -22200
rect 388908 -22342 389248 -22256
rect 388908 -22398 388981 -22342
rect 389037 -22398 389123 -22342
rect 389179 -22398 389248 -22342
rect 388908 -22484 389248 -22398
rect 388908 -22540 388981 -22484
rect 389037 -22540 389123 -22484
rect 389179 -22540 389248 -22484
rect 388908 -22626 389248 -22540
rect 388908 -22682 388981 -22626
rect 389037 -22682 389123 -22626
rect 389179 -22682 389248 -22626
rect 388908 -22768 389248 -22682
rect 388908 -22824 388981 -22768
rect 389037 -22824 389123 -22768
rect 389179 -22824 389248 -22768
rect 388908 -22910 389248 -22824
rect 388908 -22966 388981 -22910
rect 389037 -22966 389123 -22910
rect 389179 -22966 389248 -22910
rect 388908 -23052 389248 -22966
rect 388908 -23108 388981 -23052
rect 389037 -23108 389123 -23052
rect 389179 -23108 389248 -23052
rect 388908 -23194 389248 -23108
rect 388908 -23250 388981 -23194
rect 389037 -23250 389123 -23194
rect 389179 -23250 389248 -23194
rect 388908 -23336 389248 -23250
rect 388908 -23392 388981 -23336
rect 389037 -23392 389123 -23336
rect 389179 -23392 389248 -23336
rect 388908 -23478 389248 -23392
rect 388908 -23534 388981 -23478
rect 389037 -23534 389123 -23478
rect 389179 -23534 389248 -23478
rect 388908 -23620 389248 -23534
rect 388908 -23676 388981 -23620
rect 389037 -23676 389123 -23620
rect 389179 -23676 389248 -23620
rect 388908 -23762 389248 -23676
rect 388908 -23818 388981 -23762
rect 389037 -23818 389123 -23762
rect 389179 -23818 389248 -23762
rect 388908 -23904 389248 -23818
rect 388908 -23960 388981 -23904
rect 389037 -23960 389123 -23904
rect 389179 -23960 389248 -23904
rect 388908 -24046 389248 -23960
rect 388908 -24102 388981 -24046
rect 389037 -24102 389123 -24046
rect 389179 -24102 389248 -24046
rect 388908 -24188 389248 -24102
rect 388908 -24244 388981 -24188
rect 389037 -24244 389123 -24188
rect 389179 -24244 389248 -24188
rect 388908 -24330 389248 -24244
rect 388908 -24386 388981 -24330
rect 389037 -24386 389123 -24330
rect 389179 -24386 389248 -24330
rect 388908 -24472 389248 -24386
rect 388908 -24528 388981 -24472
rect 389037 -24528 389123 -24472
rect 389179 -24528 389248 -24472
rect 388908 -24614 389248 -24528
rect 388908 -24670 388981 -24614
rect 389037 -24670 389123 -24614
rect 389179 -24670 389248 -24614
rect 388908 -24756 389248 -24670
rect 388908 -24812 388981 -24756
rect 389037 -24812 389123 -24756
rect 389179 -24812 389248 -24756
rect 388908 -24898 389248 -24812
rect 388908 -24954 388981 -24898
rect 389037 -24954 389123 -24898
rect 389179 -24954 389248 -24898
rect 388908 -25040 389248 -24954
rect 388908 -25096 388981 -25040
rect 389037 -25096 389123 -25040
rect 389179 -25096 389248 -25040
rect 388908 -25182 389248 -25096
rect 388908 -25238 388981 -25182
rect 389037 -25238 389123 -25182
rect 389179 -25238 389248 -25182
rect 388908 -25324 389248 -25238
rect 388908 -25380 388981 -25324
rect 389037 -25380 389123 -25324
rect 389179 -25380 389248 -25324
rect 388908 -25466 389248 -25380
rect 388908 -25522 388981 -25466
rect 389037 -25522 389123 -25466
rect 389179 -25522 389248 -25466
rect 388908 -25532 389248 -25522
rect 389308 -13680 389648 -13670
rect 389308 -13736 389382 -13680
rect 389438 -13736 389524 -13680
rect 389580 -13736 389648 -13680
rect 389308 -13822 389648 -13736
rect 389308 -13878 389382 -13822
rect 389438 -13878 389524 -13822
rect 389580 -13878 389648 -13822
rect 389308 -13964 389648 -13878
rect 389308 -14020 389382 -13964
rect 389438 -14020 389524 -13964
rect 389580 -14020 389648 -13964
rect 389308 -14106 389648 -14020
rect 389308 -14162 389382 -14106
rect 389438 -14162 389524 -14106
rect 389580 -14162 389648 -14106
rect 389308 -14248 389648 -14162
rect 389308 -14304 389382 -14248
rect 389438 -14304 389524 -14248
rect 389580 -14304 389648 -14248
rect 389308 -14390 389648 -14304
rect 389308 -14446 389382 -14390
rect 389438 -14446 389524 -14390
rect 389580 -14446 389648 -14390
rect 389308 -14532 389648 -14446
rect 389308 -14588 389382 -14532
rect 389438 -14588 389524 -14532
rect 389580 -14588 389648 -14532
rect 389308 -14674 389648 -14588
rect 389308 -14730 389382 -14674
rect 389438 -14730 389524 -14674
rect 389580 -14730 389648 -14674
rect 389308 -14816 389648 -14730
rect 389308 -14872 389382 -14816
rect 389438 -14872 389524 -14816
rect 389580 -14872 389648 -14816
rect 389308 -14958 389648 -14872
rect 389308 -15014 389382 -14958
rect 389438 -15014 389524 -14958
rect 389580 -15014 389648 -14958
rect 389308 -15100 389648 -15014
rect 389308 -15156 389382 -15100
rect 389438 -15156 389524 -15100
rect 389580 -15156 389648 -15100
rect 389308 -15242 389648 -15156
rect 389308 -15298 389382 -15242
rect 389438 -15298 389524 -15242
rect 389580 -15298 389648 -15242
rect 389308 -15384 389648 -15298
rect 389308 -15440 389382 -15384
rect 389438 -15440 389524 -15384
rect 389580 -15440 389648 -15384
rect 389308 -15526 389648 -15440
rect 389308 -15582 389382 -15526
rect 389438 -15582 389524 -15526
rect 389580 -15582 389648 -15526
rect 389308 -15668 389648 -15582
rect 389308 -15724 389382 -15668
rect 389438 -15724 389524 -15668
rect 389580 -15724 389648 -15668
rect 389308 -15810 389648 -15724
rect 389308 -15866 389382 -15810
rect 389438 -15866 389524 -15810
rect 389580 -15866 389648 -15810
rect 389308 -15952 389648 -15866
rect 389308 -16008 389382 -15952
rect 389438 -16008 389524 -15952
rect 389580 -16008 389648 -15952
rect 389308 -16094 389648 -16008
rect 389308 -16150 389382 -16094
rect 389438 -16150 389524 -16094
rect 389580 -16150 389648 -16094
rect 389308 -16236 389648 -16150
rect 389308 -16292 389382 -16236
rect 389438 -16292 389524 -16236
rect 389580 -16292 389648 -16236
rect 389308 -16378 389648 -16292
rect 389308 -16434 389382 -16378
rect 389438 -16434 389524 -16378
rect 389580 -16434 389648 -16378
rect 389308 -16520 389648 -16434
rect 389308 -16576 389382 -16520
rect 389438 -16576 389524 -16520
rect 389580 -16576 389648 -16520
rect 389308 -16662 389648 -16576
rect 389308 -16718 389382 -16662
rect 389438 -16718 389524 -16662
rect 389580 -16718 389648 -16662
rect 389308 -16804 389648 -16718
rect 389308 -16860 389382 -16804
rect 389438 -16860 389524 -16804
rect 389580 -16860 389648 -16804
rect 389308 -16946 389648 -16860
rect 389308 -17002 389382 -16946
rect 389438 -17002 389524 -16946
rect 389580 -17002 389648 -16946
rect 389308 -17088 389648 -17002
rect 389308 -17144 389382 -17088
rect 389438 -17144 389524 -17088
rect 389580 -17144 389648 -17088
rect 389308 -17230 389648 -17144
rect 389308 -17286 389382 -17230
rect 389438 -17286 389524 -17230
rect 389580 -17286 389648 -17230
rect 389308 -17372 389648 -17286
rect 389308 -17428 389382 -17372
rect 389438 -17428 389524 -17372
rect 389580 -17428 389648 -17372
rect 389308 -17514 389648 -17428
rect 389308 -17570 389382 -17514
rect 389438 -17570 389524 -17514
rect 389580 -17570 389648 -17514
rect 389308 -17656 389648 -17570
rect 389308 -17712 389382 -17656
rect 389438 -17712 389524 -17656
rect 389580 -17712 389648 -17656
rect 389308 -17798 389648 -17712
rect 389308 -17854 389382 -17798
rect 389438 -17854 389524 -17798
rect 389580 -17854 389648 -17798
rect 389308 -17940 389648 -17854
rect 389308 -17996 389382 -17940
rect 389438 -17996 389524 -17940
rect 389580 -17996 389648 -17940
rect 389308 -18082 389648 -17996
rect 389308 -18138 389382 -18082
rect 389438 -18138 389524 -18082
rect 389580 -18138 389648 -18082
rect 389308 -18224 389648 -18138
rect 389308 -18280 389382 -18224
rect 389438 -18280 389524 -18224
rect 389580 -18280 389648 -18224
rect 389308 -18366 389648 -18280
rect 389308 -18422 389382 -18366
rect 389438 -18422 389524 -18366
rect 389580 -18422 389648 -18366
rect 389308 -18508 389648 -18422
rect 389308 -18564 389382 -18508
rect 389438 -18564 389524 -18508
rect 389580 -18564 389648 -18508
rect 389308 -18650 389648 -18564
rect 389308 -18706 389382 -18650
rect 389438 -18706 389524 -18650
rect 389580 -18706 389648 -18650
rect 389308 -18792 389648 -18706
rect 389308 -18848 389382 -18792
rect 389438 -18848 389524 -18792
rect 389580 -18848 389648 -18792
rect 389308 -18934 389648 -18848
rect 389308 -18990 389382 -18934
rect 389438 -18990 389524 -18934
rect 389580 -18990 389648 -18934
rect 389308 -19076 389648 -18990
rect 389308 -19132 389382 -19076
rect 389438 -19132 389524 -19076
rect 389580 -19132 389648 -19076
rect 389308 -19218 389648 -19132
rect 389308 -19274 389382 -19218
rect 389438 -19274 389524 -19218
rect 389580 -19274 389648 -19218
rect 389308 -19360 389648 -19274
rect 389308 -19416 389382 -19360
rect 389438 -19416 389524 -19360
rect 389580 -19416 389648 -19360
rect 389308 -19502 389648 -19416
rect 389308 -19558 389382 -19502
rect 389438 -19558 389524 -19502
rect 389580 -19558 389648 -19502
rect 389308 -19644 389648 -19558
rect 389308 -19700 389382 -19644
rect 389438 -19700 389524 -19644
rect 389580 -19700 389648 -19644
rect 389308 -19786 389648 -19700
rect 389308 -19842 389382 -19786
rect 389438 -19842 389524 -19786
rect 389580 -19842 389648 -19786
rect 389308 -19928 389648 -19842
rect 389308 -19984 389382 -19928
rect 389438 -19984 389524 -19928
rect 389580 -19984 389648 -19928
rect 389308 -20070 389648 -19984
rect 389308 -20126 389382 -20070
rect 389438 -20126 389524 -20070
rect 389580 -20126 389648 -20070
rect 389308 -20212 389648 -20126
rect 389308 -20268 389382 -20212
rect 389438 -20268 389524 -20212
rect 389580 -20268 389648 -20212
rect 389308 -20354 389648 -20268
rect 389308 -20410 389382 -20354
rect 389438 -20410 389524 -20354
rect 389580 -20410 389648 -20354
rect 389308 -20496 389648 -20410
rect 389308 -20552 389382 -20496
rect 389438 -20552 389524 -20496
rect 389580 -20552 389648 -20496
rect 389308 -20638 389648 -20552
rect 389308 -20694 389382 -20638
rect 389438 -20694 389524 -20638
rect 389580 -20694 389648 -20638
rect 389308 -20780 389648 -20694
rect 389308 -20836 389382 -20780
rect 389438 -20836 389524 -20780
rect 389580 -20836 389648 -20780
rect 389308 -20922 389648 -20836
rect 389308 -20978 389382 -20922
rect 389438 -20978 389524 -20922
rect 389580 -20978 389648 -20922
rect 389308 -21064 389648 -20978
rect 389308 -21120 389382 -21064
rect 389438 -21120 389524 -21064
rect 389580 -21120 389648 -21064
rect 389308 -21206 389648 -21120
rect 389308 -21262 389382 -21206
rect 389438 -21262 389524 -21206
rect 389580 -21262 389648 -21206
rect 389308 -21348 389648 -21262
rect 389308 -21404 389382 -21348
rect 389438 -21404 389524 -21348
rect 389580 -21404 389648 -21348
rect 389308 -21490 389648 -21404
rect 389308 -21546 389382 -21490
rect 389438 -21546 389524 -21490
rect 389580 -21546 389648 -21490
rect 389308 -21632 389648 -21546
rect 389308 -21688 389382 -21632
rect 389438 -21688 389524 -21632
rect 389580 -21688 389648 -21632
rect 389308 -21774 389648 -21688
rect 389308 -21830 389382 -21774
rect 389438 -21830 389524 -21774
rect 389580 -21830 389648 -21774
rect 389308 -21916 389648 -21830
rect 389308 -21972 389382 -21916
rect 389438 -21972 389524 -21916
rect 389580 -21972 389648 -21916
rect 389308 -22058 389648 -21972
rect 389308 -22114 389382 -22058
rect 389438 -22114 389524 -22058
rect 389580 -22114 389648 -22058
rect 389308 -22200 389648 -22114
rect 389308 -22256 389382 -22200
rect 389438 -22256 389524 -22200
rect 389580 -22256 389648 -22200
rect 389308 -22342 389648 -22256
rect 389308 -22398 389382 -22342
rect 389438 -22398 389524 -22342
rect 389580 -22398 389648 -22342
rect 389308 -22484 389648 -22398
rect 389308 -22540 389382 -22484
rect 389438 -22540 389524 -22484
rect 389580 -22540 389648 -22484
rect 389308 -22626 389648 -22540
rect 389308 -22682 389382 -22626
rect 389438 -22682 389524 -22626
rect 389580 -22682 389648 -22626
rect 389308 -22768 389648 -22682
rect 389308 -22824 389382 -22768
rect 389438 -22824 389524 -22768
rect 389580 -22824 389648 -22768
rect 389308 -22910 389648 -22824
rect 389308 -22966 389382 -22910
rect 389438 -22966 389524 -22910
rect 389580 -22966 389648 -22910
rect 389308 -23052 389648 -22966
rect 389308 -23108 389382 -23052
rect 389438 -23108 389524 -23052
rect 389580 -23108 389648 -23052
rect 389308 -23194 389648 -23108
rect 389308 -23250 389382 -23194
rect 389438 -23250 389524 -23194
rect 389580 -23250 389648 -23194
rect 389308 -23336 389648 -23250
rect 389308 -23392 389382 -23336
rect 389438 -23392 389524 -23336
rect 389580 -23392 389648 -23336
rect 389308 -23478 389648 -23392
rect 389308 -23534 389382 -23478
rect 389438 -23534 389524 -23478
rect 389580 -23534 389648 -23478
rect 389308 -23620 389648 -23534
rect 389308 -23676 389382 -23620
rect 389438 -23676 389524 -23620
rect 389580 -23676 389648 -23620
rect 389308 -23762 389648 -23676
rect 389308 -23818 389382 -23762
rect 389438 -23818 389524 -23762
rect 389580 -23818 389648 -23762
rect 389308 -23904 389648 -23818
rect 389308 -23960 389382 -23904
rect 389438 -23960 389524 -23904
rect 389580 -23960 389648 -23904
rect 389308 -24046 389648 -23960
rect 389308 -24102 389382 -24046
rect 389438 -24102 389524 -24046
rect 389580 -24102 389648 -24046
rect 389308 -24188 389648 -24102
rect 389308 -24244 389382 -24188
rect 389438 -24244 389524 -24188
rect 389580 -24244 389648 -24188
rect 389308 -24330 389648 -24244
rect 389308 -24386 389382 -24330
rect 389438 -24386 389524 -24330
rect 389580 -24386 389648 -24330
rect 389308 -24472 389648 -24386
rect 389308 -24528 389382 -24472
rect 389438 -24528 389524 -24472
rect 389580 -24528 389648 -24472
rect 389308 -24614 389648 -24528
rect 389308 -24670 389382 -24614
rect 389438 -24670 389524 -24614
rect 389580 -24670 389648 -24614
rect 389308 -24756 389648 -24670
rect 389308 -24812 389382 -24756
rect 389438 -24812 389524 -24756
rect 389580 -24812 389648 -24756
rect 389308 -24898 389648 -24812
rect 389308 -24954 389382 -24898
rect 389438 -24954 389524 -24898
rect 389580 -24954 389648 -24898
rect 389308 -25040 389648 -24954
rect 389308 -25096 389382 -25040
rect 389438 -25096 389524 -25040
rect 389580 -25096 389648 -25040
rect 389308 -25182 389648 -25096
rect 389308 -25238 389382 -25182
rect 389438 -25238 389524 -25182
rect 389580 -25238 389648 -25182
rect 389308 -25324 389648 -25238
rect 389308 -25380 389382 -25324
rect 389438 -25380 389524 -25324
rect 389580 -25380 389648 -25324
rect 389308 -25466 389648 -25380
rect 389308 -25522 389382 -25466
rect 389438 -25522 389524 -25466
rect 389580 -25522 389648 -25466
rect 389308 -25532 389648 -25522
rect 389708 -13680 390048 -13670
rect 389708 -13736 389782 -13680
rect 389838 -13736 389924 -13680
rect 389980 -13736 390048 -13680
rect 389708 -13822 390048 -13736
rect 389708 -13878 389782 -13822
rect 389838 -13878 389924 -13822
rect 389980 -13878 390048 -13822
rect 389708 -13964 390048 -13878
rect 389708 -14020 389782 -13964
rect 389838 -14020 389924 -13964
rect 389980 -14020 390048 -13964
rect 389708 -14106 390048 -14020
rect 389708 -14162 389782 -14106
rect 389838 -14162 389924 -14106
rect 389980 -14162 390048 -14106
rect 389708 -14248 390048 -14162
rect 389708 -14304 389782 -14248
rect 389838 -14304 389924 -14248
rect 389980 -14304 390048 -14248
rect 389708 -14390 390048 -14304
rect 389708 -14446 389782 -14390
rect 389838 -14446 389924 -14390
rect 389980 -14446 390048 -14390
rect 389708 -14532 390048 -14446
rect 389708 -14588 389782 -14532
rect 389838 -14588 389924 -14532
rect 389980 -14588 390048 -14532
rect 389708 -14674 390048 -14588
rect 389708 -14730 389782 -14674
rect 389838 -14730 389924 -14674
rect 389980 -14730 390048 -14674
rect 389708 -14816 390048 -14730
rect 389708 -14872 389782 -14816
rect 389838 -14872 389924 -14816
rect 389980 -14872 390048 -14816
rect 389708 -14958 390048 -14872
rect 389708 -15014 389782 -14958
rect 389838 -15014 389924 -14958
rect 389980 -15014 390048 -14958
rect 389708 -15100 390048 -15014
rect 389708 -15156 389782 -15100
rect 389838 -15156 389924 -15100
rect 389980 -15156 390048 -15100
rect 389708 -15242 390048 -15156
rect 389708 -15298 389782 -15242
rect 389838 -15298 389924 -15242
rect 389980 -15298 390048 -15242
rect 389708 -15384 390048 -15298
rect 389708 -15440 389782 -15384
rect 389838 -15440 389924 -15384
rect 389980 -15440 390048 -15384
rect 389708 -15526 390048 -15440
rect 389708 -15582 389782 -15526
rect 389838 -15582 389924 -15526
rect 389980 -15582 390048 -15526
rect 389708 -15668 390048 -15582
rect 389708 -15724 389782 -15668
rect 389838 -15724 389924 -15668
rect 389980 -15724 390048 -15668
rect 389708 -15810 390048 -15724
rect 389708 -15866 389782 -15810
rect 389838 -15866 389924 -15810
rect 389980 -15866 390048 -15810
rect 389708 -15952 390048 -15866
rect 389708 -16008 389782 -15952
rect 389838 -16008 389924 -15952
rect 389980 -16008 390048 -15952
rect 389708 -16094 390048 -16008
rect 389708 -16150 389782 -16094
rect 389838 -16150 389924 -16094
rect 389980 -16150 390048 -16094
rect 389708 -16236 390048 -16150
rect 389708 -16292 389782 -16236
rect 389838 -16292 389924 -16236
rect 389980 -16292 390048 -16236
rect 389708 -16378 390048 -16292
rect 389708 -16434 389782 -16378
rect 389838 -16434 389924 -16378
rect 389980 -16434 390048 -16378
rect 389708 -16520 390048 -16434
rect 389708 -16576 389782 -16520
rect 389838 -16576 389924 -16520
rect 389980 -16576 390048 -16520
rect 389708 -16662 390048 -16576
rect 389708 -16718 389782 -16662
rect 389838 -16718 389924 -16662
rect 389980 -16718 390048 -16662
rect 389708 -16804 390048 -16718
rect 389708 -16860 389782 -16804
rect 389838 -16860 389924 -16804
rect 389980 -16860 390048 -16804
rect 389708 -16946 390048 -16860
rect 389708 -17002 389782 -16946
rect 389838 -17002 389924 -16946
rect 389980 -17002 390048 -16946
rect 389708 -17088 390048 -17002
rect 389708 -17144 389782 -17088
rect 389838 -17144 389924 -17088
rect 389980 -17144 390048 -17088
rect 389708 -17230 390048 -17144
rect 389708 -17286 389782 -17230
rect 389838 -17286 389924 -17230
rect 389980 -17286 390048 -17230
rect 389708 -17372 390048 -17286
rect 389708 -17428 389782 -17372
rect 389838 -17428 389924 -17372
rect 389980 -17428 390048 -17372
rect 389708 -17514 390048 -17428
rect 389708 -17570 389782 -17514
rect 389838 -17570 389924 -17514
rect 389980 -17570 390048 -17514
rect 389708 -17656 390048 -17570
rect 389708 -17712 389782 -17656
rect 389838 -17712 389924 -17656
rect 389980 -17712 390048 -17656
rect 389708 -17798 390048 -17712
rect 389708 -17854 389782 -17798
rect 389838 -17854 389924 -17798
rect 389980 -17854 390048 -17798
rect 389708 -17940 390048 -17854
rect 389708 -17996 389782 -17940
rect 389838 -17996 389924 -17940
rect 389980 -17996 390048 -17940
rect 389708 -18082 390048 -17996
rect 389708 -18138 389782 -18082
rect 389838 -18138 389924 -18082
rect 389980 -18138 390048 -18082
rect 389708 -18224 390048 -18138
rect 389708 -18280 389782 -18224
rect 389838 -18280 389924 -18224
rect 389980 -18280 390048 -18224
rect 389708 -18366 390048 -18280
rect 389708 -18422 389782 -18366
rect 389838 -18422 389924 -18366
rect 389980 -18422 390048 -18366
rect 389708 -18508 390048 -18422
rect 389708 -18564 389782 -18508
rect 389838 -18564 389924 -18508
rect 389980 -18564 390048 -18508
rect 389708 -18650 390048 -18564
rect 389708 -18706 389782 -18650
rect 389838 -18706 389924 -18650
rect 389980 -18706 390048 -18650
rect 389708 -18792 390048 -18706
rect 389708 -18848 389782 -18792
rect 389838 -18848 389924 -18792
rect 389980 -18848 390048 -18792
rect 389708 -18934 390048 -18848
rect 389708 -18990 389782 -18934
rect 389838 -18990 389924 -18934
rect 389980 -18990 390048 -18934
rect 389708 -19076 390048 -18990
rect 389708 -19132 389782 -19076
rect 389838 -19132 389924 -19076
rect 389980 -19132 390048 -19076
rect 389708 -19218 390048 -19132
rect 389708 -19274 389782 -19218
rect 389838 -19274 389924 -19218
rect 389980 -19274 390048 -19218
rect 389708 -19360 390048 -19274
rect 389708 -19416 389782 -19360
rect 389838 -19416 389924 -19360
rect 389980 -19416 390048 -19360
rect 389708 -19502 390048 -19416
rect 389708 -19558 389782 -19502
rect 389838 -19558 389924 -19502
rect 389980 -19558 390048 -19502
rect 389708 -19644 390048 -19558
rect 389708 -19700 389782 -19644
rect 389838 -19700 389924 -19644
rect 389980 -19700 390048 -19644
rect 389708 -19786 390048 -19700
rect 389708 -19842 389782 -19786
rect 389838 -19842 389924 -19786
rect 389980 -19842 390048 -19786
rect 389708 -19928 390048 -19842
rect 389708 -19984 389782 -19928
rect 389838 -19984 389924 -19928
rect 389980 -19984 390048 -19928
rect 389708 -20070 390048 -19984
rect 389708 -20126 389782 -20070
rect 389838 -20126 389924 -20070
rect 389980 -20126 390048 -20070
rect 389708 -20212 390048 -20126
rect 389708 -20268 389782 -20212
rect 389838 -20268 389924 -20212
rect 389980 -20268 390048 -20212
rect 389708 -20354 390048 -20268
rect 389708 -20410 389782 -20354
rect 389838 -20410 389924 -20354
rect 389980 -20410 390048 -20354
rect 389708 -20496 390048 -20410
rect 389708 -20552 389782 -20496
rect 389838 -20552 389924 -20496
rect 389980 -20552 390048 -20496
rect 389708 -20638 390048 -20552
rect 389708 -20694 389782 -20638
rect 389838 -20694 389924 -20638
rect 389980 -20694 390048 -20638
rect 389708 -20780 390048 -20694
rect 389708 -20836 389782 -20780
rect 389838 -20836 389924 -20780
rect 389980 -20836 390048 -20780
rect 389708 -20922 390048 -20836
rect 389708 -20978 389782 -20922
rect 389838 -20978 389924 -20922
rect 389980 -20978 390048 -20922
rect 389708 -21064 390048 -20978
rect 389708 -21120 389782 -21064
rect 389838 -21120 389924 -21064
rect 389980 -21120 390048 -21064
rect 389708 -21206 390048 -21120
rect 389708 -21262 389782 -21206
rect 389838 -21262 389924 -21206
rect 389980 -21262 390048 -21206
rect 389708 -21348 390048 -21262
rect 389708 -21404 389782 -21348
rect 389838 -21404 389924 -21348
rect 389980 -21404 390048 -21348
rect 389708 -21490 390048 -21404
rect 389708 -21546 389782 -21490
rect 389838 -21546 389924 -21490
rect 389980 -21546 390048 -21490
rect 389708 -21632 390048 -21546
rect 389708 -21688 389782 -21632
rect 389838 -21688 389924 -21632
rect 389980 -21688 390048 -21632
rect 389708 -21774 390048 -21688
rect 389708 -21830 389782 -21774
rect 389838 -21830 389924 -21774
rect 389980 -21830 390048 -21774
rect 389708 -21916 390048 -21830
rect 389708 -21972 389782 -21916
rect 389838 -21972 389924 -21916
rect 389980 -21972 390048 -21916
rect 389708 -22058 390048 -21972
rect 389708 -22114 389782 -22058
rect 389838 -22114 389924 -22058
rect 389980 -22114 390048 -22058
rect 389708 -22200 390048 -22114
rect 389708 -22256 389782 -22200
rect 389838 -22256 389924 -22200
rect 389980 -22256 390048 -22200
rect 389708 -22342 390048 -22256
rect 389708 -22398 389782 -22342
rect 389838 -22398 389924 -22342
rect 389980 -22398 390048 -22342
rect 389708 -22484 390048 -22398
rect 389708 -22540 389782 -22484
rect 389838 -22540 389924 -22484
rect 389980 -22540 390048 -22484
rect 389708 -22626 390048 -22540
rect 389708 -22682 389782 -22626
rect 389838 -22682 389924 -22626
rect 389980 -22682 390048 -22626
rect 389708 -22768 390048 -22682
rect 389708 -22824 389782 -22768
rect 389838 -22824 389924 -22768
rect 389980 -22824 390048 -22768
rect 389708 -22910 390048 -22824
rect 389708 -22966 389782 -22910
rect 389838 -22966 389924 -22910
rect 389980 -22966 390048 -22910
rect 389708 -23052 390048 -22966
rect 389708 -23108 389782 -23052
rect 389838 -23108 389924 -23052
rect 389980 -23108 390048 -23052
rect 389708 -23194 390048 -23108
rect 389708 -23250 389782 -23194
rect 389838 -23250 389924 -23194
rect 389980 -23250 390048 -23194
rect 389708 -23336 390048 -23250
rect 389708 -23392 389782 -23336
rect 389838 -23392 389924 -23336
rect 389980 -23392 390048 -23336
rect 389708 -23478 390048 -23392
rect 389708 -23534 389782 -23478
rect 389838 -23534 389924 -23478
rect 389980 -23534 390048 -23478
rect 389708 -23620 390048 -23534
rect 389708 -23676 389782 -23620
rect 389838 -23676 389924 -23620
rect 389980 -23676 390048 -23620
rect 389708 -23762 390048 -23676
rect 389708 -23818 389782 -23762
rect 389838 -23818 389924 -23762
rect 389980 -23818 390048 -23762
rect 389708 -23904 390048 -23818
rect 389708 -23960 389782 -23904
rect 389838 -23960 389924 -23904
rect 389980 -23960 390048 -23904
rect 389708 -24046 390048 -23960
rect 389708 -24102 389782 -24046
rect 389838 -24102 389924 -24046
rect 389980 -24102 390048 -24046
rect 389708 -24188 390048 -24102
rect 389708 -24244 389782 -24188
rect 389838 -24244 389924 -24188
rect 389980 -24244 390048 -24188
rect 389708 -24330 390048 -24244
rect 389708 -24386 389782 -24330
rect 389838 -24386 389924 -24330
rect 389980 -24386 390048 -24330
rect 389708 -24472 390048 -24386
rect 389708 -24528 389782 -24472
rect 389838 -24528 389924 -24472
rect 389980 -24528 390048 -24472
rect 389708 -24614 390048 -24528
rect 389708 -24670 389782 -24614
rect 389838 -24670 389924 -24614
rect 389980 -24670 390048 -24614
rect 389708 -24756 390048 -24670
rect 389708 -24812 389782 -24756
rect 389838 -24812 389924 -24756
rect 389980 -24812 390048 -24756
rect 389708 -24898 390048 -24812
rect 389708 -24954 389782 -24898
rect 389838 -24954 389924 -24898
rect 389980 -24954 390048 -24898
rect 389708 -25040 390048 -24954
rect 389708 -25096 389782 -25040
rect 389838 -25096 389924 -25040
rect 389980 -25096 390048 -25040
rect 389708 -25182 390048 -25096
rect 389708 -25238 389782 -25182
rect 389838 -25238 389924 -25182
rect 389980 -25238 390048 -25182
rect 389708 -25324 390048 -25238
rect 389708 -25380 389782 -25324
rect 389838 -25380 389924 -25324
rect 389980 -25380 390048 -25324
rect 389708 -25466 390048 -25380
rect 389708 -25522 389782 -25466
rect 389838 -25522 389924 -25466
rect 389980 -25522 390048 -25466
rect 389708 -25532 390048 -25522
rect 390108 -13680 390448 -13670
rect 390108 -13736 390179 -13680
rect 390235 -13736 390321 -13680
rect 390377 -13736 390448 -13680
rect 390108 -13822 390448 -13736
rect 390108 -13878 390179 -13822
rect 390235 -13878 390321 -13822
rect 390377 -13878 390448 -13822
rect 390108 -13964 390448 -13878
rect 390108 -14020 390179 -13964
rect 390235 -14020 390321 -13964
rect 390377 -14020 390448 -13964
rect 390108 -14106 390448 -14020
rect 390108 -14162 390179 -14106
rect 390235 -14162 390321 -14106
rect 390377 -14162 390448 -14106
rect 390108 -14248 390448 -14162
rect 390108 -14304 390179 -14248
rect 390235 -14304 390321 -14248
rect 390377 -14304 390448 -14248
rect 390108 -14390 390448 -14304
rect 390108 -14446 390179 -14390
rect 390235 -14446 390321 -14390
rect 390377 -14446 390448 -14390
rect 390108 -14532 390448 -14446
rect 390108 -14588 390179 -14532
rect 390235 -14588 390321 -14532
rect 390377 -14588 390448 -14532
rect 390108 -14674 390448 -14588
rect 390108 -14730 390179 -14674
rect 390235 -14730 390321 -14674
rect 390377 -14730 390448 -14674
rect 390108 -14816 390448 -14730
rect 390108 -14872 390179 -14816
rect 390235 -14872 390321 -14816
rect 390377 -14872 390448 -14816
rect 390108 -14958 390448 -14872
rect 390108 -15014 390179 -14958
rect 390235 -15014 390321 -14958
rect 390377 -15014 390448 -14958
rect 390108 -15100 390448 -15014
rect 390108 -15156 390179 -15100
rect 390235 -15156 390321 -15100
rect 390377 -15156 390448 -15100
rect 390108 -15242 390448 -15156
rect 390108 -15298 390179 -15242
rect 390235 -15298 390321 -15242
rect 390377 -15298 390448 -15242
rect 390108 -15384 390448 -15298
rect 390108 -15440 390179 -15384
rect 390235 -15440 390321 -15384
rect 390377 -15440 390448 -15384
rect 390108 -15526 390448 -15440
rect 390108 -15582 390179 -15526
rect 390235 -15582 390321 -15526
rect 390377 -15582 390448 -15526
rect 390108 -15668 390448 -15582
rect 390108 -15724 390179 -15668
rect 390235 -15724 390321 -15668
rect 390377 -15724 390448 -15668
rect 390108 -15810 390448 -15724
rect 390108 -15866 390179 -15810
rect 390235 -15866 390321 -15810
rect 390377 -15866 390448 -15810
rect 390108 -15952 390448 -15866
rect 390108 -16008 390179 -15952
rect 390235 -16008 390321 -15952
rect 390377 -16008 390448 -15952
rect 390108 -16094 390448 -16008
rect 390108 -16150 390179 -16094
rect 390235 -16150 390321 -16094
rect 390377 -16150 390448 -16094
rect 390108 -16236 390448 -16150
rect 390108 -16292 390179 -16236
rect 390235 -16292 390321 -16236
rect 390377 -16292 390448 -16236
rect 390108 -16378 390448 -16292
rect 390108 -16434 390179 -16378
rect 390235 -16434 390321 -16378
rect 390377 -16434 390448 -16378
rect 390108 -16520 390448 -16434
rect 390108 -16576 390179 -16520
rect 390235 -16576 390321 -16520
rect 390377 -16576 390448 -16520
rect 390108 -16662 390448 -16576
rect 390108 -16718 390179 -16662
rect 390235 -16718 390321 -16662
rect 390377 -16718 390448 -16662
rect 390108 -16804 390448 -16718
rect 390108 -16860 390179 -16804
rect 390235 -16860 390321 -16804
rect 390377 -16860 390448 -16804
rect 390108 -16946 390448 -16860
rect 390108 -17002 390179 -16946
rect 390235 -17002 390321 -16946
rect 390377 -17002 390448 -16946
rect 390108 -17088 390448 -17002
rect 390108 -17144 390179 -17088
rect 390235 -17144 390321 -17088
rect 390377 -17144 390448 -17088
rect 390108 -17230 390448 -17144
rect 390108 -17286 390179 -17230
rect 390235 -17286 390321 -17230
rect 390377 -17286 390448 -17230
rect 390108 -17372 390448 -17286
rect 390108 -17428 390179 -17372
rect 390235 -17428 390321 -17372
rect 390377 -17428 390448 -17372
rect 390108 -17514 390448 -17428
rect 390108 -17570 390179 -17514
rect 390235 -17570 390321 -17514
rect 390377 -17570 390448 -17514
rect 390108 -17656 390448 -17570
rect 390108 -17712 390179 -17656
rect 390235 -17712 390321 -17656
rect 390377 -17712 390448 -17656
rect 390108 -17798 390448 -17712
rect 390108 -17854 390179 -17798
rect 390235 -17854 390321 -17798
rect 390377 -17854 390448 -17798
rect 390108 -17940 390448 -17854
rect 390108 -17996 390179 -17940
rect 390235 -17996 390321 -17940
rect 390377 -17996 390448 -17940
rect 390108 -18082 390448 -17996
rect 390108 -18138 390179 -18082
rect 390235 -18138 390321 -18082
rect 390377 -18138 390448 -18082
rect 390108 -18224 390448 -18138
rect 390108 -18280 390179 -18224
rect 390235 -18280 390321 -18224
rect 390377 -18280 390448 -18224
rect 390108 -18366 390448 -18280
rect 390108 -18422 390179 -18366
rect 390235 -18422 390321 -18366
rect 390377 -18422 390448 -18366
rect 390108 -18508 390448 -18422
rect 390108 -18564 390179 -18508
rect 390235 -18564 390321 -18508
rect 390377 -18564 390448 -18508
rect 390108 -18650 390448 -18564
rect 390108 -18706 390179 -18650
rect 390235 -18706 390321 -18650
rect 390377 -18706 390448 -18650
rect 390108 -18792 390448 -18706
rect 390108 -18848 390179 -18792
rect 390235 -18848 390321 -18792
rect 390377 -18848 390448 -18792
rect 390108 -18934 390448 -18848
rect 390108 -18990 390179 -18934
rect 390235 -18990 390321 -18934
rect 390377 -18990 390448 -18934
rect 390108 -19076 390448 -18990
rect 390108 -19132 390179 -19076
rect 390235 -19132 390321 -19076
rect 390377 -19132 390448 -19076
rect 390108 -19218 390448 -19132
rect 390108 -19274 390179 -19218
rect 390235 -19274 390321 -19218
rect 390377 -19274 390448 -19218
rect 390108 -19360 390448 -19274
rect 390108 -19416 390179 -19360
rect 390235 -19416 390321 -19360
rect 390377 -19416 390448 -19360
rect 390108 -19502 390448 -19416
rect 390108 -19558 390179 -19502
rect 390235 -19558 390321 -19502
rect 390377 -19558 390448 -19502
rect 390108 -19644 390448 -19558
rect 390108 -19700 390179 -19644
rect 390235 -19700 390321 -19644
rect 390377 -19700 390448 -19644
rect 390108 -19786 390448 -19700
rect 390108 -19842 390179 -19786
rect 390235 -19842 390321 -19786
rect 390377 -19842 390448 -19786
rect 390108 -19928 390448 -19842
rect 390108 -19984 390179 -19928
rect 390235 -19984 390321 -19928
rect 390377 -19984 390448 -19928
rect 390108 -20070 390448 -19984
rect 390108 -20126 390179 -20070
rect 390235 -20126 390321 -20070
rect 390377 -20126 390448 -20070
rect 390108 -20212 390448 -20126
rect 390108 -20268 390179 -20212
rect 390235 -20268 390321 -20212
rect 390377 -20268 390448 -20212
rect 390108 -20354 390448 -20268
rect 390108 -20410 390179 -20354
rect 390235 -20410 390321 -20354
rect 390377 -20410 390448 -20354
rect 390108 -20496 390448 -20410
rect 390108 -20552 390179 -20496
rect 390235 -20552 390321 -20496
rect 390377 -20552 390448 -20496
rect 390108 -20638 390448 -20552
rect 390108 -20694 390179 -20638
rect 390235 -20694 390321 -20638
rect 390377 -20694 390448 -20638
rect 390108 -20780 390448 -20694
rect 390108 -20836 390179 -20780
rect 390235 -20836 390321 -20780
rect 390377 -20836 390448 -20780
rect 390108 -20922 390448 -20836
rect 390108 -20978 390179 -20922
rect 390235 -20978 390321 -20922
rect 390377 -20978 390448 -20922
rect 390108 -21064 390448 -20978
rect 390108 -21120 390179 -21064
rect 390235 -21120 390321 -21064
rect 390377 -21120 390448 -21064
rect 390108 -21206 390448 -21120
rect 390108 -21262 390179 -21206
rect 390235 -21262 390321 -21206
rect 390377 -21262 390448 -21206
rect 390108 -21348 390448 -21262
rect 390108 -21404 390179 -21348
rect 390235 -21404 390321 -21348
rect 390377 -21404 390448 -21348
rect 390108 -21490 390448 -21404
rect 390108 -21546 390179 -21490
rect 390235 -21546 390321 -21490
rect 390377 -21546 390448 -21490
rect 390108 -21632 390448 -21546
rect 390108 -21688 390179 -21632
rect 390235 -21688 390321 -21632
rect 390377 -21688 390448 -21632
rect 390108 -21774 390448 -21688
rect 390108 -21830 390179 -21774
rect 390235 -21830 390321 -21774
rect 390377 -21830 390448 -21774
rect 390108 -21916 390448 -21830
rect 390108 -21972 390179 -21916
rect 390235 -21972 390321 -21916
rect 390377 -21972 390448 -21916
rect 390108 -22058 390448 -21972
rect 390108 -22114 390179 -22058
rect 390235 -22114 390321 -22058
rect 390377 -22114 390448 -22058
rect 390108 -22200 390448 -22114
rect 390108 -22256 390179 -22200
rect 390235 -22256 390321 -22200
rect 390377 -22256 390448 -22200
rect 390108 -22342 390448 -22256
rect 390108 -22398 390179 -22342
rect 390235 -22398 390321 -22342
rect 390377 -22398 390448 -22342
rect 390108 -22484 390448 -22398
rect 390108 -22540 390179 -22484
rect 390235 -22540 390321 -22484
rect 390377 -22540 390448 -22484
rect 390108 -22626 390448 -22540
rect 390108 -22682 390179 -22626
rect 390235 -22682 390321 -22626
rect 390377 -22682 390448 -22626
rect 390108 -22768 390448 -22682
rect 390108 -22824 390179 -22768
rect 390235 -22824 390321 -22768
rect 390377 -22824 390448 -22768
rect 390108 -22910 390448 -22824
rect 390108 -22966 390179 -22910
rect 390235 -22966 390321 -22910
rect 390377 -22966 390448 -22910
rect 390108 -23052 390448 -22966
rect 390108 -23108 390179 -23052
rect 390235 -23108 390321 -23052
rect 390377 -23108 390448 -23052
rect 390108 -23194 390448 -23108
rect 390108 -23250 390179 -23194
rect 390235 -23250 390321 -23194
rect 390377 -23250 390448 -23194
rect 390108 -23336 390448 -23250
rect 390108 -23392 390179 -23336
rect 390235 -23392 390321 -23336
rect 390377 -23392 390448 -23336
rect 390108 -23478 390448 -23392
rect 390108 -23534 390179 -23478
rect 390235 -23534 390321 -23478
rect 390377 -23534 390448 -23478
rect 390108 -23620 390448 -23534
rect 390108 -23676 390179 -23620
rect 390235 -23676 390321 -23620
rect 390377 -23676 390448 -23620
rect 390108 -23762 390448 -23676
rect 390108 -23818 390179 -23762
rect 390235 -23818 390321 -23762
rect 390377 -23818 390448 -23762
rect 390108 -23904 390448 -23818
rect 390108 -23960 390179 -23904
rect 390235 -23960 390321 -23904
rect 390377 -23960 390448 -23904
rect 390108 -24046 390448 -23960
rect 390108 -24102 390179 -24046
rect 390235 -24102 390321 -24046
rect 390377 -24102 390448 -24046
rect 390108 -24188 390448 -24102
rect 390108 -24244 390179 -24188
rect 390235 -24244 390321 -24188
rect 390377 -24244 390448 -24188
rect 390108 -24330 390448 -24244
rect 390108 -24386 390179 -24330
rect 390235 -24386 390321 -24330
rect 390377 -24386 390448 -24330
rect 390108 -24472 390448 -24386
rect 390108 -24528 390179 -24472
rect 390235 -24528 390321 -24472
rect 390377 -24528 390448 -24472
rect 390108 -24614 390448 -24528
rect 390108 -24670 390179 -24614
rect 390235 -24670 390321 -24614
rect 390377 -24670 390448 -24614
rect 390108 -24756 390448 -24670
rect 390108 -24812 390179 -24756
rect 390235 -24812 390321 -24756
rect 390377 -24812 390448 -24756
rect 390108 -24898 390448 -24812
rect 390108 -24954 390179 -24898
rect 390235 -24954 390321 -24898
rect 390377 -24954 390448 -24898
rect 390108 -25040 390448 -24954
rect 390108 -25096 390179 -25040
rect 390235 -25096 390321 -25040
rect 390377 -25096 390448 -25040
rect 390108 -25182 390448 -25096
rect 390108 -25238 390179 -25182
rect 390235 -25238 390321 -25182
rect 390377 -25238 390448 -25182
rect 390108 -25324 390448 -25238
rect 390108 -25380 390179 -25324
rect 390235 -25380 390321 -25324
rect 390377 -25380 390448 -25324
rect 390108 -25466 390448 -25380
rect 390108 -25522 390179 -25466
rect 390235 -25522 390321 -25466
rect 390377 -25522 390448 -25466
rect 390108 -25532 390448 -25522
rect 390508 -13680 390848 -13670
rect 390508 -13736 390576 -13680
rect 390632 -13736 390718 -13680
rect 390774 -13736 390848 -13680
rect 390508 -13822 390848 -13736
rect 390508 -13878 390576 -13822
rect 390632 -13878 390718 -13822
rect 390774 -13878 390848 -13822
rect 390508 -13964 390848 -13878
rect 390508 -14020 390576 -13964
rect 390632 -14020 390718 -13964
rect 390774 -14020 390848 -13964
rect 390508 -14106 390848 -14020
rect 390508 -14162 390576 -14106
rect 390632 -14162 390718 -14106
rect 390774 -14162 390848 -14106
rect 390508 -14248 390848 -14162
rect 390508 -14304 390576 -14248
rect 390632 -14304 390718 -14248
rect 390774 -14304 390848 -14248
rect 390508 -14390 390848 -14304
rect 390508 -14446 390576 -14390
rect 390632 -14446 390718 -14390
rect 390774 -14446 390848 -14390
rect 390508 -14532 390848 -14446
rect 390508 -14588 390576 -14532
rect 390632 -14588 390718 -14532
rect 390774 -14588 390848 -14532
rect 390508 -14674 390848 -14588
rect 390508 -14730 390576 -14674
rect 390632 -14730 390718 -14674
rect 390774 -14730 390848 -14674
rect 390508 -14816 390848 -14730
rect 390508 -14872 390576 -14816
rect 390632 -14872 390718 -14816
rect 390774 -14872 390848 -14816
rect 390508 -14958 390848 -14872
rect 390508 -15014 390576 -14958
rect 390632 -15014 390718 -14958
rect 390774 -15014 390848 -14958
rect 390508 -15100 390848 -15014
rect 390508 -15156 390576 -15100
rect 390632 -15156 390718 -15100
rect 390774 -15156 390848 -15100
rect 390508 -15242 390848 -15156
rect 390508 -15298 390576 -15242
rect 390632 -15298 390718 -15242
rect 390774 -15298 390848 -15242
rect 390508 -15384 390848 -15298
rect 390508 -15440 390576 -15384
rect 390632 -15440 390718 -15384
rect 390774 -15440 390848 -15384
rect 390508 -15526 390848 -15440
rect 390508 -15582 390576 -15526
rect 390632 -15582 390718 -15526
rect 390774 -15582 390848 -15526
rect 390508 -15668 390848 -15582
rect 390508 -15724 390576 -15668
rect 390632 -15724 390718 -15668
rect 390774 -15724 390848 -15668
rect 390508 -15810 390848 -15724
rect 390508 -15866 390576 -15810
rect 390632 -15866 390718 -15810
rect 390774 -15866 390848 -15810
rect 390508 -15952 390848 -15866
rect 390508 -16008 390576 -15952
rect 390632 -16008 390718 -15952
rect 390774 -16008 390848 -15952
rect 390508 -16094 390848 -16008
rect 390508 -16150 390576 -16094
rect 390632 -16150 390718 -16094
rect 390774 -16150 390848 -16094
rect 390508 -16236 390848 -16150
rect 390508 -16292 390576 -16236
rect 390632 -16292 390718 -16236
rect 390774 -16292 390848 -16236
rect 390508 -16378 390848 -16292
rect 390508 -16434 390576 -16378
rect 390632 -16434 390718 -16378
rect 390774 -16434 390848 -16378
rect 390508 -16520 390848 -16434
rect 390508 -16576 390576 -16520
rect 390632 -16576 390718 -16520
rect 390774 -16576 390848 -16520
rect 390508 -16662 390848 -16576
rect 390508 -16718 390576 -16662
rect 390632 -16718 390718 -16662
rect 390774 -16718 390848 -16662
rect 390508 -16804 390848 -16718
rect 390508 -16860 390576 -16804
rect 390632 -16860 390718 -16804
rect 390774 -16860 390848 -16804
rect 390508 -16946 390848 -16860
rect 390508 -17002 390576 -16946
rect 390632 -17002 390718 -16946
rect 390774 -17002 390848 -16946
rect 390508 -17088 390848 -17002
rect 390508 -17144 390576 -17088
rect 390632 -17144 390718 -17088
rect 390774 -17144 390848 -17088
rect 390508 -17230 390848 -17144
rect 390508 -17286 390576 -17230
rect 390632 -17286 390718 -17230
rect 390774 -17286 390848 -17230
rect 390508 -17372 390848 -17286
rect 390508 -17428 390576 -17372
rect 390632 -17428 390718 -17372
rect 390774 -17428 390848 -17372
rect 390508 -17514 390848 -17428
rect 390508 -17570 390576 -17514
rect 390632 -17570 390718 -17514
rect 390774 -17570 390848 -17514
rect 390508 -17656 390848 -17570
rect 390508 -17712 390576 -17656
rect 390632 -17712 390718 -17656
rect 390774 -17712 390848 -17656
rect 390508 -17798 390848 -17712
rect 390508 -17854 390576 -17798
rect 390632 -17854 390718 -17798
rect 390774 -17854 390848 -17798
rect 390508 -17940 390848 -17854
rect 390508 -17996 390576 -17940
rect 390632 -17996 390718 -17940
rect 390774 -17996 390848 -17940
rect 390508 -18082 390848 -17996
rect 390508 -18138 390576 -18082
rect 390632 -18138 390718 -18082
rect 390774 -18138 390848 -18082
rect 390508 -18224 390848 -18138
rect 390508 -18280 390576 -18224
rect 390632 -18280 390718 -18224
rect 390774 -18280 390848 -18224
rect 390508 -18366 390848 -18280
rect 390508 -18422 390576 -18366
rect 390632 -18422 390718 -18366
rect 390774 -18422 390848 -18366
rect 390508 -18508 390848 -18422
rect 390508 -18564 390576 -18508
rect 390632 -18564 390718 -18508
rect 390774 -18564 390848 -18508
rect 390508 -18650 390848 -18564
rect 390508 -18706 390576 -18650
rect 390632 -18706 390718 -18650
rect 390774 -18706 390848 -18650
rect 390508 -18792 390848 -18706
rect 390508 -18848 390576 -18792
rect 390632 -18848 390718 -18792
rect 390774 -18848 390848 -18792
rect 390508 -18934 390848 -18848
rect 390508 -18990 390576 -18934
rect 390632 -18990 390718 -18934
rect 390774 -18990 390848 -18934
rect 390508 -19076 390848 -18990
rect 390508 -19132 390576 -19076
rect 390632 -19132 390718 -19076
rect 390774 -19132 390848 -19076
rect 390508 -19218 390848 -19132
rect 390508 -19274 390576 -19218
rect 390632 -19274 390718 -19218
rect 390774 -19274 390848 -19218
rect 390508 -19360 390848 -19274
rect 390508 -19416 390576 -19360
rect 390632 -19416 390718 -19360
rect 390774 -19416 390848 -19360
rect 390508 -19502 390848 -19416
rect 390508 -19558 390576 -19502
rect 390632 -19558 390718 -19502
rect 390774 -19558 390848 -19502
rect 390508 -19644 390848 -19558
rect 390508 -19700 390576 -19644
rect 390632 -19700 390718 -19644
rect 390774 -19700 390848 -19644
rect 390508 -19786 390848 -19700
rect 390508 -19842 390576 -19786
rect 390632 -19842 390718 -19786
rect 390774 -19842 390848 -19786
rect 390508 -19928 390848 -19842
rect 390508 -19984 390576 -19928
rect 390632 -19984 390718 -19928
rect 390774 -19984 390848 -19928
rect 390508 -20070 390848 -19984
rect 390508 -20126 390576 -20070
rect 390632 -20126 390718 -20070
rect 390774 -20126 390848 -20070
rect 390508 -20212 390848 -20126
rect 390508 -20268 390576 -20212
rect 390632 -20268 390718 -20212
rect 390774 -20268 390848 -20212
rect 390508 -20354 390848 -20268
rect 390508 -20410 390576 -20354
rect 390632 -20410 390718 -20354
rect 390774 -20410 390848 -20354
rect 390508 -20496 390848 -20410
rect 390508 -20552 390576 -20496
rect 390632 -20552 390718 -20496
rect 390774 -20552 390848 -20496
rect 390508 -20638 390848 -20552
rect 390508 -20694 390576 -20638
rect 390632 -20694 390718 -20638
rect 390774 -20694 390848 -20638
rect 390508 -20780 390848 -20694
rect 390508 -20836 390576 -20780
rect 390632 -20836 390718 -20780
rect 390774 -20836 390848 -20780
rect 390508 -20922 390848 -20836
rect 390508 -20978 390576 -20922
rect 390632 -20978 390718 -20922
rect 390774 -20978 390848 -20922
rect 390508 -21064 390848 -20978
rect 390508 -21120 390576 -21064
rect 390632 -21120 390718 -21064
rect 390774 -21120 390848 -21064
rect 390508 -21206 390848 -21120
rect 390508 -21262 390576 -21206
rect 390632 -21262 390718 -21206
rect 390774 -21262 390848 -21206
rect 390508 -21348 390848 -21262
rect 390508 -21404 390576 -21348
rect 390632 -21404 390718 -21348
rect 390774 -21404 390848 -21348
rect 390508 -21490 390848 -21404
rect 390508 -21546 390576 -21490
rect 390632 -21546 390718 -21490
rect 390774 -21546 390848 -21490
rect 390508 -21632 390848 -21546
rect 390508 -21688 390576 -21632
rect 390632 -21688 390718 -21632
rect 390774 -21688 390848 -21632
rect 390508 -21774 390848 -21688
rect 390508 -21830 390576 -21774
rect 390632 -21830 390718 -21774
rect 390774 -21830 390848 -21774
rect 390508 -21916 390848 -21830
rect 390508 -21972 390576 -21916
rect 390632 -21972 390718 -21916
rect 390774 -21972 390848 -21916
rect 390508 -22058 390848 -21972
rect 390508 -22114 390576 -22058
rect 390632 -22114 390718 -22058
rect 390774 -22114 390848 -22058
rect 390508 -22200 390848 -22114
rect 390508 -22256 390576 -22200
rect 390632 -22256 390718 -22200
rect 390774 -22256 390848 -22200
rect 390508 -22342 390848 -22256
rect 390508 -22398 390576 -22342
rect 390632 -22398 390718 -22342
rect 390774 -22398 390848 -22342
rect 390508 -22484 390848 -22398
rect 390508 -22540 390576 -22484
rect 390632 -22540 390718 -22484
rect 390774 -22540 390848 -22484
rect 390508 -22626 390848 -22540
rect 390508 -22682 390576 -22626
rect 390632 -22682 390718 -22626
rect 390774 -22682 390848 -22626
rect 390508 -22768 390848 -22682
rect 390508 -22824 390576 -22768
rect 390632 -22824 390718 -22768
rect 390774 -22824 390848 -22768
rect 390508 -22910 390848 -22824
rect 390508 -22966 390576 -22910
rect 390632 -22966 390718 -22910
rect 390774 -22966 390848 -22910
rect 390508 -23052 390848 -22966
rect 390508 -23108 390576 -23052
rect 390632 -23108 390718 -23052
rect 390774 -23108 390848 -23052
rect 390508 -23194 390848 -23108
rect 390508 -23250 390576 -23194
rect 390632 -23250 390718 -23194
rect 390774 -23250 390848 -23194
rect 390508 -23336 390848 -23250
rect 390508 -23392 390576 -23336
rect 390632 -23392 390718 -23336
rect 390774 -23392 390848 -23336
rect 390508 -23478 390848 -23392
rect 390508 -23534 390576 -23478
rect 390632 -23534 390718 -23478
rect 390774 -23534 390848 -23478
rect 390508 -23620 390848 -23534
rect 390508 -23676 390576 -23620
rect 390632 -23676 390718 -23620
rect 390774 -23676 390848 -23620
rect 390508 -23762 390848 -23676
rect 390508 -23818 390576 -23762
rect 390632 -23818 390718 -23762
rect 390774 -23818 390848 -23762
rect 390508 -23904 390848 -23818
rect 390508 -23960 390576 -23904
rect 390632 -23960 390718 -23904
rect 390774 -23960 390848 -23904
rect 390508 -24046 390848 -23960
rect 390508 -24102 390576 -24046
rect 390632 -24102 390718 -24046
rect 390774 -24102 390848 -24046
rect 390508 -24188 390848 -24102
rect 390508 -24244 390576 -24188
rect 390632 -24244 390718 -24188
rect 390774 -24244 390848 -24188
rect 390508 -24330 390848 -24244
rect 390508 -24386 390576 -24330
rect 390632 -24386 390718 -24330
rect 390774 -24386 390848 -24330
rect 390508 -24472 390848 -24386
rect 390508 -24528 390576 -24472
rect 390632 -24528 390718 -24472
rect 390774 -24528 390848 -24472
rect 390508 -24614 390848 -24528
rect 390508 -24670 390576 -24614
rect 390632 -24670 390718 -24614
rect 390774 -24670 390848 -24614
rect 390508 -24756 390848 -24670
rect 390508 -24812 390576 -24756
rect 390632 -24812 390718 -24756
rect 390774 -24812 390848 -24756
rect 390508 -24898 390848 -24812
rect 390508 -24954 390576 -24898
rect 390632 -24954 390718 -24898
rect 390774 -24954 390848 -24898
rect 390508 -25040 390848 -24954
rect 390508 -25096 390576 -25040
rect 390632 -25096 390718 -25040
rect 390774 -25096 390848 -25040
rect 390508 -25182 390848 -25096
rect 390508 -25238 390576 -25182
rect 390632 -25238 390718 -25182
rect 390774 -25238 390848 -25182
rect 390508 -25324 390848 -25238
rect 390508 -25380 390576 -25324
rect 390632 -25380 390718 -25324
rect 390774 -25380 390848 -25324
rect 390508 -25466 390848 -25380
rect 390508 -25522 390576 -25466
rect 390632 -25522 390718 -25466
rect 390774 -25522 390848 -25466
rect 390508 -25532 390848 -25522
rect 390908 -13680 391248 -13670
rect 390908 -13736 390980 -13680
rect 391036 -13736 391122 -13680
rect 391178 -13736 391248 -13680
rect 390908 -13822 391248 -13736
rect 390908 -13878 390980 -13822
rect 391036 -13878 391122 -13822
rect 391178 -13878 391248 -13822
rect 390908 -13964 391248 -13878
rect 390908 -14020 390980 -13964
rect 391036 -14020 391122 -13964
rect 391178 -14020 391248 -13964
rect 390908 -14106 391248 -14020
rect 390908 -14162 390980 -14106
rect 391036 -14162 391122 -14106
rect 391178 -14162 391248 -14106
rect 390908 -14248 391248 -14162
rect 390908 -14304 390980 -14248
rect 391036 -14304 391122 -14248
rect 391178 -14304 391248 -14248
rect 390908 -14390 391248 -14304
rect 390908 -14446 390980 -14390
rect 391036 -14446 391122 -14390
rect 391178 -14446 391248 -14390
rect 390908 -14532 391248 -14446
rect 390908 -14588 390980 -14532
rect 391036 -14588 391122 -14532
rect 391178 -14588 391248 -14532
rect 390908 -14674 391248 -14588
rect 390908 -14730 390980 -14674
rect 391036 -14730 391122 -14674
rect 391178 -14730 391248 -14674
rect 390908 -14816 391248 -14730
rect 390908 -14872 390980 -14816
rect 391036 -14872 391122 -14816
rect 391178 -14872 391248 -14816
rect 390908 -14958 391248 -14872
rect 390908 -15014 390980 -14958
rect 391036 -15014 391122 -14958
rect 391178 -15014 391248 -14958
rect 390908 -15100 391248 -15014
rect 390908 -15156 390980 -15100
rect 391036 -15156 391122 -15100
rect 391178 -15156 391248 -15100
rect 390908 -15242 391248 -15156
rect 390908 -15298 390980 -15242
rect 391036 -15298 391122 -15242
rect 391178 -15298 391248 -15242
rect 390908 -15384 391248 -15298
rect 390908 -15440 390980 -15384
rect 391036 -15440 391122 -15384
rect 391178 -15440 391248 -15384
rect 390908 -15526 391248 -15440
rect 390908 -15582 390980 -15526
rect 391036 -15582 391122 -15526
rect 391178 -15582 391248 -15526
rect 390908 -15668 391248 -15582
rect 390908 -15724 390980 -15668
rect 391036 -15724 391122 -15668
rect 391178 -15724 391248 -15668
rect 390908 -15810 391248 -15724
rect 390908 -15866 390980 -15810
rect 391036 -15866 391122 -15810
rect 391178 -15866 391248 -15810
rect 390908 -15952 391248 -15866
rect 390908 -16008 390980 -15952
rect 391036 -16008 391122 -15952
rect 391178 -16008 391248 -15952
rect 390908 -16094 391248 -16008
rect 390908 -16150 390980 -16094
rect 391036 -16150 391122 -16094
rect 391178 -16150 391248 -16094
rect 390908 -16236 391248 -16150
rect 390908 -16292 390980 -16236
rect 391036 -16292 391122 -16236
rect 391178 -16292 391248 -16236
rect 390908 -16378 391248 -16292
rect 390908 -16434 390980 -16378
rect 391036 -16434 391122 -16378
rect 391178 -16434 391248 -16378
rect 390908 -16520 391248 -16434
rect 390908 -16576 390980 -16520
rect 391036 -16576 391122 -16520
rect 391178 -16576 391248 -16520
rect 390908 -16662 391248 -16576
rect 390908 -16718 390980 -16662
rect 391036 -16718 391122 -16662
rect 391178 -16718 391248 -16662
rect 390908 -16804 391248 -16718
rect 390908 -16860 390980 -16804
rect 391036 -16860 391122 -16804
rect 391178 -16860 391248 -16804
rect 390908 -16946 391248 -16860
rect 390908 -17002 390980 -16946
rect 391036 -17002 391122 -16946
rect 391178 -17002 391248 -16946
rect 390908 -17088 391248 -17002
rect 390908 -17144 390980 -17088
rect 391036 -17144 391122 -17088
rect 391178 -17144 391248 -17088
rect 390908 -17230 391248 -17144
rect 390908 -17286 390980 -17230
rect 391036 -17286 391122 -17230
rect 391178 -17286 391248 -17230
rect 390908 -17372 391248 -17286
rect 390908 -17428 390980 -17372
rect 391036 -17428 391122 -17372
rect 391178 -17428 391248 -17372
rect 390908 -17514 391248 -17428
rect 390908 -17570 390980 -17514
rect 391036 -17570 391122 -17514
rect 391178 -17570 391248 -17514
rect 390908 -17656 391248 -17570
rect 390908 -17712 390980 -17656
rect 391036 -17712 391122 -17656
rect 391178 -17712 391248 -17656
rect 390908 -17798 391248 -17712
rect 390908 -17854 390980 -17798
rect 391036 -17854 391122 -17798
rect 391178 -17854 391248 -17798
rect 390908 -17940 391248 -17854
rect 390908 -17996 390980 -17940
rect 391036 -17996 391122 -17940
rect 391178 -17996 391248 -17940
rect 390908 -18082 391248 -17996
rect 390908 -18138 390980 -18082
rect 391036 -18138 391122 -18082
rect 391178 -18138 391248 -18082
rect 390908 -18224 391248 -18138
rect 390908 -18280 390980 -18224
rect 391036 -18280 391122 -18224
rect 391178 -18280 391248 -18224
rect 390908 -18366 391248 -18280
rect 390908 -18422 390980 -18366
rect 391036 -18422 391122 -18366
rect 391178 -18422 391248 -18366
rect 390908 -18508 391248 -18422
rect 390908 -18564 390980 -18508
rect 391036 -18564 391122 -18508
rect 391178 -18564 391248 -18508
rect 390908 -18650 391248 -18564
rect 390908 -18706 390980 -18650
rect 391036 -18706 391122 -18650
rect 391178 -18706 391248 -18650
rect 390908 -18792 391248 -18706
rect 390908 -18848 390980 -18792
rect 391036 -18848 391122 -18792
rect 391178 -18848 391248 -18792
rect 390908 -18934 391248 -18848
rect 390908 -18990 390980 -18934
rect 391036 -18990 391122 -18934
rect 391178 -18990 391248 -18934
rect 390908 -19076 391248 -18990
rect 390908 -19132 390980 -19076
rect 391036 -19132 391122 -19076
rect 391178 -19132 391248 -19076
rect 390908 -19218 391248 -19132
rect 390908 -19274 390980 -19218
rect 391036 -19274 391122 -19218
rect 391178 -19274 391248 -19218
rect 390908 -19360 391248 -19274
rect 390908 -19416 390980 -19360
rect 391036 -19416 391122 -19360
rect 391178 -19416 391248 -19360
rect 390908 -19502 391248 -19416
rect 390908 -19558 390980 -19502
rect 391036 -19558 391122 -19502
rect 391178 -19558 391248 -19502
rect 390908 -19644 391248 -19558
rect 390908 -19700 390980 -19644
rect 391036 -19700 391122 -19644
rect 391178 -19700 391248 -19644
rect 390908 -19786 391248 -19700
rect 390908 -19842 390980 -19786
rect 391036 -19842 391122 -19786
rect 391178 -19842 391248 -19786
rect 390908 -19928 391248 -19842
rect 390908 -19984 390980 -19928
rect 391036 -19984 391122 -19928
rect 391178 -19984 391248 -19928
rect 390908 -20070 391248 -19984
rect 390908 -20126 390980 -20070
rect 391036 -20126 391122 -20070
rect 391178 -20126 391248 -20070
rect 390908 -20212 391248 -20126
rect 390908 -20268 390980 -20212
rect 391036 -20268 391122 -20212
rect 391178 -20268 391248 -20212
rect 390908 -20354 391248 -20268
rect 390908 -20410 390980 -20354
rect 391036 -20410 391122 -20354
rect 391178 -20410 391248 -20354
rect 390908 -20496 391248 -20410
rect 390908 -20552 390980 -20496
rect 391036 -20552 391122 -20496
rect 391178 -20552 391248 -20496
rect 390908 -20638 391248 -20552
rect 390908 -20694 390980 -20638
rect 391036 -20694 391122 -20638
rect 391178 -20694 391248 -20638
rect 390908 -20780 391248 -20694
rect 390908 -20836 390980 -20780
rect 391036 -20836 391122 -20780
rect 391178 -20836 391248 -20780
rect 390908 -20922 391248 -20836
rect 390908 -20978 390980 -20922
rect 391036 -20978 391122 -20922
rect 391178 -20978 391248 -20922
rect 390908 -21064 391248 -20978
rect 390908 -21120 390980 -21064
rect 391036 -21120 391122 -21064
rect 391178 -21120 391248 -21064
rect 390908 -21206 391248 -21120
rect 390908 -21262 390980 -21206
rect 391036 -21262 391122 -21206
rect 391178 -21262 391248 -21206
rect 390908 -21348 391248 -21262
rect 390908 -21404 390980 -21348
rect 391036 -21404 391122 -21348
rect 391178 -21404 391248 -21348
rect 390908 -21490 391248 -21404
rect 390908 -21546 390980 -21490
rect 391036 -21546 391122 -21490
rect 391178 -21546 391248 -21490
rect 390908 -21632 391248 -21546
rect 390908 -21688 390980 -21632
rect 391036 -21688 391122 -21632
rect 391178 -21688 391248 -21632
rect 390908 -21774 391248 -21688
rect 390908 -21830 390980 -21774
rect 391036 -21830 391122 -21774
rect 391178 -21830 391248 -21774
rect 390908 -21916 391248 -21830
rect 390908 -21972 390980 -21916
rect 391036 -21972 391122 -21916
rect 391178 -21972 391248 -21916
rect 390908 -22058 391248 -21972
rect 390908 -22114 390980 -22058
rect 391036 -22114 391122 -22058
rect 391178 -22114 391248 -22058
rect 390908 -22200 391248 -22114
rect 390908 -22256 390980 -22200
rect 391036 -22256 391122 -22200
rect 391178 -22256 391248 -22200
rect 390908 -22342 391248 -22256
rect 390908 -22398 390980 -22342
rect 391036 -22398 391122 -22342
rect 391178 -22398 391248 -22342
rect 390908 -22484 391248 -22398
rect 390908 -22540 390980 -22484
rect 391036 -22540 391122 -22484
rect 391178 -22540 391248 -22484
rect 390908 -22626 391248 -22540
rect 390908 -22682 390980 -22626
rect 391036 -22682 391122 -22626
rect 391178 -22682 391248 -22626
rect 390908 -22768 391248 -22682
rect 390908 -22824 390980 -22768
rect 391036 -22824 391122 -22768
rect 391178 -22824 391248 -22768
rect 390908 -22910 391248 -22824
rect 390908 -22966 390980 -22910
rect 391036 -22966 391122 -22910
rect 391178 -22966 391248 -22910
rect 390908 -23052 391248 -22966
rect 390908 -23108 390980 -23052
rect 391036 -23108 391122 -23052
rect 391178 -23108 391248 -23052
rect 390908 -23194 391248 -23108
rect 390908 -23250 390980 -23194
rect 391036 -23250 391122 -23194
rect 391178 -23250 391248 -23194
rect 390908 -23336 391248 -23250
rect 390908 -23392 390980 -23336
rect 391036 -23392 391122 -23336
rect 391178 -23392 391248 -23336
rect 390908 -23478 391248 -23392
rect 390908 -23534 390980 -23478
rect 391036 -23534 391122 -23478
rect 391178 -23534 391248 -23478
rect 390908 -23620 391248 -23534
rect 390908 -23676 390980 -23620
rect 391036 -23676 391122 -23620
rect 391178 -23676 391248 -23620
rect 390908 -23762 391248 -23676
rect 390908 -23818 390980 -23762
rect 391036 -23818 391122 -23762
rect 391178 -23818 391248 -23762
rect 390908 -23904 391248 -23818
rect 390908 -23960 390980 -23904
rect 391036 -23960 391122 -23904
rect 391178 -23960 391248 -23904
rect 390908 -24046 391248 -23960
rect 390908 -24102 390980 -24046
rect 391036 -24102 391122 -24046
rect 391178 -24102 391248 -24046
rect 390908 -24188 391248 -24102
rect 390908 -24244 390980 -24188
rect 391036 -24244 391122 -24188
rect 391178 -24244 391248 -24188
rect 390908 -24330 391248 -24244
rect 390908 -24386 390980 -24330
rect 391036 -24386 391122 -24330
rect 391178 -24386 391248 -24330
rect 390908 -24472 391248 -24386
rect 390908 -24528 390980 -24472
rect 391036 -24528 391122 -24472
rect 391178 -24528 391248 -24472
rect 390908 -24614 391248 -24528
rect 390908 -24670 390980 -24614
rect 391036 -24670 391122 -24614
rect 391178 -24670 391248 -24614
rect 390908 -24756 391248 -24670
rect 390908 -24812 390980 -24756
rect 391036 -24812 391122 -24756
rect 391178 -24812 391248 -24756
rect 390908 -24898 391248 -24812
rect 390908 -24954 390980 -24898
rect 391036 -24954 391122 -24898
rect 391178 -24954 391248 -24898
rect 390908 -25040 391248 -24954
rect 390908 -25096 390980 -25040
rect 391036 -25096 391122 -25040
rect 391178 -25096 391248 -25040
rect 390908 -25182 391248 -25096
rect 390908 -25238 390980 -25182
rect 391036 -25238 391122 -25182
rect 391178 -25238 391248 -25182
rect 390908 -25324 391248 -25238
rect 390908 -25380 390980 -25324
rect 391036 -25380 391122 -25324
rect 391178 -25380 391248 -25324
rect 390908 -25466 391248 -25380
rect 390908 -25522 390980 -25466
rect 391036 -25522 391122 -25466
rect 391178 -25522 391248 -25466
rect 390908 -25532 391248 -25522
rect 391308 -13680 391648 -13670
rect 391308 -13736 391376 -13680
rect 391432 -13736 391518 -13680
rect 391574 -13736 391648 -13680
rect 391308 -13822 391648 -13736
rect 391308 -13878 391376 -13822
rect 391432 -13878 391518 -13822
rect 391574 -13878 391648 -13822
rect 391308 -13964 391648 -13878
rect 391308 -14020 391376 -13964
rect 391432 -14020 391518 -13964
rect 391574 -14020 391648 -13964
rect 391308 -14106 391648 -14020
rect 391308 -14162 391376 -14106
rect 391432 -14162 391518 -14106
rect 391574 -14162 391648 -14106
rect 391308 -14248 391648 -14162
rect 391308 -14304 391376 -14248
rect 391432 -14304 391518 -14248
rect 391574 -14304 391648 -14248
rect 391308 -14390 391648 -14304
rect 391308 -14446 391376 -14390
rect 391432 -14446 391518 -14390
rect 391574 -14446 391648 -14390
rect 391308 -14532 391648 -14446
rect 391308 -14588 391376 -14532
rect 391432 -14588 391518 -14532
rect 391574 -14588 391648 -14532
rect 391308 -14674 391648 -14588
rect 391308 -14730 391376 -14674
rect 391432 -14730 391518 -14674
rect 391574 -14730 391648 -14674
rect 391308 -14816 391648 -14730
rect 391308 -14872 391376 -14816
rect 391432 -14872 391518 -14816
rect 391574 -14872 391648 -14816
rect 391308 -14958 391648 -14872
rect 391308 -15014 391376 -14958
rect 391432 -15014 391518 -14958
rect 391574 -15014 391648 -14958
rect 391308 -15100 391648 -15014
rect 391308 -15156 391376 -15100
rect 391432 -15156 391518 -15100
rect 391574 -15156 391648 -15100
rect 391308 -15242 391648 -15156
rect 391308 -15298 391376 -15242
rect 391432 -15298 391518 -15242
rect 391574 -15298 391648 -15242
rect 391308 -15384 391648 -15298
rect 391308 -15440 391376 -15384
rect 391432 -15440 391518 -15384
rect 391574 -15440 391648 -15384
rect 391308 -15526 391648 -15440
rect 391308 -15582 391376 -15526
rect 391432 -15582 391518 -15526
rect 391574 -15582 391648 -15526
rect 391308 -15668 391648 -15582
rect 391308 -15724 391376 -15668
rect 391432 -15724 391518 -15668
rect 391574 -15724 391648 -15668
rect 391308 -15810 391648 -15724
rect 391308 -15866 391376 -15810
rect 391432 -15866 391518 -15810
rect 391574 -15866 391648 -15810
rect 391308 -15952 391648 -15866
rect 391308 -16008 391376 -15952
rect 391432 -16008 391518 -15952
rect 391574 -16008 391648 -15952
rect 391308 -16094 391648 -16008
rect 391308 -16150 391376 -16094
rect 391432 -16150 391518 -16094
rect 391574 -16150 391648 -16094
rect 391308 -16236 391648 -16150
rect 391308 -16292 391376 -16236
rect 391432 -16292 391518 -16236
rect 391574 -16292 391648 -16236
rect 391308 -16378 391648 -16292
rect 391308 -16434 391376 -16378
rect 391432 -16434 391518 -16378
rect 391574 -16434 391648 -16378
rect 391308 -16520 391648 -16434
rect 391308 -16576 391376 -16520
rect 391432 -16576 391518 -16520
rect 391574 -16576 391648 -16520
rect 391308 -16662 391648 -16576
rect 391308 -16718 391376 -16662
rect 391432 -16718 391518 -16662
rect 391574 -16718 391648 -16662
rect 391308 -16804 391648 -16718
rect 391308 -16860 391376 -16804
rect 391432 -16860 391518 -16804
rect 391574 -16860 391648 -16804
rect 391308 -16946 391648 -16860
rect 391308 -17002 391376 -16946
rect 391432 -17002 391518 -16946
rect 391574 -17002 391648 -16946
rect 391308 -17088 391648 -17002
rect 391308 -17144 391376 -17088
rect 391432 -17144 391518 -17088
rect 391574 -17144 391648 -17088
rect 391308 -17230 391648 -17144
rect 391308 -17286 391376 -17230
rect 391432 -17286 391518 -17230
rect 391574 -17286 391648 -17230
rect 391308 -17372 391648 -17286
rect 391308 -17428 391376 -17372
rect 391432 -17428 391518 -17372
rect 391574 -17428 391648 -17372
rect 391308 -17514 391648 -17428
rect 391308 -17570 391376 -17514
rect 391432 -17570 391518 -17514
rect 391574 -17570 391648 -17514
rect 391308 -17656 391648 -17570
rect 391308 -17712 391376 -17656
rect 391432 -17712 391518 -17656
rect 391574 -17712 391648 -17656
rect 391308 -17798 391648 -17712
rect 391308 -17854 391376 -17798
rect 391432 -17854 391518 -17798
rect 391574 -17854 391648 -17798
rect 391308 -17940 391648 -17854
rect 391308 -17996 391376 -17940
rect 391432 -17996 391518 -17940
rect 391574 -17996 391648 -17940
rect 391308 -18082 391648 -17996
rect 391308 -18138 391376 -18082
rect 391432 -18138 391518 -18082
rect 391574 -18138 391648 -18082
rect 391308 -18224 391648 -18138
rect 391308 -18280 391376 -18224
rect 391432 -18280 391518 -18224
rect 391574 -18280 391648 -18224
rect 391308 -18366 391648 -18280
rect 391308 -18422 391376 -18366
rect 391432 -18422 391518 -18366
rect 391574 -18422 391648 -18366
rect 391308 -18508 391648 -18422
rect 391308 -18564 391376 -18508
rect 391432 -18564 391518 -18508
rect 391574 -18564 391648 -18508
rect 391308 -18650 391648 -18564
rect 391308 -18706 391376 -18650
rect 391432 -18706 391518 -18650
rect 391574 -18706 391648 -18650
rect 391308 -18792 391648 -18706
rect 391308 -18848 391376 -18792
rect 391432 -18848 391518 -18792
rect 391574 -18848 391648 -18792
rect 391308 -18934 391648 -18848
rect 391308 -18990 391376 -18934
rect 391432 -18990 391518 -18934
rect 391574 -18990 391648 -18934
rect 391308 -19076 391648 -18990
rect 391308 -19132 391376 -19076
rect 391432 -19132 391518 -19076
rect 391574 -19132 391648 -19076
rect 391308 -19218 391648 -19132
rect 391308 -19274 391376 -19218
rect 391432 -19274 391518 -19218
rect 391574 -19274 391648 -19218
rect 391308 -19360 391648 -19274
rect 391308 -19416 391376 -19360
rect 391432 -19416 391518 -19360
rect 391574 -19416 391648 -19360
rect 391308 -19502 391648 -19416
rect 391308 -19558 391376 -19502
rect 391432 -19558 391518 -19502
rect 391574 -19558 391648 -19502
rect 391308 -19644 391648 -19558
rect 391308 -19700 391376 -19644
rect 391432 -19700 391518 -19644
rect 391574 -19700 391648 -19644
rect 391308 -19786 391648 -19700
rect 391308 -19842 391376 -19786
rect 391432 -19842 391518 -19786
rect 391574 -19842 391648 -19786
rect 391308 -19928 391648 -19842
rect 391308 -19984 391376 -19928
rect 391432 -19984 391518 -19928
rect 391574 -19984 391648 -19928
rect 391308 -20070 391648 -19984
rect 391308 -20126 391376 -20070
rect 391432 -20126 391518 -20070
rect 391574 -20126 391648 -20070
rect 391308 -20212 391648 -20126
rect 391308 -20268 391376 -20212
rect 391432 -20268 391518 -20212
rect 391574 -20268 391648 -20212
rect 391308 -20354 391648 -20268
rect 391308 -20410 391376 -20354
rect 391432 -20410 391518 -20354
rect 391574 -20410 391648 -20354
rect 391308 -20496 391648 -20410
rect 391308 -20552 391376 -20496
rect 391432 -20552 391518 -20496
rect 391574 -20552 391648 -20496
rect 391308 -20638 391648 -20552
rect 391308 -20694 391376 -20638
rect 391432 -20694 391518 -20638
rect 391574 -20694 391648 -20638
rect 391308 -20780 391648 -20694
rect 391308 -20836 391376 -20780
rect 391432 -20836 391518 -20780
rect 391574 -20836 391648 -20780
rect 391308 -20922 391648 -20836
rect 391308 -20978 391376 -20922
rect 391432 -20978 391518 -20922
rect 391574 -20978 391648 -20922
rect 391308 -21064 391648 -20978
rect 391308 -21120 391376 -21064
rect 391432 -21120 391518 -21064
rect 391574 -21120 391648 -21064
rect 391308 -21206 391648 -21120
rect 391308 -21262 391376 -21206
rect 391432 -21262 391518 -21206
rect 391574 -21262 391648 -21206
rect 391308 -21348 391648 -21262
rect 391308 -21404 391376 -21348
rect 391432 -21404 391518 -21348
rect 391574 -21404 391648 -21348
rect 391308 -21490 391648 -21404
rect 391308 -21546 391376 -21490
rect 391432 -21546 391518 -21490
rect 391574 -21546 391648 -21490
rect 391308 -21632 391648 -21546
rect 391308 -21688 391376 -21632
rect 391432 -21688 391518 -21632
rect 391574 -21688 391648 -21632
rect 391308 -21774 391648 -21688
rect 391308 -21830 391376 -21774
rect 391432 -21830 391518 -21774
rect 391574 -21830 391648 -21774
rect 391308 -21916 391648 -21830
rect 391308 -21972 391376 -21916
rect 391432 -21972 391518 -21916
rect 391574 -21972 391648 -21916
rect 391308 -22058 391648 -21972
rect 391308 -22114 391376 -22058
rect 391432 -22114 391518 -22058
rect 391574 -22114 391648 -22058
rect 391308 -22200 391648 -22114
rect 391308 -22256 391376 -22200
rect 391432 -22256 391518 -22200
rect 391574 -22256 391648 -22200
rect 391308 -22342 391648 -22256
rect 391308 -22398 391376 -22342
rect 391432 -22398 391518 -22342
rect 391574 -22398 391648 -22342
rect 391308 -22484 391648 -22398
rect 391308 -22540 391376 -22484
rect 391432 -22540 391518 -22484
rect 391574 -22540 391648 -22484
rect 391308 -22626 391648 -22540
rect 391308 -22682 391376 -22626
rect 391432 -22682 391518 -22626
rect 391574 -22682 391648 -22626
rect 391308 -22768 391648 -22682
rect 391308 -22824 391376 -22768
rect 391432 -22824 391518 -22768
rect 391574 -22824 391648 -22768
rect 391308 -22910 391648 -22824
rect 391308 -22966 391376 -22910
rect 391432 -22966 391518 -22910
rect 391574 -22966 391648 -22910
rect 391308 -23052 391648 -22966
rect 391308 -23108 391376 -23052
rect 391432 -23108 391518 -23052
rect 391574 -23108 391648 -23052
rect 391308 -23194 391648 -23108
rect 391308 -23250 391376 -23194
rect 391432 -23250 391518 -23194
rect 391574 -23250 391648 -23194
rect 391308 -23336 391648 -23250
rect 391308 -23392 391376 -23336
rect 391432 -23392 391518 -23336
rect 391574 -23392 391648 -23336
rect 391308 -23478 391648 -23392
rect 391308 -23534 391376 -23478
rect 391432 -23534 391518 -23478
rect 391574 -23534 391648 -23478
rect 391308 -23620 391648 -23534
rect 391308 -23676 391376 -23620
rect 391432 -23676 391518 -23620
rect 391574 -23676 391648 -23620
rect 391308 -23762 391648 -23676
rect 391308 -23818 391376 -23762
rect 391432 -23818 391518 -23762
rect 391574 -23818 391648 -23762
rect 391308 -23904 391648 -23818
rect 391308 -23960 391376 -23904
rect 391432 -23960 391518 -23904
rect 391574 -23960 391648 -23904
rect 391308 -24046 391648 -23960
rect 391308 -24102 391376 -24046
rect 391432 -24102 391518 -24046
rect 391574 -24102 391648 -24046
rect 391308 -24188 391648 -24102
rect 391308 -24244 391376 -24188
rect 391432 -24244 391518 -24188
rect 391574 -24244 391648 -24188
rect 391308 -24330 391648 -24244
rect 391308 -24386 391376 -24330
rect 391432 -24386 391518 -24330
rect 391574 -24386 391648 -24330
rect 391308 -24472 391648 -24386
rect 391308 -24528 391376 -24472
rect 391432 -24528 391518 -24472
rect 391574 -24528 391648 -24472
rect 391308 -24614 391648 -24528
rect 391308 -24670 391376 -24614
rect 391432 -24670 391518 -24614
rect 391574 -24670 391648 -24614
rect 391308 -24756 391648 -24670
rect 391308 -24812 391376 -24756
rect 391432 -24812 391518 -24756
rect 391574 -24812 391648 -24756
rect 391308 -24898 391648 -24812
rect 391308 -24954 391376 -24898
rect 391432 -24954 391518 -24898
rect 391574 -24954 391648 -24898
rect 391308 -25040 391648 -24954
rect 391308 -25096 391376 -25040
rect 391432 -25096 391518 -25040
rect 391574 -25096 391648 -25040
rect 391308 -25182 391648 -25096
rect 391308 -25238 391376 -25182
rect 391432 -25238 391518 -25182
rect 391574 -25238 391648 -25182
rect 391308 -25324 391648 -25238
rect 391308 -25380 391376 -25324
rect 391432 -25380 391518 -25324
rect 391574 -25380 391648 -25324
rect 391308 -25466 391648 -25380
rect 391308 -25522 391376 -25466
rect 391432 -25522 391518 -25466
rect 391574 -25522 391648 -25466
rect 391308 -25532 391648 -25522
rect 391708 -13680 392048 -13670
rect 391708 -13736 391776 -13680
rect 391832 -13736 391918 -13680
rect 391974 -13736 392048 -13680
rect 391708 -13822 392048 -13736
rect 391708 -13878 391776 -13822
rect 391832 -13878 391918 -13822
rect 391974 -13878 392048 -13822
rect 391708 -13964 392048 -13878
rect 391708 -14020 391776 -13964
rect 391832 -14020 391918 -13964
rect 391974 -14020 392048 -13964
rect 391708 -14106 392048 -14020
rect 391708 -14162 391776 -14106
rect 391832 -14162 391918 -14106
rect 391974 -14162 392048 -14106
rect 391708 -14248 392048 -14162
rect 391708 -14304 391776 -14248
rect 391832 -14304 391918 -14248
rect 391974 -14304 392048 -14248
rect 391708 -14390 392048 -14304
rect 391708 -14446 391776 -14390
rect 391832 -14446 391918 -14390
rect 391974 -14446 392048 -14390
rect 391708 -14532 392048 -14446
rect 391708 -14588 391776 -14532
rect 391832 -14588 391918 -14532
rect 391974 -14588 392048 -14532
rect 391708 -14674 392048 -14588
rect 391708 -14730 391776 -14674
rect 391832 -14730 391918 -14674
rect 391974 -14730 392048 -14674
rect 391708 -14816 392048 -14730
rect 391708 -14872 391776 -14816
rect 391832 -14872 391918 -14816
rect 391974 -14872 392048 -14816
rect 391708 -14958 392048 -14872
rect 391708 -15014 391776 -14958
rect 391832 -15014 391918 -14958
rect 391974 -15014 392048 -14958
rect 391708 -15100 392048 -15014
rect 391708 -15156 391776 -15100
rect 391832 -15156 391918 -15100
rect 391974 -15156 392048 -15100
rect 391708 -15242 392048 -15156
rect 391708 -15298 391776 -15242
rect 391832 -15298 391918 -15242
rect 391974 -15298 392048 -15242
rect 391708 -15384 392048 -15298
rect 391708 -15440 391776 -15384
rect 391832 -15440 391918 -15384
rect 391974 -15440 392048 -15384
rect 391708 -15526 392048 -15440
rect 391708 -15582 391776 -15526
rect 391832 -15582 391918 -15526
rect 391974 -15582 392048 -15526
rect 391708 -15668 392048 -15582
rect 391708 -15724 391776 -15668
rect 391832 -15724 391918 -15668
rect 391974 -15724 392048 -15668
rect 391708 -15810 392048 -15724
rect 391708 -15866 391776 -15810
rect 391832 -15866 391918 -15810
rect 391974 -15866 392048 -15810
rect 391708 -15952 392048 -15866
rect 391708 -16008 391776 -15952
rect 391832 -16008 391918 -15952
rect 391974 -16008 392048 -15952
rect 391708 -16094 392048 -16008
rect 391708 -16150 391776 -16094
rect 391832 -16150 391918 -16094
rect 391974 -16150 392048 -16094
rect 391708 -16236 392048 -16150
rect 391708 -16292 391776 -16236
rect 391832 -16292 391918 -16236
rect 391974 -16292 392048 -16236
rect 391708 -16378 392048 -16292
rect 391708 -16434 391776 -16378
rect 391832 -16434 391918 -16378
rect 391974 -16434 392048 -16378
rect 391708 -16520 392048 -16434
rect 391708 -16576 391776 -16520
rect 391832 -16576 391918 -16520
rect 391974 -16576 392048 -16520
rect 391708 -16662 392048 -16576
rect 391708 -16718 391776 -16662
rect 391832 -16718 391918 -16662
rect 391974 -16718 392048 -16662
rect 391708 -16804 392048 -16718
rect 391708 -16860 391776 -16804
rect 391832 -16860 391918 -16804
rect 391974 -16860 392048 -16804
rect 391708 -16946 392048 -16860
rect 391708 -17002 391776 -16946
rect 391832 -17002 391918 -16946
rect 391974 -17002 392048 -16946
rect 391708 -17088 392048 -17002
rect 391708 -17144 391776 -17088
rect 391832 -17144 391918 -17088
rect 391974 -17144 392048 -17088
rect 391708 -17230 392048 -17144
rect 391708 -17286 391776 -17230
rect 391832 -17286 391918 -17230
rect 391974 -17286 392048 -17230
rect 391708 -17372 392048 -17286
rect 391708 -17428 391776 -17372
rect 391832 -17428 391918 -17372
rect 391974 -17428 392048 -17372
rect 391708 -17514 392048 -17428
rect 391708 -17570 391776 -17514
rect 391832 -17570 391918 -17514
rect 391974 -17570 392048 -17514
rect 391708 -17656 392048 -17570
rect 391708 -17712 391776 -17656
rect 391832 -17712 391918 -17656
rect 391974 -17712 392048 -17656
rect 391708 -17798 392048 -17712
rect 391708 -17854 391776 -17798
rect 391832 -17854 391918 -17798
rect 391974 -17854 392048 -17798
rect 391708 -17940 392048 -17854
rect 391708 -17996 391776 -17940
rect 391832 -17996 391918 -17940
rect 391974 -17996 392048 -17940
rect 391708 -18082 392048 -17996
rect 391708 -18138 391776 -18082
rect 391832 -18138 391918 -18082
rect 391974 -18138 392048 -18082
rect 391708 -18224 392048 -18138
rect 391708 -18280 391776 -18224
rect 391832 -18280 391918 -18224
rect 391974 -18280 392048 -18224
rect 391708 -18366 392048 -18280
rect 391708 -18422 391776 -18366
rect 391832 -18422 391918 -18366
rect 391974 -18422 392048 -18366
rect 391708 -18508 392048 -18422
rect 391708 -18564 391776 -18508
rect 391832 -18564 391918 -18508
rect 391974 -18564 392048 -18508
rect 391708 -18650 392048 -18564
rect 391708 -18706 391776 -18650
rect 391832 -18706 391918 -18650
rect 391974 -18706 392048 -18650
rect 391708 -18792 392048 -18706
rect 391708 -18848 391776 -18792
rect 391832 -18848 391918 -18792
rect 391974 -18848 392048 -18792
rect 391708 -18934 392048 -18848
rect 391708 -18990 391776 -18934
rect 391832 -18990 391918 -18934
rect 391974 -18990 392048 -18934
rect 391708 -19076 392048 -18990
rect 391708 -19132 391776 -19076
rect 391832 -19132 391918 -19076
rect 391974 -19132 392048 -19076
rect 391708 -19218 392048 -19132
rect 391708 -19274 391776 -19218
rect 391832 -19274 391918 -19218
rect 391974 -19274 392048 -19218
rect 391708 -19360 392048 -19274
rect 391708 -19416 391776 -19360
rect 391832 -19416 391918 -19360
rect 391974 -19416 392048 -19360
rect 391708 -19502 392048 -19416
rect 391708 -19558 391776 -19502
rect 391832 -19558 391918 -19502
rect 391974 -19558 392048 -19502
rect 391708 -19644 392048 -19558
rect 391708 -19700 391776 -19644
rect 391832 -19700 391918 -19644
rect 391974 -19700 392048 -19644
rect 391708 -19786 392048 -19700
rect 391708 -19842 391776 -19786
rect 391832 -19842 391918 -19786
rect 391974 -19842 392048 -19786
rect 391708 -19928 392048 -19842
rect 391708 -19984 391776 -19928
rect 391832 -19984 391918 -19928
rect 391974 -19984 392048 -19928
rect 391708 -20070 392048 -19984
rect 391708 -20126 391776 -20070
rect 391832 -20126 391918 -20070
rect 391974 -20126 392048 -20070
rect 391708 -20212 392048 -20126
rect 391708 -20268 391776 -20212
rect 391832 -20268 391918 -20212
rect 391974 -20268 392048 -20212
rect 391708 -20354 392048 -20268
rect 391708 -20410 391776 -20354
rect 391832 -20410 391918 -20354
rect 391974 -20410 392048 -20354
rect 391708 -20496 392048 -20410
rect 391708 -20552 391776 -20496
rect 391832 -20552 391918 -20496
rect 391974 -20552 392048 -20496
rect 391708 -20638 392048 -20552
rect 391708 -20694 391776 -20638
rect 391832 -20694 391918 -20638
rect 391974 -20694 392048 -20638
rect 391708 -20780 392048 -20694
rect 391708 -20836 391776 -20780
rect 391832 -20836 391918 -20780
rect 391974 -20836 392048 -20780
rect 391708 -20922 392048 -20836
rect 391708 -20978 391776 -20922
rect 391832 -20978 391918 -20922
rect 391974 -20978 392048 -20922
rect 391708 -21064 392048 -20978
rect 391708 -21120 391776 -21064
rect 391832 -21120 391918 -21064
rect 391974 -21120 392048 -21064
rect 391708 -21206 392048 -21120
rect 391708 -21262 391776 -21206
rect 391832 -21262 391918 -21206
rect 391974 -21262 392048 -21206
rect 391708 -21348 392048 -21262
rect 391708 -21404 391776 -21348
rect 391832 -21404 391918 -21348
rect 391974 -21404 392048 -21348
rect 391708 -21490 392048 -21404
rect 391708 -21546 391776 -21490
rect 391832 -21546 391918 -21490
rect 391974 -21546 392048 -21490
rect 391708 -21632 392048 -21546
rect 391708 -21688 391776 -21632
rect 391832 -21688 391918 -21632
rect 391974 -21688 392048 -21632
rect 391708 -21774 392048 -21688
rect 391708 -21830 391776 -21774
rect 391832 -21830 391918 -21774
rect 391974 -21830 392048 -21774
rect 391708 -21916 392048 -21830
rect 391708 -21972 391776 -21916
rect 391832 -21972 391918 -21916
rect 391974 -21972 392048 -21916
rect 391708 -22058 392048 -21972
rect 391708 -22114 391776 -22058
rect 391832 -22114 391918 -22058
rect 391974 -22114 392048 -22058
rect 391708 -22200 392048 -22114
rect 391708 -22256 391776 -22200
rect 391832 -22256 391918 -22200
rect 391974 -22256 392048 -22200
rect 391708 -22342 392048 -22256
rect 391708 -22398 391776 -22342
rect 391832 -22398 391918 -22342
rect 391974 -22398 392048 -22342
rect 391708 -22484 392048 -22398
rect 391708 -22540 391776 -22484
rect 391832 -22540 391918 -22484
rect 391974 -22540 392048 -22484
rect 391708 -22626 392048 -22540
rect 391708 -22682 391776 -22626
rect 391832 -22682 391918 -22626
rect 391974 -22682 392048 -22626
rect 391708 -22768 392048 -22682
rect 391708 -22824 391776 -22768
rect 391832 -22824 391918 -22768
rect 391974 -22824 392048 -22768
rect 391708 -22910 392048 -22824
rect 391708 -22966 391776 -22910
rect 391832 -22966 391918 -22910
rect 391974 -22966 392048 -22910
rect 391708 -23052 392048 -22966
rect 391708 -23108 391776 -23052
rect 391832 -23108 391918 -23052
rect 391974 -23108 392048 -23052
rect 391708 -23194 392048 -23108
rect 391708 -23250 391776 -23194
rect 391832 -23250 391918 -23194
rect 391974 -23250 392048 -23194
rect 391708 -23336 392048 -23250
rect 391708 -23392 391776 -23336
rect 391832 -23392 391918 -23336
rect 391974 -23392 392048 -23336
rect 391708 -23478 392048 -23392
rect 391708 -23534 391776 -23478
rect 391832 -23534 391918 -23478
rect 391974 -23534 392048 -23478
rect 391708 -23620 392048 -23534
rect 391708 -23676 391776 -23620
rect 391832 -23676 391918 -23620
rect 391974 -23676 392048 -23620
rect 391708 -23762 392048 -23676
rect 391708 -23818 391776 -23762
rect 391832 -23818 391918 -23762
rect 391974 -23818 392048 -23762
rect 391708 -23904 392048 -23818
rect 391708 -23960 391776 -23904
rect 391832 -23960 391918 -23904
rect 391974 -23960 392048 -23904
rect 391708 -24046 392048 -23960
rect 391708 -24102 391776 -24046
rect 391832 -24102 391918 -24046
rect 391974 -24102 392048 -24046
rect 391708 -24188 392048 -24102
rect 391708 -24244 391776 -24188
rect 391832 -24244 391918 -24188
rect 391974 -24244 392048 -24188
rect 391708 -24330 392048 -24244
rect 391708 -24386 391776 -24330
rect 391832 -24386 391918 -24330
rect 391974 -24386 392048 -24330
rect 391708 -24472 392048 -24386
rect 391708 -24528 391776 -24472
rect 391832 -24528 391918 -24472
rect 391974 -24528 392048 -24472
rect 391708 -24614 392048 -24528
rect 391708 -24670 391776 -24614
rect 391832 -24670 391918 -24614
rect 391974 -24670 392048 -24614
rect 391708 -24756 392048 -24670
rect 391708 -24812 391776 -24756
rect 391832 -24812 391918 -24756
rect 391974 -24812 392048 -24756
rect 391708 -24898 392048 -24812
rect 391708 -24954 391776 -24898
rect 391832 -24954 391918 -24898
rect 391974 -24954 392048 -24898
rect 391708 -25040 392048 -24954
rect 391708 -25096 391776 -25040
rect 391832 -25096 391918 -25040
rect 391974 -25096 392048 -25040
rect 391708 -25182 392048 -25096
rect 391708 -25238 391776 -25182
rect 391832 -25238 391918 -25182
rect 391974 -25238 392048 -25182
rect 391708 -25324 392048 -25238
rect 391708 -25380 391776 -25324
rect 391832 -25380 391918 -25324
rect 391974 -25380 392048 -25324
rect 391708 -25466 392048 -25380
rect 391708 -25522 391776 -25466
rect 391832 -25522 391918 -25466
rect 391974 -25522 392048 -25466
rect 391708 -25532 392048 -25522
rect 392108 -13680 392448 -13670
rect 392108 -13736 392173 -13680
rect 392229 -13736 392315 -13680
rect 392371 -13736 392448 -13680
rect 392108 -13822 392448 -13736
rect 392108 -13878 392173 -13822
rect 392229 -13878 392315 -13822
rect 392371 -13878 392448 -13822
rect 392108 -13964 392448 -13878
rect 392108 -14020 392173 -13964
rect 392229 -14020 392315 -13964
rect 392371 -14020 392448 -13964
rect 392108 -14106 392448 -14020
rect 392108 -14162 392173 -14106
rect 392229 -14162 392315 -14106
rect 392371 -14162 392448 -14106
rect 392108 -14248 392448 -14162
rect 392108 -14304 392173 -14248
rect 392229 -14304 392315 -14248
rect 392371 -14304 392448 -14248
rect 392108 -14390 392448 -14304
rect 392108 -14446 392173 -14390
rect 392229 -14446 392315 -14390
rect 392371 -14446 392448 -14390
rect 392108 -14532 392448 -14446
rect 392108 -14588 392173 -14532
rect 392229 -14588 392315 -14532
rect 392371 -14588 392448 -14532
rect 392108 -14674 392448 -14588
rect 392108 -14730 392173 -14674
rect 392229 -14730 392315 -14674
rect 392371 -14730 392448 -14674
rect 392108 -14816 392448 -14730
rect 392108 -14872 392173 -14816
rect 392229 -14872 392315 -14816
rect 392371 -14872 392448 -14816
rect 392108 -14958 392448 -14872
rect 392108 -15014 392173 -14958
rect 392229 -15014 392315 -14958
rect 392371 -15014 392448 -14958
rect 392108 -15100 392448 -15014
rect 392108 -15156 392173 -15100
rect 392229 -15156 392315 -15100
rect 392371 -15156 392448 -15100
rect 392108 -15242 392448 -15156
rect 392108 -15298 392173 -15242
rect 392229 -15298 392315 -15242
rect 392371 -15298 392448 -15242
rect 392108 -15384 392448 -15298
rect 392108 -15440 392173 -15384
rect 392229 -15440 392315 -15384
rect 392371 -15440 392448 -15384
rect 392108 -15526 392448 -15440
rect 392108 -15582 392173 -15526
rect 392229 -15582 392315 -15526
rect 392371 -15582 392448 -15526
rect 392108 -15668 392448 -15582
rect 392108 -15724 392173 -15668
rect 392229 -15724 392315 -15668
rect 392371 -15724 392448 -15668
rect 392108 -15810 392448 -15724
rect 392108 -15866 392173 -15810
rect 392229 -15866 392315 -15810
rect 392371 -15866 392448 -15810
rect 392108 -15952 392448 -15866
rect 392108 -16008 392173 -15952
rect 392229 -16008 392315 -15952
rect 392371 -16008 392448 -15952
rect 392108 -16094 392448 -16008
rect 392108 -16150 392173 -16094
rect 392229 -16150 392315 -16094
rect 392371 -16150 392448 -16094
rect 392108 -16236 392448 -16150
rect 392108 -16292 392173 -16236
rect 392229 -16292 392315 -16236
rect 392371 -16292 392448 -16236
rect 392108 -16378 392448 -16292
rect 392108 -16434 392173 -16378
rect 392229 -16434 392315 -16378
rect 392371 -16434 392448 -16378
rect 392108 -16520 392448 -16434
rect 392108 -16576 392173 -16520
rect 392229 -16576 392315 -16520
rect 392371 -16576 392448 -16520
rect 392108 -16662 392448 -16576
rect 392108 -16718 392173 -16662
rect 392229 -16718 392315 -16662
rect 392371 -16718 392448 -16662
rect 392108 -16804 392448 -16718
rect 392108 -16860 392173 -16804
rect 392229 -16860 392315 -16804
rect 392371 -16860 392448 -16804
rect 392108 -16946 392448 -16860
rect 392108 -17002 392173 -16946
rect 392229 -17002 392315 -16946
rect 392371 -17002 392448 -16946
rect 392108 -17088 392448 -17002
rect 392108 -17144 392173 -17088
rect 392229 -17144 392315 -17088
rect 392371 -17144 392448 -17088
rect 392108 -17230 392448 -17144
rect 392108 -17286 392173 -17230
rect 392229 -17286 392315 -17230
rect 392371 -17286 392448 -17230
rect 392108 -17372 392448 -17286
rect 392108 -17428 392173 -17372
rect 392229 -17428 392315 -17372
rect 392371 -17428 392448 -17372
rect 392108 -17514 392448 -17428
rect 392108 -17570 392173 -17514
rect 392229 -17570 392315 -17514
rect 392371 -17570 392448 -17514
rect 392108 -17656 392448 -17570
rect 392108 -17712 392173 -17656
rect 392229 -17712 392315 -17656
rect 392371 -17712 392448 -17656
rect 392108 -17798 392448 -17712
rect 392108 -17854 392173 -17798
rect 392229 -17854 392315 -17798
rect 392371 -17854 392448 -17798
rect 392108 -17940 392448 -17854
rect 392108 -17996 392173 -17940
rect 392229 -17996 392315 -17940
rect 392371 -17996 392448 -17940
rect 392108 -18082 392448 -17996
rect 392108 -18138 392173 -18082
rect 392229 -18138 392315 -18082
rect 392371 -18138 392448 -18082
rect 392108 -18224 392448 -18138
rect 392108 -18280 392173 -18224
rect 392229 -18280 392315 -18224
rect 392371 -18280 392448 -18224
rect 392108 -18366 392448 -18280
rect 392108 -18422 392173 -18366
rect 392229 -18422 392315 -18366
rect 392371 -18422 392448 -18366
rect 392108 -18508 392448 -18422
rect 392108 -18564 392173 -18508
rect 392229 -18564 392315 -18508
rect 392371 -18564 392448 -18508
rect 392108 -18650 392448 -18564
rect 392108 -18706 392173 -18650
rect 392229 -18706 392315 -18650
rect 392371 -18706 392448 -18650
rect 392108 -18792 392448 -18706
rect 392108 -18848 392173 -18792
rect 392229 -18848 392315 -18792
rect 392371 -18848 392448 -18792
rect 392108 -18934 392448 -18848
rect 392108 -18990 392173 -18934
rect 392229 -18990 392315 -18934
rect 392371 -18990 392448 -18934
rect 392108 -19076 392448 -18990
rect 392108 -19132 392173 -19076
rect 392229 -19132 392315 -19076
rect 392371 -19132 392448 -19076
rect 392108 -19218 392448 -19132
rect 392108 -19274 392173 -19218
rect 392229 -19274 392315 -19218
rect 392371 -19274 392448 -19218
rect 392108 -19360 392448 -19274
rect 392108 -19416 392173 -19360
rect 392229 -19416 392315 -19360
rect 392371 -19416 392448 -19360
rect 392108 -19502 392448 -19416
rect 392108 -19558 392173 -19502
rect 392229 -19558 392315 -19502
rect 392371 -19558 392448 -19502
rect 392108 -19644 392448 -19558
rect 392108 -19700 392173 -19644
rect 392229 -19700 392315 -19644
rect 392371 -19700 392448 -19644
rect 392108 -19786 392448 -19700
rect 392108 -19842 392173 -19786
rect 392229 -19842 392315 -19786
rect 392371 -19842 392448 -19786
rect 392108 -19928 392448 -19842
rect 392108 -19984 392173 -19928
rect 392229 -19984 392315 -19928
rect 392371 -19984 392448 -19928
rect 392108 -20070 392448 -19984
rect 392108 -20126 392173 -20070
rect 392229 -20126 392315 -20070
rect 392371 -20126 392448 -20070
rect 392108 -20212 392448 -20126
rect 392108 -20268 392173 -20212
rect 392229 -20268 392315 -20212
rect 392371 -20268 392448 -20212
rect 392108 -20354 392448 -20268
rect 392108 -20410 392173 -20354
rect 392229 -20410 392315 -20354
rect 392371 -20410 392448 -20354
rect 392108 -20496 392448 -20410
rect 392108 -20552 392173 -20496
rect 392229 -20552 392315 -20496
rect 392371 -20552 392448 -20496
rect 392108 -20638 392448 -20552
rect 392108 -20694 392173 -20638
rect 392229 -20694 392315 -20638
rect 392371 -20694 392448 -20638
rect 392108 -20780 392448 -20694
rect 392108 -20836 392173 -20780
rect 392229 -20836 392315 -20780
rect 392371 -20836 392448 -20780
rect 392108 -20922 392448 -20836
rect 392108 -20978 392173 -20922
rect 392229 -20978 392315 -20922
rect 392371 -20978 392448 -20922
rect 392108 -21064 392448 -20978
rect 392108 -21120 392173 -21064
rect 392229 -21120 392315 -21064
rect 392371 -21120 392448 -21064
rect 392108 -21206 392448 -21120
rect 392108 -21262 392173 -21206
rect 392229 -21262 392315 -21206
rect 392371 -21262 392448 -21206
rect 392108 -21348 392448 -21262
rect 392108 -21404 392173 -21348
rect 392229 -21404 392315 -21348
rect 392371 -21404 392448 -21348
rect 392108 -21490 392448 -21404
rect 392108 -21546 392173 -21490
rect 392229 -21546 392315 -21490
rect 392371 -21546 392448 -21490
rect 392108 -21632 392448 -21546
rect 392108 -21688 392173 -21632
rect 392229 -21688 392315 -21632
rect 392371 -21688 392448 -21632
rect 392108 -21774 392448 -21688
rect 392108 -21830 392173 -21774
rect 392229 -21830 392315 -21774
rect 392371 -21830 392448 -21774
rect 392108 -21916 392448 -21830
rect 392108 -21972 392173 -21916
rect 392229 -21972 392315 -21916
rect 392371 -21972 392448 -21916
rect 392108 -22058 392448 -21972
rect 392108 -22114 392173 -22058
rect 392229 -22114 392315 -22058
rect 392371 -22114 392448 -22058
rect 392108 -22200 392448 -22114
rect 392108 -22256 392173 -22200
rect 392229 -22256 392315 -22200
rect 392371 -22256 392448 -22200
rect 392108 -22342 392448 -22256
rect 392108 -22398 392173 -22342
rect 392229 -22398 392315 -22342
rect 392371 -22398 392448 -22342
rect 392108 -22484 392448 -22398
rect 392108 -22540 392173 -22484
rect 392229 -22540 392315 -22484
rect 392371 -22540 392448 -22484
rect 392108 -22626 392448 -22540
rect 392108 -22682 392173 -22626
rect 392229 -22682 392315 -22626
rect 392371 -22682 392448 -22626
rect 392108 -22768 392448 -22682
rect 392108 -22824 392173 -22768
rect 392229 -22824 392315 -22768
rect 392371 -22824 392448 -22768
rect 392108 -22910 392448 -22824
rect 392108 -22966 392173 -22910
rect 392229 -22966 392315 -22910
rect 392371 -22966 392448 -22910
rect 392108 -23052 392448 -22966
rect 392108 -23108 392173 -23052
rect 392229 -23108 392315 -23052
rect 392371 -23108 392448 -23052
rect 392108 -23194 392448 -23108
rect 392108 -23250 392173 -23194
rect 392229 -23250 392315 -23194
rect 392371 -23250 392448 -23194
rect 392108 -23336 392448 -23250
rect 392108 -23392 392173 -23336
rect 392229 -23392 392315 -23336
rect 392371 -23392 392448 -23336
rect 392108 -23478 392448 -23392
rect 392108 -23534 392173 -23478
rect 392229 -23534 392315 -23478
rect 392371 -23534 392448 -23478
rect 392108 -23620 392448 -23534
rect 392108 -23676 392173 -23620
rect 392229 -23676 392315 -23620
rect 392371 -23676 392448 -23620
rect 392108 -23762 392448 -23676
rect 392108 -23818 392173 -23762
rect 392229 -23818 392315 -23762
rect 392371 -23818 392448 -23762
rect 392108 -23904 392448 -23818
rect 392108 -23960 392173 -23904
rect 392229 -23960 392315 -23904
rect 392371 -23960 392448 -23904
rect 392108 -24046 392448 -23960
rect 392108 -24102 392173 -24046
rect 392229 -24102 392315 -24046
rect 392371 -24102 392448 -24046
rect 392108 -24188 392448 -24102
rect 392108 -24244 392173 -24188
rect 392229 -24244 392315 -24188
rect 392371 -24244 392448 -24188
rect 392108 -24330 392448 -24244
rect 392108 -24386 392173 -24330
rect 392229 -24386 392315 -24330
rect 392371 -24386 392448 -24330
rect 392108 -24472 392448 -24386
rect 392108 -24528 392173 -24472
rect 392229 -24528 392315 -24472
rect 392371 -24528 392448 -24472
rect 392108 -24614 392448 -24528
rect 392108 -24670 392173 -24614
rect 392229 -24670 392315 -24614
rect 392371 -24670 392448 -24614
rect 392108 -24756 392448 -24670
rect 392108 -24812 392173 -24756
rect 392229 -24812 392315 -24756
rect 392371 -24812 392448 -24756
rect 392108 -24898 392448 -24812
rect 392108 -24954 392173 -24898
rect 392229 -24954 392315 -24898
rect 392371 -24954 392448 -24898
rect 392108 -25040 392448 -24954
rect 392108 -25096 392173 -25040
rect 392229 -25096 392315 -25040
rect 392371 -25096 392448 -25040
rect 392108 -25182 392448 -25096
rect 392108 -25238 392173 -25182
rect 392229 -25238 392315 -25182
rect 392371 -25238 392448 -25182
rect 392108 -25324 392448 -25238
rect 392108 -25380 392173 -25324
rect 392229 -25380 392315 -25324
rect 392371 -25380 392448 -25324
rect 392108 -25466 392448 -25380
rect 392108 -25522 392173 -25466
rect 392229 -25522 392315 -25466
rect 392371 -25522 392448 -25466
rect 392108 -25532 392448 -25522
rect 392508 -13680 392848 -13670
rect 392508 -13736 392578 -13680
rect 392634 -13736 392720 -13680
rect 392776 -13736 392848 -13680
rect 392508 -13822 392848 -13736
rect 392508 -13878 392578 -13822
rect 392634 -13878 392720 -13822
rect 392776 -13878 392848 -13822
rect 392508 -13964 392848 -13878
rect 392508 -14020 392578 -13964
rect 392634 -14020 392720 -13964
rect 392776 -14020 392848 -13964
rect 392508 -14106 392848 -14020
rect 392508 -14162 392578 -14106
rect 392634 -14162 392720 -14106
rect 392776 -14162 392848 -14106
rect 392508 -14248 392848 -14162
rect 392508 -14304 392578 -14248
rect 392634 -14304 392720 -14248
rect 392776 -14304 392848 -14248
rect 392508 -14390 392848 -14304
rect 392508 -14446 392578 -14390
rect 392634 -14446 392720 -14390
rect 392776 -14446 392848 -14390
rect 392508 -14532 392848 -14446
rect 392508 -14588 392578 -14532
rect 392634 -14588 392720 -14532
rect 392776 -14588 392848 -14532
rect 392508 -14674 392848 -14588
rect 392508 -14730 392578 -14674
rect 392634 -14730 392720 -14674
rect 392776 -14730 392848 -14674
rect 392508 -14816 392848 -14730
rect 392508 -14872 392578 -14816
rect 392634 -14872 392720 -14816
rect 392776 -14872 392848 -14816
rect 392508 -14958 392848 -14872
rect 392508 -15014 392578 -14958
rect 392634 -15014 392720 -14958
rect 392776 -15014 392848 -14958
rect 392508 -15100 392848 -15014
rect 392508 -15156 392578 -15100
rect 392634 -15156 392720 -15100
rect 392776 -15156 392848 -15100
rect 392508 -15242 392848 -15156
rect 392508 -15298 392578 -15242
rect 392634 -15298 392720 -15242
rect 392776 -15298 392848 -15242
rect 392508 -15384 392848 -15298
rect 392508 -15440 392578 -15384
rect 392634 -15440 392720 -15384
rect 392776 -15440 392848 -15384
rect 392508 -15526 392848 -15440
rect 392508 -15582 392578 -15526
rect 392634 -15582 392720 -15526
rect 392776 -15582 392848 -15526
rect 392508 -15668 392848 -15582
rect 392508 -15724 392578 -15668
rect 392634 -15724 392720 -15668
rect 392776 -15724 392848 -15668
rect 392508 -15810 392848 -15724
rect 392508 -15866 392578 -15810
rect 392634 -15866 392720 -15810
rect 392776 -15866 392848 -15810
rect 392508 -15952 392848 -15866
rect 392508 -16008 392578 -15952
rect 392634 -16008 392720 -15952
rect 392776 -16008 392848 -15952
rect 392508 -16094 392848 -16008
rect 392508 -16150 392578 -16094
rect 392634 -16150 392720 -16094
rect 392776 -16150 392848 -16094
rect 392508 -16236 392848 -16150
rect 392508 -16292 392578 -16236
rect 392634 -16292 392720 -16236
rect 392776 -16292 392848 -16236
rect 392508 -16378 392848 -16292
rect 392508 -16434 392578 -16378
rect 392634 -16434 392720 -16378
rect 392776 -16434 392848 -16378
rect 392508 -16520 392848 -16434
rect 392508 -16576 392578 -16520
rect 392634 -16576 392720 -16520
rect 392776 -16576 392848 -16520
rect 392508 -16662 392848 -16576
rect 392508 -16718 392578 -16662
rect 392634 -16718 392720 -16662
rect 392776 -16718 392848 -16662
rect 392508 -16804 392848 -16718
rect 392508 -16860 392578 -16804
rect 392634 -16860 392720 -16804
rect 392776 -16860 392848 -16804
rect 392508 -16946 392848 -16860
rect 392508 -17002 392578 -16946
rect 392634 -17002 392720 -16946
rect 392776 -17002 392848 -16946
rect 392508 -17088 392848 -17002
rect 392508 -17144 392578 -17088
rect 392634 -17144 392720 -17088
rect 392776 -17144 392848 -17088
rect 392508 -17230 392848 -17144
rect 392508 -17286 392578 -17230
rect 392634 -17286 392720 -17230
rect 392776 -17286 392848 -17230
rect 392508 -17372 392848 -17286
rect 392508 -17428 392578 -17372
rect 392634 -17428 392720 -17372
rect 392776 -17428 392848 -17372
rect 392508 -17514 392848 -17428
rect 392508 -17570 392578 -17514
rect 392634 -17570 392720 -17514
rect 392776 -17570 392848 -17514
rect 392508 -17656 392848 -17570
rect 392508 -17712 392578 -17656
rect 392634 -17712 392720 -17656
rect 392776 -17712 392848 -17656
rect 392508 -17798 392848 -17712
rect 392508 -17854 392578 -17798
rect 392634 -17854 392720 -17798
rect 392776 -17854 392848 -17798
rect 392508 -17940 392848 -17854
rect 392508 -17996 392578 -17940
rect 392634 -17996 392720 -17940
rect 392776 -17996 392848 -17940
rect 392508 -18082 392848 -17996
rect 392508 -18138 392578 -18082
rect 392634 -18138 392720 -18082
rect 392776 -18138 392848 -18082
rect 392508 -18224 392848 -18138
rect 392508 -18280 392578 -18224
rect 392634 -18280 392720 -18224
rect 392776 -18280 392848 -18224
rect 392508 -18366 392848 -18280
rect 392508 -18422 392578 -18366
rect 392634 -18422 392720 -18366
rect 392776 -18422 392848 -18366
rect 392508 -18508 392848 -18422
rect 392508 -18564 392578 -18508
rect 392634 -18564 392720 -18508
rect 392776 -18564 392848 -18508
rect 392508 -18650 392848 -18564
rect 392508 -18706 392578 -18650
rect 392634 -18706 392720 -18650
rect 392776 -18706 392848 -18650
rect 392508 -18792 392848 -18706
rect 392508 -18848 392578 -18792
rect 392634 -18848 392720 -18792
rect 392776 -18848 392848 -18792
rect 392508 -18934 392848 -18848
rect 392508 -18990 392578 -18934
rect 392634 -18990 392720 -18934
rect 392776 -18990 392848 -18934
rect 392508 -19076 392848 -18990
rect 392508 -19132 392578 -19076
rect 392634 -19132 392720 -19076
rect 392776 -19132 392848 -19076
rect 392508 -19218 392848 -19132
rect 392508 -19274 392578 -19218
rect 392634 -19274 392720 -19218
rect 392776 -19274 392848 -19218
rect 392508 -19360 392848 -19274
rect 392508 -19416 392578 -19360
rect 392634 -19416 392720 -19360
rect 392776 -19416 392848 -19360
rect 392508 -19502 392848 -19416
rect 392508 -19558 392578 -19502
rect 392634 -19558 392720 -19502
rect 392776 -19558 392848 -19502
rect 392508 -19644 392848 -19558
rect 392508 -19700 392578 -19644
rect 392634 -19700 392720 -19644
rect 392776 -19700 392848 -19644
rect 392508 -19786 392848 -19700
rect 392508 -19842 392578 -19786
rect 392634 -19842 392720 -19786
rect 392776 -19842 392848 -19786
rect 392508 -19928 392848 -19842
rect 392508 -19984 392578 -19928
rect 392634 -19984 392720 -19928
rect 392776 -19984 392848 -19928
rect 392508 -20070 392848 -19984
rect 392508 -20126 392578 -20070
rect 392634 -20126 392720 -20070
rect 392776 -20126 392848 -20070
rect 392508 -20212 392848 -20126
rect 392508 -20268 392578 -20212
rect 392634 -20268 392720 -20212
rect 392776 -20268 392848 -20212
rect 392508 -20354 392848 -20268
rect 392508 -20410 392578 -20354
rect 392634 -20410 392720 -20354
rect 392776 -20410 392848 -20354
rect 392508 -20496 392848 -20410
rect 392508 -20552 392578 -20496
rect 392634 -20552 392720 -20496
rect 392776 -20552 392848 -20496
rect 392508 -20638 392848 -20552
rect 392508 -20694 392578 -20638
rect 392634 -20694 392720 -20638
rect 392776 -20694 392848 -20638
rect 392508 -20780 392848 -20694
rect 392508 -20836 392578 -20780
rect 392634 -20836 392720 -20780
rect 392776 -20836 392848 -20780
rect 392508 -20922 392848 -20836
rect 392508 -20978 392578 -20922
rect 392634 -20978 392720 -20922
rect 392776 -20978 392848 -20922
rect 392508 -21064 392848 -20978
rect 392508 -21120 392578 -21064
rect 392634 -21120 392720 -21064
rect 392776 -21120 392848 -21064
rect 392508 -21206 392848 -21120
rect 392508 -21262 392578 -21206
rect 392634 -21262 392720 -21206
rect 392776 -21262 392848 -21206
rect 392508 -21348 392848 -21262
rect 392508 -21404 392578 -21348
rect 392634 -21404 392720 -21348
rect 392776 -21404 392848 -21348
rect 392508 -21490 392848 -21404
rect 392508 -21546 392578 -21490
rect 392634 -21546 392720 -21490
rect 392776 -21546 392848 -21490
rect 392508 -21632 392848 -21546
rect 392508 -21688 392578 -21632
rect 392634 -21688 392720 -21632
rect 392776 -21688 392848 -21632
rect 392508 -21774 392848 -21688
rect 392508 -21830 392578 -21774
rect 392634 -21830 392720 -21774
rect 392776 -21830 392848 -21774
rect 392508 -21916 392848 -21830
rect 392508 -21972 392578 -21916
rect 392634 -21972 392720 -21916
rect 392776 -21972 392848 -21916
rect 392508 -22058 392848 -21972
rect 392508 -22114 392578 -22058
rect 392634 -22114 392720 -22058
rect 392776 -22114 392848 -22058
rect 392508 -22200 392848 -22114
rect 392508 -22256 392578 -22200
rect 392634 -22256 392720 -22200
rect 392776 -22256 392848 -22200
rect 392508 -22342 392848 -22256
rect 392508 -22398 392578 -22342
rect 392634 -22398 392720 -22342
rect 392776 -22398 392848 -22342
rect 392508 -22484 392848 -22398
rect 392508 -22540 392578 -22484
rect 392634 -22540 392720 -22484
rect 392776 -22540 392848 -22484
rect 392508 -22626 392848 -22540
rect 392508 -22682 392578 -22626
rect 392634 -22682 392720 -22626
rect 392776 -22682 392848 -22626
rect 392508 -22768 392848 -22682
rect 392508 -22824 392578 -22768
rect 392634 -22824 392720 -22768
rect 392776 -22824 392848 -22768
rect 392508 -22910 392848 -22824
rect 392508 -22966 392578 -22910
rect 392634 -22966 392720 -22910
rect 392776 -22966 392848 -22910
rect 392508 -23052 392848 -22966
rect 392508 -23108 392578 -23052
rect 392634 -23108 392720 -23052
rect 392776 -23108 392848 -23052
rect 392508 -23194 392848 -23108
rect 392508 -23250 392578 -23194
rect 392634 -23250 392720 -23194
rect 392776 -23250 392848 -23194
rect 392508 -23336 392848 -23250
rect 392508 -23392 392578 -23336
rect 392634 -23392 392720 -23336
rect 392776 -23392 392848 -23336
rect 392508 -23478 392848 -23392
rect 392508 -23534 392578 -23478
rect 392634 -23534 392720 -23478
rect 392776 -23534 392848 -23478
rect 392508 -23620 392848 -23534
rect 392508 -23676 392578 -23620
rect 392634 -23676 392720 -23620
rect 392776 -23676 392848 -23620
rect 392508 -23762 392848 -23676
rect 392508 -23818 392578 -23762
rect 392634 -23818 392720 -23762
rect 392776 -23818 392848 -23762
rect 392508 -23904 392848 -23818
rect 392508 -23960 392578 -23904
rect 392634 -23960 392720 -23904
rect 392776 -23960 392848 -23904
rect 392508 -24046 392848 -23960
rect 392508 -24102 392578 -24046
rect 392634 -24102 392720 -24046
rect 392776 -24102 392848 -24046
rect 392508 -24188 392848 -24102
rect 392508 -24244 392578 -24188
rect 392634 -24244 392720 -24188
rect 392776 -24244 392848 -24188
rect 392508 -24330 392848 -24244
rect 392508 -24386 392578 -24330
rect 392634 -24386 392720 -24330
rect 392776 -24386 392848 -24330
rect 392508 -24472 392848 -24386
rect 392508 -24528 392578 -24472
rect 392634 -24528 392720 -24472
rect 392776 -24528 392848 -24472
rect 392508 -24614 392848 -24528
rect 392508 -24670 392578 -24614
rect 392634 -24670 392720 -24614
rect 392776 -24670 392848 -24614
rect 392508 -24756 392848 -24670
rect 392508 -24812 392578 -24756
rect 392634 -24812 392720 -24756
rect 392776 -24812 392848 -24756
rect 392508 -24898 392848 -24812
rect 392508 -24954 392578 -24898
rect 392634 -24954 392720 -24898
rect 392776 -24954 392848 -24898
rect 392508 -25040 392848 -24954
rect 392508 -25096 392578 -25040
rect 392634 -25096 392720 -25040
rect 392776 -25096 392848 -25040
rect 392508 -25182 392848 -25096
rect 392508 -25238 392578 -25182
rect 392634 -25238 392720 -25182
rect 392776 -25238 392848 -25182
rect 392508 -25324 392848 -25238
rect 392508 -25380 392578 -25324
rect 392634 -25380 392720 -25324
rect 392776 -25380 392848 -25324
rect 392508 -25466 392848 -25380
rect 392508 -25522 392578 -25466
rect 392634 -25522 392720 -25466
rect 392776 -25522 392848 -25466
rect 392508 -25532 392848 -25522
rect 392908 -13680 393248 -13670
rect 392908 -13736 392978 -13680
rect 393034 -13736 393120 -13680
rect 393176 -13736 393248 -13680
rect 392908 -13822 393248 -13736
rect 392908 -13878 392978 -13822
rect 393034 -13878 393120 -13822
rect 393176 -13878 393248 -13822
rect 392908 -13964 393248 -13878
rect 392908 -14020 392978 -13964
rect 393034 -14020 393120 -13964
rect 393176 -14020 393248 -13964
rect 392908 -14106 393248 -14020
rect 392908 -14162 392978 -14106
rect 393034 -14162 393120 -14106
rect 393176 -14162 393248 -14106
rect 392908 -14248 393248 -14162
rect 392908 -14304 392978 -14248
rect 393034 -14304 393120 -14248
rect 393176 -14304 393248 -14248
rect 392908 -14390 393248 -14304
rect 392908 -14446 392978 -14390
rect 393034 -14446 393120 -14390
rect 393176 -14446 393248 -14390
rect 392908 -14532 393248 -14446
rect 392908 -14588 392978 -14532
rect 393034 -14588 393120 -14532
rect 393176 -14588 393248 -14532
rect 392908 -14674 393248 -14588
rect 392908 -14730 392978 -14674
rect 393034 -14730 393120 -14674
rect 393176 -14730 393248 -14674
rect 392908 -14816 393248 -14730
rect 392908 -14872 392978 -14816
rect 393034 -14872 393120 -14816
rect 393176 -14872 393248 -14816
rect 392908 -14958 393248 -14872
rect 392908 -15014 392978 -14958
rect 393034 -15014 393120 -14958
rect 393176 -15014 393248 -14958
rect 392908 -15100 393248 -15014
rect 392908 -15156 392978 -15100
rect 393034 -15156 393120 -15100
rect 393176 -15156 393248 -15100
rect 392908 -15242 393248 -15156
rect 392908 -15298 392978 -15242
rect 393034 -15298 393120 -15242
rect 393176 -15298 393248 -15242
rect 392908 -15384 393248 -15298
rect 392908 -15440 392978 -15384
rect 393034 -15440 393120 -15384
rect 393176 -15440 393248 -15384
rect 392908 -15526 393248 -15440
rect 392908 -15582 392978 -15526
rect 393034 -15582 393120 -15526
rect 393176 -15582 393248 -15526
rect 392908 -15668 393248 -15582
rect 392908 -15724 392978 -15668
rect 393034 -15724 393120 -15668
rect 393176 -15724 393248 -15668
rect 392908 -15810 393248 -15724
rect 392908 -15866 392978 -15810
rect 393034 -15866 393120 -15810
rect 393176 -15866 393248 -15810
rect 392908 -15952 393248 -15866
rect 392908 -16008 392978 -15952
rect 393034 -16008 393120 -15952
rect 393176 -16008 393248 -15952
rect 392908 -16094 393248 -16008
rect 392908 -16150 392978 -16094
rect 393034 -16150 393120 -16094
rect 393176 -16150 393248 -16094
rect 392908 -16236 393248 -16150
rect 392908 -16292 392978 -16236
rect 393034 -16292 393120 -16236
rect 393176 -16292 393248 -16236
rect 392908 -16378 393248 -16292
rect 392908 -16434 392978 -16378
rect 393034 -16434 393120 -16378
rect 393176 -16434 393248 -16378
rect 392908 -16520 393248 -16434
rect 392908 -16576 392978 -16520
rect 393034 -16576 393120 -16520
rect 393176 -16576 393248 -16520
rect 392908 -16662 393248 -16576
rect 392908 -16718 392978 -16662
rect 393034 -16718 393120 -16662
rect 393176 -16718 393248 -16662
rect 392908 -16804 393248 -16718
rect 392908 -16860 392978 -16804
rect 393034 -16860 393120 -16804
rect 393176 -16860 393248 -16804
rect 392908 -16946 393248 -16860
rect 392908 -17002 392978 -16946
rect 393034 -17002 393120 -16946
rect 393176 -17002 393248 -16946
rect 392908 -17088 393248 -17002
rect 392908 -17144 392978 -17088
rect 393034 -17144 393120 -17088
rect 393176 -17144 393248 -17088
rect 392908 -17230 393248 -17144
rect 392908 -17286 392978 -17230
rect 393034 -17286 393120 -17230
rect 393176 -17286 393248 -17230
rect 392908 -17372 393248 -17286
rect 392908 -17428 392978 -17372
rect 393034 -17428 393120 -17372
rect 393176 -17428 393248 -17372
rect 392908 -17514 393248 -17428
rect 392908 -17570 392978 -17514
rect 393034 -17570 393120 -17514
rect 393176 -17570 393248 -17514
rect 392908 -17656 393248 -17570
rect 392908 -17712 392978 -17656
rect 393034 -17712 393120 -17656
rect 393176 -17712 393248 -17656
rect 392908 -17798 393248 -17712
rect 392908 -17854 392978 -17798
rect 393034 -17854 393120 -17798
rect 393176 -17854 393248 -17798
rect 392908 -17940 393248 -17854
rect 392908 -17996 392978 -17940
rect 393034 -17996 393120 -17940
rect 393176 -17996 393248 -17940
rect 392908 -18082 393248 -17996
rect 392908 -18138 392978 -18082
rect 393034 -18138 393120 -18082
rect 393176 -18138 393248 -18082
rect 392908 -18224 393248 -18138
rect 392908 -18280 392978 -18224
rect 393034 -18280 393120 -18224
rect 393176 -18280 393248 -18224
rect 392908 -18366 393248 -18280
rect 392908 -18422 392978 -18366
rect 393034 -18422 393120 -18366
rect 393176 -18422 393248 -18366
rect 392908 -18508 393248 -18422
rect 392908 -18564 392978 -18508
rect 393034 -18564 393120 -18508
rect 393176 -18564 393248 -18508
rect 392908 -18650 393248 -18564
rect 392908 -18706 392978 -18650
rect 393034 -18706 393120 -18650
rect 393176 -18706 393248 -18650
rect 392908 -18792 393248 -18706
rect 392908 -18848 392978 -18792
rect 393034 -18848 393120 -18792
rect 393176 -18848 393248 -18792
rect 392908 -18934 393248 -18848
rect 392908 -18990 392978 -18934
rect 393034 -18990 393120 -18934
rect 393176 -18990 393248 -18934
rect 392908 -19076 393248 -18990
rect 392908 -19132 392978 -19076
rect 393034 -19132 393120 -19076
rect 393176 -19132 393248 -19076
rect 392908 -19218 393248 -19132
rect 392908 -19274 392978 -19218
rect 393034 -19274 393120 -19218
rect 393176 -19274 393248 -19218
rect 392908 -19360 393248 -19274
rect 392908 -19416 392978 -19360
rect 393034 -19416 393120 -19360
rect 393176 -19416 393248 -19360
rect 392908 -19502 393248 -19416
rect 392908 -19558 392978 -19502
rect 393034 -19558 393120 -19502
rect 393176 -19558 393248 -19502
rect 392908 -19644 393248 -19558
rect 392908 -19700 392978 -19644
rect 393034 -19700 393120 -19644
rect 393176 -19700 393248 -19644
rect 392908 -19786 393248 -19700
rect 392908 -19842 392978 -19786
rect 393034 -19842 393120 -19786
rect 393176 -19842 393248 -19786
rect 392908 -19928 393248 -19842
rect 392908 -19984 392978 -19928
rect 393034 -19984 393120 -19928
rect 393176 -19984 393248 -19928
rect 392908 -20070 393248 -19984
rect 392908 -20126 392978 -20070
rect 393034 -20126 393120 -20070
rect 393176 -20126 393248 -20070
rect 392908 -20212 393248 -20126
rect 392908 -20268 392978 -20212
rect 393034 -20268 393120 -20212
rect 393176 -20268 393248 -20212
rect 392908 -20354 393248 -20268
rect 392908 -20410 392978 -20354
rect 393034 -20410 393120 -20354
rect 393176 -20410 393248 -20354
rect 392908 -20496 393248 -20410
rect 392908 -20552 392978 -20496
rect 393034 -20552 393120 -20496
rect 393176 -20552 393248 -20496
rect 392908 -20638 393248 -20552
rect 392908 -20694 392978 -20638
rect 393034 -20694 393120 -20638
rect 393176 -20694 393248 -20638
rect 392908 -20780 393248 -20694
rect 392908 -20836 392978 -20780
rect 393034 -20836 393120 -20780
rect 393176 -20836 393248 -20780
rect 392908 -20922 393248 -20836
rect 392908 -20978 392978 -20922
rect 393034 -20978 393120 -20922
rect 393176 -20978 393248 -20922
rect 392908 -21064 393248 -20978
rect 392908 -21120 392978 -21064
rect 393034 -21120 393120 -21064
rect 393176 -21120 393248 -21064
rect 392908 -21206 393248 -21120
rect 392908 -21262 392978 -21206
rect 393034 -21262 393120 -21206
rect 393176 -21262 393248 -21206
rect 392908 -21348 393248 -21262
rect 392908 -21404 392978 -21348
rect 393034 -21404 393120 -21348
rect 393176 -21404 393248 -21348
rect 392908 -21490 393248 -21404
rect 392908 -21546 392978 -21490
rect 393034 -21546 393120 -21490
rect 393176 -21546 393248 -21490
rect 392908 -21632 393248 -21546
rect 392908 -21688 392978 -21632
rect 393034 -21688 393120 -21632
rect 393176 -21688 393248 -21632
rect 392908 -21774 393248 -21688
rect 392908 -21830 392978 -21774
rect 393034 -21830 393120 -21774
rect 393176 -21830 393248 -21774
rect 392908 -21916 393248 -21830
rect 392908 -21972 392978 -21916
rect 393034 -21972 393120 -21916
rect 393176 -21972 393248 -21916
rect 392908 -22058 393248 -21972
rect 392908 -22114 392978 -22058
rect 393034 -22114 393120 -22058
rect 393176 -22114 393248 -22058
rect 392908 -22200 393248 -22114
rect 392908 -22256 392978 -22200
rect 393034 -22256 393120 -22200
rect 393176 -22256 393248 -22200
rect 392908 -22342 393248 -22256
rect 392908 -22398 392978 -22342
rect 393034 -22398 393120 -22342
rect 393176 -22398 393248 -22342
rect 392908 -22484 393248 -22398
rect 392908 -22540 392978 -22484
rect 393034 -22540 393120 -22484
rect 393176 -22540 393248 -22484
rect 392908 -22626 393248 -22540
rect 392908 -22682 392978 -22626
rect 393034 -22682 393120 -22626
rect 393176 -22682 393248 -22626
rect 392908 -22768 393248 -22682
rect 392908 -22824 392978 -22768
rect 393034 -22824 393120 -22768
rect 393176 -22824 393248 -22768
rect 392908 -22910 393248 -22824
rect 392908 -22966 392978 -22910
rect 393034 -22966 393120 -22910
rect 393176 -22966 393248 -22910
rect 392908 -23052 393248 -22966
rect 392908 -23108 392978 -23052
rect 393034 -23108 393120 -23052
rect 393176 -23108 393248 -23052
rect 392908 -23194 393248 -23108
rect 392908 -23250 392978 -23194
rect 393034 -23250 393120 -23194
rect 393176 -23250 393248 -23194
rect 392908 -23336 393248 -23250
rect 392908 -23392 392978 -23336
rect 393034 -23392 393120 -23336
rect 393176 -23392 393248 -23336
rect 392908 -23478 393248 -23392
rect 392908 -23534 392978 -23478
rect 393034 -23534 393120 -23478
rect 393176 -23534 393248 -23478
rect 392908 -23620 393248 -23534
rect 392908 -23676 392978 -23620
rect 393034 -23676 393120 -23620
rect 393176 -23676 393248 -23620
rect 392908 -23762 393248 -23676
rect 392908 -23818 392978 -23762
rect 393034 -23818 393120 -23762
rect 393176 -23818 393248 -23762
rect 392908 -23904 393248 -23818
rect 392908 -23960 392978 -23904
rect 393034 -23960 393120 -23904
rect 393176 -23960 393248 -23904
rect 392908 -24046 393248 -23960
rect 392908 -24102 392978 -24046
rect 393034 -24102 393120 -24046
rect 393176 -24102 393248 -24046
rect 392908 -24188 393248 -24102
rect 392908 -24244 392978 -24188
rect 393034 -24244 393120 -24188
rect 393176 -24244 393248 -24188
rect 392908 -24330 393248 -24244
rect 392908 -24386 392978 -24330
rect 393034 -24386 393120 -24330
rect 393176 -24386 393248 -24330
rect 392908 -24472 393248 -24386
rect 392908 -24528 392978 -24472
rect 393034 -24528 393120 -24472
rect 393176 -24528 393248 -24472
rect 392908 -24614 393248 -24528
rect 392908 -24670 392978 -24614
rect 393034 -24670 393120 -24614
rect 393176 -24670 393248 -24614
rect 392908 -24756 393248 -24670
rect 392908 -24812 392978 -24756
rect 393034 -24812 393120 -24756
rect 393176 -24812 393248 -24756
rect 392908 -24898 393248 -24812
rect 392908 -24954 392978 -24898
rect 393034 -24954 393120 -24898
rect 393176 -24954 393248 -24898
rect 392908 -25040 393248 -24954
rect 392908 -25096 392978 -25040
rect 393034 -25096 393120 -25040
rect 393176 -25096 393248 -25040
rect 392908 -25182 393248 -25096
rect 392908 -25238 392978 -25182
rect 393034 -25238 393120 -25182
rect 393176 -25238 393248 -25182
rect 392908 -25324 393248 -25238
rect 392908 -25380 392978 -25324
rect 393034 -25380 393120 -25324
rect 393176 -25380 393248 -25324
rect 392908 -25466 393248 -25380
rect 392908 -25522 392978 -25466
rect 393034 -25522 393120 -25466
rect 393176 -25522 393248 -25466
rect 392908 -25532 393248 -25522
rect 393308 -13680 393648 -13670
rect 393308 -13736 393383 -13680
rect 393439 -13736 393525 -13680
rect 393581 -13736 393648 -13680
rect 393308 -13822 393648 -13736
rect 393308 -13878 393383 -13822
rect 393439 -13878 393525 -13822
rect 393581 -13878 393648 -13822
rect 393308 -13964 393648 -13878
rect 393308 -14020 393383 -13964
rect 393439 -14020 393525 -13964
rect 393581 -14020 393648 -13964
rect 393308 -14106 393648 -14020
rect 393308 -14162 393383 -14106
rect 393439 -14162 393525 -14106
rect 393581 -14162 393648 -14106
rect 393308 -14248 393648 -14162
rect 393308 -14304 393383 -14248
rect 393439 -14304 393525 -14248
rect 393581 -14304 393648 -14248
rect 393308 -14390 393648 -14304
rect 393308 -14446 393383 -14390
rect 393439 -14446 393525 -14390
rect 393581 -14446 393648 -14390
rect 393308 -14532 393648 -14446
rect 393308 -14588 393383 -14532
rect 393439 -14588 393525 -14532
rect 393581 -14588 393648 -14532
rect 393308 -14674 393648 -14588
rect 393308 -14730 393383 -14674
rect 393439 -14730 393525 -14674
rect 393581 -14730 393648 -14674
rect 393308 -14816 393648 -14730
rect 393308 -14872 393383 -14816
rect 393439 -14872 393525 -14816
rect 393581 -14872 393648 -14816
rect 393308 -14958 393648 -14872
rect 393308 -15014 393383 -14958
rect 393439 -15014 393525 -14958
rect 393581 -15014 393648 -14958
rect 393308 -15100 393648 -15014
rect 393308 -15156 393383 -15100
rect 393439 -15156 393525 -15100
rect 393581 -15156 393648 -15100
rect 393308 -15242 393648 -15156
rect 393308 -15298 393383 -15242
rect 393439 -15298 393525 -15242
rect 393581 -15298 393648 -15242
rect 393308 -15384 393648 -15298
rect 393308 -15440 393383 -15384
rect 393439 -15440 393525 -15384
rect 393581 -15440 393648 -15384
rect 393308 -15526 393648 -15440
rect 393308 -15582 393383 -15526
rect 393439 -15582 393525 -15526
rect 393581 -15582 393648 -15526
rect 393308 -15668 393648 -15582
rect 393308 -15724 393383 -15668
rect 393439 -15724 393525 -15668
rect 393581 -15724 393648 -15668
rect 393308 -15810 393648 -15724
rect 393308 -15866 393383 -15810
rect 393439 -15866 393525 -15810
rect 393581 -15866 393648 -15810
rect 393308 -15952 393648 -15866
rect 393308 -16008 393383 -15952
rect 393439 -16008 393525 -15952
rect 393581 -16008 393648 -15952
rect 393308 -16094 393648 -16008
rect 393308 -16150 393383 -16094
rect 393439 -16150 393525 -16094
rect 393581 -16150 393648 -16094
rect 393308 -16236 393648 -16150
rect 393308 -16292 393383 -16236
rect 393439 -16292 393525 -16236
rect 393581 -16292 393648 -16236
rect 393308 -16378 393648 -16292
rect 393308 -16434 393383 -16378
rect 393439 -16434 393525 -16378
rect 393581 -16434 393648 -16378
rect 393308 -16520 393648 -16434
rect 393308 -16576 393383 -16520
rect 393439 -16576 393525 -16520
rect 393581 -16576 393648 -16520
rect 393308 -16662 393648 -16576
rect 393308 -16718 393383 -16662
rect 393439 -16718 393525 -16662
rect 393581 -16718 393648 -16662
rect 393308 -16804 393648 -16718
rect 393308 -16860 393383 -16804
rect 393439 -16860 393525 -16804
rect 393581 -16860 393648 -16804
rect 393308 -16946 393648 -16860
rect 393308 -17002 393383 -16946
rect 393439 -17002 393525 -16946
rect 393581 -17002 393648 -16946
rect 393308 -17088 393648 -17002
rect 393308 -17144 393383 -17088
rect 393439 -17144 393525 -17088
rect 393581 -17144 393648 -17088
rect 393308 -17230 393648 -17144
rect 393308 -17286 393383 -17230
rect 393439 -17286 393525 -17230
rect 393581 -17286 393648 -17230
rect 393308 -17372 393648 -17286
rect 393308 -17428 393383 -17372
rect 393439 -17428 393525 -17372
rect 393581 -17428 393648 -17372
rect 393308 -17514 393648 -17428
rect 393308 -17570 393383 -17514
rect 393439 -17570 393525 -17514
rect 393581 -17570 393648 -17514
rect 393308 -17656 393648 -17570
rect 393308 -17712 393383 -17656
rect 393439 -17712 393525 -17656
rect 393581 -17712 393648 -17656
rect 393308 -17798 393648 -17712
rect 393308 -17854 393383 -17798
rect 393439 -17854 393525 -17798
rect 393581 -17854 393648 -17798
rect 393308 -17940 393648 -17854
rect 393308 -17996 393383 -17940
rect 393439 -17996 393525 -17940
rect 393581 -17996 393648 -17940
rect 393308 -18082 393648 -17996
rect 393308 -18138 393383 -18082
rect 393439 -18138 393525 -18082
rect 393581 -18138 393648 -18082
rect 393308 -18224 393648 -18138
rect 393308 -18280 393383 -18224
rect 393439 -18280 393525 -18224
rect 393581 -18280 393648 -18224
rect 393308 -18366 393648 -18280
rect 393308 -18422 393383 -18366
rect 393439 -18422 393525 -18366
rect 393581 -18422 393648 -18366
rect 393308 -18508 393648 -18422
rect 393308 -18564 393383 -18508
rect 393439 -18564 393525 -18508
rect 393581 -18564 393648 -18508
rect 393308 -18650 393648 -18564
rect 393308 -18706 393383 -18650
rect 393439 -18706 393525 -18650
rect 393581 -18706 393648 -18650
rect 393308 -18792 393648 -18706
rect 393308 -18848 393383 -18792
rect 393439 -18848 393525 -18792
rect 393581 -18848 393648 -18792
rect 393308 -18934 393648 -18848
rect 393308 -18990 393383 -18934
rect 393439 -18990 393525 -18934
rect 393581 -18990 393648 -18934
rect 393308 -19076 393648 -18990
rect 393308 -19132 393383 -19076
rect 393439 -19132 393525 -19076
rect 393581 -19132 393648 -19076
rect 393308 -19218 393648 -19132
rect 393308 -19274 393383 -19218
rect 393439 -19274 393525 -19218
rect 393581 -19274 393648 -19218
rect 393308 -19360 393648 -19274
rect 393308 -19416 393383 -19360
rect 393439 -19416 393525 -19360
rect 393581 -19416 393648 -19360
rect 393308 -19502 393648 -19416
rect 393308 -19558 393383 -19502
rect 393439 -19558 393525 -19502
rect 393581 -19558 393648 -19502
rect 393308 -19644 393648 -19558
rect 393308 -19700 393383 -19644
rect 393439 -19700 393525 -19644
rect 393581 -19700 393648 -19644
rect 393308 -19786 393648 -19700
rect 393308 -19842 393383 -19786
rect 393439 -19842 393525 -19786
rect 393581 -19842 393648 -19786
rect 393308 -19928 393648 -19842
rect 393308 -19984 393383 -19928
rect 393439 -19984 393525 -19928
rect 393581 -19984 393648 -19928
rect 393308 -20070 393648 -19984
rect 393308 -20126 393383 -20070
rect 393439 -20126 393525 -20070
rect 393581 -20126 393648 -20070
rect 393308 -20212 393648 -20126
rect 393308 -20268 393383 -20212
rect 393439 -20268 393525 -20212
rect 393581 -20268 393648 -20212
rect 393308 -20354 393648 -20268
rect 393308 -20410 393383 -20354
rect 393439 -20410 393525 -20354
rect 393581 -20410 393648 -20354
rect 393308 -20496 393648 -20410
rect 393308 -20552 393383 -20496
rect 393439 -20552 393525 -20496
rect 393581 -20552 393648 -20496
rect 393308 -20638 393648 -20552
rect 393308 -20694 393383 -20638
rect 393439 -20694 393525 -20638
rect 393581 -20694 393648 -20638
rect 393308 -20780 393648 -20694
rect 393308 -20836 393383 -20780
rect 393439 -20836 393525 -20780
rect 393581 -20836 393648 -20780
rect 393308 -20922 393648 -20836
rect 393308 -20978 393383 -20922
rect 393439 -20978 393525 -20922
rect 393581 -20978 393648 -20922
rect 393308 -21064 393648 -20978
rect 393308 -21120 393383 -21064
rect 393439 -21120 393525 -21064
rect 393581 -21120 393648 -21064
rect 393308 -21206 393648 -21120
rect 393308 -21262 393383 -21206
rect 393439 -21262 393525 -21206
rect 393581 -21262 393648 -21206
rect 393308 -21348 393648 -21262
rect 393308 -21404 393383 -21348
rect 393439 -21404 393525 -21348
rect 393581 -21404 393648 -21348
rect 393308 -21490 393648 -21404
rect 393308 -21546 393383 -21490
rect 393439 -21546 393525 -21490
rect 393581 -21546 393648 -21490
rect 393308 -21632 393648 -21546
rect 393308 -21688 393383 -21632
rect 393439 -21688 393525 -21632
rect 393581 -21688 393648 -21632
rect 393308 -21774 393648 -21688
rect 393308 -21830 393383 -21774
rect 393439 -21830 393525 -21774
rect 393581 -21830 393648 -21774
rect 393308 -21916 393648 -21830
rect 393308 -21972 393383 -21916
rect 393439 -21972 393525 -21916
rect 393581 -21972 393648 -21916
rect 393308 -22058 393648 -21972
rect 393308 -22114 393383 -22058
rect 393439 -22114 393525 -22058
rect 393581 -22114 393648 -22058
rect 393308 -22200 393648 -22114
rect 393308 -22256 393383 -22200
rect 393439 -22256 393525 -22200
rect 393581 -22256 393648 -22200
rect 393308 -22342 393648 -22256
rect 393308 -22398 393383 -22342
rect 393439 -22398 393525 -22342
rect 393581 -22398 393648 -22342
rect 393308 -22484 393648 -22398
rect 393308 -22540 393383 -22484
rect 393439 -22540 393525 -22484
rect 393581 -22540 393648 -22484
rect 393308 -22626 393648 -22540
rect 393308 -22682 393383 -22626
rect 393439 -22682 393525 -22626
rect 393581 -22682 393648 -22626
rect 393308 -22768 393648 -22682
rect 393308 -22824 393383 -22768
rect 393439 -22824 393525 -22768
rect 393581 -22824 393648 -22768
rect 393308 -22910 393648 -22824
rect 393308 -22966 393383 -22910
rect 393439 -22966 393525 -22910
rect 393581 -22966 393648 -22910
rect 393308 -23052 393648 -22966
rect 393308 -23108 393383 -23052
rect 393439 -23108 393525 -23052
rect 393581 -23108 393648 -23052
rect 393308 -23194 393648 -23108
rect 393308 -23250 393383 -23194
rect 393439 -23250 393525 -23194
rect 393581 -23250 393648 -23194
rect 393308 -23336 393648 -23250
rect 393308 -23392 393383 -23336
rect 393439 -23392 393525 -23336
rect 393581 -23392 393648 -23336
rect 393308 -23478 393648 -23392
rect 393308 -23534 393383 -23478
rect 393439 -23534 393525 -23478
rect 393581 -23534 393648 -23478
rect 393308 -23620 393648 -23534
rect 393308 -23676 393383 -23620
rect 393439 -23676 393525 -23620
rect 393581 -23676 393648 -23620
rect 393308 -23762 393648 -23676
rect 393308 -23818 393383 -23762
rect 393439 -23818 393525 -23762
rect 393581 -23818 393648 -23762
rect 393308 -23904 393648 -23818
rect 393308 -23960 393383 -23904
rect 393439 -23960 393525 -23904
rect 393581 -23960 393648 -23904
rect 393308 -24046 393648 -23960
rect 393308 -24102 393383 -24046
rect 393439 -24102 393525 -24046
rect 393581 -24102 393648 -24046
rect 393308 -24188 393648 -24102
rect 393308 -24244 393383 -24188
rect 393439 -24244 393525 -24188
rect 393581 -24244 393648 -24188
rect 393308 -24330 393648 -24244
rect 393308 -24386 393383 -24330
rect 393439 -24386 393525 -24330
rect 393581 -24386 393648 -24330
rect 393308 -24472 393648 -24386
rect 393308 -24528 393383 -24472
rect 393439 -24528 393525 -24472
rect 393581 -24528 393648 -24472
rect 393308 -24614 393648 -24528
rect 393308 -24670 393383 -24614
rect 393439 -24670 393525 -24614
rect 393581 -24670 393648 -24614
rect 393308 -24756 393648 -24670
rect 393308 -24812 393383 -24756
rect 393439 -24812 393525 -24756
rect 393581 -24812 393648 -24756
rect 393308 -24898 393648 -24812
rect 393308 -24954 393383 -24898
rect 393439 -24954 393525 -24898
rect 393581 -24954 393648 -24898
rect 393308 -25040 393648 -24954
rect 393308 -25096 393383 -25040
rect 393439 -25096 393525 -25040
rect 393581 -25096 393648 -25040
rect 393308 -25182 393648 -25096
rect 393308 -25238 393383 -25182
rect 393439 -25238 393525 -25182
rect 393581 -25238 393648 -25182
rect 393308 -25324 393648 -25238
rect 393308 -25380 393383 -25324
rect 393439 -25380 393525 -25324
rect 393581 -25380 393648 -25324
rect 393308 -25466 393648 -25380
rect 393308 -25522 393383 -25466
rect 393439 -25522 393525 -25466
rect 393581 -25522 393648 -25466
rect 393308 -25532 393648 -25522
rect 393708 -13680 394048 -13670
rect 393708 -13736 393780 -13680
rect 393836 -13736 393922 -13680
rect 393978 -13736 394048 -13680
rect 393708 -13822 394048 -13736
rect 393708 -13878 393780 -13822
rect 393836 -13878 393922 -13822
rect 393978 -13878 394048 -13822
rect 393708 -13964 394048 -13878
rect 393708 -14020 393780 -13964
rect 393836 -14020 393922 -13964
rect 393978 -14020 394048 -13964
rect 393708 -14106 394048 -14020
rect 393708 -14162 393780 -14106
rect 393836 -14162 393922 -14106
rect 393978 -14162 394048 -14106
rect 393708 -14248 394048 -14162
rect 393708 -14304 393780 -14248
rect 393836 -14304 393922 -14248
rect 393978 -14304 394048 -14248
rect 393708 -14390 394048 -14304
rect 393708 -14446 393780 -14390
rect 393836 -14446 393922 -14390
rect 393978 -14446 394048 -14390
rect 393708 -14532 394048 -14446
rect 393708 -14588 393780 -14532
rect 393836 -14588 393922 -14532
rect 393978 -14588 394048 -14532
rect 393708 -14674 394048 -14588
rect 393708 -14730 393780 -14674
rect 393836 -14730 393922 -14674
rect 393978 -14730 394048 -14674
rect 393708 -14816 394048 -14730
rect 393708 -14872 393780 -14816
rect 393836 -14872 393922 -14816
rect 393978 -14872 394048 -14816
rect 393708 -14958 394048 -14872
rect 393708 -15014 393780 -14958
rect 393836 -15014 393922 -14958
rect 393978 -15014 394048 -14958
rect 393708 -15100 394048 -15014
rect 393708 -15156 393780 -15100
rect 393836 -15156 393922 -15100
rect 393978 -15156 394048 -15100
rect 393708 -15242 394048 -15156
rect 393708 -15298 393780 -15242
rect 393836 -15298 393922 -15242
rect 393978 -15298 394048 -15242
rect 393708 -15384 394048 -15298
rect 393708 -15440 393780 -15384
rect 393836 -15440 393922 -15384
rect 393978 -15440 394048 -15384
rect 393708 -15526 394048 -15440
rect 393708 -15582 393780 -15526
rect 393836 -15582 393922 -15526
rect 393978 -15582 394048 -15526
rect 393708 -15668 394048 -15582
rect 393708 -15724 393780 -15668
rect 393836 -15724 393922 -15668
rect 393978 -15724 394048 -15668
rect 393708 -15810 394048 -15724
rect 393708 -15866 393780 -15810
rect 393836 -15866 393922 -15810
rect 393978 -15866 394048 -15810
rect 393708 -15952 394048 -15866
rect 393708 -16008 393780 -15952
rect 393836 -16008 393922 -15952
rect 393978 -16008 394048 -15952
rect 393708 -16094 394048 -16008
rect 393708 -16150 393780 -16094
rect 393836 -16150 393922 -16094
rect 393978 -16150 394048 -16094
rect 393708 -16236 394048 -16150
rect 393708 -16292 393780 -16236
rect 393836 -16292 393922 -16236
rect 393978 -16292 394048 -16236
rect 393708 -16378 394048 -16292
rect 393708 -16434 393780 -16378
rect 393836 -16434 393922 -16378
rect 393978 -16434 394048 -16378
rect 393708 -16520 394048 -16434
rect 393708 -16576 393780 -16520
rect 393836 -16576 393922 -16520
rect 393978 -16576 394048 -16520
rect 393708 -16662 394048 -16576
rect 393708 -16718 393780 -16662
rect 393836 -16718 393922 -16662
rect 393978 -16718 394048 -16662
rect 393708 -16804 394048 -16718
rect 393708 -16860 393780 -16804
rect 393836 -16860 393922 -16804
rect 393978 -16860 394048 -16804
rect 393708 -16946 394048 -16860
rect 393708 -17002 393780 -16946
rect 393836 -17002 393922 -16946
rect 393978 -17002 394048 -16946
rect 393708 -17088 394048 -17002
rect 393708 -17144 393780 -17088
rect 393836 -17144 393922 -17088
rect 393978 -17144 394048 -17088
rect 393708 -17230 394048 -17144
rect 393708 -17286 393780 -17230
rect 393836 -17286 393922 -17230
rect 393978 -17286 394048 -17230
rect 393708 -17372 394048 -17286
rect 393708 -17428 393780 -17372
rect 393836 -17428 393922 -17372
rect 393978 -17428 394048 -17372
rect 393708 -17514 394048 -17428
rect 393708 -17570 393780 -17514
rect 393836 -17570 393922 -17514
rect 393978 -17570 394048 -17514
rect 393708 -17656 394048 -17570
rect 393708 -17712 393780 -17656
rect 393836 -17712 393922 -17656
rect 393978 -17712 394048 -17656
rect 393708 -17798 394048 -17712
rect 393708 -17854 393780 -17798
rect 393836 -17854 393922 -17798
rect 393978 -17854 394048 -17798
rect 393708 -17940 394048 -17854
rect 393708 -17996 393780 -17940
rect 393836 -17996 393922 -17940
rect 393978 -17996 394048 -17940
rect 393708 -18082 394048 -17996
rect 393708 -18138 393780 -18082
rect 393836 -18138 393922 -18082
rect 393978 -18138 394048 -18082
rect 393708 -18224 394048 -18138
rect 393708 -18280 393780 -18224
rect 393836 -18280 393922 -18224
rect 393978 -18280 394048 -18224
rect 393708 -18366 394048 -18280
rect 393708 -18422 393780 -18366
rect 393836 -18422 393922 -18366
rect 393978 -18422 394048 -18366
rect 393708 -18508 394048 -18422
rect 393708 -18564 393780 -18508
rect 393836 -18564 393922 -18508
rect 393978 -18564 394048 -18508
rect 393708 -18650 394048 -18564
rect 393708 -18706 393780 -18650
rect 393836 -18706 393922 -18650
rect 393978 -18706 394048 -18650
rect 393708 -18792 394048 -18706
rect 393708 -18848 393780 -18792
rect 393836 -18848 393922 -18792
rect 393978 -18848 394048 -18792
rect 393708 -18934 394048 -18848
rect 393708 -18990 393780 -18934
rect 393836 -18990 393922 -18934
rect 393978 -18990 394048 -18934
rect 393708 -19076 394048 -18990
rect 393708 -19132 393780 -19076
rect 393836 -19132 393922 -19076
rect 393978 -19132 394048 -19076
rect 393708 -19218 394048 -19132
rect 393708 -19274 393780 -19218
rect 393836 -19274 393922 -19218
rect 393978 -19274 394048 -19218
rect 393708 -19360 394048 -19274
rect 393708 -19416 393780 -19360
rect 393836 -19416 393922 -19360
rect 393978 -19416 394048 -19360
rect 393708 -19502 394048 -19416
rect 393708 -19558 393780 -19502
rect 393836 -19558 393922 -19502
rect 393978 -19558 394048 -19502
rect 393708 -19644 394048 -19558
rect 393708 -19700 393780 -19644
rect 393836 -19700 393922 -19644
rect 393978 -19700 394048 -19644
rect 393708 -19786 394048 -19700
rect 393708 -19842 393780 -19786
rect 393836 -19842 393922 -19786
rect 393978 -19842 394048 -19786
rect 393708 -19928 394048 -19842
rect 393708 -19984 393780 -19928
rect 393836 -19984 393922 -19928
rect 393978 -19984 394048 -19928
rect 393708 -20070 394048 -19984
rect 393708 -20126 393780 -20070
rect 393836 -20126 393922 -20070
rect 393978 -20126 394048 -20070
rect 393708 -20212 394048 -20126
rect 393708 -20268 393780 -20212
rect 393836 -20268 393922 -20212
rect 393978 -20268 394048 -20212
rect 393708 -20354 394048 -20268
rect 393708 -20410 393780 -20354
rect 393836 -20410 393922 -20354
rect 393978 -20410 394048 -20354
rect 393708 -20496 394048 -20410
rect 393708 -20552 393780 -20496
rect 393836 -20552 393922 -20496
rect 393978 -20552 394048 -20496
rect 393708 -20638 394048 -20552
rect 393708 -20694 393780 -20638
rect 393836 -20694 393922 -20638
rect 393978 -20694 394048 -20638
rect 393708 -20780 394048 -20694
rect 393708 -20836 393780 -20780
rect 393836 -20836 393922 -20780
rect 393978 -20836 394048 -20780
rect 393708 -20922 394048 -20836
rect 393708 -20978 393780 -20922
rect 393836 -20978 393922 -20922
rect 393978 -20978 394048 -20922
rect 393708 -21064 394048 -20978
rect 393708 -21120 393780 -21064
rect 393836 -21120 393922 -21064
rect 393978 -21120 394048 -21064
rect 393708 -21206 394048 -21120
rect 393708 -21262 393780 -21206
rect 393836 -21262 393922 -21206
rect 393978 -21262 394048 -21206
rect 393708 -21348 394048 -21262
rect 393708 -21404 393780 -21348
rect 393836 -21404 393922 -21348
rect 393978 -21404 394048 -21348
rect 393708 -21490 394048 -21404
rect 393708 -21546 393780 -21490
rect 393836 -21546 393922 -21490
rect 393978 -21546 394048 -21490
rect 393708 -21632 394048 -21546
rect 393708 -21688 393780 -21632
rect 393836 -21688 393922 -21632
rect 393978 -21688 394048 -21632
rect 393708 -21774 394048 -21688
rect 393708 -21830 393780 -21774
rect 393836 -21830 393922 -21774
rect 393978 -21830 394048 -21774
rect 393708 -21916 394048 -21830
rect 393708 -21972 393780 -21916
rect 393836 -21972 393922 -21916
rect 393978 -21972 394048 -21916
rect 393708 -22058 394048 -21972
rect 393708 -22114 393780 -22058
rect 393836 -22114 393922 -22058
rect 393978 -22114 394048 -22058
rect 393708 -22200 394048 -22114
rect 393708 -22256 393780 -22200
rect 393836 -22256 393922 -22200
rect 393978 -22256 394048 -22200
rect 393708 -22342 394048 -22256
rect 393708 -22398 393780 -22342
rect 393836 -22398 393922 -22342
rect 393978 -22398 394048 -22342
rect 393708 -22484 394048 -22398
rect 393708 -22540 393780 -22484
rect 393836 -22540 393922 -22484
rect 393978 -22540 394048 -22484
rect 393708 -22626 394048 -22540
rect 393708 -22682 393780 -22626
rect 393836 -22682 393922 -22626
rect 393978 -22682 394048 -22626
rect 393708 -22768 394048 -22682
rect 393708 -22824 393780 -22768
rect 393836 -22824 393922 -22768
rect 393978 -22824 394048 -22768
rect 393708 -22910 394048 -22824
rect 393708 -22966 393780 -22910
rect 393836 -22966 393922 -22910
rect 393978 -22966 394048 -22910
rect 393708 -23052 394048 -22966
rect 393708 -23108 393780 -23052
rect 393836 -23108 393922 -23052
rect 393978 -23108 394048 -23052
rect 393708 -23194 394048 -23108
rect 393708 -23250 393780 -23194
rect 393836 -23250 393922 -23194
rect 393978 -23250 394048 -23194
rect 393708 -23336 394048 -23250
rect 393708 -23392 393780 -23336
rect 393836 -23392 393922 -23336
rect 393978 -23392 394048 -23336
rect 393708 -23478 394048 -23392
rect 393708 -23534 393780 -23478
rect 393836 -23534 393922 -23478
rect 393978 -23534 394048 -23478
rect 393708 -23620 394048 -23534
rect 393708 -23676 393780 -23620
rect 393836 -23676 393922 -23620
rect 393978 -23676 394048 -23620
rect 393708 -23762 394048 -23676
rect 393708 -23818 393780 -23762
rect 393836 -23818 393922 -23762
rect 393978 -23818 394048 -23762
rect 393708 -23904 394048 -23818
rect 393708 -23960 393780 -23904
rect 393836 -23960 393922 -23904
rect 393978 -23960 394048 -23904
rect 393708 -24046 394048 -23960
rect 393708 -24102 393780 -24046
rect 393836 -24102 393922 -24046
rect 393978 -24102 394048 -24046
rect 393708 -24188 394048 -24102
rect 393708 -24244 393780 -24188
rect 393836 -24244 393922 -24188
rect 393978 -24244 394048 -24188
rect 393708 -24330 394048 -24244
rect 393708 -24386 393780 -24330
rect 393836 -24386 393922 -24330
rect 393978 -24386 394048 -24330
rect 393708 -24472 394048 -24386
rect 393708 -24528 393780 -24472
rect 393836 -24528 393922 -24472
rect 393978 -24528 394048 -24472
rect 393708 -24614 394048 -24528
rect 393708 -24670 393780 -24614
rect 393836 -24670 393922 -24614
rect 393978 -24670 394048 -24614
rect 393708 -24756 394048 -24670
rect 393708 -24812 393780 -24756
rect 393836 -24812 393922 -24756
rect 393978 -24812 394048 -24756
rect 393708 -24898 394048 -24812
rect 393708 -24954 393780 -24898
rect 393836 -24954 393922 -24898
rect 393978 -24954 394048 -24898
rect 393708 -25040 394048 -24954
rect 393708 -25096 393780 -25040
rect 393836 -25096 393922 -25040
rect 393978 -25096 394048 -25040
rect 393708 -25182 394048 -25096
rect 393708 -25238 393780 -25182
rect 393836 -25238 393922 -25182
rect 393978 -25238 394048 -25182
rect 393708 -25324 394048 -25238
rect 393708 -25380 393780 -25324
rect 393836 -25380 393922 -25324
rect 393978 -25380 394048 -25324
rect 393708 -25466 394048 -25380
rect 393708 -25522 393780 -25466
rect 393836 -25522 393922 -25466
rect 393978 -25522 394048 -25466
rect 393708 -25532 394048 -25522
rect 394108 -13680 394448 -13670
rect 394108 -13736 394177 -13680
rect 394233 -13736 394319 -13680
rect 394375 -13736 394448 -13680
rect 394108 -13822 394448 -13736
rect 394108 -13878 394177 -13822
rect 394233 -13878 394319 -13822
rect 394375 -13878 394448 -13822
rect 394108 -13964 394448 -13878
rect 394108 -14020 394177 -13964
rect 394233 -14020 394319 -13964
rect 394375 -14020 394448 -13964
rect 394108 -14106 394448 -14020
rect 394108 -14162 394177 -14106
rect 394233 -14162 394319 -14106
rect 394375 -14162 394448 -14106
rect 394108 -14248 394448 -14162
rect 394108 -14304 394177 -14248
rect 394233 -14304 394319 -14248
rect 394375 -14304 394448 -14248
rect 394108 -14390 394448 -14304
rect 394108 -14446 394177 -14390
rect 394233 -14446 394319 -14390
rect 394375 -14446 394448 -14390
rect 394108 -14532 394448 -14446
rect 394108 -14588 394177 -14532
rect 394233 -14588 394319 -14532
rect 394375 -14588 394448 -14532
rect 394108 -14674 394448 -14588
rect 394108 -14730 394177 -14674
rect 394233 -14730 394319 -14674
rect 394375 -14730 394448 -14674
rect 394108 -14816 394448 -14730
rect 394108 -14872 394177 -14816
rect 394233 -14872 394319 -14816
rect 394375 -14872 394448 -14816
rect 394108 -14958 394448 -14872
rect 394108 -15014 394177 -14958
rect 394233 -15014 394319 -14958
rect 394375 -15014 394448 -14958
rect 394108 -15100 394448 -15014
rect 394108 -15156 394177 -15100
rect 394233 -15156 394319 -15100
rect 394375 -15156 394448 -15100
rect 394108 -15242 394448 -15156
rect 394108 -15298 394177 -15242
rect 394233 -15298 394319 -15242
rect 394375 -15298 394448 -15242
rect 394108 -15384 394448 -15298
rect 394108 -15440 394177 -15384
rect 394233 -15440 394319 -15384
rect 394375 -15440 394448 -15384
rect 394108 -15526 394448 -15440
rect 394108 -15582 394177 -15526
rect 394233 -15582 394319 -15526
rect 394375 -15582 394448 -15526
rect 394108 -15668 394448 -15582
rect 394108 -15724 394177 -15668
rect 394233 -15724 394319 -15668
rect 394375 -15724 394448 -15668
rect 394108 -15810 394448 -15724
rect 394108 -15866 394177 -15810
rect 394233 -15866 394319 -15810
rect 394375 -15866 394448 -15810
rect 394108 -15952 394448 -15866
rect 394108 -16008 394177 -15952
rect 394233 -16008 394319 -15952
rect 394375 -16008 394448 -15952
rect 394108 -16094 394448 -16008
rect 394108 -16150 394177 -16094
rect 394233 -16150 394319 -16094
rect 394375 -16150 394448 -16094
rect 394108 -16236 394448 -16150
rect 394108 -16292 394177 -16236
rect 394233 -16292 394319 -16236
rect 394375 -16292 394448 -16236
rect 394108 -16378 394448 -16292
rect 394108 -16434 394177 -16378
rect 394233 -16434 394319 -16378
rect 394375 -16434 394448 -16378
rect 394108 -16520 394448 -16434
rect 394108 -16576 394177 -16520
rect 394233 -16576 394319 -16520
rect 394375 -16576 394448 -16520
rect 394108 -16662 394448 -16576
rect 394108 -16718 394177 -16662
rect 394233 -16718 394319 -16662
rect 394375 -16718 394448 -16662
rect 394108 -16804 394448 -16718
rect 394108 -16860 394177 -16804
rect 394233 -16860 394319 -16804
rect 394375 -16860 394448 -16804
rect 394108 -16946 394448 -16860
rect 394108 -17002 394177 -16946
rect 394233 -17002 394319 -16946
rect 394375 -17002 394448 -16946
rect 394108 -17088 394448 -17002
rect 394108 -17144 394177 -17088
rect 394233 -17144 394319 -17088
rect 394375 -17144 394448 -17088
rect 394108 -17230 394448 -17144
rect 394108 -17286 394177 -17230
rect 394233 -17286 394319 -17230
rect 394375 -17286 394448 -17230
rect 394108 -17372 394448 -17286
rect 394108 -17428 394177 -17372
rect 394233 -17428 394319 -17372
rect 394375 -17428 394448 -17372
rect 394108 -17514 394448 -17428
rect 394108 -17570 394177 -17514
rect 394233 -17570 394319 -17514
rect 394375 -17570 394448 -17514
rect 394108 -17656 394448 -17570
rect 394108 -17712 394177 -17656
rect 394233 -17712 394319 -17656
rect 394375 -17712 394448 -17656
rect 394108 -17798 394448 -17712
rect 394108 -17854 394177 -17798
rect 394233 -17854 394319 -17798
rect 394375 -17854 394448 -17798
rect 394108 -17940 394448 -17854
rect 394108 -17996 394177 -17940
rect 394233 -17996 394319 -17940
rect 394375 -17996 394448 -17940
rect 394108 -18082 394448 -17996
rect 394108 -18138 394177 -18082
rect 394233 -18138 394319 -18082
rect 394375 -18138 394448 -18082
rect 394108 -18224 394448 -18138
rect 394108 -18280 394177 -18224
rect 394233 -18280 394319 -18224
rect 394375 -18280 394448 -18224
rect 394108 -18366 394448 -18280
rect 394108 -18422 394177 -18366
rect 394233 -18422 394319 -18366
rect 394375 -18422 394448 -18366
rect 394108 -18508 394448 -18422
rect 394108 -18564 394177 -18508
rect 394233 -18564 394319 -18508
rect 394375 -18564 394448 -18508
rect 394108 -18650 394448 -18564
rect 394108 -18706 394177 -18650
rect 394233 -18706 394319 -18650
rect 394375 -18706 394448 -18650
rect 394108 -18792 394448 -18706
rect 394108 -18848 394177 -18792
rect 394233 -18848 394319 -18792
rect 394375 -18848 394448 -18792
rect 394108 -18934 394448 -18848
rect 394108 -18990 394177 -18934
rect 394233 -18990 394319 -18934
rect 394375 -18990 394448 -18934
rect 394108 -19076 394448 -18990
rect 394108 -19132 394177 -19076
rect 394233 -19132 394319 -19076
rect 394375 -19132 394448 -19076
rect 394108 -19218 394448 -19132
rect 394108 -19274 394177 -19218
rect 394233 -19274 394319 -19218
rect 394375 -19274 394448 -19218
rect 394108 -19360 394448 -19274
rect 394108 -19416 394177 -19360
rect 394233 -19416 394319 -19360
rect 394375 -19416 394448 -19360
rect 394108 -19502 394448 -19416
rect 394108 -19558 394177 -19502
rect 394233 -19558 394319 -19502
rect 394375 -19558 394448 -19502
rect 394108 -19644 394448 -19558
rect 394108 -19700 394177 -19644
rect 394233 -19700 394319 -19644
rect 394375 -19700 394448 -19644
rect 394108 -19786 394448 -19700
rect 394108 -19842 394177 -19786
rect 394233 -19842 394319 -19786
rect 394375 -19842 394448 -19786
rect 394108 -19928 394448 -19842
rect 394108 -19984 394177 -19928
rect 394233 -19984 394319 -19928
rect 394375 -19984 394448 -19928
rect 394108 -20070 394448 -19984
rect 394108 -20126 394177 -20070
rect 394233 -20126 394319 -20070
rect 394375 -20126 394448 -20070
rect 394108 -20212 394448 -20126
rect 394108 -20268 394177 -20212
rect 394233 -20268 394319 -20212
rect 394375 -20268 394448 -20212
rect 394108 -20354 394448 -20268
rect 394108 -20410 394177 -20354
rect 394233 -20410 394319 -20354
rect 394375 -20410 394448 -20354
rect 394108 -20496 394448 -20410
rect 394108 -20552 394177 -20496
rect 394233 -20552 394319 -20496
rect 394375 -20552 394448 -20496
rect 394108 -20638 394448 -20552
rect 394108 -20694 394177 -20638
rect 394233 -20694 394319 -20638
rect 394375 -20694 394448 -20638
rect 394108 -20780 394448 -20694
rect 394108 -20836 394177 -20780
rect 394233 -20836 394319 -20780
rect 394375 -20836 394448 -20780
rect 394108 -20922 394448 -20836
rect 394108 -20978 394177 -20922
rect 394233 -20978 394319 -20922
rect 394375 -20978 394448 -20922
rect 394108 -21064 394448 -20978
rect 394108 -21120 394177 -21064
rect 394233 -21120 394319 -21064
rect 394375 -21120 394448 -21064
rect 394108 -21206 394448 -21120
rect 394108 -21262 394177 -21206
rect 394233 -21262 394319 -21206
rect 394375 -21262 394448 -21206
rect 394108 -21348 394448 -21262
rect 394108 -21404 394177 -21348
rect 394233 -21404 394319 -21348
rect 394375 -21404 394448 -21348
rect 394108 -21490 394448 -21404
rect 394108 -21546 394177 -21490
rect 394233 -21546 394319 -21490
rect 394375 -21546 394448 -21490
rect 394108 -21632 394448 -21546
rect 394108 -21688 394177 -21632
rect 394233 -21688 394319 -21632
rect 394375 -21688 394448 -21632
rect 394108 -21774 394448 -21688
rect 394108 -21830 394177 -21774
rect 394233 -21830 394319 -21774
rect 394375 -21830 394448 -21774
rect 394108 -21916 394448 -21830
rect 394108 -21972 394177 -21916
rect 394233 -21972 394319 -21916
rect 394375 -21972 394448 -21916
rect 394108 -22058 394448 -21972
rect 394108 -22114 394177 -22058
rect 394233 -22114 394319 -22058
rect 394375 -22114 394448 -22058
rect 394108 -22200 394448 -22114
rect 394108 -22256 394177 -22200
rect 394233 -22256 394319 -22200
rect 394375 -22256 394448 -22200
rect 394108 -22342 394448 -22256
rect 394108 -22398 394177 -22342
rect 394233 -22398 394319 -22342
rect 394375 -22398 394448 -22342
rect 394108 -22484 394448 -22398
rect 394108 -22540 394177 -22484
rect 394233 -22540 394319 -22484
rect 394375 -22540 394448 -22484
rect 394108 -22626 394448 -22540
rect 394108 -22682 394177 -22626
rect 394233 -22682 394319 -22626
rect 394375 -22682 394448 -22626
rect 394108 -22768 394448 -22682
rect 394108 -22824 394177 -22768
rect 394233 -22824 394319 -22768
rect 394375 -22824 394448 -22768
rect 394108 -22910 394448 -22824
rect 394108 -22966 394177 -22910
rect 394233 -22966 394319 -22910
rect 394375 -22966 394448 -22910
rect 394108 -23052 394448 -22966
rect 394108 -23108 394177 -23052
rect 394233 -23108 394319 -23052
rect 394375 -23108 394448 -23052
rect 394108 -23194 394448 -23108
rect 394108 -23250 394177 -23194
rect 394233 -23250 394319 -23194
rect 394375 -23250 394448 -23194
rect 394108 -23336 394448 -23250
rect 394108 -23392 394177 -23336
rect 394233 -23392 394319 -23336
rect 394375 -23392 394448 -23336
rect 394108 -23478 394448 -23392
rect 394108 -23534 394177 -23478
rect 394233 -23534 394319 -23478
rect 394375 -23534 394448 -23478
rect 394108 -23620 394448 -23534
rect 394108 -23676 394177 -23620
rect 394233 -23676 394319 -23620
rect 394375 -23676 394448 -23620
rect 394108 -23762 394448 -23676
rect 394108 -23818 394177 -23762
rect 394233 -23818 394319 -23762
rect 394375 -23818 394448 -23762
rect 394108 -23904 394448 -23818
rect 394108 -23960 394177 -23904
rect 394233 -23960 394319 -23904
rect 394375 -23960 394448 -23904
rect 394108 -24046 394448 -23960
rect 394108 -24102 394177 -24046
rect 394233 -24102 394319 -24046
rect 394375 -24102 394448 -24046
rect 394108 -24188 394448 -24102
rect 394108 -24244 394177 -24188
rect 394233 -24244 394319 -24188
rect 394375 -24244 394448 -24188
rect 394108 -24330 394448 -24244
rect 394108 -24386 394177 -24330
rect 394233 -24386 394319 -24330
rect 394375 -24386 394448 -24330
rect 394108 -24472 394448 -24386
rect 394108 -24528 394177 -24472
rect 394233 -24528 394319 -24472
rect 394375 -24528 394448 -24472
rect 394108 -24614 394448 -24528
rect 394108 -24670 394177 -24614
rect 394233 -24670 394319 -24614
rect 394375 -24670 394448 -24614
rect 394108 -24756 394448 -24670
rect 394108 -24812 394177 -24756
rect 394233 -24812 394319 -24756
rect 394375 -24812 394448 -24756
rect 394108 -24898 394448 -24812
rect 394108 -24954 394177 -24898
rect 394233 -24954 394319 -24898
rect 394375 -24954 394448 -24898
rect 394108 -25040 394448 -24954
rect 394108 -25096 394177 -25040
rect 394233 -25096 394319 -25040
rect 394375 -25096 394448 -25040
rect 394108 -25182 394448 -25096
rect 394108 -25238 394177 -25182
rect 394233 -25238 394319 -25182
rect 394375 -25238 394448 -25182
rect 394108 -25324 394448 -25238
rect 394108 -25380 394177 -25324
rect 394233 -25380 394319 -25324
rect 394375 -25380 394448 -25324
rect 394108 -25466 394448 -25380
rect 394108 -25522 394177 -25466
rect 394233 -25522 394319 -25466
rect 394375 -25522 394448 -25466
rect 394108 -25532 394448 -25522
rect 394508 -13680 394848 -13670
rect 394508 -13736 394580 -13680
rect 394636 -13736 394722 -13680
rect 394778 -13736 394848 -13680
rect 394508 -13822 394848 -13736
rect 394508 -13878 394580 -13822
rect 394636 -13878 394722 -13822
rect 394778 -13878 394848 -13822
rect 394508 -13964 394848 -13878
rect 394508 -14020 394580 -13964
rect 394636 -14020 394722 -13964
rect 394778 -14020 394848 -13964
rect 394508 -14106 394848 -14020
rect 394508 -14162 394580 -14106
rect 394636 -14162 394722 -14106
rect 394778 -14162 394848 -14106
rect 394508 -14248 394848 -14162
rect 394508 -14304 394580 -14248
rect 394636 -14304 394722 -14248
rect 394778 -14304 394848 -14248
rect 394508 -14390 394848 -14304
rect 394508 -14446 394580 -14390
rect 394636 -14446 394722 -14390
rect 394778 -14446 394848 -14390
rect 394508 -14532 394848 -14446
rect 394508 -14588 394580 -14532
rect 394636 -14588 394722 -14532
rect 394778 -14588 394848 -14532
rect 394508 -14674 394848 -14588
rect 394508 -14730 394580 -14674
rect 394636 -14730 394722 -14674
rect 394778 -14730 394848 -14674
rect 394508 -14816 394848 -14730
rect 394508 -14872 394580 -14816
rect 394636 -14872 394722 -14816
rect 394778 -14872 394848 -14816
rect 394508 -14958 394848 -14872
rect 394508 -15014 394580 -14958
rect 394636 -15014 394722 -14958
rect 394778 -15014 394848 -14958
rect 394508 -15100 394848 -15014
rect 394508 -15156 394580 -15100
rect 394636 -15156 394722 -15100
rect 394778 -15156 394848 -15100
rect 394508 -15242 394848 -15156
rect 394508 -15298 394580 -15242
rect 394636 -15298 394722 -15242
rect 394778 -15298 394848 -15242
rect 394508 -15384 394848 -15298
rect 394508 -15440 394580 -15384
rect 394636 -15440 394722 -15384
rect 394778 -15440 394848 -15384
rect 394508 -15526 394848 -15440
rect 394508 -15582 394580 -15526
rect 394636 -15582 394722 -15526
rect 394778 -15582 394848 -15526
rect 394508 -15668 394848 -15582
rect 394508 -15724 394580 -15668
rect 394636 -15724 394722 -15668
rect 394778 -15724 394848 -15668
rect 394508 -15810 394848 -15724
rect 394508 -15866 394580 -15810
rect 394636 -15866 394722 -15810
rect 394778 -15866 394848 -15810
rect 394508 -15952 394848 -15866
rect 394508 -16008 394580 -15952
rect 394636 -16008 394722 -15952
rect 394778 -16008 394848 -15952
rect 394508 -16094 394848 -16008
rect 394508 -16150 394580 -16094
rect 394636 -16150 394722 -16094
rect 394778 -16150 394848 -16094
rect 394508 -16236 394848 -16150
rect 394508 -16292 394580 -16236
rect 394636 -16292 394722 -16236
rect 394778 -16292 394848 -16236
rect 394508 -16378 394848 -16292
rect 394508 -16434 394580 -16378
rect 394636 -16434 394722 -16378
rect 394778 -16434 394848 -16378
rect 394508 -16520 394848 -16434
rect 394508 -16576 394580 -16520
rect 394636 -16576 394722 -16520
rect 394778 -16576 394848 -16520
rect 394508 -16662 394848 -16576
rect 394508 -16718 394580 -16662
rect 394636 -16718 394722 -16662
rect 394778 -16718 394848 -16662
rect 394508 -16804 394848 -16718
rect 394508 -16860 394580 -16804
rect 394636 -16860 394722 -16804
rect 394778 -16860 394848 -16804
rect 394508 -16946 394848 -16860
rect 394508 -17002 394580 -16946
rect 394636 -17002 394722 -16946
rect 394778 -17002 394848 -16946
rect 394508 -17088 394848 -17002
rect 394508 -17144 394580 -17088
rect 394636 -17144 394722 -17088
rect 394778 -17144 394848 -17088
rect 394508 -17230 394848 -17144
rect 394508 -17286 394580 -17230
rect 394636 -17286 394722 -17230
rect 394778 -17286 394848 -17230
rect 394508 -17372 394848 -17286
rect 394508 -17428 394580 -17372
rect 394636 -17428 394722 -17372
rect 394778 -17428 394848 -17372
rect 394508 -17514 394848 -17428
rect 394508 -17570 394580 -17514
rect 394636 -17570 394722 -17514
rect 394778 -17570 394848 -17514
rect 394508 -17656 394848 -17570
rect 394508 -17712 394580 -17656
rect 394636 -17712 394722 -17656
rect 394778 -17712 394848 -17656
rect 394508 -17798 394848 -17712
rect 394508 -17854 394580 -17798
rect 394636 -17854 394722 -17798
rect 394778 -17854 394848 -17798
rect 394508 -17940 394848 -17854
rect 394508 -17996 394580 -17940
rect 394636 -17996 394722 -17940
rect 394778 -17996 394848 -17940
rect 394508 -18082 394848 -17996
rect 394508 -18138 394580 -18082
rect 394636 -18138 394722 -18082
rect 394778 -18138 394848 -18082
rect 394508 -18224 394848 -18138
rect 394508 -18280 394580 -18224
rect 394636 -18280 394722 -18224
rect 394778 -18280 394848 -18224
rect 394508 -18366 394848 -18280
rect 394508 -18422 394580 -18366
rect 394636 -18422 394722 -18366
rect 394778 -18422 394848 -18366
rect 394508 -18508 394848 -18422
rect 394508 -18564 394580 -18508
rect 394636 -18564 394722 -18508
rect 394778 -18564 394848 -18508
rect 394508 -18650 394848 -18564
rect 394508 -18706 394580 -18650
rect 394636 -18706 394722 -18650
rect 394778 -18706 394848 -18650
rect 394508 -18792 394848 -18706
rect 394508 -18848 394580 -18792
rect 394636 -18848 394722 -18792
rect 394778 -18848 394848 -18792
rect 394508 -18934 394848 -18848
rect 394508 -18990 394580 -18934
rect 394636 -18990 394722 -18934
rect 394778 -18990 394848 -18934
rect 394508 -19076 394848 -18990
rect 394508 -19132 394580 -19076
rect 394636 -19132 394722 -19076
rect 394778 -19132 394848 -19076
rect 394508 -19218 394848 -19132
rect 394508 -19274 394580 -19218
rect 394636 -19274 394722 -19218
rect 394778 -19274 394848 -19218
rect 394508 -19360 394848 -19274
rect 394508 -19416 394580 -19360
rect 394636 -19416 394722 -19360
rect 394778 -19416 394848 -19360
rect 394508 -19502 394848 -19416
rect 394508 -19558 394580 -19502
rect 394636 -19558 394722 -19502
rect 394778 -19558 394848 -19502
rect 394508 -19644 394848 -19558
rect 394508 -19700 394580 -19644
rect 394636 -19700 394722 -19644
rect 394778 -19700 394848 -19644
rect 394508 -19786 394848 -19700
rect 394508 -19842 394580 -19786
rect 394636 -19842 394722 -19786
rect 394778 -19842 394848 -19786
rect 394508 -19928 394848 -19842
rect 394508 -19984 394580 -19928
rect 394636 -19984 394722 -19928
rect 394778 -19984 394848 -19928
rect 394508 -20070 394848 -19984
rect 394508 -20126 394580 -20070
rect 394636 -20126 394722 -20070
rect 394778 -20126 394848 -20070
rect 394508 -20212 394848 -20126
rect 394508 -20268 394580 -20212
rect 394636 -20268 394722 -20212
rect 394778 -20268 394848 -20212
rect 394508 -20354 394848 -20268
rect 394508 -20410 394580 -20354
rect 394636 -20410 394722 -20354
rect 394778 -20410 394848 -20354
rect 394508 -20496 394848 -20410
rect 394508 -20552 394580 -20496
rect 394636 -20552 394722 -20496
rect 394778 -20552 394848 -20496
rect 394508 -20638 394848 -20552
rect 394508 -20694 394580 -20638
rect 394636 -20694 394722 -20638
rect 394778 -20694 394848 -20638
rect 394508 -20780 394848 -20694
rect 394508 -20836 394580 -20780
rect 394636 -20836 394722 -20780
rect 394778 -20836 394848 -20780
rect 394508 -20922 394848 -20836
rect 394508 -20978 394580 -20922
rect 394636 -20978 394722 -20922
rect 394778 -20978 394848 -20922
rect 394508 -21064 394848 -20978
rect 394508 -21120 394580 -21064
rect 394636 -21120 394722 -21064
rect 394778 -21120 394848 -21064
rect 394508 -21206 394848 -21120
rect 394508 -21262 394580 -21206
rect 394636 -21262 394722 -21206
rect 394778 -21262 394848 -21206
rect 394508 -21348 394848 -21262
rect 394508 -21404 394580 -21348
rect 394636 -21404 394722 -21348
rect 394778 -21404 394848 -21348
rect 394508 -21490 394848 -21404
rect 394508 -21546 394580 -21490
rect 394636 -21546 394722 -21490
rect 394778 -21546 394848 -21490
rect 394508 -21632 394848 -21546
rect 394508 -21688 394580 -21632
rect 394636 -21688 394722 -21632
rect 394778 -21688 394848 -21632
rect 394508 -21774 394848 -21688
rect 394508 -21830 394580 -21774
rect 394636 -21830 394722 -21774
rect 394778 -21830 394848 -21774
rect 394508 -21916 394848 -21830
rect 394508 -21972 394580 -21916
rect 394636 -21972 394722 -21916
rect 394778 -21972 394848 -21916
rect 394508 -22058 394848 -21972
rect 394508 -22114 394580 -22058
rect 394636 -22114 394722 -22058
rect 394778 -22114 394848 -22058
rect 394508 -22200 394848 -22114
rect 394508 -22256 394580 -22200
rect 394636 -22256 394722 -22200
rect 394778 -22256 394848 -22200
rect 394508 -22342 394848 -22256
rect 394508 -22398 394580 -22342
rect 394636 -22398 394722 -22342
rect 394778 -22398 394848 -22342
rect 394508 -22484 394848 -22398
rect 394508 -22540 394580 -22484
rect 394636 -22540 394722 -22484
rect 394778 -22540 394848 -22484
rect 394508 -22626 394848 -22540
rect 394508 -22682 394580 -22626
rect 394636 -22682 394722 -22626
rect 394778 -22682 394848 -22626
rect 394508 -22768 394848 -22682
rect 394508 -22824 394580 -22768
rect 394636 -22824 394722 -22768
rect 394778 -22824 394848 -22768
rect 394508 -22910 394848 -22824
rect 394508 -22966 394580 -22910
rect 394636 -22966 394722 -22910
rect 394778 -22966 394848 -22910
rect 394508 -23052 394848 -22966
rect 394508 -23108 394580 -23052
rect 394636 -23108 394722 -23052
rect 394778 -23108 394848 -23052
rect 394508 -23194 394848 -23108
rect 394508 -23250 394580 -23194
rect 394636 -23250 394722 -23194
rect 394778 -23250 394848 -23194
rect 394508 -23336 394848 -23250
rect 394508 -23392 394580 -23336
rect 394636 -23392 394722 -23336
rect 394778 -23392 394848 -23336
rect 394508 -23478 394848 -23392
rect 394508 -23534 394580 -23478
rect 394636 -23534 394722 -23478
rect 394778 -23534 394848 -23478
rect 394508 -23620 394848 -23534
rect 394508 -23676 394580 -23620
rect 394636 -23676 394722 -23620
rect 394778 -23676 394848 -23620
rect 394508 -23762 394848 -23676
rect 394508 -23818 394580 -23762
rect 394636 -23818 394722 -23762
rect 394778 -23818 394848 -23762
rect 394508 -23904 394848 -23818
rect 394508 -23960 394580 -23904
rect 394636 -23960 394722 -23904
rect 394778 -23960 394848 -23904
rect 394508 -24046 394848 -23960
rect 394508 -24102 394580 -24046
rect 394636 -24102 394722 -24046
rect 394778 -24102 394848 -24046
rect 394508 -24188 394848 -24102
rect 394508 -24244 394580 -24188
rect 394636 -24244 394722 -24188
rect 394778 -24244 394848 -24188
rect 394508 -24330 394848 -24244
rect 394508 -24386 394580 -24330
rect 394636 -24386 394722 -24330
rect 394778 -24386 394848 -24330
rect 394508 -24472 394848 -24386
rect 394508 -24528 394580 -24472
rect 394636 -24528 394722 -24472
rect 394778 -24528 394848 -24472
rect 394508 -24614 394848 -24528
rect 394508 -24670 394580 -24614
rect 394636 -24670 394722 -24614
rect 394778 -24670 394848 -24614
rect 394508 -24756 394848 -24670
rect 394508 -24812 394580 -24756
rect 394636 -24812 394722 -24756
rect 394778 -24812 394848 -24756
rect 394508 -24898 394848 -24812
rect 394508 -24954 394580 -24898
rect 394636 -24954 394722 -24898
rect 394778 -24954 394848 -24898
rect 394508 -25040 394848 -24954
rect 394508 -25096 394580 -25040
rect 394636 -25096 394722 -25040
rect 394778 -25096 394848 -25040
rect 394508 -25182 394848 -25096
rect 394508 -25238 394580 -25182
rect 394636 -25238 394722 -25182
rect 394778 -25238 394848 -25182
rect 394508 -25324 394848 -25238
rect 394508 -25380 394580 -25324
rect 394636 -25380 394722 -25324
rect 394778 -25380 394848 -25324
rect 394508 -25466 394848 -25380
rect 394508 -25522 394580 -25466
rect 394636 -25522 394722 -25466
rect 394778 -25522 394848 -25466
rect 394508 -25532 394848 -25522
rect 394908 -13680 395248 -13670
rect 394908 -13736 394982 -13680
rect 395038 -13736 395124 -13680
rect 395180 -13736 395248 -13680
rect 394908 -13822 395248 -13736
rect 394908 -13878 394982 -13822
rect 395038 -13878 395124 -13822
rect 395180 -13878 395248 -13822
rect 394908 -13964 395248 -13878
rect 394908 -14020 394982 -13964
rect 395038 -14020 395124 -13964
rect 395180 -14020 395248 -13964
rect 394908 -14106 395248 -14020
rect 394908 -14162 394982 -14106
rect 395038 -14162 395124 -14106
rect 395180 -14162 395248 -14106
rect 394908 -14248 395248 -14162
rect 394908 -14304 394982 -14248
rect 395038 -14304 395124 -14248
rect 395180 -14304 395248 -14248
rect 394908 -14390 395248 -14304
rect 394908 -14446 394982 -14390
rect 395038 -14446 395124 -14390
rect 395180 -14446 395248 -14390
rect 394908 -14532 395248 -14446
rect 394908 -14588 394982 -14532
rect 395038 -14588 395124 -14532
rect 395180 -14588 395248 -14532
rect 394908 -14674 395248 -14588
rect 394908 -14730 394982 -14674
rect 395038 -14730 395124 -14674
rect 395180 -14730 395248 -14674
rect 394908 -14816 395248 -14730
rect 394908 -14872 394982 -14816
rect 395038 -14872 395124 -14816
rect 395180 -14872 395248 -14816
rect 394908 -14958 395248 -14872
rect 394908 -15014 394982 -14958
rect 395038 -15014 395124 -14958
rect 395180 -15014 395248 -14958
rect 394908 -15100 395248 -15014
rect 394908 -15156 394982 -15100
rect 395038 -15156 395124 -15100
rect 395180 -15156 395248 -15100
rect 394908 -15242 395248 -15156
rect 394908 -15298 394982 -15242
rect 395038 -15298 395124 -15242
rect 395180 -15298 395248 -15242
rect 394908 -15384 395248 -15298
rect 394908 -15440 394982 -15384
rect 395038 -15440 395124 -15384
rect 395180 -15440 395248 -15384
rect 394908 -15526 395248 -15440
rect 394908 -15582 394982 -15526
rect 395038 -15582 395124 -15526
rect 395180 -15582 395248 -15526
rect 394908 -15668 395248 -15582
rect 394908 -15724 394982 -15668
rect 395038 -15724 395124 -15668
rect 395180 -15724 395248 -15668
rect 394908 -15810 395248 -15724
rect 394908 -15866 394982 -15810
rect 395038 -15866 395124 -15810
rect 395180 -15866 395248 -15810
rect 394908 -15952 395248 -15866
rect 394908 -16008 394982 -15952
rect 395038 -16008 395124 -15952
rect 395180 -16008 395248 -15952
rect 394908 -16094 395248 -16008
rect 394908 -16150 394982 -16094
rect 395038 -16150 395124 -16094
rect 395180 -16150 395248 -16094
rect 394908 -16236 395248 -16150
rect 394908 -16292 394982 -16236
rect 395038 -16292 395124 -16236
rect 395180 -16292 395248 -16236
rect 394908 -16378 395248 -16292
rect 394908 -16434 394982 -16378
rect 395038 -16434 395124 -16378
rect 395180 -16434 395248 -16378
rect 394908 -16520 395248 -16434
rect 394908 -16576 394982 -16520
rect 395038 -16576 395124 -16520
rect 395180 -16576 395248 -16520
rect 394908 -16662 395248 -16576
rect 394908 -16718 394982 -16662
rect 395038 -16718 395124 -16662
rect 395180 -16718 395248 -16662
rect 394908 -16804 395248 -16718
rect 394908 -16860 394982 -16804
rect 395038 -16860 395124 -16804
rect 395180 -16860 395248 -16804
rect 394908 -16946 395248 -16860
rect 394908 -17002 394982 -16946
rect 395038 -17002 395124 -16946
rect 395180 -17002 395248 -16946
rect 394908 -17088 395248 -17002
rect 394908 -17144 394982 -17088
rect 395038 -17144 395124 -17088
rect 395180 -17144 395248 -17088
rect 394908 -17230 395248 -17144
rect 394908 -17286 394982 -17230
rect 395038 -17286 395124 -17230
rect 395180 -17286 395248 -17230
rect 394908 -17372 395248 -17286
rect 394908 -17428 394982 -17372
rect 395038 -17428 395124 -17372
rect 395180 -17428 395248 -17372
rect 394908 -17514 395248 -17428
rect 394908 -17570 394982 -17514
rect 395038 -17570 395124 -17514
rect 395180 -17570 395248 -17514
rect 394908 -17656 395248 -17570
rect 394908 -17712 394982 -17656
rect 395038 -17712 395124 -17656
rect 395180 -17712 395248 -17656
rect 394908 -17798 395248 -17712
rect 394908 -17854 394982 -17798
rect 395038 -17854 395124 -17798
rect 395180 -17854 395248 -17798
rect 394908 -17940 395248 -17854
rect 394908 -17996 394982 -17940
rect 395038 -17996 395124 -17940
rect 395180 -17996 395248 -17940
rect 394908 -18082 395248 -17996
rect 394908 -18138 394982 -18082
rect 395038 -18138 395124 -18082
rect 395180 -18138 395248 -18082
rect 394908 -18224 395248 -18138
rect 394908 -18280 394982 -18224
rect 395038 -18280 395124 -18224
rect 395180 -18280 395248 -18224
rect 394908 -18366 395248 -18280
rect 394908 -18422 394982 -18366
rect 395038 -18422 395124 -18366
rect 395180 -18422 395248 -18366
rect 394908 -18508 395248 -18422
rect 394908 -18564 394982 -18508
rect 395038 -18564 395124 -18508
rect 395180 -18564 395248 -18508
rect 394908 -18650 395248 -18564
rect 394908 -18706 394982 -18650
rect 395038 -18706 395124 -18650
rect 395180 -18706 395248 -18650
rect 394908 -18792 395248 -18706
rect 394908 -18848 394982 -18792
rect 395038 -18848 395124 -18792
rect 395180 -18848 395248 -18792
rect 394908 -18934 395248 -18848
rect 394908 -18990 394982 -18934
rect 395038 -18990 395124 -18934
rect 395180 -18990 395248 -18934
rect 394908 -19076 395248 -18990
rect 394908 -19132 394982 -19076
rect 395038 -19132 395124 -19076
rect 395180 -19132 395248 -19076
rect 394908 -19218 395248 -19132
rect 394908 -19274 394982 -19218
rect 395038 -19274 395124 -19218
rect 395180 -19274 395248 -19218
rect 394908 -19360 395248 -19274
rect 394908 -19416 394982 -19360
rect 395038 -19416 395124 -19360
rect 395180 -19416 395248 -19360
rect 394908 -19502 395248 -19416
rect 394908 -19558 394982 -19502
rect 395038 -19558 395124 -19502
rect 395180 -19558 395248 -19502
rect 394908 -19644 395248 -19558
rect 394908 -19700 394982 -19644
rect 395038 -19700 395124 -19644
rect 395180 -19700 395248 -19644
rect 394908 -19786 395248 -19700
rect 394908 -19842 394982 -19786
rect 395038 -19842 395124 -19786
rect 395180 -19842 395248 -19786
rect 394908 -19928 395248 -19842
rect 394908 -19984 394982 -19928
rect 395038 -19984 395124 -19928
rect 395180 -19984 395248 -19928
rect 394908 -20070 395248 -19984
rect 394908 -20126 394982 -20070
rect 395038 -20126 395124 -20070
rect 395180 -20126 395248 -20070
rect 394908 -20212 395248 -20126
rect 394908 -20268 394982 -20212
rect 395038 -20268 395124 -20212
rect 395180 -20268 395248 -20212
rect 394908 -20354 395248 -20268
rect 394908 -20410 394982 -20354
rect 395038 -20410 395124 -20354
rect 395180 -20410 395248 -20354
rect 394908 -20496 395248 -20410
rect 394908 -20552 394982 -20496
rect 395038 -20552 395124 -20496
rect 395180 -20552 395248 -20496
rect 394908 -20638 395248 -20552
rect 394908 -20694 394982 -20638
rect 395038 -20694 395124 -20638
rect 395180 -20694 395248 -20638
rect 394908 -20780 395248 -20694
rect 394908 -20836 394982 -20780
rect 395038 -20836 395124 -20780
rect 395180 -20836 395248 -20780
rect 394908 -20922 395248 -20836
rect 394908 -20978 394982 -20922
rect 395038 -20978 395124 -20922
rect 395180 -20978 395248 -20922
rect 394908 -21064 395248 -20978
rect 394908 -21120 394982 -21064
rect 395038 -21120 395124 -21064
rect 395180 -21120 395248 -21064
rect 394908 -21206 395248 -21120
rect 394908 -21262 394982 -21206
rect 395038 -21262 395124 -21206
rect 395180 -21262 395248 -21206
rect 394908 -21348 395248 -21262
rect 394908 -21404 394982 -21348
rect 395038 -21404 395124 -21348
rect 395180 -21404 395248 -21348
rect 394908 -21490 395248 -21404
rect 394908 -21546 394982 -21490
rect 395038 -21546 395124 -21490
rect 395180 -21546 395248 -21490
rect 394908 -21632 395248 -21546
rect 394908 -21688 394982 -21632
rect 395038 -21688 395124 -21632
rect 395180 -21688 395248 -21632
rect 394908 -21774 395248 -21688
rect 394908 -21830 394982 -21774
rect 395038 -21830 395124 -21774
rect 395180 -21830 395248 -21774
rect 394908 -21916 395248 -21830
rect 394908 -21972 394982 -21916
rect 395038 -21972 395124 -21916
rect 395180 -21972 395248 -21916
rect 394908 -22058 395248 -21972
rect 394908 -22114 394982 -22058
rect 395038 -22114 395124 -22058
rect 395180 -22114 395248 -22058
rect 394908 -22200 395248 -22114
rect 394908 -22256 394982 -22200
rect 395038 -22256 395124 -22200
rect 395180 -22256 395248 -22200
rect 394908 -22342 395248 -22256
rect 394908 -22398 394982 -22342
rect 395038 -22398 395124 -22342
rect 395180 -22398 395248 -22342
rect 394908 -22484 395248 -22398
rect 394908 -22540 394982 -22484
rect 395038 -22540 395124 -22484
rect 395180 -22540 395248 -22484
rect 394908 -22626 395248 -22540
rect 394908 -22682 394982 -22626
rect 395038 -22682 395124 -22626
rect 395180 -22682 395248 -22626
rect 394908 -22768 395248 -22682
rect 394908 -22824 394982 -22768
rect 395038 -22824 395124 -22768
rect 395180 -22824 395248 -22768
rect 394908 -22910 395248 -22824
rect 394908 -22966 394982 -22910
rect 395038 -22966 395124 -22910
rect 395180 -22966 395248 -22910
rect 394908 -23052 395248 -22966
rect 394908 -23108 394982 -23052
rect 395038 -23108 395124 -23052
rect 395180 -23108 395248 -23052
rect 394908 -23194 395248 -23108
rect 394908 -23250 394982 -23194
rect 395038 -23250 395124 -23194
rect 395180 -23250 395248 -23194
rect 394908 -23336 395248 -23250
rect 394908 -23392 394982 -23336
rect 395038 -23392 395124 -23336
rect 395180 -23392 395248 -23336
rect 394908 -23478 395248 -23392
rect 394908 -23534 394982 -23478
rect 395038 -23534 395124 -23478
rect 395180 -23534 395248 -23478
rect 394908 -23620 395248 -23534
rect 394908 -23676 394982 -23620
rect 395038 -23676 395124 -23620
rect 395180 -23676 395248 -23620
rect 394908 -23762 395248 -23676
rect 394908 -23818 394982 -23762
rect 395038 -23818 395124 -23762
rect 395180 -23818 395248 -23762
rect 394908 -23904 395248 -23818
rect 394908 -23960 394982 -23904
rect 395038 -23960 395124 -23904
rect 395180 -23960 395248 -23904
rect 394908 -24046 395248 -23960
rect 394908 -24102 394982 -24046
rect 395038 -24102 395124 -24046
rect 395180 -24102 395248 -24046
rect 394908 -24188 395248 -24102
rect 394908 -24244 394982 -24188
rect 395038 -24244 395124 -24188
rect 395180 -24244 395248 -24188
rect 394908 -24330 395248 -24244
rect 394908 -24386 394982 -24330
rect 395038 -24386 395124 -24330
rect 395180 -24386 395248 -24330
rect 394908 -24472 395248 -24386
rect 394908 -24528 394982 -24472
rect 395038 -24528 395124 -24472
rect 395180 -24528 395248 -24472
rect 394908 -24614 395248 -24528
rect 394908 -24670 394982 -24614
rect 395038 -24670 395124 -24614
rect 395180 -24670 395248 -24614
rect 394908 -24756 395248 -24670
rect 394908 -24812 394982 -24756
rect 395038 -24812 395124 -24756
rect 395180 -24812 395248 -24756
rect 394908 -24898 395248 -24812
rect 394908 -24954 394982 -24898
rect 395038 -24954 395124 -24898
rect 395180 -24954 395248 -24898
rect 394908 -25040 395248 -24954
rect 394908 -25096 394982 -25040
rect 395038 -25096 395124 -25040
rect 395180 -25096 395248 -25040
rect 394908 -25182 395248 -25096
rect 394908 -25238 394982 -25182
rect 395038 -25238 395124 -25182
rect 395180 -25238 395248 -25182
rect 394908 -25324 395248 -25238
rect 394908 -25380 394982 -25324
rect 395038 -25380 395124 -25324
rect 395180 -25380 395248 -25324
rect 394908 -25466 395248 -25380
rect 394908 -25522 394982 -25466
rect 395038 -25522 395124 -25466
rect 395180 -25522 395248 -25466
rect 394908 -25532 395248 -25522
rect 395308 -13680 395648 -13670
rect 395308 -13736 395385 -13680
rect 395441 -13736 395527 -13680
rect 395583 -13736 395648 -13680
rect 395308 -13822 395648 -13736
rect 395308 -13878 395385 -13822
rect 395441 -13878 395527 -13822
rect 395583 -13878 395648 -13822
rect 395308 -13964 395648 -13878
rect 395308 -14020 395385 -13964
rect 395441 -14020 395527 -13964
rect 395583 -14020 395648 -13964
rect 395308 -14106 395648 -14020
rect 395308 -14162 395385 -14106
rect 395441 -14162 395527 -14106
rect 395583 -14162 395648 -14106
rect 395308 -14248 395648 -14162
rect 395308 -14304 395385 -14248
rect 395441 -14304 395527 -14248
rect 395583 -14304 395648 -14248
rect 395308 -14390 395648 -14304
rect 395308 -14446 395385 -14390
rect 395441 -14446 395527 -14390
rect 395583 -14446 395648 -14390
rect 395308 -14532 395648 -14446
rect 395308 -14588 395385 -14532
rect 395441 -14588 395527 -14532
rect 395583 -14588 395648 -14532
rect 395308 -14674 395648 -14588
rect 395308 -14730 395385 -14674
rect 395441 -14730 395527 -14674
rect 395583 -14730 395648 -14674
rect 395308 -14816 395648 -14730
rect 395308 -14872 395385 -14816
rect 395441 -14872 395527 -14816
rect 395583 -14872 395648 -14816
rect 395308 -14958 395648 -14872
rect 395308 -15014 395385 -14958
rect 395441 -15014 395527 -14958
rect 395583 -15014 395648 -14958
rect 395308 -15100 395648 -15014
rect 395308 -15156 395385 -15100
rect 395441 -15156 395527 -15100
rect 395583 -15156 395648 -15100
rect 395308 -15242 395648 -15156
rect 395308 -15298 395385 -15242
rect 395441 -15298 395527 -15242
rect 395583 -15298 395648 -15242
rect 395308 -15384 395648 -15298
rect 395308 -15440 395385 -15384
rect 395441 -15440 395527 -15384
rect 395583 -15440 395648 -15384
rect 395308 -15526 395648 -15440
rect 395308 -15582 395385 -15526
rect 395441 -15582 395527 -15526
rect 395583 -15582 395648 -15526
rect 395308 -15668 395648 -15582
rect 395308 -15724 395385 -15668
rect 395441 -15724 395527 -15668
rect 395583 -15724 395648 -15668
rect 395308 -15810 395648 -15724
rect 395308 -15866 395385 -15810
rect 395441 -15866 395527 -15810
rect 395583 -15866 395648 -15810
rect 395308 -15952 395648 -15866
rect 395308 -16008 395385 -15952
rect 395441 -16008 395527 -15952
rect 395583 -16008 395648 -15952
rect 395308 -16094 395648 -16008
rect 395308 -16150 395385 -16094
rect 395441 -16150 395527 -16094
rect 395583 -16150 395648 -16094
rect 395308 -16236 395648 -16150
rect 395308 -16292 395385 -16236
rect 395441 -16292 395527 -16236
rect 395583 -16292 395648 -16236
rect 395308 -16378 395648 -16292
rect 395308 -16434 395385 -16378
rect 395441 -16434 395527 -16378
rect 395583 -16434 395648 -16378
rect 395308 -16520 395648 -16434
rect 395308 -16576 395385 -16520
rect 395441 -16576 395527 -16520
rect 395583 -16576 395648 -16520
rect 395308 -16662 395648 -16576
rect 395308 -16718 395385 -16662
rect 395441 -16718 395527 -16662
rect 395583 -16718 395648 -16662
rect 395308 -16804 395648 -16718
rect 395308 -16860 395385 -16804
rect 395441 -16860 395527 -16804
rect 395583 -16860 395648 -16804
rect 395308 -16946 395648 -16860
rect 395308 -17002 395385 -16946
rect 395441 -17002 395527 -16946
rect 395583 -17002 395648 -16946
rect 395308 -17088 395648 -17002
rect 395308 -17144 395385 -17088
rect 395441 -17144 395527 -17088
rect 395583 -17144 395648 -17088
rect 395308 -17230 395648 -17144
rect 395308 -17286 395385 -17230
rect 395441 -17286 395527 -17230
rect 395583 -17286 395648 -17230
rect 395308 -17372 395648 -17286
rect 395308 -17428 395385 -17372
rect 395441 -17428 395527 -17372
rect 395583 -17428 395648 -17372
rect 395308 -17514 395648 -17428
rect 395308 -17570 395385 -17514
rect 395441 -17570 395527 -17514
rect 395583 -17570 395648 -17514
rect 395308 -17656 395648 -17570
rect 395308 -17712 395385 -17656
rect 395441 -17712 395527 -17656
rect 395583 -17712 395648 -17656
rect 395308 -17798 395648 -17712
rect 395308 -17854 395385 -17798
rect 395441 -17854 395527 -17798
rect 395583 -17854 395648 -17798
rect 395308 -17940 395648 -17854
rect 395308 -17996 395385 -17940
rect 395441 -17996 395527 -17940
rect 395583 -17996 395648 -17940
rect 395308 -18082 395648 -17996
rect 395308 -18138 395385 -18082
rect 395441 -18138 395527 -18082
rect 395583 -18138 395648 -18082
rect 395308 -18224 395648 -18138
rect 395308 -18280 395385 -18224
rect 395441 -18280 395527 -18224
rect 395583 -18280 395648 -18224
rect 395308 -18366 395648 -18280
rect 395308 -18422 395385 -18366
rect 395441 -18422 395527 -18366
rect 395583 -18422 395648 -18366
rect 395308 -18508 395648 -18422
rect 395308 -18564 395385 -18508
rect 395441 -18564 395527 -18508
rect 395583 -18564 395648 -18508
rect 395308 -18650 395648 -18564
rect 395308 -18706 395385 -18650
rect 395441 -18706 395527 -18650
rect 395583 -18706 395648 -18650
rect 395308 -18792 395648 -18706
rect 395308 -18848 395385 -18792
rect 395441 -18848 395527 -18792
rect 395583 -18848 395648 -18792
rect 395308 -18934 395648 -18848
rect 395308 -18990 395385 -18934
rect 395441 -18990 395527 -18934
rect 395583 -18990 395648 -18934
rect 395308 -19076 395648 -18990
rect 395308 -19132 395385 -19076
rect 395441 -19132 395527 -19076
rect 395583 -19132 395648 -19076
rect 395308 -19218 395648 -19132
rect 395308 -19274 395385 -19218
rect 395441 -19274 395527 -19218
rect 395583 -19274 395648 -19218
rect 395308 -19360 395648 -19274
rect 395308 -19416 395385 -19360
rect 395441 -19416 395527 -19360
rect 395583 -19416 395648 -19360
rect 395308 -19502 395648 -19416
rect 395308 -19558 395385 -19502
rect 395441 -19558 395527 -19502
rect 395583 -19558 395648 -19502
rect 395308 -19644 395648 -19558
rect 395308 -19700 395385 -19644
rect 395441 -19700 395527 -19644
rect 395583 -19700 395648 -19644
rect 395308 -19786 395648 -19700
rect 395308 -19842 395385 -19786
rect 395441 -19842 395527 -19786
rect 395583 -19842 395648 -19786
rect 395308 -19928 395648 -19842
rect 395308 -19984 395385 -19928
rect 395441 -19984 395527 -19928
rect 395583 -19984 395648 -19928
rect 395308 -20070 395648 -19984
rect 395308 -20126 395385 -20070
rect 395441 -20126 395527 -20070
rect 395583 -20126 395648 -20070
rect 395308 -20212 395648 -20126
rect 395308 -20268 395385 -20212
rect 395441 -20268 395527 -20212
rect 395583 -20268 395648 -20212
rect 395308 -20354 395648 -20268
rect 395308 -20410 395385 -20354
rect 395441 -20410 395527 -20354
rect 395583 -20410 395648 -20354
rect 395308 -20496 395648 -20410
rect 395308 -20552 395385 -20496
rect 395441 -20552 395527 -20496
rect 395583 -20552 395648 -20496
rect 395308 -20638 395648 -20552
rect 395308 -20694 395385 -20638
rect 395441 -20694 395527 -20638
rect 395583 -20694 395648 -20638
rect 395308 -20780 395648 -20694
rect 395308 -20836 395385 -20780
rect 395441 -20836 395527 -20780
rect 395583 -20836 395648 -20780
rect 395308 -20922 395648 -20836
rect 395308 -20978 395385 -20922
rect 395441 -20978 395527 -20922
rect 395583 -20978 395648 -20922
rect 395308 -21064 395648 -20978
rect 395308 -21120 395385 -21064
rect 395441 -21120 395527 -21064
rect 395583 -21120 395648 -21064
rect 395308 -21206 395648 -21120
rect 395308 -21262 395385 -21206
rect 395441 -21262 395527 -21206
rect 395583 -21262 395648 -21206
rect 395308 -21348 395648 -21262
rect 395308 -21404 395385 -21348
rect 395441 -21404 395527 -21348
rect 395583 -21404 395648 -21348
rect 395308 -21490 395648 -21404
rect 395308 -21546 395385 -21490
rect 395441 -21546 395527 -21490
rect 395583 -21546 395648 -21490
rect 395308 -21632 395648 -21546
rect 395308 -21688 395385 -21632
rect 395441 -21688 395527 -21632
rect 395583 -21688 395648 -21632
rect 395308 -21774 395648 -21688
rect 395308 -21830 395385 -21774
rect 395441 -21830 395527 -21774
rect 395583 -21830 395648 -21774
rect 395308 -21916 395648 -21830
rect 395308 -21972 395385 -21916
rect 395441 -21972 395527 -21916
rect 395583 -21972 395648 -21916
rect 395308 -22058 395648 -21972
rect 395308 -22114 395385 -22058
rect 395441 -22114 395527 -22058
rect 395583 -22114 395648 -22058
rect 395308 -22200 395648 -22114
rect 395308 -22256 395385 -22200
rect 395441 -22256 395527 -22200
rect 395583 -22256 395648 -22200
rect 395308 -22342 395648 -22256
rect 395308 -22398 395385 -22342
rect 395441 -22398 395527 -22342
rect 395583 -22398 395648 -22342
rect 395308 -22484 395648 -22398
rect 395308 -22540 395385 -22484
rect 395441 -22540 395527 -22484
rect 395583 -22540 395648 -22484
rect 395308 -22626 395648 -22540
rect 395308 -22682 395385 -22626
rect 395441 -22682 395527 -22626
rect 395583 -22682 395648 -22626
rect 395308 -22768 395648 -22682
rect 395308 -22824 395385 -22768
rect 395441 -22824 395527 -22768
rect 395583 -22824 395648 -22768
rect 395308 -22910 395648 -22824
rect 395308 -22966 395385 -22910
rect 395441 -22966 395527 -22910
rect 395583 -22966 395648 -22910
rect 395308 -23052 395648 -22966
rect 395308 -23108 395385 -23052
rect 395441 -23108 395527 -23052
rect 395583 -23108 395648 -23052
rect 395308 -23194 395648 -23108
rect 395308 -23250 395385 -23194
rect 395441 -23250 395527 -23194
rect 395583 -23250 395648 -23194
rect 395308 -23336 395648 -23250
rect 395308 -23392 395385 -23336
rect 395441 -23392 395527 -23336
rect 395583 -23392 395648 -23336
rect 395308 -23478 395648 -23392
rect 395308 -23534 395385 -23478
rect 395441 -23534 395527 -23478
rect 395583 -23534 395648 -23478
rect 395308 -23620 395648 -23534
rect 395308 -23676 395385 -23620
rect 395441 -23676 395527 -23620
rect 395583 -23676 395648 -23620
rect 395308 -23762 395648 -23676
rect 395308 -23818 395385 -23762
rect 395441 -23818 395527 -23762
rect 395583 -23818 395648 -23762
rect 395308 -23904 395648 -23818
rect 395308 -23960 395385 -23904
rect 395441 -23960 395527 -23904
rect 395583 -23960 395648 -23904
rect 395308 -24046 395648 -23960
rect 395308 -24102 395385 -24046
rect 395441 -24102 395527 -24046
rect 395583 -24102 395648 -24046
rect 395308 -24188 395648 -24102
rect 395308 -24244 395385 -24188
rect 395441 -24244 395527 -24188
rect 395583 -24244 395648 -24188
rect 395308 -24330 395648 -24244
rect 395308 -24386 395385 -24330
rect 395441 -24386 395527 -24330
rect 395583 -24386 395648 -24330
rect 395308 -24472 395648 -24386
rect 395308 -24528 395385 -24472
rect 395441 -24528 395527 -24472
rect 395583 -24528 395648 -24472
rect 395308 -24614 395648 -24528
rect 395308 -24670 395385 -24614
rect 395441 -24670 395527 -24614
rect 395583 -24670 395648 -24614
rect 395308 -24756 395648 -24670
rect 395308 -24812 395385 -24756
rect 395441 -24812 395527 -24756
rect 395583 -24812 395648 -24756
rect 395308 -24898 395648 -24812
rect 395308 -24954 395385 -24898
rect 395441 -24954 395527 -24898
rect 395583 -24954 395648 -24898
rect 395308 -25040 395648 -24954
rect 395308 -25096 395385 -25040
rect 395441 -25096 395527 -25040
rect 395583 -25096 395648 -25040
rect 395308 -25182 395648 -25096
rect 395308 -25238 395385 -25182
rect 395441 -25238 395527 -25182
rect 395583 -25238 395648 -25182
rect 395308 -25324 395648 -25238
rect 395308 -25380 395385 -25324
rect 395441 -25380 395527 -25324
rect 395583 -25380 395648 -25324
rect 395308 -25466 395648 -25380
rect 395308 -25522 395385 -25466
rect 395441 -25522 395527 -25466
rect 395583 -25522 395648 -25466
rect 395308 -25532 395648 -25522
rect 395708 -13680 396048 -13670
rect 395708 -13736 395779 -13680
rect 395835 -13736 395921 -13680
rect 395977 -13736 396048 -13680
rect 395708 -13822 396048 -13736
rect 395708 -13878 395779 -13822
rect 395835 -13878 395921 -13822
rect 395977 -13878 396048 -13822
rect 395708 -13964 396048 -13878
rect 395708 -14020 395779 -13964
rect 395835 -14020 395921 -13964
rect 395977 -14020 396048 -13964
rect 395708 -14106 396048 -14020
rect 395708 -14162 395779 -14106
rect 395835 -14162 395921 -14106
rect 395977 -14162 396048 -14106
rect 395708 -14248 396048 -14162
rect 395708 -14304 395779 -14248
rect 395835 -14304 395921 -14248
rect 395977 -14304 396048 -14248
rect 395708 -14390 396048 -14304
rect 395708 -14446 395779 -14390
rect 395835 -14446 395921 -14390
rect 395977 -14446 396048 -14390
rect 395708 -14532 396048 -14446
rect 395708 -14588 395779 -14532
rect 395835 -14588 395921 -14532
rect 395977 -14588 396048 -14532
rect 395708 -14674 396048 -14588
rect 395708 -14730 395779 -14674
rect 395835 -14730 395921 -14674
rect 395977 -14730 396048 -14674
rect 395708 -14816 396048 -14730
rect 395708 -14872 395779 -14816
rect 395835 -14872 395921 -14816
rect 395977 -14872 396048 -14816
rect 395708 -14958 396048 -14872
rect 395708 -15014 395779 -14958
rect 395835 -15014 395921 -14958
rect 395977 -15014 396048 -14958
rect 395708 -15100 396048 -15014
rect 395708 -15156 395779 -15100
rect 395835 -15156 395921 -15100
rect 395977 -15156 396048 -15100
rect 395708 -15242 396048 -15156
rect 395708 -15298 395779 -15242
rect 395835 -15298 395921 -15242
rect 395977 -15298 396048 -15242
rect 395708 -15384 396048 -15298
rect 395708 -15440 395779 -15384
rect 395835 -15440 395921 -15384
rect 395977 -15440 396048 -15384
rect 395708 -15526 396048 -15440
rect 395708 -15582 395779 -15526
rect 395835 -15582 395921 -15526
rect 395977 -15582 396048 -15526
rect 395708 -15668 396048 -15582
rect 395708 -15724 395779 -15668
rect 395835 -15724 395921 -15668
rect 395977 -15724 396048 -15668
rect 395708 -15810 396048 -15724
rect 395708 -15866 395779 -15810
rect 395835 -15866 395921 -15810
rect 395977 -15866 396048 -15810
rect 395708 -15952 396048 -15866
rect 395708 -16008 395779 -15952
rect 395835 -16008 395921 -15952
rect 395977 -16008 396048 -15952
rect 395708 -16094 396048 -16008
rect 395708 -16150 395779 -16094
rect 395835 -16150 395921 -16094
rect 395977 -16150 396048 -16094
rect 395708 -16236 396048 -16150
rect 395708 -16292 395779 -16236
rect 395835 -16292 395921 -16236
rect 395977 -16292 396048 -16236
rect 395708 -16378 396048 -16292
rect 395708 -16434 395779 -16378
rect 395835 -16434 395921 -16378
rect 395977 -16434 396048 -16378
rect 395708 -16520 396048 -16434
rect 395708 -16576 395779 -16520
rect 395835 -16576 395921 -16520
rect 395977 -16576 396048 -16520
rect 395708 -16662 396048 -16576
rect 395708 -16718 395779 -16662
rect 395835 -16718 395921 -16662
rect 395977 -16718 396048 -16662
rect 395708 -16804 396048 -16718
rect 395708 -16860 395779 -16804
rect 395835 -16860 395921 -16804
rect 395977 -16860 396048 -16804
rect 395708 -16946 396048 -16860
rect 395708 -17002 395779 -16946
rect 395835 -17002 395921 -16946
rect 395977 -17002 396048 -16946
rect 395708 -17088 396048 -17002
rect 395708 -17144 395779 -17088
rect 395835 -17144 395921 -17088
rect 395977 -17144 396048 -17088
rect 395708 -17230 396048 -17144
rect 395708 -17286 395779 -17230
rect 395835 -17286 395921 -17230
rect 395977 -17286 396048 -17230
rect 395708 -17372 396048 -17286
rect 395708 -17428 395779 -17372
rect 395835 -17428 395921 -17372
rect 395977 -17428 396048 -17372
rect 395708 -17514 396048 -17428
rect 395708 -17570 395779 -17514
rect 395835 -17570 395921 -17514
rect 395977 -17570 396048 -17514
rect 395708 -17656 396048 -17570
rect 395708 -17712 395779 -17656
rect 395835 -17712 395921 -17656
rect 395977 -17712 396048 -17656
rect 395708 -17798 396048 -17712
rect 395708 -17854 395779 -17798
rect 395835 -17854 395921 -17798
rect 395977 -17854 396048 -17798
rect 395708 -17940 396048 -17854
rect 395708 -17996 395779 -17940
rect 395835 -17996 395921 -17940
rect 395977 -17996 396048 -17940
rect 395708 -18082 396048 -17996
rect 395708 -18138 395779 -18082
rect 395835 -18138 395921 -18082
rect 395977 -18138 396048 -18082
rect 395708 -18224 396048 -18138
rect 395708 -18280 395779 -18224
rect 395835 -18280 395921 -18224
rect 395977 -18280 396048 -18224
rect 395708 -18366 396048 -18280
rect 395708 -18422 395779 -18366
rect 395835 -18422 395921 -18366
rect 395977 -18422 396048 -18366
rect 395708 -18508 396048 -18422
rect 395708 -18564 395779 -18508
rect 395835 -18564 395921 -18508
rect 395977 -18564 396048 -18508
rect 395708 -18650 396048 -18564
rect 395708 -18706 395779 -18650
rect 395835 -18706 395921 -18650
rect 395977 -18706 396048 -18650
rect 395708 -18792 396048 -18706
rect 395708 -18848 395779 -18792
rect 395835 -18848 395921 -18792
rect 395977 -18848 396048 -18792
rect 395708 -18934 396048 -18848
rect 395708 -18990 395779 -18934
rect 395835 -18990 395921 -18934
rect 395977 -18990 396048 -18934
rect 395708 -19076 396048 -18990
rect 395708 -19132 395779 -19076
rect 395835 -19132 395921 -19076
rect 395977 -19132 396048 -19076
rect 395708 -19218 396048 -19132
rect 395708 -19274 395779 -19218
rect 395835 -19274 395921 -19218
rect 395977 -19274 396048 -19218
rect 395708 -19360 396048 -19274
rect 395708 -19416 395779 -19360
rect 395835 -19416 395921 -19360
rect 395977 -19416 396048 -19360
rect 395708 -19502 396048 -19416
rect 395708 -19558 395779 -19502
rect 395835 -19558 395921 -19502
rect 395977 -19558 396048 -19502
rect 395708 -19644 396048 -19558
rect 395708 -19700 395779 -19644
rect 395835 -19700 395921 -19644
rect 395977 -19700 396048 -19644
rect 395708 -19786 396048 -19700
rect 395708 -19842 395779 -19786
rect 395835 -19842 395921 -19786
rect 395977 -19842 396048 -19786
rect 395708 -19928 396048 -19842
rect 395708 -19984 395779 -19928
rect 395835 -19984 395921 -19928
rect 395977 -19984 396048 -19928
rect 395708 -20070 396048 -19984
rect 395708 -20126 395779 -20070
rect 395835 -20126 395921 -20070
rect 395977 -20126 396048 -20070
rect 395708 -20212 396048 -20126
rect 395708 -20268 395779 -20212
rect 395835 -20268 395921 -20212
rect 395977 -20268 396048 -20212
rect 395708 -20354 396048 -20268
rect 395708 -20410 395779 -20354
rect 395835 -20410 395921 -20354
rect 395977 -20410 396048 -20354
rect 395708 -20496 396048 -20410
rect 395708 -20552 395779 -20496
rect 395835 -20552 395921 -20496
rect 395977 -20552 396048 -20496
rect 395708 -20638 396048 -20552
rect 395708 -20694 395779 -20638
rect 395835 -20694 395921 -20638
rect 395977 -20694 396048 -20638
rect 395708 -20780 396048 -20694
rect 395708 -20836 395779 -20780
rect 395835 -20836 395921 -20780
rect 395977 -20836 396048 -20780
rect 395708 -20922 396048 -20836
rect 395708 -20978 395779 -20922
rect 395835 -20978 395921 -20922
rect 395977 -20978 396048 -20922
rect 395708 -21064 396048 -20978
rect 395708 -21120 395779 -21064
rect 395835 -21120 395921 -21064
rect 395977 -21120 396048 -21064
rect 395708 -21206 396048 -21120
rect 395708 -21262 395779 -21206
rect 395835 -21262 395921 -21206
rect 395977 -21262 396048 -21206
rect 395708 -21348 396048 -21262
rect 395708 -21404 395779 -21348
rect 395835 -21404 395921 -21348
rect 395977 -21404 396048 -21348
rect 395708 -21490 396048 -21404
rect 395708 -21546 395779 -21490
rect 395835 -21546 395921 -21490
rect 395977 -21546 396048 -21490
rect 395708 -21632 396048 -21546
rect 395708 -21688 395779 -21632
rect 395835 -21688 395921 -21632
rect 395977 -21688 396048 -21632
rect 395708 -21774 396048 -21688
rect 395708 -21830 395779 -21774
rect 395835 -21830 395921 -21774
rect 395977 -21830 396048 -21774
rect 395708 -21916 396048 -21830
rect 395708 -21972 395779 -21916
rect 395835 -21972 395921 -21916
rect 395977 -21972 396048 -21916
rect 395708 -22058 396048 -21972
rect 395708 -22114 395779 -22058
rect 395835 -22114 395921 -22058
rect 395977 -22114 396048 -22058
rect 395708 -22200 396048 -22114
rect 395708 -22256 395779 -22200
rect 395835 -22256 395921 -22200
rect 395977 -22256 396048 -22200
rect 395708 -22342 396048 -22256
rect 395708 -22398 395779 -22342
rect 395835 -22398 395921 -22342
rect 395977 -22398 396048 -22342
rect 395708 -22484 396048 -22398
rect 395708 -22540 395779 -22484
rect 395835 -22540 395921 -22484
rect 395977 -22540 396048 -22484
rect 395708 -22626 396048 -22540
rect 395708 -22682 395779 -22626
rect 395835 -22682 395921 -22626
rect 395977 -22682 396048 -22626
rect 395708 -22768 396048 -22682
rect 395708 -22824 395779 -22768
rect 395835 -22824 395921 -22768
rect 395977 -22824 396048 -22768
rect 395708 -22910 396048 -22824
rect 395708 -22966 395779 -22910
rect 395835 -22966 395921 -22910
rect 395977 -22966 396048 -22910
rect 395708 -23052 396048 -22966
rect 395708 -23108 395779 -23052
rect 395835 -23108 395921 -23052
rect 395977 -23108 396048 -23052
rect 395708 -23194 396048 -23108
rect 395708 -23250 395779 -23194
rect 395835 -23250 395921 -23194
rect 395977 -23250 396048 -23194
rect 395708 -23336 396048 -23250
rect 395708 -23392 395779 -23336
rect 395835 -23392 395921 -23336
rect 395977 -23392 396048 -23336
rect 395708 -23478 396048 -23392
rect 395708 -23534 395779 -23478
rect 395835 -23534 395921 -23478
rect 395977 -23534 396048 -23478
rect 395708 -23620 396048 -23534
rect 395708 -23676 395779 -23620
rect 395835 -23676 395921 -23620
rect 395977 -23676 396048 -23620
rect 395708 -23762 396048 -23676
rect 395708 -23818 395779 -23762
rect 395835 -23818 395921 -23762
rect 395977 -23818 396048 -23762
rect 395708 -23904 396048 -23818
rect 395708 -23960 395779 -23904
rect 395835 -23960 395921 -23904
rect 395977 -23960 396048 -23904
rect 395708 -24046 396048 -23960
rect 395708 -24102 395779 -24046
rect 395835 -24102 395921 -24046
rect 395977 -24102 396048 -24046
rect 395708 -24188 396048 -24102
rect 395708 -24244 395779 -24188
rect 395835 -24244 395921 -24188
rect 395977 -24244 396048 -24188
rect 395708 -24330 396048 -24244
rect 395708 -24386 395779 -24330
rect 395835 -24386 395921 -24330
rect 395977 -24386 396048 -24330
rect 395708 -24472 396048 -24386
rect 395708 -24528 395779 -24472
rect 395835 -24528 395921 -24472
rect 395977 -24528 396048 -24472
rect 395708 -24614 396048 -24528
rect 395708 -24670 395779 -24614
rect 395835 -24670 395921 -24614
rect 395977 -24670 396048 -24614
rect 395708 -24756 396048 -24670
rect 395708 -24812 395779 -24756
rect 395835 -24812 395921 -24756
rect 395977 -24812 396048 -24756
rect 395708 -24898 396048 -24812
rect 395708 -24954 395779 -24898
rect 395835 -24954 395921 -24898
rect 395977 -24954 396048 -24898
rect 395708 -25040 396048 -24954
rect 395708 -25096 395779 -25040
rect 395835 -25096 395921 -25040
rect 395977 -25096 396048 -25040
rect 395708 -25182 396048 -25096
rect 395708 -25238 395779 -25182
rect 395835 -25238 395921 -25182
rect 395977 -25238 396048 -25182
rect 395708 -25324 396048 -25238
rect 395708 -25380 395779 -25324
rect 395835 -25380 395921 -25324
rect 395977 -25380 396048 -25324
rect 395708 -25466 396048 -25380
rect 395708 -25522 395779 -25466
rect 395835 -25522 395921 -25466
rect 395977 -25522 396048 -25466
rect 395708 -25532 396048 -25522
rect 396108 -13680 396448 -13670
rect 396108 -13736 396180 -13680
rect 396236 -13736 396322 -13680
rect 396378 -13736 396448 -13680
rect 396108 -13822 396448 -13736
rect 396108 -13878 396180 -13822
rect 396236 -13878 396322 -13822
rect 396378 -13878 396448 -13822
rect 396108 -13964 396448 -13878
rect 396108 -14020 396180 -13964
rect 396236 -14020 396322 -13964
rect 396378 -14020 396448 -13964
rect 396108 -14106 396448 -14020
rect 396108 -14162 396180 -14106
rect 396236 -14162 396322 -14106
rect 396378 -14162 396448 -14106
rect 396108 -14248 396448 -14162
rect 396108 -14304 396180 -14248
rect 396236 -14304 396322 -14248
rect 396378 -14304 396448 -14248
rect 396108 -14390 396448 -14304
rect 396108 -14446 396180 -14390
rect 396236 -14446 396322 -14390
rect 396378 -14446 396448 -14390
rect 396108 -14532 396448 -14446
rect 396108 -14588 396180 -14532
rect 396236 -14588 396322 -14532
rect 396378 -14588 396448 -14532
rect 396108 -14674 396448 -14588
rect 396108 -14730 396180 -14674
rect 396236 -14730 396322 -14674
rect 396378 -14730 396448 -14674
rect 396108 -14816 396448 -14730
rect 396108 -14872 396180 -14816
rect 396236 -14872 396322 -14816
rect 396378 -14872 396448 -14816
rect 396108 -14958 396448 -14872
rect 396108 -15014 396180 -14958
rect 396236 -15014 396322 -14958
rect 396378 -15014 396448 -14958
rect 396108 -15100 396448 -15014
rect 396108 -15156 396180 -15100
rect 396236 -15156 396322 -15100
rect 396378 -15156 396448 -15100
rect 396108 -15242 396448 -15156
rect 396108 -15298 396180 -15242
rect 396236 -15298 396322 -15242
rect 396378 -15298 396448 -15242
rect 396108 -15384 396448 -15298
rect 396108 -15440 396180 -15384
rect 396236 -15440 396322 -15384
rect 396378 -15440 396448 -15384
rect 396108 -15526 396448 -15440
rect 396108 -15582 396180 -15526
rect 396236 -15582 396322 -15526
rect 396378 -15582 396448 -15526
rect 396108 -15668 396448 -15582
rect 396108 -15724 396180 -15668
rect 396236 -15724 396322 -15668
rect 396378 -15724 396448 -15668
rect 396108 -15810 396448 -15724
rect 396108 -15866 396180 -15810
rect 396236 -15866 396322 -15810
rect 396378 -15866 396448 -15810
rect 396108 -15952 396448 -15866
rect 396108 -16008 396180 -15952
rect 396236 -16008 396322 -15952
rect 396378 -16008 396448 -15952
rect 396108 -16094 396448 -16008
rect 396108 -16150 396180 -16094
rect 396236 -16150 396322 -16094
rect 396378 -16150 396448 -16094
rect 396108 -16236 396448 -16150
rect 396108 -16292 396180 -16236
rect 396236 -16292 396322 -16236
rect 396378 -16292 396448 -16236
rect 396108 -16378 396448 -16292
rect 396108 -16434 396180 -16378
rect 396236 -16434 396322 -16378
rect 396378 -16434 396448 -16378
rect 396108 -16520 396448 -16434
rect 396108 -16576 396180 -16520
rect 396236 -16576 396322 -16520
rect 396378 -16576 396448 -16520
rect 396108 -16662 396448 -16576
rect 396108 -16718 396180 -16662
rect 396236 -16718 396322 -16662
rect 396378 -16718 396448 -16662
rect 396108 -16804 396448 -16718
rect 396108 -16860 396180 -16804
rect 396236 -16860 396322 -16804
rect 396378 -16860 396448 -16804
rect 396108 -16946 396448 -16860
rect 396108 -17002 396180 -16946
rect 396236 -17002 396322 -16946
rect 396378 -17002 396448 -16946
rect 396108 -17088 396448 -17002
rect 396108 -17144 396180 -17088
rect 396236 -17144 396322 -17088
rect 396378 -17144 396448 -17088
rect 396108 -17230 396448 -17144
rect 396108 -17286 396180 -17230
rect 396236 -17286 396322 -17230
rect 396378 -17286 396448 -17230
rect 396108 -17372 396448 -17286
rect 396108 -17428 396180 -17372
rect 396236 -17428 396322 -17372
rect 396378 -17428 396448 -17372
rect 396108 -17514 396448 -17428
rect 396108 -17570 396180 -17514
rect 396236 -17570 396322 -17514
rect 396378 -17570 396448 -17514
rect 396108 -17656 396448 -17570
rect 396108 -17712 396180 -17656
rect 396236 -17712 396322 -17656
rect 396378 -17712 396448 -17656
rect 396108 -17798 396448 -17712
rect 396108 -17854 396180 -17798
rect 396236 -17854 396322 -17798
rect 396378 -17854 396448 -17798
rect 396108 -17940 396448 -17854
rect 396108 -17996 396180 -17940
rect 396236 -17996 396322 -17940
rect 396378 -17996 396448 -17940
rect 396108 -18082 396448 -17996
rect 396108 -18138 396180 -18082
rect 396236 -18138 396322 -18082
rect 396378 -18138 396448 -18082
rect 396108 -18224 396448 -18138
rect 396108 -18280 396180 -18224
rect 396236 -18280 396322 -18224
rect 396378 -18280 396448 -18224
rect 396108 -18366 396448 -18280
rect 396108 -18422 396180 -18366
rect 396236 -18422 396322 -18366
rect 396378 -18422 396448 -18366
rect 396108 -18508 396448 -18422
rect 396108 -18564 396180 -18508
rect 396236 -18564 396322 -18508
rect 396378 -18564 396448 -18508
rect 396108 -18650 396448 -18564
rect 396108 -18706 396180 -18650
rect 396236 -18706 396322 -18650
rect 396378 -18706 396448 -18650
rect 396108 -18792 396448 -18706
rect 396108 -18848 396180 -18792
rect 396236 -18848 396322 -18792
rect 396378 -18848 396448 -18792
rect 396108 -18934 396448 -18848
rect 396108 -18990 396180 -18934
rect 396236 -18990 396322 -18934
rect 396378 -18990 396448 -18934
rect 396108 -19076 396448 -18990
rect 396108 -19132 396180 -19076
rect 396236 -19132 396322 -19076
rect 396378 -19132 396448 -19076
rect 396108 -19218 396448 -19132
rect 396108 -19274 396180 -19218
rect 396236 -19274 396322 -19218
rect 396378 -19274 396448 -19218
rect 396108 -19360 396448 -19274
rect 396108 -19416 396180 -19360
rect 396236 -19416 396322 -19360
rect 396378 -19416 396448 -19360
rect 396108 -19502 396448 -19416
rect 396108 -19558 396180 -19502
rect 396236 -19558 396322 -19502
rect 396378 -19558 396448 -19502
rect 396108 -19644 396448 -19558
rect 396108 -19700 396180 -19644
rect 396236 -19700 396322 -19644
rect 396378 -19700 396448 -19644
rect 396108 -19786 396448 -19700
rect 396108 -19842 396180 -19786
rect 396236 -19842 396322 -19786
rect 396378 -19842 396448 -19786
rect 396108 -19928 396448 -19842
rect 396108 -19984 396180 -19928
rect 396236 -19984 396322 -19928
rect 396378 -19984 396448 -19928
rect 396108 -20070 396448 -19984
rect 396108 -20126 396180 -20070
rect 396236 -20126 396322 -20070
rect 396378 -20126 396448 -20070
rect 396108 -20212 396448 -20126
rect 396108 -20268 396180 -20212
rect 396236 -20268 396322 -20212
rect 396378 -20268 396448 -20212
rect 396108 -20354 396448 -20268
rect 396108 -20410 396180 -20354
rect 396236 -20410 396322 -20354
rect 396378 -20410 396448 -20354
rect 396108 -20496 396448 -20410
rect 396108 -20552 396180 -20496
rect 396236 -20552 396322 -20496
rect 396378 -20552 396448 -20496
rect 396108 -20638 396448 -20552
rect 396108 -20694 396180 -20638
rect 396236 -20694 396322 -20638
rect 396378 -20694 396448 -20638
rect 396108 -20780 396448 -20694
rect 396108 -20836 396180 -20780
rect 396236 -20836 396322 -20780
rect 396378 -20836 396448 -20780
rect 396108 -20922 396448 -20836
rect 396108 -20978 396180 -20922
rect 396236 -20978 396322 -20922
rect 396378 -20978 396448 -20922
rect 396108 -21064 396448 -20978
rect 396108 -21120 396180 -21064
rect 396236 -21120 396322 -21064
rect 396378 -21120 396448 -21064
rect 396108 -21206 396448 -21120
rect 396108 -21262 396180 -21206
rect 396236 -21262 396322 -21206
rect 396378 -21262 396448 -21206
rect 396108 -21348 396448 -21262
rect 396108 -21404 396180 -21348
rect 396236 -21404 396322 -21348
rect 396378 -21404 396448 -21348
rect 396108 -21490 396448 -21404
rect 396108 -21546 396180 -21490
rect 396236 -21546 396322 -21490
rect 396378 -21546 396448 -21490
rect 396108 -21632 396448 -21546
rect 396108 -21688 396180 -21632
rect 396236 -21688 396322 -21632
rect 396378 -21688 396448 -21632
rect 396108 -21774 396448 -21688
rect 396108 -21830 396180 -21774
rect 396236 -21830 396322 -21774
rect 396378 -21830 396448 -21774
rect 396108 -21916 396448 -21830
rect 396108 -21972 396180 -21916
rect 396236 -21972 396322 -21916
rect 396378 -21972 396448 -21916
rect 396108 -22058 396448 -21972
rect 396108 -22114 396180 -22058
rect 396236 -22114 396322 -22058
rect 396378 -22114 396448 -22058
rect 396108 -22200 396448 -22114
rect 396108 -22256 396180 -22200
rect 396236 -22256 396322 -22200
rect 396378 -22256 396448 -22200
rect 396108 -22342 396448 -22256
rect 396108 -22398 396180 -22342
rect 396236 -22398 396322 -22342
rect 396378 -22398 396448 -22342
rect 396108 -22484 396448 -22398
rect 396108 -22540 396180 -22484
rect 396236 -22540 396322 -22484
rect 396378 -22540 396448 -22484
rect 396108 -22626 396448 -22540
rect 396108 -22682 396180 -22626
rect 396236 -22682 396322 -22626
rect 396378 -22682 396448 -22626
rect 396108 -22768 396448 -22682
rect 396108 -22824 396180 -22768
rect 396236 -22824 396322 -22768
rect 396378 -22824 396448 -22768
rect 396108 -22910 396448 -22824
rect 396108 -22966 396180 -22910
rect 396236 -22966 396322 -22910
rect 396378 -22966 396448 -22910
rect 396108 -23052 396448 -22966
rect 396108 -23108 396180 -23052
rect 396236 -23108 396322 -23052
rect 396378 -23108 396448 -23052
rect 396108 -23194 396448 -23108
rect 396108 -23250 396180 -23194
rect 396236 -23250 396322 -23194
rect 396378 -23250 396448 -23194
rect 396108 -23336 396448 -23250
rect 396108 -23392 396180 -23336
rect 396236 -23392 396322 -23336
rect 396378 -23392 396448 -23336
rect 396108 -23478 396448 -23392
rect 396108 -23534 396180 -23478
rect 396236 -23534 396322 -23478
rect 396378 -23534 396448 -23478
rect 396108 -23620 396448 -23534
rect 396108 -23676 396180 -23620
rect 396236 -23676 396322 -23620
rect 396378 -23676 396448 -23620
rect 396108 -23762 396448 -23676
rect 396108 -23818 396180 -23762
rect 396236 -23818 396322 -23762
rect 396378 -23818 396448 -23762
rect 396108 -23904 396448 -23818
rect 396108 -23960 396180 -23904
rect 396236 -23960 396322 -23904
rect 396378 -23960 396448 -23904
rect 396108 -24046 396448 -23960
rect 396108 -24102 396180 -24046
rect 396236 -24102 396322 -24046
rect 396378 -24102 396448 -24046
rect 396108 -24188 396448 -24102
rect 396108 -24244 396180 -24188
rect 396236 -24244 396322 -24188
rect 396378 -24244 396448 -24188
rect 396108 -24330 396448 -24244
rect 396108 -24386 396180 -24330
rect 396236 -24386 396322 -24330
rect 396378 -24386 396448 -24330
rect 396108 -24472 396448 -24386
rect 396108 -24528 396180 -24472
rect 396236 -24528 396322 -24472
rect 396378 -24528 396448 -24472
rect 396108 -24614 396448 -24528
rect 396108 -24670 396180 -24614
rect 396236 -24670 396322 -24614
rect 396378 -24670 396448 -24614
rect 396108 -24756 396448 -24670
rect 396108 -24812 396180 -24756
rect 396236 -24812 396322 -24756
rect 396378 -24812 396448 -24756
rect 396108 -24898 396448 -24812
rect 396108 -24954 396180 -24898
rect 396236 -24954 396322 -24898
rect 396378 -24954 396448 -24898
rect 396108 -25040 396448 -24954
rect 396108 -25096 396180 -25040
rect 396236 -25096 396322 -25040
rect 396378 -25096 396448 -25040
rect 396108 -25182 396448 -25096
rect 396108 -25238 396180 -25182
rect 396236 -25238 396322 -25182
rect 396378 -25238 396448 -25182
rect 396108 -25324 396448 -25238
rect 396108 -25380 396180 -25324
rect 396236 -25380 396322 -25324
rect 396378 -25380 396448 -25324
rect 396108 -25466 396448 -25380
rect 396108 -25522 396180 -25466
rect 396236 -25522 396322 -25466
rect 396378 -25522 396448 -25466
rect 396108 -25532 396448 -25522
rect 396508 -13680 396848 -13670
rect 396508 -13736 396580 -13680
rect 396636 -13736 396722 -13680
rect 396778 -13736 396848 -13680
rect 396508 -13822 396848 -13736
rect 396508 -13878 396580 -13822
rect 396636 -13878 396722 -13822
rect 396778 -13878 396848 -13822
rect 396508 -13964 396848 -13878
rect 396508 -14020 396580 -13964
rect 396636 -14020 396722 -13964
rect 396778 -14020 396848 -13964
rect 396508 -14106 396848 -14020
rect 396508 -14162 396580 -14106
rect 396636 -14162 396722 -14106
rect 396778 -14162 396848 -14106
rect 396508 -14248 396848 -14162
rect 396508 -14304 396580 -14248
rect 396636 -14304 396722 -14248
rect 396778 -14304 396848 -14248
rect 396508 -14390 396848 -14304
rect 396508 -14446 396580 -14390
rect 396636 -14446 396722 -14390
rect 396778 -14446 396848 -14390
rect 396508 -14532 396848 -14446
rect 396508 -14588 396580 -14532
rect 396636 -14588 396722 -14532
rect 396778 -14588 396848 -14532
rect 396508 -14674 396848 -14588
rect 396508 -14730 396580 -14674
rect 396636 -14730 396722 -14674
rect 396778 -14730 396848 -14674
rect 396508 -14816 396848 -14730
rect 396508 -14872 396580 -14816
rect 396636 -14872 396722 -14816
rect 396778 -14872 396848 -14816
rect 396508 -14958 396848 -14872
rect 396508 -15014 396580 -14958
rect 396636 -15014 396722 -14958
rect 396778 -15014 396848 -14958
rect 396508 -15100 396848 -15014
rect 396508 -15156 396580 -15100
rect 396636 -15156 396722 -15100
rect 396778 -15156 396848 -15100
rect 396508 -15242 396848 -15156
rect 396508 -15298 396580 -15242
rect 396636 -15298 396722 -15242
rect 396778 -15298 396848 -15242
rect 396508 -15384 396848 -15298
rect 396508 -15440 396580 -15384
rect 396636 -15440 396722 -15384
rect 396778 -15440 396848 -15384
rect 396508 -15526 396848 -15440
rect 396508 -15582 396580 -15526
rect 396636 -15582 396722 -15526
rect 396778 -15582 396848 -15526
rect 396508 -15668 396848 -15582
rect 396508 -15724 396580 -15668
rect 396636 -15724 396722 -15668
rect 396778 -15724 396848 -15668
rect 396508 -15810 396848 -15724
rect 396508 -15866 396580 -15810
rect 396636 -15866 396722 -15810
rect 396778 -15866 396848 -15810
rect 396508 -15952 396848 -15866
rect 396508 -16008 396580 -15952
rect 396636 -16008 396722 -15952
rect 396778 -16008 396848 -15952
rect 396508 -16094 396848 -16008
rect 396508 -16150 396580 -16094
rect 396636 -16150 396722 -16094
rect 396778 -16150 396848 -16094
rect 396508 -16236 396848 -16150
rect 396508 -16292 396580 -16236
rect 396636 -16292 396722 -16236
rect 396778 -16292 396848 -16236
rect 396508 -16378 396848 -16292
rect 396508 -16434 396580 -16378
rect 396636 -16434 396722 -16378
rect 396778 -16434 396848 -16378
rect 396508 -16520 396848 -16434
rect 396508 -16576 396580 -16520
rect 396636 -16576 396722 -16520
rect 396778 -16576 396848 -16520
rect 396508 -16662 396848 -16576
rect 396508 -16718 396580 -16662
rect 396636 -16718 396722 -16662
rect 396778 -16718 396848 -16662
rect 396508 -16804 396848 -16718
rect 396508 -16860 396580 -16804
rect 396636 -16860 396722 -16804
rect 396778 -16860 396848 -16804
rect 396508 -16946 396848 -16860
rect 396508 -17002 396580 -16946
rect 396636 -17002 396722 -16946
rect 396778 -17002 396848 -16946
rect 396508 -17088 396848 -17002
rect 396508 -17144 396580 -17088
rect 396636 -17144 396722 -17088
rect 396778 -17144 396848 -17088
rect 396508 -17230 396848 -17144
rect 396508 -17286 396580 -17230
rect 396636 -17286 396722 -17230
rect 396778 -17286 396848 -17230
rect 396508 -17372 396848 -17286
rect 396508 -17428 396580 -17372
rect 396636 -17428 396722 -17372
rect 396778 -17428 396848 -17372
rect 396508 -17514 396848 -17428
rect 396508 -17570 396580 -17514
rect 396636 -17570 396722 -17514
rect 396778 -17570 396848 -17514
rect 396508 -17656 396848 -17570
rect 396508 -17712 396580 -17656
rect 396636 -17712 396722 -17656
rect 396778 -17712 396848 -17656
rect 396508 -17798 396848 -17712
rect 396508 -17854 396580 -17798
rect 396636 -17854 396722 -17798
rect 396778 -17854 396848 -17798
rect 396508 -17940 396848 -17854
rect 396508 -17996 396580 -17940
rect 396636 -17996 396722 -17940
rect 396778 -17996 396848 -17940
rect 396508 -18082 396848 -17996
rect 396508 -18138 396580 -18082
rect 396636 -18138 396722 -18082
rect 396778 -18138 396848 -18082
rect 396508 -18224 396848 -18138
rect 396508 -18280 396580 -18224
rect 396636 -18280 396722 -18224
rect 396778 -18280 396848 -18224
rect 396508 -18366 396848 -18280
rect 396508 -18422 396580 -18366
rect 396636 -18422 396722 -18366
rect 396778 -18422 396848 -18366
rect 396508 -18508 396848 -18422
rect 396508 -18564 396580 -18508
rect 396636 -18564 396722 -18508
rect 396778 -18564 396848 -18508
rect 396508 -18650 396848 -18564
rect 396508 -18706 396580 -18650
rect 396636 -18706 396722 -18650
rect 396778 -18706 396848 -18650
rect 396508 -18792 396848 -18706
rect 396508 -18848 396580 -18792
rect 396636 -18848 396722 -18792
rect 396778 -18848 396848 -18792
rect 396508 -18934 396848 -18848
rect 396508 -18990 396580 -18934
rect 396636 -18990 396722 -18934
rect 396778 -18990 396848 -18934
rect 396508 -19076 396848 -18990
rect 396508 -19132 396580 -19076
rect 396636 -19132 396722 -19076
rect 396778 -19132 396848 -19076
rect 396508 -19218 396848 -19132
rect 396508 -19274 396580 -19218
rect 396636 -19274 396722 -19218
rect 396778 -19274 396848 -19218
rect 396508 -19360 396848 -19274
rect 396508 -19416 396580 -19360
rect 396636 -19416 396722 -19360
rect 396778 -19416 396848 -19360
rect 396508 -19502 396848 -19416
rect 396508 -19558 396580 -19502
rect 396636 -19558 396722 -19502
rect 396778 -19558 396848 -19502
rect 396508 -19644 396848 -19558
rect 396508 -19700 396580 -19644
rect 396636 -19700 396722 -19644
rect 396778 -19700 396848 -19644
rect 396508 -19786 396848 -19700
rect 396508 -19842 396580 -19786
rect 396636 -19842 396722 -19786
rect 396778 -19842 396848 -19786
rect 396508 -19928 396848 -19842
rect 396508 -19984 396580 -19928
rect 396636 -19984 396722 -19928
rect 396778 -19984 396848 -19928
rect 396508 -20070 396848 -19984
rect 396508 -20126 396580 -20070
rect 396636 -20126 396722 -20070
rect 396778 -20126 396848 -20070
rect 396508 -20212 396848 -20126
rect 396508 -20268 396580 -20212
rect 396636 -20268 396722 -20212
rect 396778 -20268 396848 -20212
rect 396508 -20354 396848 -20268
rect 396508 -20410 396580 -20354
rect 396636 -20410 396722 -20354
rect 396778 -20410 396848 -20354
rect 396508 -20496 396848 -20410
rect 396508 -20552 396580 -20496
rect 396636 -20552 396722 -20496
rect 396778 -20552 396848 -20496
rect 396508 -20638 396848 -20552
rect 396508 -20694 396580 -20638
rect 396636 -20694 396722 -20638
rect 396778 -20694 396848 -20638
rect 396508 -20780 396848 -20694
rect 396508 -20836 396580 -20780
rect 396636 -20836 396722 -20780
rect 396778 -20836 396848 -20780
rect 396508 -20922 396848 -20836
rect 396508 -20978 396580 -20922
rect 396636 -20978 396722 -20922
rect 396778 -20978 396848 -20922
rect 396508 -21064 396848 -20978
rect 396508 -21120 396580 -21064
rect 396636 -21120 396722 -21064
rect 396778 -21120 396848 -21064
rect 396508 -21206 396848 -21120
rect 396508 -21262 396580 -21206
rect 396636 -21262 396722 -21206
rect 396778 -21262 396848 -21206
rect 396508 -21348 396848 -21262
rect 396508 -21404 396580 -21348
rect 396636 -21404 396722 -21348
rect 396778 -21404 396848 -21348
rect 396508 -21490 396848 -21404
rect 396508 -21546 396580 -21490
rect 396636 -21546 396722 -21490
rect 396778 -21546 396848 -21490
rect 396508 -21632 396848 -21546
rect 396508 -21688 396580 -21632
rect 396636 -21688 396722 -21632
rect 396778 -21688 396848 -21632
rect 396508 -21774 396848 -21688
rect 396508 -21830 396580 -21774
rect 396636 -21830 396722 -21774
rect 396778 -21830 396848 -21774
rect 396508 -21916 396848 -21830
rect 396508 -21972 396580 -21916
rect 396636 -21972 396722 -21916
rect 396778 -21972 396848 -21916
rect 396508 -22058 396848 -21972
rect 396508 -22114 396580 -22058
rect 396636 -22114 396722 -22058
rect 396778 -22114 396848 -22058
rect 396508 -22200 396848 -22114
rect 396508 -22256 396580 -22200
rect 396636 -22256 396722 -22200
rect 396778 -22256 396848 -22200
rect 396508 -22342 396848 -22256
rect 396508 -22398 396580 -22342
rect 396636 -22398 396722 -22342
rect 396778 -22398 396848 -22342
rect 396508 -22484 396848 -22398
rect 396508 -22540 396580 -22484
rect 396636 -22540 396722 -22484
rect 396778 -22540 396848 -22484
rect 396508 -22626 396848 -22540
rect 396508 -22682 396580 -22626
rect 396636 -22682 396722 -22626
rect 396778 -22682 396848 -22626
rect 396508 -22768 396848 -22682
rect 396508 -22824 396580 -22768
rect 396636 -22824 396722 -22768
rect 396778 -22824 396848 -22768
rect 396508 -22910 396848 -22824
rect 396508 -22966 396580 -22910
rect 396636 -22966 396722 -22910
rect 396778 -22966 396848 -22910
rect 396508 -23052 396848 -22966
rect 396508 -23108 396580 -23052
rect 396636 -23108 396722 -23052
rect 396778 -23108 396848 -23052
rect 396508 -23194 396848 -23108
rect 396508 -23250 396580 -23194
rect 396636 -23250 396722 -23194
rect 396778 -23250 396848 -23194
rect 396508 -23336 396848 -23250
rect 396508 -23392 396580 -23336
rect 396636 -23392 396722 -23336
rect 396778 -23392 396848 -23336
rect 396508 -23478 396848 -23392
rect 396508 -23534 396580 -23478
rect 396636 -23534 396722 -23478
rect 396778 -23534 396848 -23478
rect 396508 -23620 396848 -23534
rect 396508 -23676 396580 -23620
rect 396636 -23676 396722 -23620
rect 396778 -23676 396848 -23620
rect 396508 -23762 396848 -23676
rect 396508 -23818 396580 -23762
rect 396636 -23818 396722 -23762
rect 396778 -23818 396848 -23762
rect 396508 -23904 396848 -23818
rect 396508 -23960 396580 -23904
rect 396636 -23960 396722 -23904
rect 396778 -23960 396848 -23904
rect 396508 -24046 396848 -23960
rect 396508 -24102 396580 -24046
rect 396636 -24102 396722 -24046
rect 396778 -24102 396848 -24046
rect 396508 -24188 396848 -24102
rect 396508 -24244 396580 -24188
rect 396636 -24244 396722 -24188
rect 396778 -24244 396848 -24188
rect 396508 -24330 396848 -24244
rect 396508 -24386 396580 -24330
rect 396636 -24386 396722 -24330
rect 396778 -24386 396848 -24330
rect 396508 -24472 396848 -24386
rect 396508 -24528 396580 -24472
rect 396636 -24528 396722 -24472
rect 396778 -24528 396848 -24472
rect 396508 -24614 396848 -24528
rect 396508 -24670 396580 -24614
rect 396636 -24670 396722 -24614
rect 396778 -24670 396848 -24614
rect 396508 -24756 396848 -24670
rect 396508 -24812 396580 -24756
rect 396636 -24812 396722 -24756
rect 396778 -24812 396848 -24756
rect 396508 -24898 396848 -24812
rect 396508 -24954 396580 -24898
rect 396636 -24954 396722 -24898
rect 396778 -24954 396848 -24898
rect 396508 -25040 396848 -24954
rect 396508 -25096 396580 -25040
rect 396636 -25096 396722 -25040
rect 396778 -25096 396848 -25040
rect 396508 -25182 396848 -25096
rect 396508 -25238 396580 -25182
rect 396636 -25238 396722 -25182
rect 396778 -25238 396848 -25182
rect 396508 -25324 396848 -25238
rect 396508 -25380 396580 -25324
rect 396636 -25380 396722 -25324
rect 396778 -25380 396848 -25324
rect 396508 -25466 396848 -25380
rect 396508 -25522 396580 -25466
rect 396636 -25522 396722 -25466
rect 396778 -25522 396848 -25466
rect 396508 -25532 396848 -25522
rect 396908 -13680 397248 -13670
rect 396908 -13736 396977 -13680
rect 397033 -13736 397119 -13680
rect 397175 -13736 397248 -13680
rect 396908 -13822 397248 -13736
rect 396908 -13878 396977 -13822
rect 397033 -13878 397119 -13822
rect 397175 -13878 397248 -13822
rect 396908 -13964 397248 -13878
rect 396908 -14020 396977 -13964
rect 397033 -14020 397119 -13964
rect 397175 -14020 397248 -13964
rect 396908 -14106 397248 -14020
rect 396908 -14162 396977 -14106
rect 397033 -14162 397119 -14106
rect 397175 -14162 397248 -14106
rect 396908 -14248 397248 -14162
rect 396908 -14304 396977 -14248
rect 397033 -14304 397119 -14248
rect 397175 -14304 397248 -14248
rect 396908 -14390 397248 -14304
rect 396908 -14446 396977 -14390
rect 397033 -14446 397119 -14390
rect 397175 -14446 397248 -14390
rect 396908 -14532 397248 -14446
rect 396908 -14588 396977 -14532
rect 397033 -14588 397119 -14532
rect 397175 -14588 397248 -14532
rect 396908 -14674 397248 -14588
rect 396908 -14730 396977 -14674
rect 397033 -14730 397119 -14674
rect 397175 -14730 397248 -14674
rect 396908 -14816 397248 -14730
rect 396908 -14872 396977 -14816
rect 397033 -14872 397119 -14816
rect 397175 -14872 397248 -14816
rect 396908 -14958 397248 -14872
rect 396908 -15014 396977 -14958
rect 397033 -15014 397119 -14958
rect 397175 -15014 397248 -14958
rect 396908 -15100 397248 -15014
rect 396908 -15156 396977 -15100
rect 397033 -15156 397119 -15100
rect 397175 -15156 397248 -15100
rect 396908 -15242 397248 -15156
rect 396908 -15298 396977 -15242
rect 397033 -15298 397119 -15242
rect 397175 -15298 397248 -15242
rect 396908 -15384 397248 -15298
rect 396908 -15440 396977 -15384
rect 397033 -15440 397119 -15384
rect 397175 -15440 397248 -15384
rect 396908 -15526 397248 -15440
rect 396908 -15582 396977 -15526
rect 397033 -15582 397119 -15526
rect 397175 -15582 397248 -15526
rect 396908 -15668 397248 -15582
rect 396908 -15724 396977 -15668
rect 397033 -15724 397119 -15668
rect 397175 -15724 397248 -15668
rect 396908 -15810 397248 -15724
rect 396908 -15866 396977 -15810
rect 397033 -15866 397119 -15810
rect 397175 -15866 397248 -15810
rect 396908 -15952 397248 -15866
rect 396908 -16008 396977 -15952
rect 397033 -16008 397119 -15952
rect 397175 -16008 397248 -15952
rect 396908 -16094 397248 -16008
rect 396908 -16150 396977 -16094
rect 397033 -16150 397119 -16094
rect 397175 -16150 397248 -16094
rect 396908 -16236 397248 -16150
rect 396908 -16292 396977 -16236
rect 397033 -16292 397119 -16236
rect 397175 -16292 397248 -16236
rect 396908 -16378 397248 -16292
rect 396908 -16434 396977 -16378
rect 397033 -16434 397119 -16378
rect 397175 -16434 397248 -16378
rect 396908 -16520 397248 -16434
rect 396908 -16576 396977 -16520
rect 397033 -16576 397119 -16520
rect 397175 -16576 397248 -16520
rect 396908 -16662 397248 -16576
rect 396908 -16718 396977 -16662
rect 397033 -16718 397119 -16662
rect 397175 -16718 397248 -16662
rect 396908 -16804 397248 -16718
rect 396908 -16860 396977 -16804
rect 397033 -16860 397119 -16804
rect 397175 -16860 397248 -16804
rect 396908 -16946 397248 -16860
rect 396908 -17002 396977 -16946
rect 397033 -17002 397119 -16946
rect 397175 -17002 397248 -16946
rect 396908 -17088 397248 -17002
rect 396908 -17144 396977 -17088
rect 397033 -17144 397119 -17088
rect 397175 -17144 397248 -17088
rect 396908 -17230 397248 -17144
rect 396908 -17286 396977 -17230
rect 397033 -17286 397119 -17230
rect 397175 -17286 397248 -17230
rect 396908 -17372 397248 -17286
rect 396908 -17428 396977 -17372
rect 397033 -17428 397119 -17372
rect 397175 -17428 397248 -17372
rect 396908 -17514 397248 -17428
rect 396908 -17570 396977 -17514
rect 397033 -17570 397119 -17514
rect 397175 -17570 397248 -17514
rect 396908 -17656 397248 -17570
rect 396908 -17712 396977 -17656
rect 397033 -17712 397119 -17656
rect 397175 -17712 397248 -17656
rect 396908 -17798 397248 -17712
rect 396908 -17854 396977 -17798
rect 397033 -17854 397119 -17798
rect 397175 -17854 397248 -17798
rect 396908 -17940 397248 -17854
rect 396908 -17996 396977 -17940
rect 397033 -17996 397119 -17940
rect 397175 -17996 397248 -17940
rect 396908 -18082 397248 -17996
rect 396908 -18138 396977 -18082
rect 397033 -18138 397119 -18082
rect 397175 -18138 397248 -18082
rect 396908 -18224 397248 -18138
rect 396908 -18280 396977 -18224
rect 397033 -18280 397119 -18224
rect 397175 -18280 397248 -18224
rect 396908 -18366 397248 -18280
rect 396908 -18422 396977 -18366
rect 397033 -18422 397119 -18366
rect 397175 -18422 397248 -18366
rect 396908 -18508 397248 -18422
rect 396908 -18564 396977 -18508
rect 397033 -18564 397119 -18508
rect 397175 -18564 397248 -18508
rect 396908 -18650 397248 -18564
rect 396908 -18706 396977 -18650
rect 397033 -18706 397119 -18650
rect 397175 -18706 397248 -18650
rect 396908 -18792 397248 -18706
rect 396908 -18848 396977 -18792
rect 397033 -18848 397119 -18792
rect 397175 -18848 397248 -18792
rect 396908 -18934 397248 -18848
rect 396908 -18990 396977 -18934
rect 397033 -18990 397119 -18934
rect 397175 -18990 397248 -18934
rect 396908 -19076 397248 -18990
rect 396908 -19132 396977 -19076
rect 397033 -19132 397119 -19076
rect 397175 -19132 397248 -19076
rect 396908 -19218 397248 -19132
rect 396908 -19274 396977 -19218
rect 397033 -19274 397119 -19218
rect 397175 -19274 397248 -19218
rect 396908 -19360 397248 -19274
rect 396908 -19416 396977 -19360
rect 397033 -19416 397119 -19360
rect 397175 -19416 397248 -19360
rect 396908 -19502 397248 -19416
rect 396908 -19558 396977 -19502
rect 397033 -19558 397119 -19502
rect 397175 -19558 397248 -19502
rect 396908 -19644 397248 -19558
rect 396908 -19700 396977 -19644
rect 397033 -19700 397119 -19644
rect 397175 -19700 397248 -19644
rect 396908 -19786 397248 -19700
rect 396908 -19842 396977 -19786
rect 397033 -19842 397119 -19786
rect 397175 -19842 397248 -19786
rect 396908 -19928 397248 -19842
rect 396908 -19984 396977 -19928
rect 397033 -19984 397119 -19928
rect 397175 -19984 397248 -19928
rect 396908 -20070 397248 -19984
rect 396908 -20126 396977 -20070
rect 397033 -20126 397119 -20070
rect 397175 -20126 397248 -20070
rect 396908 -20212 397248 -20126
rect 396908 -20268 396977 -20212
rect 397033 -20268 397119 -20212
rect 397175 -20268 397248 -20212
rect 396908 -20354 397248 -20268
rect 396908 -20410 396977 -20354
rect 397033 -20410 397119 -20354
rect 397175 -20410 397248 -20354
rect 396908 -20496 397248 -20410
rect 396908 -20552 396977 -20496
rect 397033 -20552 397119 -20496
rect 397175 -20552 397248 -20496
rect 396908 -20638 397248 -20552
rect 396908 -20694 396977 -20638
rect 397033 -20694 397119 -20638
rect 397175 -20694 397248 -20638
rect 396908 -20780 397248 -20694
rect 396908 -20836 396977 -20780
rect 397033 -20836 397119 -20780
rect 397175 -20836 397248 -20780
rect 396908 -20922 397248 -20836
rect 396908 -20978 396977 -20922
rect 397033 -20978 397119 -20922
rect 397175 -20978 397248 -20922
rect 396908 -21064 397248 -20978
rect 396908 -21120 396977 -21064
rect 397033 -21120 397119 -21064
rect 397175 -21120 397248 -21064
rect 396908 -21206 397248 -21120
rect 396908 -21262 396977 -21206
rect 397033 -21262 397119 -21206
rect 397175 -21262 397248 -21206
rect 396908 -21348 397248 -21262
rect 396908 -21404 396977 -21348
rect 397033 -21404 397119 -21348
rect 397175 -21404 397248 -21348
rect 396908 -21490 397248 -21404
rect 396908 -21546 396977 -21490
rect 397033 -21546 397119 -21490
rect 397175 -21546 397248 -21490
rect 396908 -21632 397248 -21546
rect 396908 -21688 396977 -21632
rect 397033 -21688 397119 -21632
rect 397175 -21688 397248 -21632
rect 396908 -21774 397248 -21688
rect 396908 -21830 396977 -21774
rect 397033 -21830 397119 -21774
rect 397175 -21830 397248 -21774
rect 396908 -21916 397248 -21830
rect 396908 -21972 396977 -21916
rect 397033 -21972 397119 -21916
rect 397175 -21972 397248 -21916
rect 396908 -22058 397248 -21972
rect 396908 -22114 396977 -22058
rect 397033 -22114 397119 -22058
rect 397175 -22114 397248 -22058
rect 396908 -22200 397248 -22114
rect 396908 -22256 396977 -22200
rect 397033 -22256 397119 -22200
rect 397175 -22256 397248 -22200
rect 396908 -22342 397248 -22256
rect 396908 -22398 396977 -22342
rect 397033 -22398 397119 -22342
rect 397175 -22398 397248 -22342
rect 396908 -22484 397248 -22398
rect 396908 -22540 396977 -22484
rect 397033 -22540 397119 -22484
rect 397175 -22540 397248 -22484
rect 396908 -22626 397248 -22540
rect 396908 -22682 396977 -22626
rect 397033 -22682 397119 -22626
rect 397175 -22682 397248 -22626
rect 396908 -22768 397248 -22682
rect 396908 -22824 396977 -22768
rect 397033 -22824 397119 -22768
rect 397175 -22824 397248 -22768
rect 396908 -22910 397248 -22824
rect 396908 -22966 396977 -22910
rect 397033 -22966 397119 -22910
rect 397175 -22966 397248 -22910
rect 396908 -23052 397248 -22966
rect 396908 -23108 396977 -23052
rect 397033 -23108 397119 -23052
rect 397175 -23108 397248 -23052
rect 396908 -23194 397248 -23108
rect 396908 -23250 396977 -23194
rect 397033 -23250 397119 -23194
rect 397175 -23250 397248 -23194
rect 396908 -23336 397248 -23250
rect 396908 -23392 396977 -23336
rect 397033 -23392 397119 -23336
rect 397175 -23392 397248 -23336
rect 396908 -23478 397248 -23392
rect 396908 -23534 396977 -23478
rect 397033 -23534 397119 -23478
rect 397175 -23534 397248 -23478
rect 396908 -23620 397248 -23534
rect 396908 -23676 396977 -23620
rect 397033 -23676 397119 -23620
rect 397175 -23676 397248 -23620
rect 396908 -23762 397248 -23676
rect 396908 -23818 396977 -23762
rect 397033 -23818 397119 -23762
rect 397175 -23818 397248 -23762
rect 396908 -23904 397248 -23818
rect 396908 -23960 396977 -23904
rect 397033 -23960 397119 -23904
rect 397175 -23960 397248 -23904
rect 396908 -24046 397248 -23960
rect 396908 -24102 396977 -24046
rect 397033 -24102 397119 -24046
rect 397175 -24102 397248 -24046
rect 396908 -24188 397248 -24102
rect 396908 -24244 396977 -24188
rect 397033 -24244 397119 -24188
rect 397175 -24244 397248 -24188
rect 396908 -24330 397248 -24244
rect 396908 -24386 396977 -24330
rect 397033 -24386 397119 -24330
rect 397175 -24386 397248 -24330
rect 396908 -24472 397248 -24386
rect 396908 -24528 396977 -24472
rect 397033 -24528 397119 -24472
rect 397175 -24528 397248 -24472
rect 396908 -24614 397248 -24528
rect 396908 -24670 396977 -24614
rect 397033 -24670 397119 -24614
rect 397175 -24670 397248 -24614
rect 396908 -24756 397248 -24670
rect 396908 -24812 396977 -24756
rect 397033 -24812 397119 -24756
rect 397175 -24812 397248 -24756
rect 396908 -24898 397248 -24812
rect 396908 -24954 396977 -24898
rect 397033 -24954 397119 -24898
rect 397175 -24954 397248 -24898
rect 396908 -25040 397248 -24954
rect 396908 -25096 396977 -25040
rect 397033 -25096 397119 -25040
rect 397175 -25096 397248 -25040
rect 396908 -25182 397248 -25096
rect 396908 -25238 396977 -25182
rect 397033 -25238 397119 -25182
rect 397175 -25238 397248 -25182
rect 396908 -25324 397248 -25238
rect 396908 -25380 396977 -25324
rect 397033 -25380 397119 -25324
rect 397175 -25380 397248 -25324
rect 396908 -25466 397248 -25380
rect 396908 -25522 396977 -25466
rect 397033 -25522 397119 -25466
rect 397175 -25522 397248 -25466
rect 396908 -25532 397248 -25522
rect 397308 -13680 397648 -13670
rect 397308 -13736 397374 -13680
rect 397430 -13736 397516 -13680
rect 397572 -13736 397648 -13680
rect 397308 -13822 397648 -13736
rect 397308 -13878 397374 -13822
rect 397430 -13878 397516 -13822
rect 397572 -13878 397648 -13822
rect 397308 -13964 397648 -13878
rect 397308 -14020 397374 -13964
rect 397430 -14020 397516 -13964
rect 397572 -14020 397648 -13964
rect 397308 -14106 397648 -14020
rect 397308 -14162 397374 -14106
rect 397430 -14162 397516 -14106
rect 397572 -14162 397648 -14106
rect 397308 -14248 397648 -14162
rect 397308 -14304 397374 -14248
rect 397430 -14304 397516 -14248
rect 397572 -14304 397648 -14248
rect 397308 -14390 397648 -14304
rect 397308 -14446 397374 -14390
rect 397430 -14446 397516 -14390
rect 397572 -14446 397648 -14390
rect 397308 -14532 397648 -14446
rect 397308 -14588 397374 -14532
rect 397430 -14588 397516 -14532
rect 397572 -14588 397648 -14532
rect 397308 -14674 397648 -14588
rect 397308 -14730 397374 -14674
rect 397430 -14730 397516 -14674
rect 397572 -14730 397648 -14674
rect 397308 -14816 397648 -14730
rect 397308 -14872 397374 -14816
rect 397430 -14872 397516 -14816
rect 397572 -14872 397648 -14816
rect 397308 -14958 397648 -14872
rect 397308 -15014 397374 -14958
rect 397430 -15014 397516 -14958
rect 397572 -15014 397648 -14958
rect 397308 -15100 397648 -15014
rect 397308 -15156 397374 -15100
rect 397430 -15156 397516 -15100
rect 397572 -15156 397648 -15100
rect 397308 -15242 397648 -15156
rect 397308 -15298 397374 -15242
rect 397430 -15298 397516 -15242
rect 397572 -15298 397648 -15242
rect 397308 -15384 397648 -15298
rect 397308 -15440 397374 -15384
rect 397430 -15440 397516 -15384
rect 397572 -15440 397648 -15384
rect 397308 -15526 397648 -15440
rect 397308 -15582 397374 -15526
rect 397430 -15582 397516 -15526
rect 397572 -15582 397648 -15526
rect 397308 -15668 397648 -15582
rect 397308 -15724 397374 -15668
rect 397430 -15724 397516 -15668
rect 397572 -15724 397648 -15668
rect 397308 -15810 397648 -15724
rect 397308 -15866 397374 -15810
rect 397430 -15866 397516 -15810
rect 397572 -15866 397648 -15810
rect 397308 -15952 397648 -15866
rect 397308 -16008 397374 -15952
rect 397430 -16008 397516 -15952
rect 397572 -16008 397648 -15952
rect 397308 -16094 397648 -16008
rect 397308 -16150 397374 -16094
rect 397430 -16150 397516 -16094
rect 397572 -16150 397648 -16094
rect 397308 -16236 397648 -16150
rect 397308 -16292 397374 -16236
rect 397430 -16292 397516 -16236
rect 397572 -16292 397648 -16236
rect 397308 -16378 397648 -16292
rect 397308 -16434 397374 -16378
rect 397430 -16434 397516 -16378
rect 397572 -16434 397648 -16378
rect 397308 -16520 397648 -16434
rect 397308 -16576 397374 -16520
rect 397430 -16576 397516 -16520
rect 397572 -16576 397648 -16520
rect 397308 -16662 397648 -16576
rect 397308 -16718 397374 -16662
rect 397430 -16718 397516 -16662
rect 397572 -16718 397648 -16662
rect 397308 -16804 397648 -16718
rect 397308 -16860 397374 -16804
rect 397430 -16860 397516 -16804
rect 397572 -16860 397648 -16804
rect 397308 -16946 397648 -16860
rect 397308 -17002 397374 -16946
rect 397430 -17002 397516 -16946
rect 397572 -17002 397648 -16946
rect 397308 -17088 397648 -17002
rect 397308 -17144 397374 -17088
rect 397430 -17144 397516 -17088
rect 397572 -17144 397648 -17088
rect 397308 -17230 397648 -17144
rect 397308 -17286 397374 -17230
rect 397430 -17286 397516 -17230
rect 397572 -17286 397648 -17230
rect 397308 -17372 397648 -17286
rect 397308 -17428 397374 -17372
rect 397430 -17428 397516 -17372
rect 397572 -17428 397648 -17372
rect 397308 -17514 397648 -17428
rect 397308 -17570 397374 -17514
rect 397430 -17570 397516 -17514
rect 397572 -17570 397648 -17514
rect 397308 -17656 397648 -17570
rect 397308 -17712 397374 -17656
rect 397430 -17712 397516 -17656
rect 397572 -17712 397648 -17656
rect 397308 -17798 397648 -17712
rect 397308 -17854 397374 -17798
rect 397430 -17854 397516 -17798
rect 397572 -17854 397648 -17798
rect 397308 -17940 397648 -17854
rect 397308 -17996 397374 -17940
rect 397430 -17996 397516 -17940
rect 397572 -17996 397648 -17940
rect 397308 -18082 397648 -17996
rect 397308 -18138 397374 -18082
rect 397430 -18138 397516 -18082
rect 397572 -18138 397648 -18082
rect 397308 -18224 397648 -18138
rect 397308 -18280 397374 -18224
rect 397430 -18280 397516 -18224
rect 397572 -18280 397648 -18224
rect 397308 -18366 397648 -18280
rect 397308 -18422 397374 -18366
rect 397430 -18422 397516 -18366
rect 397572 -18422 397648 -18366
rect 397308 -18508 397648 -18422
rect 397308 -18564 397374 -18508
rect 397430 -18564 397516 -18508
rect 397572 -18564 397648 -18508
rect 397308 -18650 397648 -18564
rect 397308 -18706 397374 -18650
rect 397430 -18706 397516 -18650
rect 397572 -18706 397648 -18650
rect 397308 -18792 397648 -18706
rect 397308 -18848 397374 -18792
rect 397430 -18848 397516 -18792
rect 397572 -18848 397648 -18792
rect 397308 -18934 397648 -18848
rect 397308 -18990 397374 -18934
rect 397430 -18990 397516 -18934
rect 397572 -18990 397648 -18934
rect 397308 -19076 397648 -18990
rect 397308 -19132 397374 -19076
rect 397430 -19132 397516 -19076
rect 397572 -19132 397648 -19076
rect 397308 -19218 397648 -19132
rect 397308 -19274 397374 -19218
rect 397430 -19274 397516 -19218
rect 397572 -19274 397648 -19218
rect 397308 -19360 397648 -19274
rect 397308 -19416 397374 -19360
rect 397430 -19416 397516 -19360
rect 397572 -19416 397648 -19360
rect 397308 -19502 397648 -19416
rect 397308 -19558 397374 -19502
rect 397430 -19558 397516 -19502
rect 397572 -19558 397648 -19502
rect 397308 -19644 397648 -19558
rect 397308 -19700 397374 -19644
rect 397430 -19700 397516 -19644
rect 397572 -19700 397648 -19644
rect 397308 -19786 397648 -19700
rect 397308 -19842 397374 -19786
rect 397430 -19842 397516 -19786
rect 397572 -19842 397648 -19786
rect 397308 -19928 397648 -19842
rect 397308 -19984 397374 -19928
rect 397430 -19984 397516 -19928
rect 397572 -19984 397648 -19928
rect 397308 -20070 397648 -19984
rect 397308 -20126 397374 -20070
rect 397430 -20126 397516 -20070
rect 397572 -20126 397648 -20070
rect 397308 -20212 397648 -20126
rect 397308 -20268 397374 -20212
rect 397430 -20268 397516 -20212
rect 397572 -20268 397648 -20212
rect 397308 -20354 397648 -20268
rect 397308 -20410 397374 -20354
rect 397430 -20410 397516 -20354
rect 397572 -20410 397648 -20354
rect 397308 -20496 397648 -20410
rect 397308 -20552 397374 -20496
rect 397430 -20552 397516 -20496
rect 397572 -20552 397648 -20496
rect 397308 -20638 397648 -20552
rect 397308 -20694 397374 -20638
rect 397430 -20694 397516 -20638
rect 397572 -20694 397648 -20638
rect 397308 -20780 397648 -20694
rect 397308 -20836 397374 -20780
rect 397430 -20836 397516 -20780
rect 397572 -20836 397648 -20780
rect 397308 -20922 397648 -20836
rect 397308 -20978 397374 -20922
rect 397430 -20978 397516 -20922
rect 397572 -20978 397648 -20922
rect 397308 -21064 397648 -20978
rect 397308 -21120 397374 -21064
rect 397430 -21120 397516 -21064
rect 397572 -21120 397648 -21064
rect 397308 -21206 397648 -21120
rect 397308 -21262 397374 -21206
rect 397430 -21262 397516 -21206
rect 397572 -21262 397648 -21206
rect 397308 -21348 397648 -21262
rect 397308 -21404 397374 -21348
rect 397430 -21404 397516 -21348
rect 397572 -21404 397648 -21348
rect 397308 -21490 397648 -21404
rect 397308 -21546 397374 -21490
rect 397430 -21546 397516 -21490
rect 397572 -21546 397648 -21490
rect 397308 -21632 397648 -21546
rect 397308 -21688 397374 -21632
rect 397430 -21688 397516 -21632
rect 397572 -21688 397648 -21632
rect 397308 -21774 397648 -21688
rect 397308 -21830 397374 -21774
rect 397430 -21830 397516 -21774
rect 397572 -21830 397648 -21774
rect 397308 -21916 397648 -21830
rect 397308 -21972 397374 -21916
rect 397430 -21972 397516 -21916
rect 397572 -21972 397648 -21916
rect 397308 -22058 397648 -21972
rect 397308 -22114 397374 -22058
rect 397430 -22114 397516 -22058
rect 397572 -22114 397648 -22058
rect 397308 -22200 397648 -22114
rect 397308 -22256 397374 -22200
rect 397430 -22256 397516 -22200
rect 397572 -22256 397648 -22200
rect 397308 -22342 397648 -22256
rect 397308 -22398 397374 -22342
rect 397430 -22398 397516 -22342
rect 397572 -22398 397648 -22342
rect 397308 -22484 397648 -22398
rect 397308 -22540 397374 -22484
rect 397430 -22540 397516 -22484
rect 397572 -22540 397648 -22484
rect 397308 -22626 397648 -22540
rect 397308 -22682 397374 -22626
rect 397430 -22682 397516 -22626
rect 397572 -22682 397648 -22626
rect 397308 -22768 397648 -22682
rect 397308 -22824 397374 -22768
rect 397430 -22824 397516 -22768
rect 397572 -22824 397648 -22768
rect 397308 -22910 397648 -22824
rect 397308 -22966 397374 -22910
rect 397430 -22966 397516 -22910
rect 397572 -22966 397648 -22910
rect 397308 -23052 397648 -22966
rect 397308 -23108 397374 -23052
rect 397430 -23108 397516 -23052
rect 397572 -23108 397648 -23052
rect 397308 -23194 397648 -23108
rect 397308 -23250 397374 -23194
rect 397430 -23250 397516 -23194
rect 397572 -23250 397648 -23194
rect 397308 -23336 397648 -23250
rect 397308 -23392 397374 -23336
rect 397430 -23392 397516 -23336
rect 397572 -23392 397648 -23336
rect 397308 -23478 397648 -23392
rect 397308 -23534 397374 -23478
rect 397430 -23534 397516 -23478
rect 397572 -23534 397648 -23478
rect 397308 -23620 397648 -23534
rect 397308 -23676 397374 -23620
rect 397430 -23676 397516 -23620
rect 397572 -23676 397648 -23620
rect 397308 -23762 397648 -23676
rect 397308 -23818 397374 -23762
rect 397430 -23818 397516 -23762
rect 397572 -23818 397648 -23762
rect 397308 -23904 397648 -23818
rect 397308 -23960 397374 -23904
rect 397430 -23960 397516 -23904
rect 397572 -23960 397648 -23904
rect 397308 -24046 397648 -23960
rect 397308 -24102 397374 -24046
rect 397430 -24102 397516 -24046
rect 397572 -24102 397648 -24046
rect 397308 -24188 397648 -24102
rect 397308 -24244 397374 -24188
rect 397430 -24244 397516 -24188
rect 397572 -24244 397648 -24188
rect 397308 -24330 397648 -24244
rect 397308 -24386 397374 -24330
rect 397430 -24386 397516 -24330
rect 397572 -24386 397648 -24330
rect 397308 -24472 397648 -24386
rect 397308 -24528 397374 -24472
rect 397430 -24528 397516 -24472
rect 397572 -24528 397648 -24472
rect 397308 -24614 397648 -24528
rect 397308 -24670 397374 -24614
rect 397430 -24670 397516 -24614
rect 397572 -24670 397648 -24614
rect 397308 -24756 397648 -24670
rect 397308 -24812 397374 -24756
rect 397430 -24812 397516 -24756
rect 397572 -24812 397648 -24756
rect 397308 -24898 397648 -24812
rect 397308 -24954 397374 -24898
rect 397430 -24954 397516 -24898
rect 397572 -24954 397648 -24898
rect 397308 -25040 397648 -24954
rect 397308 -25096 397374 -25040
rect 397430 -25096 397516 -25040
rect 397572 -25096 397648 -25040
rect 397308 -25182 397648 -25096
rect 397308 -25238 397374 -25182
rect 397430 -25238 397516 -25182
rect 397572 -25238 397648 -25182
rect 397308 -25324 397648 -25238
rect 397308 -25380 397374 -25324
rect 397430 -25380 397516 -25324
rect 397572 -25380 397648 -25324
rect 397308 -25466 397648 -25380
rect 397308 -25522 397374 -25466
rect 397430 -25522 397516 -25466
rect 397572 -25522 397648 -25466
rect 397308 -25532 397648 -25522
rect 397708 -13680 398048 -13670
rect 397708 -13736 397778 -13680
rect 397834 -13736 397920 -13680
rect 397976 -13736 398048 -13680
rect 397708 -13822 398048 -13736
rect 397708 -13878 397778 -13822
rect 397834 -13878 397920 -13822
rect 397976 -13878 398048 -13822
rect 397708 -13964 398048 -13878
rect 397708 -14020 397778 -13964
rect 397834 -14020 397920 -13964
rect 397976 -14020 398048 -13964
rect 397708 -14106 398048 -14020
rect 397708 -14162 397778 -14106
rect 397834 -14162 397920 -14106
rect 397976 -14162 398048 -14106
rect 397708 -14248 398048 -14162
rect 397708 -14304 397778 -14248
rect 397834 -14304 397920 -14248
rect 397976 -14304 398048 -14248
rect 397708 -14390 398048 -14304
rect 397708 -14446 397778 -14390
rect 397834 -14446 397920 -14390
rect 397976 -14446 398048 -14390
rect 397708 -14532 398048 -14446
rect 397708 -14588 397778 -14532
rect 397834 -14588 397920 -14532
rect 397976 -14588 398048 -14532
rect 397708 -14674 398048 -14588
rect 397708 -14730 397778 -14674
rect 397834 -14730 397920 -14674
rect 397976 -14730 398048 -14674
rect 397708 -14816 398048 -14730
rect 397708 -14872 397778 -14816
rect 397834 -14872 397920 -14816
rect 397976 -14872 398048 -14816
rect 397708 -14958 398048 -14872
rect 397708 -15014 397778 -14958
rect 397834 -15014 397920 -14958
rect 397976 -15014 398048 -14958
rect 397708 -15100 398048 -15014
rect 397708 -15156 397778 -15100
rect 397834 -15156 397920 -15100
rect 397976 -15156 398048 -15100
rect 397708 -15242 398048 -15156
rect 397708 -15298 397778 -15242
rect 397834 -15298 397920 -15242
rect 397976 -15298 398048 -15242
rect 397708 -15384 398048 -15298
rect 397708 -15440 397778 -15384
rect 397834 -15440 397920 -15384
rect 397976 -15440 398048 -15384
rect 397708 -15526 398048 -15440
rect 397708 -15582 397778 -15526
rect 397834 -15582 397920 -15526
rect 397976 -15582 398048 -15526
rect 397708 -15668 398048 -15582
rect 397708 -15724 397778 -15668
rect 397834 -15724 397920 -15668
rect 397976 -15724 398048 -15668
rect 397708 -15810 398048 -15724
rect 397708 -15866 397778 -15810
rect 397834 -15866 397920 -15810
rect 397976 -15866 398048 -15810
rect 397708 -15952 398048 -15866
rect 397708 -16008 397778 -15952
rect 397834 -16008 397920 -15952
rect 397976 -16008 398048 -15952
rect 397708 -16094 398048 -16008
rect 397708 -16150 397778 -16094
rect 397834 -16150 397920 -16094
rect 397976 -16150 398048 -16094
rect 397708 -16236 398048 -16150
rect 397708 -16292 397778 -16236
rect 397834 -16292 397920 -16236
rect 397976 -16292 398048 -16236
rect 397708 -16378 398048 -16292
rect 397708 -16434 397778 -16378
rect 397834 -16434 397920 -16378
rect 397976 -16434 398048 -16378
rect 397708 -16520 398048 -16434
rect 397708 -16576 397778 -16520
rect 397834 -16576 397920 -16520
rect 397976 -16576 398048 -16520
rect 397708 -16662 398048 -16576
rect 397708 -16718 397778 -16662
rect 397834 -16718 397920 -16662
rect 397976 -16718 398048 -16662
rect 397708 -16804 398048 -16718
rect 397708 -16860 397778 -16804
rect 397834 -16860 397920 -16804
rect 397976 -16860 398048 -16804
rect 397708 -16946 398048 -16860
rect 397708 -17002 397778 -16946
rect 397834 -17002 397920 -16946
rect 397976 -17002 398048 -16946
rect 397708 -17088 398048 -17002
rect 397708 -17144 397778 -17088
rect 397834 -17144 397920 -17088
rect 397976 -17144 398048 -17088
rect 397708 -17230 398048 -17144
rect 397708 -17286 397778 -17230
rect 397834 -17286 397920 -17230
rect 397976 -17286 398048 -17230
rect 397708 -17372 398048 -17286
rect 397708 -17428 397778 -17372
rect 397834 -17428 397920 -17372
rect 397976 -17428 398048 -17372
rect 397708 -17514 398048 -17428
rect 397708 -17570 397778 -17514
rect 397834 -17570 397920 -17514
rect 397976 -17570 398048 -17514
rect 397708 -17656 398048 -17570
rect 397708 -17712 397778 -17656
rect 397834 -17712 397920 -17656
rect 397976 -17712 398048 -17656
rect 397708 -17798 398048 -17712
rect 397708 -17854 397778 -17798
rect 397834 -17854 397920 -17798
rect 397976 -17854 398048 -17798
rect 397708 -17940 398048 -17854
rect 397708 -17996 397778 -17940
rect 397834 -17996 397920 -17940
rect 397976 -17996 398048 -17940
rect 397708 -18082 398048 -17996
rect 397708 -18138 397778 -18082
rect 397834 -18138 397920 -18082
rect 397976 -18138 398048 -18082
rect 397708 -18224 398048 -18138
rect 397708 -18280 397778 -18224
rect 397834 -18280 397920 -18224
rect 397976 -18280 398048 -18224
rect 397708 -18366 398048 -18280
rect 397708 -18422 397778 -18366
rect 397834 -18422 397920 -18366
rect 397976 -18422 398048 -18366
rect 397708 -18508 398048 -18422
rect 397708 -18564 397778 -18508
rect 397834 -18564 397920 -18508
rect 397976 -18564 398048 -18508
rect 397708 -18650 398048 -18564
rect 397708 -18706 397778 -18650
rect 397834 -18706 397920 -18650
rect 397976 -18706 398048 -18650
rect 397708 -18792 398048 -18706
rect 397708 -18848 397778 -18792
rect 397834 -18848 397920 -18792
rect 397976 -18848 398048 -18792
rect 397708 -18934 398048 -18848
rect 397708 -18990 397778 -18934
rect 397834 -18990 397920 -18934
rect 397976 -18990 398048 -18934
rect 397708 -19076 398048 -18990
rect 397708 -19132 397778 -19076
rect 397834 -19132 397920 -19076
rect 397976 -19132 398048 -19076
rect 397708 -19218 398048 -19132
rect 397708 -19274 397778 -19218
rect 397834 -19274 397920 -19218
rect 397976 -19274 398048 -19218
rect 397708 -19360 398048 -19274
rect 397708 -19416 397778 -19360
rect 397834 -19416 397920 -19360
rect 397976 -19416 398048 -19360
rect 397708 -19502 398048 -19416
rect 397708 -19558 397778 -19502
rect 397834 -19558 397920 -19502
rect 397976 -19558 398048 -19502
rect 397708 -19644 398048 -19558
rect 397708 -19700 397778 -19644
rect 397834 -19700 397920 -19644
rect 397976 -19700 398048 -19644
rect 397708 -19786 398048 -19700
rect 397708 -19842 397778 -19786
rect 397834 -19842 397920 -19786
rect 397976 -19842 398048 -19786
rect 397708 -19928 398048 -19842
rect 397708 -19984 397778 -19928
rect 397834 -19984 397920 -19928
rect 397976 -19984 398048 -19928
rect 397708 -20070 398048 -19984
rect 397708 -20126 397778 -20070
rect 397834 -20126 397920 -20070
rect 397976 -20126 398048 -20070
rect 397708 -20212 398048 -20126
rect 397708 -20268 397778 -20212
rect 397834 -20268 397920 -20212
rect 397976 -20268 398048 -20212
rect 397708 -20354 398048 -20268
rect 397708 -20410 397778 -20354
rect 397834 -20410 397920 -20354
rect 397976 -20410 398048 -20354
rect 397708 -20496 398048 -20410
rect 397708 -20552 397778 -20496
rect 397834 -20552 397920 -20496
rect 397976 -20552 398048 -20496
rect 397708 -20638 398048 -20552
rect 397708 -20694 397778 -20638
rect 397834 -20694 397920 -20638
rect 397976 -20694 398048 -20638
rect 397708 -20780 398048 -20694
rect 397708 -20836 397778 -20780
rect 397834 -20836 397920 -20780
rect 397976 -20836 398048 -20780
rect 397708 -20922 398048 -20836
rect 397708 -20978 397778 -20922
rect 397834 -20978 397920 -20922
rect 397976 -20978 398048 -20922
rect 397708 -21064 398048 -20978
rect 397708 -21120 397778 -21064
rect 397834 -21120 397920 -21064
rect 397976 -21120 398048 -21064
rect 397708 -21206 398048 -21120
rect 397708 -21262 397778 -21206
rect 397834 -21262 397920 -21206
rect 397976 -21262 398048 -21206
rect 397708 -21348 398048 -21262
rect 397708 -21404 397778 -21348
rect 397834 -21404 397920 -21348
rect 397976 -21404 398048 -21348
rect 397708 -21490 398048 -21404
rect 397708 -21546 397778 -21490
rect 397834 -21546 397920 -21490
rect 397976 -21546 398048 -21490
rect 397708 -21632 398048 -21546
rect 397708 -21688 397778 -21632
rect 397834 -21688 397920 -21632
rect 397976 -21688 398048 -21632
rect 397708 -21774 398048 -21688
rect 397708 -21830 397778 -21774
rect 397834 -21830 397920 -21774
rect 397976 -21830 398048 -21774
rect 397708 -21916 398048 -21830
rect 397708 -21972 397778 -21916
rect 397834 -21972 397920 -21916
rect 397976 -21972 398048 -21916
rect 397708 -22058 398048 -21972
rect 397708 -22114 397778 -22058
rect 397834 -22114 397920 -22058
rect 397976 -22114 398048 -22058
rect 397708 -22200 398048 -22114
rect 397708 -22256 397778 -22200
rect 397834 -22256 397920 -22200
rect 397976 -22256 398048 -22200
rect 397708 -22342 398048 -22256
rect 397708 -22398 397778 -22342
rect 397834 -22398 397920 -22342
rect 397976 -22398 398048 -22342
rect 397708 -22484 398048 -22398
rect 397708 -22540 397778 -22484
rect 397834 -22540 397920 -22484
rect 397976 -22540 398048 -22484
rect 397708 -22626 398048 -22540
rect 397708 -22682 397778 -22626
rect 397834 -22682 397920 -22626
rect 397976 -22682 398048 -22626
rect 397708 -22768 398048 -22682
rect 397708 -22824 397778 -22768
rect 397834 -22824 397920 -22768
rect 397976 -22824 398048 -22768
rect 397708 -22910 398048 -22824
rect 397708 -22966 397778 -22910
rect 397834 -22966 397920 -22910
rect 397976 -22966 398048 -22910
rect 397708 -23052 398048 -22966
rect 397708 -23108 397778 -23052
rect 397834 -23108 397920 -23052
rect 397976 -23108 398048 -23052
rect 397708 -23194 398048 -23108
rect 397708 -23250 397778 -23194
rect 397834 -23250 397920 -23194
rect 397976 -23250 398048 -23194
rect 397708 -23336 398048 -23250
rect 397708 -23392 397778 -23336
rect 397834 -23392 397920 -23336
rect 397976 -23392 398048 -23336
rect 397708 -23478 398048 -23392
rect 397708 -23534 397778 -23478
rect 397834 -23534 397920 -23478
rect 397976 -23534 398048 -23478
rect 397708 -23620 398048 -23534
rect 397708 -23676 397778 -23620
rect 397834 -23676 397920 -23620
rect 397976 -23676 398048 -23620
rect 397708 -23762 398048 -23676
rect 397708 -23818 397778 -23762
rect 397834 -23818 397920 -23762
rect 397976 -23818 398048 -23762
rect 397708 -23904 398048 -23818
rect 397708 -23960 397778 -23904
rect 397834 -23960 397920 -23904
rect 397976 -23960 398048 -23904
rect 397708 -24046 398048 -23960
rect 397708 -24102 397778 -24046
rect 397834 -24102 397920 -24046
rect 397976 -24102 398048 -24046
rect 397708 -24188 398048 -24102
rect 397708 -24244 397778 -24188
rect 397834 -24244 397920 -24188
rect 397976 -24244 398048 -24188
rect 397708 -24330 398048 -24244
rect 397708 -24386 397778 -24330
rect 397834 -24386 397920 -24330
rect 397976 -24386 398048 -24330
rect 397708 -24472 398048 -24386
rect 397708 -24528 397778 -24472
rect 397834 -24528 397920 -24472
rect 397976 -24528 398048 -24472
rect 397708 -24614 398048 -24528
rect 397708 -24670 397778 -24614
rect 397834 -24670 397920 -24614
rect 397976 -24670 398048 -24614
rect 397708 -24756 398048 -24670
rect 397708 -24812 397778 -24756
rect 397834 -24812 397920 -24756
rect 397976 -24812 398048 -24756
rect 397708 -24898 398048 -24812
rect 397708 -24954 397778 -24898
rect 397834 -24954 397920 -24898
rect 397976 -24954 398048 -24898
rect 397708 -25040 398048 -24954
rect 397708 -25096 397778 -25040
rect 397834 -25096 397920 -25040
rect 397976 -25096 398048 -25040
rect 397708 -25182 398048 -25096
rect 397708 -25238 397778 -25182
rect 397834 -25238 397920 -25182
rect 397976 -25238 398048 -25182
rect 397708 -25324 398048 -25238
rect 397708 -25380 397778 -25324
rect 397834 -25380 397920 -25324
rect 397976 -25380 398048 -25324
rect 397708 -25466 398048 -25380
rect 397708 -25522 397778 -25466
rect 397834 -25522 397920 -25466
rect 397976 -25522 398048 -25466
rect 397708 -25532 398048 -25522
rect 398108 -13680 398448 -13670
rect 398108 -13736 398174 -13680
rect 398230 -13736 398316 -13680
rect 398372 -13736 398448 -13680
rect 398108 -13822 398448 -13736
rect 398108 -13878 398174 -13822
rect 398230 -13878 398316 -13822
rect 398372 -13878 398448 -13822
rect 398108 -13964 398448 -13878
rect 398108 -14020 398174 -13964
rect 398230 -14020 398316 -13964
rect 398372 -14020 398448 -13964
rect 398108 -14106 398448 -14020
rect 398108 -14162 398174 -14106
rect 398230 -14162 398316 -14106
rect 398372 -14162 398448 -14106
rect 398108 -14248 398448 -14162
rect 398108 -14304 398174 -14248
rect 398230 -14304 398316 -14248
rect 398372 -14304 398448 -14248
rect 398108 -14390 398448 -14304
rect 398108 -14446 398174 -14390
rect 398230 -14446 398316 -14390
rect 398372 -14446 398448 -14390
rect 398108 -14532 398448 -14446
rect 398108 -14588 398174 -14532
rect 398230 -14588 398316 -14532
rect 398372 -14588 398448 -14532
rect 398108 -14674 398448 -14588
rect 398108 -14730 398174 -14674
rect 398230 -14730 398316 -14674
rect 398372 -14730 398448 -14674
rect 398108 -14816 398448 -14730
rect 398108 -14872 398174 -14816
rect 398230 -14872 398316 -14816
rect 398372 -14872 398448 -14816
rect 398108 -14958 398448 -14872
rect 398108 -15014 398174 -14958
rect 398230 -15014 398316 -14958
rect 398372 -15014 398448 -14958
rect 398108 -15100 398448 -15014
rect 398108 -15156 398174 -15100
rect 398230 -15156 398316 -15100
rect 398372 -15156 398448 -15100
rect 398108 -15242 398448 -15156
rect 398108 -15298 398174 -15242
rect 398230 -15298 398316 -15242
rect 398372 -15298 398448 -15242
rect 398108 -15384 398448 -15298
rect 398108 -15440 398174 -15384
rect 398230 -15440 398316 -15384
rect 398372 -15440 398448 -15384
rect 398108 -15526 398448 -15440
rect 398108 -15582 398174 -15526
rect 398230 -15582 398316 -15526
rect 398372 -15582 398448 -15526
rect 398108 -15668 398448 -15582
rect 398108 -15724 398174 -15668
rect 398230 -15724 398316 -15668
rect 398372 -15724 398448 -15668
rect 398108 -15810 398448 -15724
rect 398108 -15866 398174 -15810
rect 398230 -15866 398316 -15810
rect 398372 -15866 398448 -15810
rect 398108 -15952 398448 -15866
rect 398108 -16008 398174 -15952
rect 398230 -16008 398316 -15952
rect 398372 -16008 398448 -15952
rect 398108 -16094 398448 -16008
rect 398108 -16150 398174 -16094
rect 398230 -16150 398316 -16094
rect 398372 -16150 398448 -16094
rect 398108 -16236 398448 -16150
rect 398108 -16292 398174 -16236
rect 398230 -16292 398316 -16236
rect 398372 -16292 398448 -16236
rect 398108 -16378 398448 -16292
rect 398108 -16434 398174 -16378
rect 398230 -16434 398316 -16378
rect 398372 -16434 398448 -16378
rect 398108 -16520 398448 -16434
rect 398108 -16576 398174 -16520
rect 398230 -16576 398316 -16520
rect 398372 -16576 398448 -16520
rect 398108 -16662 398448 -16576
rect 398108 -16718 398174 -16662
rect 398230 -16718 398316 -16662
rect 398372 -16718 398448 -16662
rect 398108 -16804 398448 -16718
rect 398108 -16860 398174 -16804
rect 398230 -16860 398316 -16804
rect 398372 -16860 398448 -16804
rect 398108 -16946 398448 -16860
rect 398108 -17002 398174 -16946
rect 398230 -17002 398316 -16946
rect 398372 -17002 398448 -16946
rect 398108 -17088 398448 -17002
rect 398108 -17144 398174 -17088
rect 398230 -17144 398316 -17088
rect 398372 -17144 398448 -17088
rect 398108 -17230 398448 -17144
rect 398108 -17286 398174 -17230
rect 398230 -17286 398316 -17230
rect 398372 -17286 398448 -17230
rect 398108 -17372 398448 -17286
rect 398108 -17428 398174 -17372
rect 398230 -17428 398316 -17372
rect 398372 -17428 398448 -17372
rect 398108 -17514 398448 -17428
rect 398108 -17570 398174 -17514
rect 398230 -17570 398316 -17514
rect 398372 -17570 398448 -17514
rect 398108 -17656 398448 -17570
rect 398108 -17712 398174 -17656
rect 398230 -17712 398316 -17656
rect 398372 -17712 398448 -17656
rect 398108 -17798 398448 -17712
rect 398108 -17854 398174 -17798
rect 398230 -17854 398316 -17798
rect 398372 -17854 398448 -17798
rect 398108 -17940 398448 -17854
rect 398108 -17996 398174 -17940
rect 398230 -17996 398316 -17940
rect 398372 -17996 398448 -17940
rect 398108 -18082 398448 -17996
rect 398108 -18138 398174 -18082
rect 398230 -18138 398316 -18082
rect 398372 -18138 398448 -18082
rect 398108 -18224 398448 -18138
rect 398108 -18280 398174 -18224
rect 398230 -18280 398316 -18224
rect 398372 -18280 398448 -18224
rect 398108 -18366 398448 -18280
rect 398108 -18422 398174 -18366
rect 398230 -18422 398316 -18366
rect 398372 -18422 398448 -18366
rect 398108 -18508 398448 -18422
rect 398108 -18564 398174 -18508
rect 398230 -18564 398316 -18508
rect 398372 -18564 398448 -18508
rect 398108 -18650 398448 -18564
rect 398108 -18706 398174 -18650
rect 398230 -18706 398316 -18650
rect 398372 -18706 398448 -18650
rect 398108 -18792 398448 -18706
rect 398108 -18848 398174 -18792
rect 398230 -18848 398316 -18792
rect 398372 -18848 398448 -18792
rect 398108 -18934 398448 -18848
rect 398108 -18990 398174 -18934
rect 398230 -18990 398316 -18934
rect 398372 -18990 398448 -18934
rect 398108 -19076 398448 -18990
rect 398108 -19132 398174 -19076
rect 398230 -19132 398316 -19076
rect 398372 -19132 398448 -19076
rect 398108 -19218 398448 -19132
rect 398108 -19274 398174 -19218
rect 398230 -19274 398316 -19218
rect 398372 -19274 398448 -19218
rect 398108 -19360 398448 -19274
rect 398108 -19416 398174 -19360
rect 398230 -19416 398316 -19360
rect 398372 -19416 398448 -19360
rect 398108 -19502 398448 -19416
rect 398108 -19558 398174 -19502
rect 398230 -19558 398316 -19502
rect 398372 -19558 398448 -19502
rect 398108 -19644 398448 -19558
rect 398108 -19700 398174 -19644
rect 398230 -19700 398316 -19644
rect 398372 -19700 398448 -19644
rect 398108 -19786 398448 -19700
rect 398108 -19842 398174 -19786
rect 398230 -19842 398316 -19786
rect 398372 -19842 398448 -19786
rect 398108 -19928 398448 -19842
rect 398108 -19984 398174 -19928
rect 398230 -19984 398316 -19928
rect 398372 -19984 398448 -19928
rect 398108 -20070 398448 -19984
rect 398108 -20126 398174 -20070
rect 398230 -20126 398316 -20070
rect 398372 -20126 398448 -20070
rect 398108 -20212 398448 -20126
rect 398108 -20268 398174 -20212
rect 398230 -20268 398316 -20212
rect 398372 -20268 398448 -20212
rect 398108 -20354 398448 -20268
rect 398108 -20410 398174 -20354
rect 398230 -20410 398316 -20354
rect 398372 -20410 398448 -20354
rect 398108 -20496 398448 -20410
rect 398108 -20552 398174 -20496
rect 398230 -20552 398316 -20496
rect 398372 -20552 398448 -20496
rect 398108 -20638 398448 -20552
rect 398108 -20694 398174 -20638
rect 398230 -20694 398316 -20638
rect 398372 -20694 398448 -20638
rect 398108 -20780 398448 -20694
rect 398108 -20836 398174 -20780
rect 398230 -20836 398316 -20780
rect 398372 -20836 398448 -20780
rect 398108 -20922 398448 -20836
rect 398108 -20978 398174 -20922
rect 398230 -20978 398316 -20922
rect 398372 -20978 398448 -20922
rect 398108 -21064 398448 -20978
rect 398108 -21120 398174 -21064
rect 398230 -21120 398316 -21064
rect 398372 -21120 398448 -21064
rect 398108 -21206 398448 -21120
rect 398108 -21262 398174 -21206
rect 398230 -21262 398316 -21206
rect 398372 -21262 398448 -21206
rect 398108 -21348 398448 -21262
rect 398108 -21404 398174 -21348
rect 398230 -21404 398316 -21348
rect 398372 -21404 398448 -21348
rect 398108 -21490 398448 -21404
rect 398108 -21546 398174 -21490
rect 398230 -21546 398316 -21490
rect 398372 -21546 398448 -21490
rect 398108 -21632 398448 -21546
rect 398108 -21688 398174 -21632
rect 398230 -21688 398316 -21632
rect 398372 -21688 398448 -21632
rect 398108 -21774 398448 -21688
rect 398108 -21830 398174 -21774
rect 398230 -21830 398316 -21774
rect 398372 -21830 398448 -21774
rect 398108 -21916 398448 -21830
rect 398108 -21972 398174 -21916
rect 398230 -21972 398316 -21916
rect 398372 -21972 398448 -21916
rect 398108 -22058 398448 -21972
rect 398108 -22114 398174 -22058
rect 398230 -22114 398316 -22058
rect 398372 -22114 398448 -22058
rect 398108 -22200 398448 -22114
rect 398108 -22256 398174 -22200
rect 398230 -22256 398316 -22200
rect 398372 -22256 398448 -22200
rect 398108 -22342 398448 -22256
rect 398108 -22398 398174 -22342
rect 398230 -22398 398316 -22342
rect 398372 -22398 398448 -22342
rect 398108 -22484 398448 -22398
rect 398108 -22540 398174 -22484
rect 398230 -22540 398316 -22484
rect 398372 -22540 398448 -22484
rect 398108 -22626 398448 -22540
rect 398108 -22682 398174 -22626
rect 398230 -22682 398316 -22626
rect 398372 -22682 398448 -22626
rect 398108 -22768 398448 -22682
rect 398108 -22824 398174 -22768
rect 398230 -22824 398316 -22768
rect 398372 -22824 398448 -22768
rect 398108 -22910 398448 -22824
rect 398108 -22966 398174 -22910
rect 398230 -22966 398316 -22910
rect 398372 -22966 398448 -22910
rect 398108 -23052 398448 -22966
rect 398108 -23108 398174 -23052
rect 398230 -23108 398316 -23052
rect 398372 -23108 398448 -23052
rect 398108 -23194 398448 -23108
rect 398108 -23250 398174 -23194
rect 398230 -23250 398316 -23194
rect 398372 -23250 398448 -23194
rect 398108 -23336 398448 -23250
rect 398108 -23392 398174 -23336
rect 398230 -23392 398316 -23336
rect 398372 -23392 398448 -23336
rect 398108 -23478 398448 -23392
rect 398108 -23534 398174 -23478
rect 398230 -23534 398316 -23478
rect 398372 -23534 398448 -23478
rect 398108 -23620 398448 -23534
rect 398108 -23676 398174 -23620
rect 398230 -23676 398316 -23620
rect 398372 -23676 398448 -23620
rect 398108 -23762 398448 -23676
rect 398108 -23818 398174 -23762
rect 398230 -23818 398316 -23762
rect 398372 -23818 398448 -23762
rect 398108 -23904 398448 -23818
rect 398108 -23960 398174 -23904
rect 398230 -23960 398316 -23904
rect 398372 -23960 398448 -23904
rect 398108 -24046 398448 -23960
rect 398108 -24102 398174 -24046
rect 398230 -24102 398316 -24046
rect 398372 -24102 398448 -24046
rect 398108 -24188 398448 -24102
rect 398108 -24244 398174 -24188
rect 398230 -24244 398316 -24188
rect 398372 -24244 398448 -24188
rect 398108 -24330 398448 -24244
rect 398108 -24386 398174 -24330
rect 398230 -24386 398316 -24330
rect 398372 -24386 398448 -24330
rect 398108 -24472 398448 -24386
rect 398108 -24528 398174 -24472
rect 398230 -24528 398316 -24472
rect 398372 -24528 398448 -24472
rect 398108 -24614 398448 -24528
rect 398108 -24670 398174 -24614
rect 398230 -24670 398316 -24614
rect 398372 -24670 398448 -24614
rect 398108 -24756 398448 -24670
rect 398108 -24812 398174 -24756
rect 398230 -24812 398316 -24756
rect 398372 -24812 398448 -24756
rect 398108 -24898 398448 -24812
rect 398108 -24954 398174 -24898
rect 398230 -24954 398316 -24898
rect 398372 -24954 398448 -24898
rect 398108 -25040 398448 -24954
rect 398108 -25096 398174 -25040
rect 398230 -25096 398316 -25040
rect 398372 -25096 398448 -25040
rect 398108 -25182 398448 -25096
rect 398108 -25238 398174 -25182
rect 398230 -25238 398316 -25182
rect 398372 -25238 398448 -25182
rect 398108 -25324 398448 -25238
rect 398108 -25380 398174 -25324
rect 398230 -25380 398316 -25324
rect 398372 -25380 398448 -25324
rect 398108 -25466 398448 -25380
rect 398108 -25522 398174 -25466
rect 398230 -25522 398316 -25466
rect 398372 -25522 398448 -25466
rect 398108 -25532 398448 -25522
rect 398508 -13680 398848 -13670
rect 398508 -13736 398574 -13680
rect 398630 -13736 398716 -13680
rect 398772 -13736 398848 -13680
rect 398508 -13822 398848 -13736
rect 398508 -13878 398574 -13822
rect 398630 -13878 398716 -13822
rect 398772 -13878 398848 -13822
rect 398508 -13964 398848 -13878
rect 398508 -14020 398574 -13964
rect 398630 -14020 398716 -13964
rect 398772 -14020 398848 -13964
rect 398508 -14106 398848 -14020
rect 398508 -14162 398574 -14106
rect 398630 -14162 398716 -14106
rect 398772 -14162 398848 -14106
rect 398508 -14248 398848 -14162
rect 398508 -14304 398574 -14248
rect 398630 -14304 398716 -14248
rect 398772 -14304 398848 -14248
rect 398508 -14390 398848 -14304
rect 398508 -14446 398574 -14390
rect 398630 -14446 398716 -14390
rect 398772 -14446 398848 -14390
rect 398508 -14532 398848 -14446
rect 398508 -14588 398574 -14532
rect 398630 -14588 398716 -14532
rect 398772 -14588 398848 -14532
rect 398508 -14674 398848 -14588
rect 398508 -14730 398574 -14674
rect 398630 -14730 398716 -14674
rect 398772 -14730 398848 -14674
rect 398508 -14816 398848 -14730
rect 398508 -14872 398574 -14816
rect 398630 -14872 398716 -14816
rect 398772 -14872 398848 -14816
rect 398508 -14958 398848 -14872
rect 398508 -15014 398574 -14958
rect 398630 -15014 398716 -14958
rect 398772 -15014 398848 -14958
rect 398508 -15100 398848 -15014
rect 398508 -15156 398574 -15100
rect 398630 -15156 398716 -15100
rect 398772 -15156 398848 -15100
rect 398508 -15242 398848 -15156
rect 398508 -15298 398574 -15242
rect 398630 -15298 398716 -15242
rect 398772 -15298 398848 -15242
rect 398508 -15384 398848 -15298
rect 398508 -15440 398574 -15384
rect 398630 -15440 398716 -15384
rect 398772 -15440 398848 -15384
rect 398508 -15526 398848 -15440
rect 398508 -15582 398574 -15526
rect 398630 -15582 398716 -15526
rect 398772 -15582 398848 -15526
rect 398508 -15668 398848 -15582
rect 398508 -15724 398574 -15668
rect 398630 -15724 398716 -15668
rect 398772 -15724 398848 -15668
rect 398508 -15810 398848 -15724
rect 398508 -15866 398574 -15810
rect 398630 -15866 398716 -15810
rect 398772 -15866 398848 -15810
rect 398508 -15952 398848 -15866
rect 398508 -16008 398574 -15952
rect 398630 -16008 398716 -15952
rect 398772 -16008 398848 -15952
rect 398508 -16094 398848 -16008
rect 398508 -16150 398574 -16094
rect 398630 -16150 398716 -16094
rect 398772 -16150 398848 -16094
rect 398508 -16236 398848 -16150
rect 398508 -16292 398574 -16236
rect 398630 -16292 398716 -16236
rect 398772 -16292 398848 -16236
rect 398508 -16378 398848 -16292
rect 398508 -16434 398574 -16378
rect 398630 -16434 398716 -16378
rect 398772 -16434 398848 -16378
rect 398508 -16520 398848 -16434
rect 398508 -16576 398574 -16520
rect 398630 -16576 398716 -16520
rect 398772 -16576 398848 -16520
rect 398508 -16662 398848 -16576
rect 398508 -16718 398574 -16662
rect 398630 -16718 398716 -16662
rect 398772 -16718 398848 -16662
rect 398508 -16804 398848 -16718
rect 398508 -16860 398574 -16804
rect 398630 -16860 398716 -16804
rect 398772 -16860 398848 -16804
rect 398508 -16946 398848 -16860
rect 398508 -17002 398574 -16946
rect 398630 -17002 398716 -16946
rect 398772 -17002 398848 -16946
rect 398508 -17088 398848 -17002
rect 398508 -17144 398574 -17088
rect 398630 -17144 398716 -17088
rect 398772 -17144 398848 -17088
rect 398508 -17230 398848 -17144
rect 398508 -17286 398574 -17230
rect 398630 -17286 398716 -17230
rect 398772 -17286 398848 -17230
rect 398508 -17372 398848 -17286
rect 398508 -17428 398574 -17372
rect 398630 -17428 398716 -17372
rect 398772 -17428 398848 -17372
rect 398508 -17514 398848 -17428
rect 398508 -17570 398574 -17514
rect 398630 -17570 398716 -17514
rect 398772 -17570 398848 -17514
rect 398508 -17656 398848 -17570
rect 398508 -17712 398574 -17656
rect 398630 -17712 398716 -17656
rect 398772 -17712 398848 -17656
rect 398508 -17798 398848 -17712
rect 398508 -17854 398574 -17798
rect 398630 -17854 398716 -17798
rect 398772 -17854 398848 -17798
rect 398508 -17940 398848 -17854
rect 398508 -17996 398574 -17940
rect 398630 -17996 398716 -17940
rect 398772 -17996 398848 -17940
rect 398508 -18082 398848 -17996
rect 398508 -18138 398574 -18082
rect 398630 -18138 398716 -18082
rect 398772 -18138 398848 -18082
rect 398508 -18224 398848 -18138
rect 398508 -18280 398574 -18224
rect 398630 -18280 398716 -18224
rect 398772 -18280 398848 -18224
rect 398508 -18366 398848 -18280
rect 398508 -18422 398574 -18366
rect 398630 -18422 398716 -18366
rect 398772 -18422 398848 -18366
rect 398508 -18508 398848 -18422
rect 398508 -18564 398574 -18508
rect 398630 -18564 398716 -18508
rect 398772 -18564 398848 -18508
rect 398508 -18650 398848 -18564
rect 398508 -18706 398574 -18650
rect 398630 -18706 398716 -18650
rect 398772 -18706 398848 -18650
rect 398508 -18792 398848 -18706
rect 398508 -18848 398574 -18792
rect 398630 -18848 398716 -18792
rect 398772 -18848 398848 -18792
rect 398508 -18934 398848 -18848
rect 398508 -18990 398574 -18934
rect 398630 -18990 398716 -18934
rect 398772 -18990 398848 -18934
rect 398508 -19076 398848 -18990
rect 398508 -19132 398574 -19076
rect 398630 -19132 398716 -19076
rect 398772 -19132 398848 -19076
rect 398508 -19218 398848 -19132
rect 398508 -19274 398574 -19218
rect 398630 -19274 398716 -19218
rect 398772 -19274 398848 -19218
rect 398508 -19360 398848 -19274
rect 398508 -19416 398574 -19360
rect 398630 -19416 398716 -19360
rect 398772 -19416 398848 -19360
rect 398508 -19502 398848 -19416
rect 398508 -19558 398574 -19502
rect 398630 -19558 398716 -19502
rect 398772 -19558 398848 -19502
rect 398508 -19644 398848 -19558
rect 398508 -19700 398574 -19644
rect 398630 -19700 398716 -19644
rect 398772 -19700 398848 -19644
rect 398508 -19786 398848 -19700
rect 398508 -19842 398574 -19786
rect 398630 -19842 398716 -19786
rect 398772 -19842 398848 -19786
rect 398508 -19928 398848 -19842
rect 398508 -19984 398574 -19928
rect 398630 -19984 398716 -19928
rect 398772 -19984 398848 -19928
rect 398508 -20070 398848 -19984
rect 398508 -20126 398574 -20070
rect 398630 -20126 398716 -20070
rect 398772 -20126 398848 -20070
rect 398508 -20212 398848 -20126
rect 398508 -20268 398574 -20212
rect 398630 -20268 398716 -20212
rect 398772 -20268 398848 -20212
rect 398508 -20354 398848 -20268
rect 398508 -20410 398574 -20354
rect 398630 -20410 398716 -20354
rect 398772 -20410 398848 -20354
rect 398508 -20496 398848 -20410
rect 398508 -20552 398574 -20496
rect 398630 -20552 398716 -20496
rect 398772 -20552 398848 -20496
rect 398508 -20638 398848 -20552
rect 398508 -20694 398574 -20638
rect 398630 -20694 398716 -20638
rect 398772 -20694 398848 -20638
rect 398508 -20780 398848 -20694
rect 398508 -20836 398574 -20780
rect 398630 -20836 398716 -20780
rect 398772 -20836 398848 -20780
rect 398508 -20922 398848 -20836
rect 398508 -20978 398574 -20922
rect 398630 -20978 398716 -20922
rect 398772 -20978 398848 -20922
rect 398508 -21064 398848 -20978
rect 398508 -21120 398574 -21064
rect 398630 -21120 398716 -21064
rect 398772 -21120 398848 -21064
rect 398508 -21206 398848 -21120
rect 398508 -21262 398574 -21206
rect 398630 -21262 398716 -21206
rect 398772 -21262 398848 -21206
rect 398508 -21348 398848 -21262
rect 398508 -21404 398574 -21348
rect 398630 -21404 398716 -21348
rect 398772 -21404 398848 -21348
rect 398508 -21490 398848 -21404
rect 398508 -21546 398574 -21490
rect 398630 -21546 398716 -21490
rect 398772 -21546 398848 -21490
rect 398508 -21632 398848 -21546
rect 398508 -21688 398574 -21632
rect 398630 -21688 398716 -21632
rect 398772 -21688 398848 -21632
rect 398508 -21774 398848 -21688
rect 398508 -21830 398574 -21774
rect 398630 -21830 398716 -21774
rect 398772 -21830 398848 -21774
rect 398508 -21916 398848 -21830
rect 398508 -21972 398574 -21916
rect 398630 -21972 398716 -21916
rect 398772 -21972 398848 -21916
rect 398508 -22058 398848 -21972
rect 398508 -22114 398574 -22058
rect 398630 -22114 398716 -22058
rect 398772 -22114 398848 -22058
rect 398508 -22200 398848 -22114
rect 398508 -22256 398574 -22200
rect 398630 -22256 398716 -22200
rect 398772 -22256 398848 -22200
rect 398508 -22342 398848 -22256
rect 398508 -22398 398574 -22342
rect 398630 -22398 398716 -22342
rect 398772 -22398 398848 -22342
rect 398508 -22484 398848 -22398
rect 398508 -22540 398574 -22484
rect 398630 -22540 398716 -22484
rect 398772 -22540 398848 -22484
rect 398508 -22626 398848 -22540
rect 398508 -22682 398574 -22626
rect 398630 -22682 398716 -22626
rect 398772 -22682 398848 -22626
rect 398508 -22768 398848 -22682
rect 398508 -22824 398574 -22768
rect 398630 -22824 398716 -22768
rect 398772 -22824 398848 -22768
rect 398508 -22910 398848 -22824
rect 398508 -22966 398574 -22910
rect 398630 -22966 398716 -22910
rect 398772 -22966 398848 -22910
rect 398508 -23052 398848 -22966
rect 398508 -23108 398574 -23052
rect 398630 -23108 398716 -23052
rect 398772 -23108 398848 -23052
rect 398508 -23194 398848 -23108
rect 398508 -23250 398574 -23194
rect 398630 -23250 398716 -23194
rect 398772 -23250 398848 -23194
rect 398508 -23336 398848 -23250
rect 398508 -23392 398574 -23336
rect 398630 -23392 398716 -23336
rect 398772 -23392 398848 -23336
rect 398508 -23478 398848 -23392
rect 398508 -23534 398574 -23478
rect 398630 -23534 398716 -23478
rect 398772 -23534 398848 -23478
rect 398508 -23620 398848 -23534
rect 398508 -23676 398574 -23620
rect 398630 -23676 398716 -23620
rect 398772 -23676 398848 -23620
rect 398508 -23762 398848 -23676
rect 398508 -23818 398574 -23762
rect 398630 -23818 398716 -23762
rect 398772 -23818 398848 -23762
rect 398508 -23904 398848 -23818
rect 398508 -23960 398574 -23904
rect 398630 -23960 398716 -23904
rect 398772 -23960 398848 -23904
rect 398508 -24046 398848 -23960
rect 398508 -24102 398574 -24046
rect 398630 -24102 398716 -24046
rect 398772 -24102 398848 -24046
rect 398508 -24188 398848 -24102
rect 398508 -24244 398574 -24188
rect 398630 -24244 398716 -24188
rect 398772 -24244 398848 -24188
rect 398508 -24330 398848 -24244
rect 398508 -24386 398574 -24330
rect 398630 -24386 398716 -24330
rect 398772 -24386 398848 -24330
rect 398508 -24472 398848 -24386
rect 398508 -24528 398574 -24472
rect 398630 -24528 398716 -24472
rect 398772 -24528 398848 -24472
rect 398508 -24614 398848 -24528
rect 398508 -24670 398574 -24614
rect 398630 -24670 398716 -24614
rect 398772 -24670 398848 -24614
rect 398508 -24756 398848 -24670
rect 398508 -24812 398574 -24756
rect 398630 -24812 398716 -24756
rect 398772 -24812 398848 -24756
rect 398508 -24898 398848 -24812
rect 398508 -24954 398574 -24898
rect 398630 -24954 398716 -24898
rect 398772 -24954 398848 -24898
rect 398508 -25040 398848 -24954
rect 398508 -25096 398574 -25040
rect 398630 -25096 398716 -25040
rect 398772 -25096 398848 -25040
rect 398508 -25182 398848 -25096
rect 398508 -25238 398574 -25182
rect 398630 -25238 398716 -25182
rect 398772 -25238 398848 -25182
rect 398508 -25324 398848 -25238
rect 398508 -25380 398574 -25324
rect 398630 -25380 398716 -25324
rect 398772 -25380 398848 -25324
rect 398508 -25466 398848 -25380
rect 398508 -25522 398574 -25466
rect 398630 -25522 398716 -25466
rect 398772 -25522 398848 -25466
rect 398508 -25532 398848 -25522
rect 398908 -13680 399248 -13670
rect 398908 -13736 398971 -13680
rect 399027 -13736 399113 -13680
rect 399169 -13736 399248 -13680
rect 398908 -13822 399248 -13736
rect 398908 -13878 398971 -13822
rect 399027 -13878 399113 -13822
rect 399169 -13878 399248 -13822
rect 398908 -13964 399248 -13878
rect 398908 -14020 398971 -13964
rect 399027 -14020 399113 -13964
rect 399169 -14020 399248 -13964
rect 398908 -14106 399248 -14020
rect 398908 -14162 398971 -14106
rect 399027 -14162 399113 -14106
rect 399169 -14162 399248 -14106
rect 398908 -14248 399248 -14162
rect 398908 -14304 398971 -14248
rect 399027 -14304 399113 -14248
rect 399169 -14304 399248 -14248
rect 398908 -14390 399248 -14304
rect 398908 -14446 398971 -14390
rect 399027 -14446 399113 -14390
rect 399169 -14446 399248 -14390
rect 398908 -14532 399248 -14446
rect 398908 -14588 398971 -14532
rect 399027 -14588 399113 -14532
rect 399169 -14588 399248 -14532
rect 398908 -14674 399248 -14588
rect 398908 -14730 398971 -14674
rect 399027 -14730 399113 -14674
rect 399169 -14730 399248 -14674
rect 398908 -14816 399248 -14730
rect 398908 -14872 398971 -14816
rect 399027 -14872 399113 -14816
rect 399169 -14872 399248 -14816
rect 398908 -14958 399248 -14872
rect 398908 -15014 398971 -14958
rect 399027 -15014 399113 -14958
rect 399169 -15014 399248 -14958
rect 398908 -15100 399248 -15014
rect 398908 -15156 398971 -15100
rect 399027 -15156 399113 -15100
rect 399169 -15156 399248 -15100
rect 398908 -15242 399248 -15156
rect 398908 -15298 398971 -15242
rect 399027 -15298 399113 -15242
rect 399169 -15298 399248 -15242
rect 398908 -15384 399248 -15298
rect 398908 -15440 398971 -15384
rect 399027 -15440 399113 -15384
rect 399169 -15440 399248 -15384
rect 398908 -15526 399248 -15440
rect 398908 -15582 398971 -15526
rect 399027 -15582 399113 -15526
rect 399169 -15582 399248 -15526
rect 398908 -15668 399248 -15582
rect 398908 -15724 398971 -15668
rect 399027 -15724 399113 -15668
rect 399169 -15724 399248 -15668
rect 398908 -15810 399248 -15724
rect 398908 -15866 398971 -15810
rect 399027 -15866 399113 -15810
rect 399169 -15866 399248 -15810
rect 398908 -15952 399248 -15866
rect 398908 -16008 398971 -15952
rect 399027 -16008 399113 -15952
rect 399169 -16008 399248 -15952
rect 398908 -16094 399248 -16008
rect 398908 -16150 398971 -16094
rect 399027 -16150 399113 -16094
rect 399169 -16150 399248 -16094
rect 398908 -16236 399248 -16150
rect 398908 -16292 398971 -16236
rect 399027 -16292 399113 -16236
rect 399169 -16292 399248 -16236
rect 398908 -16378 399248 -16292
rect 398908 -16434 398971 -16378
rect 399027 -16434 399113 -16378
rect 399169 -16434 399248 -16378
rect 398908 -16520 399248 -16434
rect 398908 -16576 398971 -16520
rect 399027 -16576 399113 -16520
rect 399169 -16576 399248 -16520
rect 398908 -16662 399248 -16576
rect 398908 -16718 398971 -16662
rect 399027 -16718 399113 -16662
rect 399169 -16718 399248 -16662
rect 398908 -16804 399248 -16718
rect 398908 -16860 398971 -16804
rect 399027 -16860 399113 -16804
rect 399169 -16860 399248 -16804
rect 398908 -16946 399248 -16860
rect 398908 -17002 398971 -16946
rect 399027 -17002 399113 -16946
rect 399169 -17002 399248 -16946
rect 398908 -17088 399248 -17002
rect 398908 -17144 398971 -17088
rect 399027 -17144 399113 -17088
rect 399169 -17144 399248 -17088
rect 398908 -17230 399248 -17144
rect 398908 -17286 398971 -17230
rect 399027 -17286 399113 -17230
rect 399169 -17286 399248 -17230
rect 398908 -17372 399248 -17286
rect 398908 -17428 398971 -17372
rect 399027 -17428 399113 -17372
rect 399169 -17428 399248 -17372
rect 398908 -17514 399248 -17428
rect 398908 -17570 398971 -17514
rect 399027 -17570 399113 -17514
rect 399169 -17570 399248 -17514
rect 398908 -17656 399248 -17570
rect 398908 -17712 398971 -17656
rect 399027 -17712 399113 -17656
rect 399169 -17712 399248 -17656
rect 398908 -17798 399248 -17712
rect 398908 -17854 398971 -17798
rect 399027 -17854 399113 -17798
rect 399169 -17854 399248 -17798
rect 398908 -17940 399248 -17854
rect 398908 -17996 398971 -17940
rect 399027 -17996 399113 -17940
rect 399169 -17996 399248 -17940
rect 398908 -18082 399248 -17996
rect 398908 -18138 398971 -18082
rect 399027 -18138 399113 -18082
rect 399169 -18138 399248 -18082
rect 398908 -18224 399248 -18138
rect 398908 -18280 398971 -18224
rect 399027 -18280 399113 -18224
rect 399169 -18280 399248 -18224
rect 398908 -18366 399248 -18280
rect 398908 -18422 398971 -18366
rect 399027 -18422 399113 -18366
rect 399169 -18422 399248 -18366
rect 398908 -18508 399248 -18422
rect 398908 -18564 398971 -18508
rect 399027 -18564 399113 -18508
rect 399169 -18564 399248 -18508
rect 398908 -18650 399248 -18564
rect 398908 -18706 398971 -18650
rect 399027 -18706 399113 -18650
rect 399169 -18706 399248 -18650
rect 398908 -18792 399248 -18706
rect 398908 -18848 398971 -18792
rect 399027 -18848 399113 -18792
rect 399169 -18848 399248 -18792
rect 398908 -18934 399248 -18848
rect 398908 -18990 398971 -18934
rect 399027 -18990 399113 -18934
rect 399169 -18990 399248 -18934
rect 398908 -19076 399248 -18990
rect 398908 -19132 398971 -19076
rect 399027 -19132 399113 -19076
rect 399169 -19132 399248 -19076
rect 398908 -19218 399248 -19132
rect 398908 -19274 398971 -19218
rect 399027 -19274 399113 -19218
rect 399169 -19274 399248 -19218
rect 398908 -19360 399248 -19274
rect 398908 -19416 398971 -19360
rect 399027 -19416 399113 -19360
rect 399169 -19416 399248 -19360
rect 398908 -19502 399248 -19416
rect 398908 -19558 398971 -19502
rect 399027 -19558 399113 -19502
rect 399169 -19558 399248 -19502
rect 398908 -19644 399248 -19558
rect 398908 -19700 398971 -19644
rect 399027 -19700 399113 -19644
rect 399169 -19700 399248 -19644
rect 398908 -19786 399248 -19700
rect 398908 -19842 398971 -19786
rect 399027 -19842 399113 -19786
rect 399169 -19842 399248 -19786
rect 398908 -19928 399248 -19842
rect 398908 -19984 398971 -19928
rect 399027 -19984 399113 -19928
rect 399169 -19984 399248 -19928
rect 398908 -20070 399248 -19984
rect 398908 -20126 398971 -20070
rect 399027 -20126 399113 -20070
rect 399169 -20126 399248 -20070
rect 398908 -20212 399248 -20126
rect 398908 -20268 398971 -20212
rect 399027 -20268 399113 -20212
rect 399169 -20268 399248 -20212
rect 398908 -20354 399248 -20268
rect 398908 -20410 398971 -20354
rect 399027 -20410 399113 -20354
rect 399169 -20410 399248 -20354
rect 398908 -20496 399248 -20410
rect 398908 -20552 398971 -20496
rect 399027 -20552 399113 -20496
rect 399169 -20552 399248 -20496
rect 398908 -20638 399248 -20552
rect 398908 -20694 398971 -20638
rect 399027 -20694 399113 -20638
rect 399169 -20694 399248 -20638
rect 398908 -20780 399248 -20694
rect 398908 -20836 398971 -20780
rect 399027 -20836 399113 -20780
rect 399169 -20836 399248 -20780
rect 398908 -20922 399248 -20836
rect 398908 -20978 398971 -20922
rect 399027 -20978 399113 -20922
rect 399169 -20978 399248 -20922
rect 398908 -21064 399248 -20978
rect 398908 -21120 398971 -21064
rect 399027 -21120 399113 -21064
rect 399169 -21120 399248 -21064
rect 398908 -21206 399248 -21120
rect 398908 -21262 398971 -21206
rect 399027 -21262 399113 -21206
rect 399169 -21262 399248 -21206
rect 398908 -21348 399248 -21262
rect 398908 -21404 398971 -21348
rect 399027 -21404 399113 -21348
rect 399169 -21404 399248 -21348
rect 398908 -21490 399248 -21404
rect 398908 -21546 398971 -21490
rect 399027 -21546 399113 -21490
rect 399169 -21546 399248 -21490
rect 398908 -21632 399248 -21546
rect 398908 -21688 398971 -21632
rect 399027 -21688 399113 -21632
rect 399169 -21688 399248 -21632
rect 398908 -21774 399248 -21688
rect 398908 -21830 398971 -21774
rect 399027 -21830 399113 -21774
rect 399169 -21830 399248 -21774
rect 398908 -21916 399248 -21830
rect 398908 -21972 398971 -21916
rect 399027 -21972 399113 -21916
rect 399169 -21972 399248 -21916
rect 398908 -22058 399248 -21972
rect 398908 -22114 398971 -22058
rect 399027 -22114 399113 -22058
rect 399169 -22114 399248 -22058
rect 398908 -22200 399248 -22114
rect 398908 -22256 398971 -22200
rect 399027 -22256 399113 -22200
rect 399169 -22256 399248 -22200
rect 398908 -22342 399248 -22256
rect 398908 -22398 398971 -22342
rect 399027 -22398 399113 -22342
rect 399169 -22398 399248 -22342
rect 398908 -22484 399248 -22398
rect 398908 -22540 398971 -22484
rect 399027 -22540 399113 -22484
rect 399169 -22540 399248 -22484
rect 398908 -22626 399248 -22540
rect 398908 -22682 398971 -22626
rect 399027 -22682 399113 -22626
rect 399169 -22682 399248 -22626
rect 398908 -22768 399248 -22682
rect 398908 -22824 398971 -22768
rect 399027 -22824 399113 -22768
rect 399169 -22824 399248 -22768
rect 398908 -22910 399248 -22824
rect 398908 -22966 398971 -22910
rect 399027 -22966 399113 -22910
rect 399169 -22966 399248 -22910
rect 398908 -23052 399248 -22966
rect 398908 -23108 398971 -23052
rect 399027 -23108 399113 -23052
rect 399169 -23108 399248 -23052
rect 398908 -23194 399248 -23108
rect 398908 -23250 398971 -23194
rect 399027 -23250 399113 -23194
rect 399169 -23250 399248 -23194
rect 398908 -23336 399248 -23250
rect 398908 -23392 398971 -23336
rect 399027 -23392 399113 -23336
rect 399169 -23392 399248 -23336
rect 398908 -23478 399248 -23392
rect 398908 -23534 398971 -23478
rect 399027 -23534 399113 -23478
rect 399169 -23534 399248 -23478
rect 398908 -23620 399248 -23534
rect 398908 -23676 398971 -23620
rect 399027 -23676 399113 -23620
rect 399169 -23676 399248 -23620
rect 398908 -23762 399248 -23676
rect 398908 -23818 398971 -23762
rect 399027 -23818 399113 -23762
rect 399169 -23818 399248 -23762
rect 398908 -23904 399248 -23818
rect 398908 -23960 398971 -23904
rect 399027 -23960 399113 -23904
rect 399169 -23960 399248 -23904
rect 398908 -24046 399248 -23960
rect 398908 -24102 398971 -24046
rect 399027 -24102 399113 -24046
rect 399169 -24102 399248 -24046
rect 398908 -24188 399248 -24102
rect 398908 -24244 398971 -24188
rect 399027 -24244 399113 -24188
rect 399169 -24244 399248 -24188
rect 398908 -24330 399248 -24244
rect 398908 -24386 398971 -24330
rect 399027 -24386 399113 -24330
rect 399169 -24386 399248 -24330
rect 398908 -24472 399248 -24386
rect 398908 -24528 398971 -24472
rect 399027 -24528 399113 -24472
rect 399169 -24528 399248 -24472
rect 398908 -24614 399248 -24528
rect 398908 -24670 398971 -24614
rect 399027 -24670 399113 -24614
rect 399169 -24670 399248 -24614
rect 398908 -24756 399248 -24670
rect 398908 -24812 398971 -24756
rect 399027 -24812 399113 -24756
rect 399169 -24812 399248 -24756
rect 398908 -24898 399248 -24812
rect 398908 -24954 398971 -24898
rect 399027 -24954 399113 -24898
rect 399169 -24954 399248 -24898
rect 398908 -25040 399248 -24954
rect 398908 -25096 398971 -25040
rect 399027 -25096 399113 -25040
rect 399169 -25096 399248 -25040
rect 398908 -25182 399248 -25096
rect 398908 -25238 398971 -25182
rect 399027 -25238 399113 -25182
rect 399169 -25238 399248 -25182
rect 398908 -25324 399248 -25238
rect 398908 -25380 398971 -25324
rect 399027 -25380 399113 -25324
rect 399169 -25380 399248 -25324
rect 398908 -25466 399248 -25380
rect 398908 -25522 398971 -25466
rect 399027 -25522 399113 -25466
rect 399169 -25522 399248 -25466
rect 398908 -25532 399248 -25522
rect 399308 -13680 399648 -13670
rect 399308 -13736 399376 -13680
rect 399432 -13736 399518 -13680
rect 399574 -13736 399648 -13680
rect 399308 -13822 399648 -13736
rect 399308 -13878 399376 -13822
rect 399432 -13878 399518 -13822
rect 399574 -13878 399648 -13822
rect 399308 -13964 399648 -13878
rect 399308 -14020 399376 -13964
rect 399432 -14020 399518 -13964
rect 399574 -14020 399648 -13964
rect 399308 -14106 399648 -14020
rect 399308 -14162 399376 -14106
rect 399432 -14162 399518 -14106
rect 399574 -14162 399648 -14106
rect 399308 -14248 399648 -14162
rect 399308 -14304 399376 -14248
rect 399432 -14304 399518 -14248
rect 399574 -14304 399648 -14248
rect 399308 -14390 399648 -14304
rect 399308 -14446 399376 -14390
rect 399432 -14446 399518 -14390
rect 399574 -14446 399648 -14390
rect 399308 -14532 399648 -14446
rect 399308 -14588 399376 -14532
rect 399432 -14588 399518 -14532
rect 399574 -14588 399648 -14532
rect 399308 -14674 399648 -14588
rect 399308 -14730 399376 -14674
rect 399432 -14730 399518 -14674
rect 399574 -14730 399648 -14674
rect 399308 -14816 399648 -14730
rect 399308 -14872 399376 -14816
rect 399432 -14872 399518 -14816
rect 399574 -14872 399648 -14816
rect 399308 -14958 399648 -14872
rect 399308 -15014 399376 -14958
rect 399432 -15014 399518 -14958
rect 399574 -15014 399648 -14958
rect 399308 -15100 399648 -15014
rect 399308 -15156 399376 -15100
rect 399432 -15156 399518 -15100
rect 399574 -15156 399648 -15100
rect 399308 -15242 399648 -15156
rect 399308 -15298 399376 -15242
rect 399432 -15298 399518 -15242
rect 399574 -15298 399648 -15242
rect 399308 -15384 399648 -15298
rect 399308 -15440 399376 -15384
rect 399432 -15440 399518 -15384
rect 399574 -15440 399648 -15384
rect 399308 -15526 399648 -15440
rect 399308 -15582 399376 -15526
rect 399432 -15582 399518 -15526
rect 399574 -15582 399648 -15526
rect 399308 -15668 399648 -15582
rect 399308 -15724 399376 -15668
rect 399432 -15724 399518 -15668
rect 399574 -15724 399648 -15668
rect 399308 -15810 399648 -15724
rect 399308 -15866 399376 -15810
rect 399432 -15866 399518 -15810
rect 399574 -15866 399648 -15810
rect 399308 -15952 399648 -15866
rect 399308 -16008 399376 -15952
rect 399432 -16008 399518 -15952
rect 399574 -16008 399648 -15952
rect 399308 -16094 399648 -16008
rect 399308 -16150 399376 -16094
rect 399432 -16150 399518 -16094
rect 399574 -16150 399648 -16094
rect 399308 -16236 399648 -16150
rect 399308 -16292 399376 -16236
rect 399432 -16292 399518 -16236
rect 399574 -16292 399648 -16236
rect 399308 -16378 399648 -16292
rect 399308 -16434 399376 -16378
rect 399432 -16434 399518 -16378
rect 399574 -16434 399648 -16378
rect 399308 -16520 399648 -16434
rect 399308 -16576 399376 -16520
rect 399432 -16576 399518 -16520
rect 399574 -16576 399648 -16520
rect 399308 -16662 399648 -16576
rect 399308 -16718 399376 -16662
rect 399432 -16718 399518 -16662
rect 399574 -16718 399648 -16662
rect 399308 -16804 399648 -16718
rect 399308 -16860 399376 -16804
rect 399432 -16860 399518 -16804
rect 399574 -16860 399648 -16804
rect 399308 -16946 399648 -16860
rect 399308 -17002 399376 -16946
rect 399432 -17002 399518 -16946
rect 399574 -17002 399648 -16946
rect 399308 -17088 399648 -17002
rect 399308 -17144 399376 -17088
rect 399432 -17144 399518 -17088
rect 399574 -17144 399648 -17088
rect 399308 -17230 399648 -17144
rect 399308 -17286 399376 -17230
rect 399432 -17286 399518 -17230
rect 399574 -17286 399648 -17230
rect 399308 -17372 399648 -17286
rect 399308 -17428 399376 -17372
rect 399432 -17428 399518 -17372
rect 399574 -17428 399648 -17372
rect 399308 -17514 399648 -17428
rect 399308 -17570 399376 -17514
rect 399432 -17570 399518 -17514
rect 399574 -17570 399648 -17514
rect 399308 -17656 399648 -17570
rect 399308 -17712 399376 -17656
rect 399432 -17712 399518 -17656
rect 399574 -17712 399648 -17656
rect 399308 -17798 399648 -17712
rect 399308 -17854 399376 -17798
rect 399432 -17854 399518 -17798
rect 399574 -17854 399648 -17798
rect 399308 -17940 399648 -17854
rect 399308 -17996 399376 -17940
rect 399432 -17996 399518 -17940
rect 399574 -17996 399648 -17940
rect 399308 -18082 399648 -17996
rect 399308 -18138 399376 -18082
rect 399432 -18138 399518 -18082
rect 399574 -18138 399648 -18082
rect 399308 -18224 399648 -18138
rect 399308 -18280 399376 -18224
rect 399432 -18280 399518 -18224
rect 399574 -18280 399648 -18224
rect 399308 -18366 399648 -18280
rect 399308 -18422 399376 -18366
rect 399432 -18422 399518 -18366
rect 399574 -18422 399648 -18366
rect 399308 -18508 399648 -18422
rect 399308 -18564 399376 -18508
rect 399432 -18564 399518 -18508
rect 399574 -18564 399648 -18508
rect 399308 -18650 399648 -18564
rect 399308 -18706 399376 -18650
rect 399432 -18706 399518 -18650
rect 399574 -18706 399648 -18650
rect 399308 -18792 399648 -18706
rect 399308 -18848 399376 -18792
rect 399432 -18848 399518 -18792
rect 399574 -18848 399648 -18792
rect 399308 -18934 399648 -18848
rect 399308 -18990 399376 -18934
rect 399432 -18990 399518 -18934
rect 399574 -18990 399648 -18934
rect 399308 -19076 399648 -18990
rect 399308 -19132 399376 -19076
rect 399432 -19132 399518 -19076
rect 399574 -19132 399648 -19076
rect 399308 -19218 399648 -19132
rect 399308 -19274 399376 -19218
rect 399432 -19274 399518 -19218
rect 399574 -19274 399648 -19218
rect 399308 -19360 399648 -19274
rect 399308 -19416 399376 -19360
rect 399432 -19416 399518 -19360
rect 399574 -19416 399648 -19360
rect 399308 -19502 399648 -19416
rect 399308 -19558 399376 -19502
rect 399432 -19558 399518 -19502
rect 399574 -19558 399648 -19502
rect 399308 -19644 399648 -19558
rect 399308 -19700 399376 -19644
rect 399432 -19700 399518 -19644
rect 399574 -19700 399648 -19644
rect 399308 -19786 399648 -19700
rect 399308 -19842 399376 -19786
rect 399432 -19842 399518 -19786
rect 399574 -19842 399648 -19786
rect 399308 -19928 399648 -19842
rect 399308 -19984 399376 -19928
rect 399432 -19984 399518 -19928
rect 399574 -19984 399648 -19928
rect 399308 -20070 399648 -19984
rect 399308 -20126 399376 -20070
rect 399432 -20126 399518 -20070
rect 399574 -20126 399648 -20070
rect 399308 -20212 399648 -20126
rect 399308 -20268 399376 -20212
rect 399432 -20268 399518 -20212
rect 399574 -20268 399648 -20212
rect 399308 -20354 399648 -20268
rect 399308 -20410 399376 -20354
rect 399432 -20410 399518 -20354
rect 399574 -20410 399648 -20354
rect 399308 -20496 399648 -20410
rect 399308 -20552 399376 -20496
rect 399432 -20552 399518 -20496
rect 399574 -20552 399648 -20496
rect 399308 -20638 399648 -20552
rect 399308 -20694 399376 -20638
rect 399432 -20694 399518 -20638
rect 399574 -20694 399648 -20638
rect 399308 -20780 399648 -20694
rect 399308 -20836 399376 -20780
rect 399432 -20836 399518 -20780
rect 399574 -20836 399648 -20780
rect 399308 -20922 399648 -20836
rect 399308 -20978 399376 -20922
rect 399432 -20978 399518 -20922
rect 399574 -20978 399648 -20922
rect 399308 -21064 399648 -20978
rect 399308 -21120 399376 -21064
rect 399432 -21120 399518 -21064
rect 399574 -21120 399648 -21064
rect 399308 -21206 399648 -21120
rect 399308 -21262 399376 -21206
rect 399432 -21262 399518 -21206
rect 399574 -21262 399648 -21206
rect 399308 -21348 399648 -21262
rect 399308 -21404 399376 -21348
rect 399432 -21404 399518 -21348
rect 399574 -21404 399648 -21348
rect 399308 -21490 399648 -21404
rect 399308 -21546 399376 -21490
rect 399432 -21546 399518 -21490
rect 399574 -21546 399648 -21490
rect 399308 -21632 399648 -21546
rect 399308 -21688 399376 -21632
rect 399432 -21688 399518 -21632
rect 399574 -21688 399648 -21632
rect 399308 -21774 399648 -21688
rect 399308 -21830 399376 -21774
rect 399432 -21830 399518 -21774
rect 399574 -21830 399648 -21774
rect 399308 -21916 399648 -21830
rect 399308 -21972 399376 -21916
rect 399432 -21972 399518 -21916
rect 399574 -21972 399648 -21916
rect 399308 -22058 399648 -21972
rect 399308 -22114 399376 -22058
rect 399432 -22114 399518 -22058
rect 399574 -22114 399648 -22058
rect 399308 -22200 399648 -22114
rect 399308 -22256 399376 -22200
rect 399432 -22256 399518 -22200
rect 399574 -22256 399648 -22200
rect 399308 -22342 399648 -22256
rect 399308 -22398 399376 -22342
rect 399432 -22398 399518 -22342
rect 399574 -22398 399648 -22342
rect 399308 -22484 399648 -22398
rect 399308 -22540 399376 -22484
rect 399432 -22540 399518 -22484
rect 399574 -22540 399648 -22484
rect 399308 -22626 399648 -22540
rect 399308 -22682 399376 -22626
rect 399432 -22682 399518 -22626
rect 399574 -22682 399648 -22626
rect 399308 -22768 399648 -22682
rect 399308 -22824 399376 -22768
rect 399432 -22824 399518 -22768
rect 399574 -22824 399648 -22768
rect 399308 -22910 399648 -22824
rect 399308 -22966 399376 -22910
rect 399432 -22966 399518 -22910
rect 399574 -22966 399648 -22910
rect 399308 -23052 399648 -22966
rect 399308 -23108 399376 -23052
rect 399432 -23108 399518 -23052
rect 399574 -23108 399648 -23052
rect 399308 -23194 399648 -23108
rect 399308 -23250 399376 -23194
rect 399432 -23250 399518 -23194
rect 399574 -23250 399648 -23194
rect 399308 -23336 399648 -23250
rect 399308 -23392 399376 -23336
rect 399432 -23392 399518 -23336
rect 399574 -23392 399648 -23336
rect 399308 -23478 399648 -23392
rect 399308 -23534 399376 -23478
rect 399432 -23534 399518 -23478
rect 399574 -23534 399648 -23478
rect 399308 -23620 399648 -23534
rect 399308 -23676 399376 -23620
rect 399432 -23676 399518 -23620
rect 399574 -23676 399648 -23620
rect 399308 -23762 399648 -23676
rect 399308 -23818 399376 -23762
rect 399432 -23818 399518 -23762
rect 399574 -23818 399648 -23762
rect 399308 -23904 399648 -23818
rect 399308 -23960 399376 -23904
rect 399432 -23960 399518 -23904
rect 399574 -23960 399648 -23904
rect 399308 -24046 399648 -23960
rect 399308 -24102 399376 -24046
rect 399432 -24102 399518 -24046
rect 399574 -24102 399648 -24046
rect 399308 -24188 399648 -24102
rect 399308 -24244 399376 -24188
rect 399432 -24244 399518 -24188
rect 399574 -24244 399648 -24188
rect 399308 -24330 399648 -24244
rect 399308 -24386 399376 -24330
rect 399432 -24386 399518 -24330
rect 399574 -24386 399648 -24330
rect 399308 -24472 399648 -24386
rect 399308 -24528 399376 -24472
rect 399432 -24528 399518 -24472
rect 399574 -24528 399648 -24472
rect 399308 -24614 399648 -24528
rect 399308 -24670 399376 -24614
rect 399432 -24670 399518 -24614
rect 399574 -24670 399648 -24614
rect 399308 -24756 399648 -24670
rect 399308 -24812 399376 -24756
rect 399432 -24812 399518 -24756
rect 399574 -24812 399648 -24756
rect 399308 -24898 399648 -24812
rect 399308 -24954 399376 -24898
rect 399432 -24954 399518 -24898
rect 399574 -24954 399648 -24898
rect 399308 -25040 399648 -24954
rect 399308 -25096 399376 -25040
rect 399432 -25096 399518 -25040
rect 399574 -25096 399648 -25040
rect 399308 -25182 399648 -25096
rect 399308 -25238 399376 -25182
rect 399432 -25238 399518 -25182
rect 399574 -25238 399648 -25182
rect 399308 -25324 399648 -25238
rect 399308 -25380 399376 -25324
rect 399432 -25380 399518 -25324
rect 399574 -25380 399648 -25324
rect 399308 -25466 399648 -25380
rect 399308 -25522 399376 -25466
rect 399432 -25522 399518 -25466
rect 399574 -25522 399648 -25466
rect 399308 -25532 399648 -25522
rect 399708 -13680 400048 -13670
rect 399708 -13736 399776 -13680
rect 399832 -13736 399918 -13680
rect 399974 -13736 400048 -13680
rect 399708 -13822 400048 -13736
rect 399708 -13878 399776 -13822
rect 399832 -13878 399918 -13822
rect 399974 -13878 400048 -13822
rect 399708 -13964 400048 -13878
rect 399708 -14020 399776 -13964
rect 399832 -14020 399918 -13964
rect 399974 -14020 400048 -13964
rect 399708 -14106 400048 -14020
rect 399708 -14162 399776 -14106
rect 399832 -14162 399918 -14106
rect 399974 -14162 400048 -14106
rect 399708 -14248 400048 -14162
rect 399708 -14304 399776 -14248
rect 399832 -14304 399918 -14248
rect 399974 -14304 400048 -14248
rect 399708 -14390 400048 -14304
rect 399708 -14446 399776 -14390
rect 399832 -14446 399918 -14390
rect 399974 -14446 400048 -14390
rect 399708 -14532 400048 -14446
rect 399708 -14588 399776 -14532
rect 399832 -14588 399918 -14532
rect 399974 -14588 400048 -14532
rect 399708 -14674 400048 -14588
rect 399708 -14730 399776 -14674
rect 399832 -14730 399918 -14674
rect 399974 -14730 400048 -14674
rect 399708 -14816 400048 -14730
rect 399708 -14872 399776 -14816
rect 399832 -14872 399918 -14816
rect 399974 -14872 400048 -14816
rect 399708 -14958 400048 -14872
rect 399708 -15014 399776 -14958
rect 399832 -15014 399918 -14958
rect 399974 -15014 400048 -14958
rect 399708 -15100 400048 -15014
rect 399708 -15156 399776 -15100
rect 399832 -15156 399918 -15100
rect 399974 -15156 400048 -15100
rect 399708 -15242 400048 -15156
rect 399708 -15298 399776 -15242
rect 399832 -15298 399918 -15242
rect 399974 -15298 400048 -15242
rect 399708 -15384 400048 -15298
rect 399708 -15440 399776 -15384
rect 399832 -15440 399918 -15384
rect 399974 -15440 400048 -15384
rect 399708 -15526 400048 -15440
rect 399708 -15582 399776 -15526
rect 399832 -15582 399918 -15526
rect 399974 -15582 400048 -15526
rect 399708 -15668 400048 -15582
rect 399708 -15724 399776 -15668
rect 399832 -15724 399918 -15668
rect 399974 -15724 400048 -15668
rect 399708 -15810 400048 -15724
rect 399708 -15866 399776 -15810
rect 399832 -15866 399918 -15810
rect 399974 -15866 400048 -15810
rect 399708 -15952 400048 -15866
rect 399708 -16008 399776 -15952
rect 399832 -16008 399918 -15952
rect 399974 -16008 400048 -15952
rect 399708 -16094 400048 -16008
rect 399708 -16150 399776 -16094
rect 399832 -16150 399918 -16094
rect 399974 -16150 400048 -16094
rect 399708 -16236 400048 -16150
rect 399708 -16292 399776 -16236
rect 399832 -16292 399918 -16236
rect 399974 -16292 400048 -16236
rect 399708 -16378 400048 -16292
rect 399708 -16434 399776 -16378
rect 399832 -16434 399918 -16378
rect 399974 -16434 400048 -16378
rect 399708 -16520 400048 -16434
rect 399708 -16576 399776 -16520
rect 399832 -16576 399918 -16520
rect 399974 -16576 400048 -16520
rect 399708 -16662 400048 -16576
rect 399708 -16718 399776 -16662
rect 399832 -16718 399918 -16662
rect 399974 -16718 400048 -16662
rect 399708 -16804 400048 -16718
rect 399708 -16860 399776 -16804
rect 399832 -16860 399918 -16804
rect 399974 -16860 400048 -16804
rect 399708 -16946 400048 -16860
rect 399708 -17002 399776 -16946
rect 399832 -17002 399918 -16946
rect 399974 -17002 400048 -16946
rect 399708 -17088 400048 -17002
rect 399708 -17144 399776 -17088
rect 399832 -17144 399918 -17088
rect 399974 -17144 400048 -17088
rect 399708 -17230 400048 -17144
rect 399708 -17286 399776 -17230
rect 399832 -17286 399918 -17230
rect 399974 -17286 400048 -17230
rect 399708 -17372 400048 -17286
rect 399708 -17428 399776 -17372
rect 399832 -17428 399918 -17372
rect 399974 -17428 400048 -17372
rect 399708 -17514 400048 -17428
rect 399708 -17570 399776 -17514
rect 399832 -17570 399918 -17514
rect 399974 -17570 400048 -17514
rect 399708 -17656 400048 -17570
rect 399708 -17712 399776 -17656
rect 399832 -17712 399918 -17656
rect 399974 -17712 400048 -17656
rect 399708 -17798 400048 -17712
rect 399708 -17854 399776 -17798
rect 399832 -17854 399918 -17798
rect 399974 -17854 400048 -17798
rect 399708 -17940 400048 -17854
rect 399708 -17996 399776 -17940
rect 399832 -17996 399918 -17940
rect 399974 -17996 400048 -17940
rect 399708 -18082 400048 -17996
rect 399708 -18138 399776 -18082
rect 399832 -18138 399918 -18082
rect 399974 -18138 400048 -18082
rect 399708 -18224 400048 -18138
rect 399708 -18280 399776 -18224
rect 399832 -18280 399918 -18224
rect 399974 -18280 400048 -18224
rect 399708 -18366 400048 -18280
rect 399708 -18422 399776 -18366
rect 399832 -18422 399918 -18366
rect 399974 -18422 400048 -18366
rect 399708 -18508 400048 -18422
rect 399708 -18564 399776 -18508
rect 399832 -18564 399918 -18508
rect 399974 -18564 400048 -18508
rect 399708 -18650 400048 -18564
rect 399708 -18706 399776 -18650
rect 399832 -18706 399918 -18650
rect 399974 -18706 400048 -18650
rect 399708 -18792 400048 -18706
rect 399708 -18848 399776 -18792
rect 399832 -18848 399918 -18792
rect 399974 -18848 400048 -18792
rect 399708 -18934 400048 -18848
rect 399708 -18990 399776 -18934
rect 399832 -18990 399918 -18934
rect 399974 -18990 400048 -18934
rect 399708 -19076 400048 -18990
rect 399708 -19132 399776 -19076
rect 399832 -19132 399918 -19076
rect 399974 -19132 400048 -19076
rect 399708 -19218 400048 -19132
rect 399708 -19274 399776 -19218
rect 399832 -19274 399918 -19218
rect 399974 -19274 400048 -19218
rect 399708 -19360 400048 -19274
rect 399708 -19416 399776 -19360
rect 399832 -19416 399918 -19360
rect 399974 -19416 400048 -19360
rect 399708 -19502 400048 -19416
rect 399708 -19558 399776 -19502
rect 399832 -19558 399918 -19502
rect 399974 -19558 400048 -19502
rect 399708 -19644 400048 -19558
rect 399708 -19700 399776 -19644
rect 399832 -19700 399918 -19644
rect 399974 -19700 400048 -19644
rect 399708 -19786 400048 -19700
rect 399708 -19842 399776 -19786
rect 399832 -19842 399918 -19786
rect 399974 -19842 400048 -19786
rect 399708 -19928 400048 -19842
rect 399708 -19984 399776 -19928
rect 399832 -19984 399918 -19928
rect 399974 -19984 400048 -19928
rect 399708 -20070 400048 -19984
rect 399708 -20126 399776 -20070
rect 399832 -20126 399918 -20070
rect 399974 -20126 400048 -20070
rect 399708 -20212 400048 -20126
rect 399708 -20268 399776 -20212
rect 399832 -20268 399918 -20212
rect 399974 -20268 400048 -20212
rect 399708 -20354 400048 -20268
rect 399708 -20410 399776 -20354
rect 399832 -20410 399918 -20354
rect 399974 -20410 400048 -20354
rect 399708 -20496 400048 -20410
rect 399708 -20552 399776 -20496
rect 399832 -20552 399918 -20496
rect 399974 -20552 400048 -20496
rect 399708 -20638 400048 -20552
rect 399708 -20694 399776 -20638
rect 399832 -20694 399918 -20638
rect 399974 -20694 400048 -20638
rect 399708 -20780 400048 -20694
rect 399708 -20836 399776 -20780
rect 399832 -20836 399918 -20780
rect 399974 -20836 400048 -20780
rect 399708 -20922 400048 -20836
rect 399708 -20978 399776 -20922
rect 399832 -20978 399918 -20922
rect 399974 -20978 400048 -20922
rect 399708 -21064 400048 -20978
rect 399708 -21120 399776 -21064
rect 399832 -21120 399918 -21064
rect 399974 -21120 400048 -21064
rect 399708 -21206 400048 -21120
rect 399708 -21262 399776 -21206
rect 399832 -21262 399918 -21206
rect 399974 -21262 400048 -21206
rect 399708 -21348 400048 -21262
rect 399708 -21404 399776 -21348
rect 399832 -21404 399918 -21348
rect 399974 -21404 400048 -21348
rect 399708 -21490 400048 -21404
rect 399708 -21546 399776 -21490
rect 399832 -21546 399918 -21490
rect 399974 -21546 400048 -21490
rect 399708 -21632 400048 -21546
rect 399708 -21688 399776 -21632
rect 399832 -21688 399918 -21632
rect 399974 -21688 400048 -21632
rect 399708 -21774 400048 -21688
rect 399708 -21830 399776 -21774
rect 399832 -21830 399918 -21774
rect 399974 -21830 400048 -21774
rect 399708 -21916 400048 -21830
rect 399708 -21972 399776 -21916
rect 399832 -21972 399918 -21916
rect 399974 -21972 400048 -21916
rect 399708 -22058 400048 -21972
rect 399708 -22114 399776 -22058
rect 399832 -22114 399918 -22058
rect 399974 -22114 400048 -22058
rect 399708 -22200 400048 -22114
rect 399708 -22256 399776 -22200
rect 399832 -22256 399918 -22200
rect 399974 -22256 400048 -22200
rect 399708 -22342 400048 -22256
rect 399708 -22398 399776 -22342
rect 399832 -22398 399918 -22342
rect 399974 -22398 400048 -22342
rect 399708 -22484 400048 -22398
rect 399708 -22540 399776 -22484
rect 399832 -22540 399918 -22484
rect 399974 -22540 400048 -22484
rect 399708 -22626 400048 -22540
rect 399708 -22682 399776 -22626
rect 399832 -22682 399918 -22626
rect 399974 -22682 400048 -22626
rect 399708 -22768 400048 -22682
rect 399708 -22824 399776 -22768
rect 399832 -22824 399918 -22768
rect 399974 -22824 400048 -22768
rect 399708 -22910 400048 -22824
rect 399708 -22966 399776 -22910
rect 399832 -22966 399918 -22910
rect 399974 -22966 400048 -22910
rect 399708 -23052 400048 -22966
rect 399708 -23108 399776 -23052
rect 399832 -23108 399918 -23052
rect 399974 -23108 400048 -23052
rect 399708 -23194 400048 -23108
rect 399708 -23250 399776 -23194
rect 399832 -23250 399918 -23194
rect 399974 -23250 400048 -23194
rect 399708 -23336 400048 -23250
rect 399708 -23392 399776 -23336
rect 399832 -23392 399918 -23336
rect 399974 -23392 400048 -23336
rect 399708 -23478 400048 -23392
rect 399708 -23534 399776 -23478
rect 399832 -23534 399918 -23478
rect 399974 -23534 400048 -23478
rect 399708 -23620 400048 -23534
rect 399708 -23676 399776 -23620
rect 399832 -23676 399918 -23620
rect 399974 -23676 400048 -23620
rect 399708 -23762 400048 -23676
rect 399708 -23818 399776 -23762
rect 399832 -23818 399918 -23762
rect 399974 -23818 400048 -23762
rect 399708 -23904 400048 -23818
rect 399708 -23960 399776 -23904
rect 399832 -23960 399918 -23904
rect 399974 -23960 400048 -23904
rect 399708 -24046 400048 -23960
rect 399708 -24102 399776 -24046
rect 399832 -24102 399918 -24046
rect 399974 -24102 400048 -24046
rect 399708 -24188 400048 -24102
rect 399708 -24244 399776 -24188
rect 399832 -24244 399918 -24188
rect 399974 -24244 400048 -24188
rect 399708 -24330 400048 -24244
rect 399708 -24386 399776 -24330
rect 399832 -24386 399918 -24330
rect 399974 -24386 400048 -24330
rect 399708 -24472 400048 -24386
rect 399708 -24528 399776 -24472
rect 399832 -24528 399918 -24472
rect 399974 -24528 400048 -24472
rect 399708 -24614 400048 -24528
rect 399708 -24670 399776 -24614
rect 399832 -24670 399918 -24614
rect 399974 -24670 400048 -24614
rect 399708 -24756 400048 -24670
rect 399708 -24812 399776 -24756
rect 399832 -24812 399918 -24756
rect 399974 -24812 400048 -24756
rect 399708 -24898 400048 -24812
rect 399708 -24954 399776 -24898
rect 399832 -24954 399918 -24898
rect 399974 -24954 400048 -24898
rect 399708 -25040 400048 -24954
rect 399708 -25096 399776 -25040
rect 399832 -25096 399918 -25040
rect 399974 -25096 400048 -25040
rect 399708 -25182 400048 -25096
rect 399708 -25238 399776 -25182
rect 399832 -25238 399918 -25182
rect 399974 -25238 400048 -25182
rect 399708 -25324 400048 -25238
rect 399708 -25380 399776 -25324
rect 399832 -25380 399918 -25324
rect 399974 -25380 400048 -25324
rect 399708 -25466 400048 -25380
rect 399708 -25522 399776 -25466
rect 399832 -25522 399918 -25466
rect 399974 -25522 400048 -25466
rect 399708 -25532 400048 -25522
rect 400108 -13680 400448 -13670
rect 400108 -13736 400181 -13680
rect 400237 -13736 400323 -13680
rect 400379 -13736 400448 -13680
rect 400108 -13822 400448 -13736
rect 400108 -13878 400181 -13822
rect 400237 -13878 400323 -13822
rect 400379 -13878 400448 -13822
rect 400108 -13964 400448 -13878
rect 400108 -14020 400181 -13964
rect 400237 -14020 400323 -13964
rect 400379 -14020 400448 -13964
rect 400108 -14106 400448 -14020
rect 400108 -14162 400181 -14106
rect 400237 -14162 400323 -14106
rect 400379 -14162 400448 -14106
rect 400108 -14248 400448 -14162
rect 400108 -14304 400181 -14248
rect 400237 -14304 400323 -14248
rect 400379 -14304 400448 -14248
rect 400108 -14390 400448 -14304
rect 400108 -14446 400181 -14390
rect 400237 -14446 400323 -14390
rect 400379 -14446 400448 -14390
rect 400108 -14532 400448 -14446
rect 400108 -14588 400181 -14532
rect 400237 -14588 400323 -14532
rect 400379 -14588 400448 -14532
rect 400108 -14674 400448 -14588
rect 400108 -14730 400181 -14674
rect 400237 -14730 400323 -14674
rect 400379 -14730 400448 -14674
rect 400108 -14816 400448 -14730
rect 400108 -14872 400181 -14816
rect 400237 -14872 400323 -14816
rect 400379 -14872 400448 -14816
rect 400108 -14958 400448 -14872
rect 400108 -15014 400181 -14958
rect 400237 -15014 400323 -14958
rect 400379 -15014 400448 -14958
rect 400108 -15100 400448 -15014
rect 400108 -15156 400181 -15100
rect 400237 -15156 400323 -15100
rect 400379 -15156 400448 -15100
rect 400108 -15242 400448 -15156
rect 400108 -15298 400181 -15242
rect 400237 -15298 400323 -15242
rect 400379 -15298 400448 -15242
rect 400108 -15384 400448 -15298
rect 400108 -15440 400181 -15384
rect 400237 -15440 400323 -15384
rect 400379 -15440 400448 -15384
rect 400108 -15526 400448 -15440
rect 400108 -15582 400181 -15526
rect 400237 -15582 400323 -15526
rect 400379 -15582 400448 -15526
rect 400108 -15668 400448 -15582
rect 400108 -15724 400181 -15668
rect 400237 -15724 400323 -15668
rect 400379 -15724 400448 -15668
rect 400108 -15810 400448 -15724
rect 400108 -15866 400181 -15810
rect 400237 -15866 400323 -15810
rect 400379 -15866 400448 -15810
rect 400108 -15952 400448 -15866
rect 400108 -16008 400181 -15952
rect 400237 -16008 400323 -15952
rect 400379 -16008 400448 -15952
rect 400108 -16094 400448 -16008
rect 400108 -16150 400181 -16094
rect 400237 -16150 400323 -16094
rect 400379 -16150 400448 -16094
rect 400108 -16236 400448 -16150
rect 400108 -16292 400181 -16236
rect 400237 -16292 400323 -16236
rect 400379 -16292 400448 -16236
rect 400108 -16378 400448 -16292
rect 400108 -16434 400181 -16378
rect 400237 -16434 400323 -16378
rect 400379 -16434 400448 -16378
rect 400108 -16520 400448 -16434
rect 400108 -16576 400181 -16520
rect 400237 -16576 400323 -16520
rect 400379 -16576 400448 -16520
rect 400108 -16662 400448 -16576
rect 400108 -16718 400181 -16662
rect 400237 -16718 400323 -16662
rect 400379 -16718 400448 -16662
rect 400108 -16804 400448 -16718
rect 400108 -16860 400181 -16804
rect 400237 -16860 400323 -16804
rect 400379 -16860 400448 -16804
rect 400108 -16946 400448 -16860
rect 400108 -17002 400181 -16946
rect 400237 -17002 400323 -16946
rect 400379 -17002 400448 -16946
rect 400108 -17088 400448 -17002
rect 400108 -17144 400181 -17088
rect 400237 -17144 400323 -17088
rect 400379 -17144 400448 -17088
rect 400108 -17230 400448 -17144
rect 400108 -17286 400181 -17230
rect 400237 -17286 400323 -17230
rect 400379 -17286 400448 -17230
rect 400108 -17372 400448 -17286
rect 400108 -17428 400181 -17372
rect 400237 -17428 400323 -17372
rect 400379 -17428 400448 -17372
rect 400108 -17514 400448 -17428
rect 400108 -17570 400181 -17514
rect 400237 -17570 400323 -17514
rect 400379 -17570 400448 -17514
rect 400108 -17656 400448 -17570
rect 400108 -17712 400181 -17656
rect 400237 -17712 400323 -17656
rect 400379 -17712 400448 -17656
rect 400108 -17798 400448 -17712
rect 400108 -17854 400181 -17798
rect 400237 -17854 400323 -17798
rect 400379 -17854 400448 -17798
rect 400108 -17940 400448 -17854
rect 400108 -17996 400181 -17940
rect 400237 -17996 400323 -17940
rect 400379 -17996 400448 -17940
rect 400108 -18082 400448 -17996
rect 400108 -18138 400181 -18082
rect 400237 -18138 400323 -18082
rect 400379 -18138 400448 -18082
rect 400108 -18224 400448 -18138
rect 400108 -18280 400181 -18224
rect 400237 -18280 400323 -18224
rect 400379 -18280 400448 -18224
rect 400108 -18366 400448 -18280
rect 400108 -18422 400181 -18366
rect 400237 -18422 400323 -18366
rect 400379 -18422 400448 -18366
rect 400108 -18508 400448 -18422
rect 400108 -18564 400181 -18508
rect 400237 -18564 400323 -18508
rect 400379 -18564 400448 -18508
rect 400108 -18650 400448 -18564
rect 400108 -18706 400181 -18650
rect 400237 -18706 400323 -18650
rect 400379 -18706 400448 -18650
rect 400108 -18792 400448 -18706
rect 400108 -18848 400181 -18792
rect 400237 -18848 400323 -18792
rect 400379 -18848 400448 -18792
rect 400108 -18934 400448 -18848
rect 400108 -18990 400181 -18934
rect 400237 -18990 400323 -18934
rect 400379 -18990 400448 -18934
rect 400108 -19076 400448 -18990
rect 400108 -19132 400181 -19076
rect 400237 -19132 400323 -19076
rect 400379 -19132 400448 -19076
rect 400108 -19218 400448 -19132
rect 400108 -19274 400181 -19218
rect 400237 -19274 400323 -19218
rect 400379 -19274 400448 -19218
rect 400108 -19360 400448 -19274
rect 400108 -19416 400181 -19360
rect 400237 -19416 400323 -19360
rect 400379 -19416 400448 -19360
rect 400108 -19502 400448 -19416
rect 400108 -19558 400181 -19502
rect 400237 -19558 400323 -19502
rect 400379 -19558 400448 -19502
rect 400108 -19644 400448 -19558
rect 400108 -19700 400181 -19644
rect 400237 -19700 400323 -19644
rect 400379 -19700 400448 -19644
rect 400108 -19786 400448 -19700
rect 400108 -19842 400181 -19786
rect 400237 -19842 400323 -19786
rect 400379 -19842 400448 -19786
rect 400108 -19928 400448 -19842
rect 400108 -19984 400181 -19928
rect 400237 -19984 400323 -19928
rect 400379 -19984 400448 -19928
rect 400108 -20070 400448 -19984
rect 400108 -20126 400181 -20070
rect 400237 -20126 400323 -20070
rect 400379 -20126 400448 -20070
rect 400108 -20212 400448 -20126
rect 400108 -20268 400181 -20212
rect 400237 -20268 400323 -20212
rect 400379 -20268 400448 -20212
rect 400108 -20354 400448 -20268
rect 400108 -20410 400181 -20354
rect 400237 -20410 400323 -20354
rect 400379 -20410 400448 -20354
rect 400108 -20496 400448 -20410
rect 400108 -20552 400181 -20496
rect 400237 -20552 400323 -20496
rect 400379 -20552 400448 -20496
rect 400108 -20638 400448 -20552
rect 400108 -20694 400181 -20638
rect 400237 -20694 400323 -20638
rect 400379 -20694 400448 -20638
rect 400108 -20780 400448 -20694
rect 400108 -20836 400181 -20780
rect 400237 -20836 400323 -20780
rect 400379 -20836 400448 -20780
rect 400108 -20922 400448 -20836
rect 400108 -20978 400181 -20922
rect 400237 -20978 400323 -20922
rect 400379 -20978 400448 -20922
rect 400108 -21064 400448 -20978
rect 400108 -21120 400181 -21064
rect 400237 -21120 400323 -21064
rect 400379 -21120 400448 -21064
rect 400108 -21206 400448 -21120
rect 400108 -21262 400181 -21206
rect 400237 -21262 400323 -21206
rect 400379 -21262 400448 -21206
rect 400108 -21348 400448 -21262
rect 400108 -21404 400181 -21348
rect 400237 -21404 400323 -21348
rect 400379 -21404 400448 -21348
rect 400108 -21490 400448 -21404
rect 400108 -21546 400181 -21490
rect 400237 -21546 400323 -21490
rect 400379 -21546 400448 -21490
rect 400108 -21632 400448 -21546
rect 400108 -21688 400181 -21632
rect 400237 -21688 400323 -21632
rect 400379 -21688 400448 -21632
rect 400108 -21774 400448 -21688
rect 400108 -21830 400181 -21774
rect 400237 -21830 400323 -21774
rect 400379 -21830 400448 -21774
rect 400108 -21916 400448 -21830
rect 400108 -21972 400181 -21916
rect 400237 -21972 400323 -21916
rect 400379 -21972 400448 -21916
rect 400108 -22058 400448 -21972
rect 400108 -22114 400181 -22058
rect 400237 -22114 400323 -22058
rect 400379 -22114 400448 -22058
rect 400108 -22200 400448 -22114
rect 400108 -22256 400181 -22200
rect 400237 -22256 400323 -22200
rect 400379 -22256 400448 -22200
rect 400108 -22342 400448 -22256
rect 400108 -22398 400181 -22342
rect 400237 -22398 400323 -22342
rect 400379 -22398 400448 -22342
rect 400108 -22484 400448 -22398
rect 400108 -22540 400181 -22484
rect 400237 -22540 400323 -22484
rect 400379 -22540 400448 -22484
rect 400108 -22626 400448 -22540
rect 400108 -22682 400181 -22626
rect 400237 -22682 400323 -22626
rect 400379 -22682 400448 -22626
rect 400108 -22768 400448 -22682
rect 400108 -22824 400181 -22768
rect 400237 -22824 400323 -22768
rect 400379 -22824 400448 -22768
rect 400108 -22910 400448 -22824
rect 400108 -22966 400181 -22910
rect 400237 -22966 400323 -22910
rect 400379 -22966 400448 -22910
rect 400108 -23052 400448 -22966
rect 400108 -23108 400181 -23052
rect 400237 -23108 400323 -23052
rect 400379 -23108 400448 -23052
rect 400108 -23194 400448 -23108
rect 400108 -23250 400181 -23194
rect 400237 -23250 400323 -23194
rect 400379 -23250 400448 -23194
rect 400108 -23336 400448 -23250
rect 400108 -23392 400181 -23336
rect 400237 -23392 400323 -23336
rect 400379 -23392 400448 -23336
rect 400108 -23478 400448 -23392
rect 400108 -23534 400181 -23478
rect 400237 -23534 400323 -23478
rect 400379 -23534 400448 -23478
rect 400108 -23620 400448 -23534
rect 400108 -23676 400181 -23620
rect 400237 -23676 400323 -23620
rect 400379 -23676 400448 -23620
rect 400108 -23762 400448 -23676
rect 400108 -23818 400181 -23762
rect 400237 -23818 400323 -23762
rect 400379 -23818 400448 -23762
rect 400108 -23904 400448 -23818
rect 400108 -23960 400181 -23904
rect 400237 -23960 400323 -23904
rect 400379 -23960 400448 -23904
rect 400108 -24046 400448 -23960
rect 400108 -24102 400181 -24046
rect 400237 -24102 400323 -24046
rect 400379 -24102 400448 -24046
rect 400108 -24188 400448 -24102
rect 400108 -24244 400181 -24188
rect 400237 -24244 400323 -24188
rect 400379 -24244 400448 -24188
rect 400108 -24330 400448 -24244
rect 400108 -24386 400181 -24330
rect 400237 -24386 400323 -24330
rect 400379 -24386 400448 -24330
rect 400108 -24472 400448 -24386
rect 400108 -24528 400181 -24472
rect 400237 -24528 400323 -24472
rect 400379 -24528 400448 -24472
rect 400108 -24614 400448 -24528
rect 400108 -24670 400181 -24614
rect 400237 -24670 400323 -24614
rect 400379 -24670 400448 -24614
rect 400108 -24756 400448 -24670
rect 400108 -24812 400181 -24756
rect 400237 -24812 400323 -24756
rect 400379 -24812 400448 -24756
rect 400108 -24898 400448 -24812
rect 400108 -24954 400181 -24898
rect 400237 -24954 400323 -24898
rect 400379 -24954 400448 -24898
rect 400108 -25040 400448 -24954
rect 400108 -25096 400181 -25040
rect 400237 -25096 400323 -25040
rect 400379 -25096 400448 -25040
rect 400108 -25182 400448 -25096
rect 400108 -25238 400181 -25182
rect 400237 -25238 400323 -25182
rect 400379 -25238 400448 -25182
rect 400108 -25324 400448 -25238
rect 400108 -25380 400181 -25324
rect 400237 -25380 400323 -25324
rect 400379 -25380 400448 -25324
rect 400108 -25466 400448 -25380
rect 400108 -25522 400181 -25466
rect 400237 -25522 400323 -25466
rect 400379 -25522 400448 -25466
rect 400108 -25532 400448 -25522
rect 400640 -13688 400766 -13670
rect 400822 -13688 400890 -13632
rect 400946 -13688 401014 -13632
rect 401070 -13688 401138 -13632
rect 401194 -13688 401262 -13632
rect 401318 -13688 401440 -13632
rect 400640 -13756 401440 -13688
rect 400640 -13812 400766 -13756
rect 400822 -13812 400890 -13756
rect 400946 -13812 401014 -13756
rect 401070 -13812 401138 -13756
rect 401194 -13812 401262 -13756
rect 401318 -13812 401440 -13756
rect 400640 -13880 401440 -13812
rect 400640 -13936 400766 -13880
rect 400822 -13936 400890 -13880
rect 400946 -13936 401014 -13880
rect 401070 -13936 401138 -13880
rect 401194 -13936 401262 -13880
rect 401318 -13936 401440 -13880
rect 400640 -14004 401440 -13936
rect 400640 -14060 400766 -14004
rect 400822 -14060 400890 -14004
rect 400946 -14060 401014 -14004
rect 401070 -14060 401138 -14004
rect 401194 -14060 401262 -14004
rect 401318 -14060 401440 -14004
rect 400640 -14128 401440 -14060
rect 400640 -14184 400766 -14128
rect 400822 -14184 400890 -14128
rect 400946 -14184 401014 -14128
rect 401070 -14184 401138 -14128
rect 401194 -14184 401262 -14128
rect 401318 -14184 401440 -14128
rect 400640 -14252 401440 -14184
rect 400640 -14308 400766 -14252
rect 400822 -14308 400890 -14252
rect 400946 -14308 401014 -14252
rect 401070 -14308 401138 -14252
rect 401194 -14308 401262 -14252
rect 401318 -14308 401440 -14252
rect 400640 -14376 401440 -14308
rect 400640 -14432 400766 -14376
rect 400822 -14432 400890 -14376
rect 400946 -14432 401014 -14376
rect 401070 -14432 401138 -14376
rect 401194 -14432 401262 -14376
rect 401318 -14432 401440 -14376
rect 400640 -14500 401440 -14432
rect 400640 -14556 400766 -14500
rect 400822 -14556 400890 -14500
rect 400946 -14556 401014 -14500
rect 401070 -14556 401138 -14500
rect 401194 -14556 401262 -14500
rect 401318 -14556 401440 -14500
rect 400640 -14624 401440 -14556
rect 400640 -14680 400766 -14624
rect 400822 -14680 400890 -14624
rect 400946 -14680 401014 -14624
rect 401070 -14680 401138 -14624
rect 401194 -14680 401262 -14624
rect 401318 -14680 401440 -14624
rect 400640 -14748 401440 -14680
rect 400640 -14804 400766 -14748
rect 400822 -14804 400890 -14748
rect 400946 -14804 401014 -14748
rect 401070 -14804 401138 -14748
rect 401194 -14804 401262 -14748
rect 401318 -14804 401440 -14748
rect 400640 -14872 401440 -14804
rect 400640 -14928 400766 -14872
rect 400822 -14928 400890 -14872
rect 400946 -14928 401014 -14872
rect 401070 -14928 401138 -14872
rect 401194 -14928 401262 -14872
rect 401318 -14928 401440 -14872
rect 400640 -14996 401440 -14928
rect 400640 -15052 400766 -14996
rect 400822 -15052 400890 -14996
rect 400946 -15052 401014 -14996
rect 401070 -15052 401138 -14996
rect 401194 -15052 401262 -14996
rect 401318 -15052 401440 -14996
rect 400640 -15120 401440 -15052
rect 400640 -15176 400766 -15120
rect 400822 -15176 400890 -15120
rect 400946 -15176 401014 -15120
rect 401070 -15176 401138 -15120
rect 401194 -15176 401262 -15120
rect 401318 -15176 401440 -15120
rect 400640 -15244 401440 -15176
rect 400640 -15300 400766 -15244
rect 400822 -15300 400890 -15244
rect 400946 -15300 401014 -15244
rect 401070 -15300 401138 -15244
rect 401194 -15300 401262 -15244
rect 401318 -15300 401440 -15244
rect 400640 -15368 401440 -15300
rect 400640 -15424 400766 -15368
rect 400822 -15424 400890 -15368
rect 400946 -15424 401014 -15368
rect 401070 -15424 401138 -15368
rect 401194 -15424 401262 -15368
rect 401318 -15424 401440 -15368
rect 400640 -15492 401440 -15424
rect 400640 -15548 400766 -15492
rect 400822 -15548 400890 -15492
rect 400946 -15548 401014 -15492
rect 401070 -15548 401138 -15492
rect 401194 -15548 401262 -15492
rect 401318 -15548 401440 -15492
rect 400640 -15616 401440 -15548
rect 400640 -15672 400766 -15616
rect 400822 -15672 400890 -15616
rect 400946 -15672 401014 -15616
rect 401070 -15672 401138 -15616
rect 401194 -15672 401262 -15616
rect 401318 -15672 401440 -15616
rect 400640 -15740 401440 -15672
rect 400640 -15796 400766 -15740
rect 400822 -15796 400890 -15740
rect 400946 -15796 401014 -15740
rect 401070 -15796 401138 -15740
rect 401194 -15796 401262 -15740
rect 401318 -15796 401440 -15740
rect 400640 -15864 401440 -15796
rect 400640 -15920 400766 -15864
rect 400822 -15920 400890 -15864
rect 400946 -15920 401014 -15864
rect 401070 -15920 401138 -15864
rect 401194 -15920 401262 -15864
rect 401318 -15920 401440 -15864
rect 400640 -15988 401440 -15920
rect 400640 -16044 400766 -15988
rect 400822 -16044 400890 -15988
rect 400946 -16044 401014 -15988
rect 401070 -16044 401138 -15988
rect 401194 -16044 401262 -15988
rect 401318 -16044 401440 -15988
rect 400640 -16112 401440 -16044
rect 400640 -16168 400766 -16112
rect 400822 -16168 400890 -16112
rect 400946 -16168 401014 -16112
rect 401070 -16168 401138 -16112
rect 401194 -16168 401262 -16112
rect 401318 -16168 401440 -16112
rect 400640 -16236 401440 -16168
rect 400640 -16292 400766 -16236
rect 400822 -16292 400890 -16236
rect 400946 -16292 401014 -16236
rect 401070 -16292 401138 -16236
rect 401194 -16292 401262 -16236
rect 401318 -16292 401440 -16236
rect 400640 -16360 401440 -16292
rect 400640 -16416 400766 -16360
rect 400822 -16416 400890 -16360
rect 400946 -16416 401014 -16360
rect 401070 -16416 401138 -16360
rect 401194 -16416 401262 -16360
rect 401318 -16416 401440 -16360
rect 400640 -16484 401440 -16416
rect 400640 -16540 400766 -16484
rect 400822 -16540 400890 -16484
rect 400946 -16540 401014 -16484
rect 401070 -16540 401138 -16484
rect 401194 -16540 401262 -16484
rect 401318 -16540 401440 -16484
rect 400640 -16608 401440 -16540
rect 400640 -16664 400766 -16608
rect 400822 -16664 400890 -16608
rect 400946 -16664 401014 -16608
rect 401070 -16664 401138 -16608
rect 401194 -16664 401262 -16608
rect 401318 -16664 401440 -16608
rect 400640 -16732 401440 -16664
rect 400640 -16788 400766 -16732
rect 400822 -16788 400890 -16732
rect 400946 -16788 401014 -16732
rect 401070 -16788 401138 -16732
rect 401194 -16788 401262 -16732
rect 401318 -16788 401440 -16732
rect 400640 -16856 401440 -16788
rect 400640 -16912 400766 -16856
rect 400822 -16912 400890 -16856
rect 400946 -16912 401014 -16856
rect 401070 -16912 401138 -16856
rect 401194 -16912 401262 -16856
rect 401318 -16912 401440 -16856
rect 400640 -16980 401440 -16912
rect 400640 -17036 400766 -16980
rect 400822 -17036 400890 -16980
rect 400946 -17036 401014 -16980
rect 401070 -17036 401138 -16980
rect 401194 -17036 401262 -16980
rect 401318 -17036 401440 -16980
rect 400640 -17104 401440 -17036
rect 400640 -17160 400766 -17104
rect 400822 -17160 400890 -17104
rect 400946 -17160 401014 -17104
rect 401070 -17160 401138 -17104
rect 401194 -17160 401262 -17104
rect 401318 -17160 401440 -17104
rect 400640 -17228 401440 -17160
rect 400640 -17284 400766 -17228
rect 400822 -17284 400890 -17228
rect 400946 -17284 401014 -17228
rect 401070 -17284 401138 -17228
rect 401194 -17284 401262 -17228
rect 401318 -17284 401440 -17228
rect 400640 -17352 401440 -17284
rect 400640 -17408 400766 -17352
rect 400822 -17408 400890 -17352
rect 400946 -17408 401014 -17352
rect 401070 -17408 401138 -17352
rect 401194 -17408 401262 -17352
rect 401318 -17408 401440 -17352
rect 400640 -17476 401440 -17408
rect 400640 -17532 400766 -17476
rect 400822 -17532 400890 -17476
rect 400946 -17532 401014 -17476
rect 401070 -17532 401138 -17476
rect 401194 -17532 401262 -17476
rect 401318 -17532 401440 -17476
rect 400640 -17600 401440 -17532
rect 400640 -17656 400766 -17600
rect 400822 -17656 400890 -17600
rect 400946 -17656 401014 -17600
rect 401070 -17656 401138 -17600
rect 401194 -17656 401262 -17600
rect 401318 -17656 401440 -17600
rect 400640 -17724 401440 -17656
rect 400640 -17780 400766 -17724
rect 400822 -17780 400890 -17724
rect 400946 -17780 401014 -17724
rect 401070 -17780 401138 -17724
rect 401194 -17780 401262 -17724
rect 401318 -17780 401440 -17724
rect 400640 -17848 401440 -17780
rect 400640 -17904 400766 -17848
rect 400822 -17904 400890 -17848
rect 400946 -17904 401014 -17848
rect 401070 -17904 401138 -17848
rect 401194 -17904 401262 -17848
rect 401318 -17904 401440 -17848
rect 400640 -17972 401440 -17904
rect 400640 -18028 400766 -17972
rect 400822 -18028 400890 -17972
rect 400946 -18028 401014 -17972
rect 401070 -18028 401138 -17972
rect 401194 -18028 401262 -17972
rect 401318 -18028 401440 -17972
rect 400640 -18096 401440 -18028
rect 400640 -18152 400766 -18096
rect 400822 -18152 400890 -18096
rect 400946 -18152 401014 -18096
rect 401070 -18152 401138 -18096
rect 401194 -18152 401262 -18096
rect 401318 -18152 401440 -18096
rect 400640 -18220 401440 -18152
rect 400640 -18276 400766 -18220
rect 400822 -18276 400890 -18220
rect 400946 -18276 401014 -18220
rect 401070 -18276 401138 -18220
rect 401194 -18276 401262 -18220
rect 401318 -18276 401440 -18220
rect 400640 -18344 401440 -18276
rect 400640 -18400 400766 -18344
rect 400822 -18400 400890 -18344
rect 400946 -18400 401014 -18344
rect 401070 -18400 401138 -18344
rect 401194 -18400 401262 -18344
rect 401318 -18400 401440 -18344
rect 400640 -18468 401440 -18400
rect 400640 -18524 400766 -18468
rect 400822 -18524 400890 -18468
rect 400946 -18524 401014 -18468
rect 401070 -18524 401138 -18468
rect 401194 -18524 401262 -18468
rect 401318 -18524 401440 -18468
rect 400640 -18592 401440 -18524
rect 400640 -18648 400766 -18592
rect 400822 -18648 400890 -18592
rect 400946 -18648 401014 -18592
rect 401070 -18648 401138 -18592
rect 401194 -18648 401262 -18592
rect 401318 -18648 401440 -18592
rect 400640 -18716 401440 -18648
rect 400640 -18772 400766 -18716
rect 400822 -18772 400890 -18716
rect 400946 -18772 401014 -18716
rect 401070 -18772 401138 -18716
rect 401194 -18772 401262 -18716
rect 401318 -18772 401440 -18716
rect 400640 -18840 401440 -18772
rect 400640 -18896 400766 -18840
rect 400822 -18896 400890 -18840
rect 400946 -18896 401014 -18840
rect 401070 -18896 401138 -18840
rect 401194 -18896 401262 -18840
rect 401318 -18896 401440 -18840
rect 400640 -18964 401440 -18896
rect 400640 -19020 400766 -18964
rect 400822 -19020 400890 -18964
rect 400946 -19020 401014 -18964
rect 401070 -19020 401138 -18964
rect 401194 -19020 401262 -18964
rect 401318 -19020 401440 -18964
rect 400640 -19088 401440 -19020
rect 400640 -19144 400766 -19088
rect 400822 -19144 400890 -19088
rect 400946 -19144 401014 -19088
rect 401070 -19144 401138 -19088
rect 401194 -19144 401262 -19088
rect 401318 -19144 401440 -19088
rect 400640 -19212 401440 -19144
rect 400640 -19268 400766 -19212
rect 400822 -19268 400890 -19212
rect 400946 -19268 401014 -19212
rect 401070 -19268 401138 -19212
rect 401194 -19268 401262 -19212
rect 401318 -19268 401440 -19212
rect 400640 -19336 401440 -19268
rect 400640 -19392 400766 -19336
rect 400822 -19392 400890 -19336
rect 400946 -19392 401014 -19336
rect 401070 -19392 401138 -19336
rect 401194 -19392 401262 -19336
rect 401318 -19392 401440 -19336
rect 400640 -19460 401440 -19392
rect 400640 -19516 400766 -19460
rect 400822 -19516 400890 -19460
rect 400946 -19516 401014 -19460
rect 401070 -19516 401138 -19460
rect 401194 -19516 401262 -19460
rect 401318 -19516 401440 -19460
rect 400640 -19584 401440 -19516
rect 400640 -19640 400766 -19584
rect 400822 -19640 400890 -19584
rect 400946 -19640 401014 -19584
rect 401070 -19640 401138 -19584
rect 401194 -19640 401262 -19584
rect 401318 -19640 401440 -19584
rect 400640 -19708 401440 -19640
rect 400640 -19764 400766 -19708
rect 400822 -19764 400890 -19708
rect 400946 -19764 401014 -19708
rect 401070 -19764 401138 -19708
rect 401194 -19764 401262 -19708
rect 401318 -19764 401440 -19708
rect 400640 -19832 401440 -19764
rect 400640 -19888 400766 -19832
rect 400822 -19888 400890 -19832
rect 400946 -19888 401014 -19832
rect 401070 -19888 401138 -19832
rect 401194 -19888 401262 -19832
rect 401318 -19888 401440 -19832
rect 400640 -19956 401440 -19888
rect 400640 -20012 400766 -19956
rect 400822 -20012 400890 -19956
rect 400946 -20012 401014 -19956
rect 401070 -20012 401138 -19956
rect 401194 -20012 401262 -19956
rect 401318 -20012 401440 -19956
rect 400640 -20080 401440 -20012
rect 400640 -20136 400766 -20080
rect 400822 -20136 400890 -20080
rect 400946 -20136 401014 -20080
rect 401070 -20136 401138 -20080
rect 401194 -20136 401262 -20080
rect 401318 -20136 401440 -20080
rect 400640 -20204 401440 -20136
rect 400640 -20260 400766 -20204
rect 400822 -20260 400890 -20204
rect 400946 -20260 401014 -20204
rect 401070 -20260 401138 -20204
rect 401194 -20260 401262 -20204
rect 401318 -20260 401440 -20204
rect 400640 -20328 401440 -20260
rect 400640 -20384 400766 -20328
rect 400822 -20384 400890 -20328
rect 400946 -20384 401014 -20328
rect 401070 -20384 401138 -20328
rect 401194 -20384 401262 -20328
rect 401318 -20384 401440 -20328
rect 400640 -20452 401440 -20384
rect 400640 -20508 400766 -20452
rect 400822 -20508 400890 -20452
rect 400946 -20508 401014 -20452
rect 401070 -20508 401138 -20452
rect 401194 -20508 401262 -20452
rect 401318 -20508 401440 -20452
rect 400640 -20576 401440 -20508
rect 400640 -20632 400766 -20576
rect 400822 -20632 400890 -20576
rect 400946 -20632 401014 -20576
rect 401070 -20632 401138 -20576
rect 401194 -20632 401262 -20576
rect 401318 -20632 401440 -20576
rect 400640 -20700 401440 -20632
rect 400640 -20756 400766 -20700
rect 400822 -20756 400890 -20700
rect 400946 -20756 401014 -20700
rect 401070 -20756 401138 -20700
rect 401194 -20756 401262 -20700
rect 401318 -20756 401440 -20700
rect 400640 -20824 401440 -20756
rect 400640 -20880 400766 -20824
rect 400822 -20880 400890 -20824
rect 400946 -20880 401014 -20824
rect 401070 -20880 401138 -20824
rect 401194 -20880 401262 -20824
rect 401318 -20880 401440 -20824
rect 400640 -20948 401440 -20880
rect 400640 -21004 400766 -20948
rect 400822 -21004 400890 -20948
rect 400946 -21004 401014 -20948
rect 401070 -21004 401138 -20948
rect 401194 -21004 401262 -20948
rect 401318 -21004 401440 -20948
rect 400640 -21072 401440 -21004
rect 400640 -21128 400766 -21072
rect 400822 -21128 400890 -21072
rect 400946 -21128 401014 -21072
rect 401070 -21128 401138 -21072
rect 401194 -21128 401262 -21072
rect 401318 -21128 401440 -21072
rect 400640 -21196 401440 -21128
rect 400640 -21252 400766 -21196
rect 400822 -21252 400890 -21196
rect 400946 -21252 401014 -21196
rect 401070 -21252 401138 -21196
rect 401194 -21252 401262 -21196
rect 401318 -21252 401440 -21196
rect 400640 -21320 401440 -21252
rect 400640 -21376 400766 -21320
rect 400822 -21376 400890 -21320
rect 400946 -21376 401014 -21320
rect 401070 -21376 401138 -21320
rect 401194 -21376 401262 -21320
rect 401318 -21376 401440 -21320
rect 400640 -21444 401440 -21376
rect 400640 -21500 400766 -21444
rect 400822 -21500 400890 -21444
rect 400946 -21500 401014 -21444
rect 401070 -21500 401138 -21444
rect 401194 -21500 401262 -21444
rect 401318 -21500 401440 -21444
rect 400640 -21568 401440 -21500
rect 400640 -21624 400766 -21568
rect 400822 -21624 400890 -21568
rect 400946 -21624 401014 -21568
rect 401070 -21624 401138 -21568
rect 401194 -21624 401262 -21568
rect 401318 -21624 401440 -21568
rect 400640 -21692 401440 -21624
rect 400640 -21748 400766 -21692
rect 400822 -21748 400890 -21692
rect 400946 -21748 401014 -21692
rect 401070 -21748 401138 -21692
rect 401194 -21748 401262 -21692
rect 401318 -21748 401440 -21692
rect 400640 -21816 401440 -21748
rect 400640 -21872 400766 -21816
rect 400822 -21872 400890 -21816
rect 400946 -21872 401014 -21816
rect 401070 -21872 401138 -21816
rect 401194 -21872 401262 -21816
rect 401318 -21872 401440 -21816
rect 400640 -21940 401440 -21872
rect 400640 -21996 400766 -21940
rect 400822 -21996 400890 -21940
rect 400946 -21996 401014 -21940
rect 401070 -21996 401138 -21940
rect 401194 -21996 401262 -21940
rect 401318 -21996 401440 -21940
rect 400640 -22064 401440 -21996
rect 400640 -22120 400766 -22064
rect 400822 -22120 400890 -22064
rect 400946 -22120 401014 -22064
rect 401070 -22120 401138 -22064
rect 401194 -22120 401262 -22064
rect 401318 -22120 401440 -22064
rect 400640 -22188 401440 -22120
rect 400640 -22244 400766 -22188
rect 400822 -22244 400890 -22188
rect 400946 -22244 401014 -22188
rect 401070 -22244 401138 -22188
rect 401194 -22244 401262 -22188
rect 401318 -22244 401440 -22188
rect 400640 -22312 401440 -22244
rect 400640 -22368 400766 -22312
rect 400822 -22368 400890 -22312
rect 400946 -22368 401014 -22312
rect 401070 -22368 401138 -22312
rect 401194 -22368 401262 -22312
rect 401318 -22368 401440 -22312
rect 400640 -22436 401440 -22368
rect 400640 -22492 400766 -22436
rect 400822 -22492 400890 -22436
rect 400946 -22492 401014 -22436
rect 401070 -22492 401138 -22436
rect 401194 -22492 401262 -22436
rect 401318 -22492 401440 -22436
rect 400640 -22560 401440 -22492
rect 400640 -22616 400766 -22560
rect 400822 -22616 400890 -22560
rect 400946 -22616 401014 -22560
rect 401070 -22616 401138 -22560
rect 401194 -22616 401262 -22560
rect 401318 -22616 401440 -22560
rect 400640 -22684 401440 -22616
rect 400640 -22740 400766 -22684
rect 400822 -22740 400890 -22684
rect 400946 -22740 401014 -22684
rect 401070 -22740 401138 -22684
rect 401194 -22740 401262 -22684
rect 401318 -22740 401440 -22684
rect 400640 -22808 401440 -22740
rect 400640 -22864 400766 -22808
rect 400822 -22864 400890 -22808
rect 400946 -22864 401014 -22808
rect 401070 -22864 401138 -22808
rect 401194 -22864 401262 -22808
rect 401318 -22864 401440 -22808
rect 400640 -22932 401440 -22864
rect 400640 -22988 400766 -22932
rect 400822 -22988 400890 -22932
rect 400946 -22988 401014 -22932
rect 401070 -22988 401138 -22932
rect 401194 -22988 401262 -22932
rect 401318 -22988 401440 -22932
rect 400640 -23056 401440 -22988
rect 400640 -23112 400766 -23056
rect 400822 -23112 400890 -23056
rect 400946 -23112 401014 -23056
rect 401070 -23112 401138 -23056
rect 401194 -23112 401262 -23056
rect 401318 -23112 401440 -23056
rect 400640 -23180 401440 -23112
rect 400640 -23236 400766 -23180
rect 400822 -23236 400890 -23180
rect 400946 -23236 401014 -23180
rect 401070 -23236 401138 -23180
rect 401194 -23236 401262 -23180
rect 401318 -23236 401440 -23180
rect 400640 -23304 401440 -23236
rect 400640 -23360 400766 -23304
rect 400822 -23360 400890 -23304
rect 400946 -23360 401014 -23304
rect 401070 -23360 401138 -23304
rect 401194 -23360 401262 -23304
rect 401318 -23360 401440 -23304
rect 400640 -23428 401440 -23360
rect 400640 -23484 400766 -23428
rect 400822 -23484 400890 -23428
rect 400946 -23484 401014 -23428
rect 401070 -23484 401138 -23428
rect 401194 -23484 401262 -23428
rect 401318 -23484 401440 -23428
rect 400640 -23552 401440 -23484
rect 400640 -23608 400766 -23552
rect 400822 -23608 400890 -23552
rect 400946 -23608 401014 -23552
rect 401070 -23608 401138 -23552
rect 401194 -23608 401262 -23552
rect 401318 -23608 401440 -23552
rect 400640 -23676 401440 -23608
rect 400640 -23732 400766 -23676
rect 400822 -23732 400890 -23676
rect 400946 -23732 401014 -23676
rect 401070 -23732 401138 -23676
rect 401194 -23732 401262 -23676
rect 401318 -23732 401440 -23676
rect 400640 -23800 401440 -23732
rect 400640 -23856 400766 -23800
rect 400822 -23856 400890 -23800
rect 400946 -23856 401014 -23800
rect 401070 -23856 401138 -23800
rect 401194 -23856 401262 -23800
rect 401318 -23856 401440 -23800
rect 400640 -23924 401440 -23856
rect 400640 -23980 400766 -23924
rect 400822 -23980 400890 -23924
rect 400946 -23980 401014 -23924
rect 401070 -23980 401138 -23924
rect 401194 -23980 401262 -23924
rect 401318 -23980 401440 -23924
rect 400640 -24048 401440 -23980
rect 400640 -24104 400766 -24048
rect 400822 -24104 400890 -24048
rect 400946 -24104 401014 -24048
rect 401070 -24104 401138 -24048
rect 401194 -24104 401262 -24048
rect 401318 -24104 401440 -24048
rect 400640 -24172 401440 -24104
rect 400640 -24228 400766 -24172
rect 400822 -24228 400890 -24172
rect 400946 -24228 401014 -24172
rect 401070 -24228 401138 -24172
rect 401194 -24228 401262 -24172
rect 401318 -24228 401440 -24172
rect 400640 -24296 401440 -24228
rect 400640 -24352 400766 -24296
rect 400822 -24352 400890 -24296
rect 400946 -24352 401014 -24296
rect 401070 -24352 401138 -24296
rect 401194 -24352 401262 -24296
rect 401318 -24352 401440 -24296
rect 400640 -24420 401440 -24352
rect 400640 -24476 400766 -24420
rect 400822 -24476 400890 -24420
rect 400946 -24476 401014 -24420
rect 401070 -24476 401138 -24420
rect 401194 -24476 401262 -24420
rect 401318 -24476 401440 -24420
rect 400640 -24544 401440 -24476
rect 400640 -24600 400766 -24544
rect 400822 -24600 400890 -24544
rect 400946 -24600 401014 -24544
rect 401070 -24600 401138 -24544
rect 401194 -24600 401262 -24544
rect 401318 -24600 401440 -24544
rect 400640 -24668 401440 -24600
rect 400640 -24724 400766 -24668
rect 400822 -24724 400890 -24668
rect 400946 -24724 401014 -24668
rect 401070 -24724 401138 -24668
rect 401194 -24724 401262 -24668
rect 401318 -24724 401440 -24668
rect 400640 -24792 401440 -24724
rect 400640 -24848 400766 -24792
rect 400822 -24848 400890 -24792
rect 400946 -24848 401014 -24792
rect 401070 -24848 401138 -24792
rect 401194 -24848 401262 -24792
rect 401318 -24848 401440 -24792
rect 400640 -24916 401440 -24848
rect 400640 -24972 400766 -24916
rect 400822 -24972 400890 -24916
rect 400946 -24972 401014 -24916
rect 401070 -24972 401138 -24916
rect 401194 -24972 401262 -24916
rect 401318 -24972 401440 -24916
rect 400640 -25040 401440 -24972
rect 400640 -25096 400766 -25040
rect 400822 -25096 400890 -25040
rect 400946 -25096 401014 -25040
rect 401070 -25096 401138 -25040
rect 401194 -25096 401262 -25040
rect 401318 -25096 401440 -25040
rect 400640 -25164 401440 -25096
rect 400640 -25220 400766 -25164
rect 400822 -25220 400890 -25164
rect 400946 -25220 401014 -25164
rect 401070 -25220 401138 -25164
rect 401194 -25220 401262 -25164
rect 401318 -25220 401440 -25164
rect 400640 -25288 401440 -25220
rect 400640 -25344 400766 -25288
rect 400822 -25344 400890 -25288
rect 400946 -25344 401014 -25288
rect 401070 -25344 401138 -25288
rect 401194 -25344 401262 -25288
rect 401318 -25344 401440 -25288
rect 400640 -25412 401440 -25344
rect 400640 -25468 400766 -25412
rect 400822 -25468 400890 -25412
rect 400946 -25468 401014 -25412
rect 401070 -25468 401138 -25412
rect 401194 -25468 401262 -25412
rect 401318 -25468 401440 -25412
rect 400640 -25532 401440 -25468
rect 387840 -25536 401440 -25532
rect 387840 -25592 387954 -25536
rect 388010 -25592 388078 -25536
rect 388134 -25592 388202 -25536
rect 388258 -25592 388326 -25536
rect 388382 -25592 388450 -25536
rect 388506 -25592 400766 -25536
rect 400822 -25592 400890 -25536
rect 400946 -25592 401014 -25536
rect 401070 -25592 401138 -25536
rect 401194 -25592 401262 -25536
rect 401318 -25592 401440 -25536
rect 387840 -25660 401440 -25592
rect 387840 -25716 387954 -25660
rect 388010 -25716 388078 -25660
rect 388134 -25716 388202 -25660
rect 388258 -25716 388326 -25660
rect 388382 -25716 388450 -25660
rect 388506 -25688 400766 -25660
rect 388506 -25716 388655 -25688
rect 387840 -25744 388655 -25716
rect 388711 -25744 388797 -25688
rect 388853 -25744 388939 -25688
rect 388995 -25744 389081 -25688
rect 389137 -25744 389223 -25688
rect 389279 -25744 389365 -25688
rect 389421 -25744 389507 -25688
rect 389563 -25744 389649 -25688
rect 389705 -25744 389791 -25688
rect 389847 -25744 389933 -25688
rect 389989 -25744 390075 -25688
rect 390131 -25744 390217 -25688
rect 390273 -25744 390359 -25688
rect 390415 -25744 390501 -25688
rect 390557 -25744 390643 -25688
rect 390699 -25744 390785 -25688
rect 390841 -25744 390927 -25688
rect 390983 -25744 391069 -25688
rect 391125 -25744 391211 -25688
rect 391267 -25744 391353 -25688
rect 391409 -25744 391495 -25688
rect 391551 -25744 391637 -25688
rect 391693 -25744 391779 -25688
rect 391835 -25744 391921 -25688
rect 391977 -25744 392063 -25688
rect 392119 -25744 392205 -25688
rect 392261 -25744 392347 -25688
rect 392403 -25744 392489 -25688
rect 392545 -25744 392631 -25688
rect 392687 -25744 392773 -25688
rect 392829 -25744 392915 -25688
rect 392971 -25744 393057 -25688
rect 393113 -25744 393199 -25688
rect 393255 -25744 393341 -25688
rect 393397 -25744 393483 -25688
rect 393539 -25744 393625 -25688
rect 393681 -25744 393767 -25688
rect 393823 -25744 393909 -25688
rect 393965 -25744 394051 -25688
rect 394107 -25744 394193 -25688
rect 394249 -25744 394335 -25688
rect 394391 -25744 394477 -25688
rect 394533 -25744 394619 -25688
rect 394675 -25744 394761 -25688
rect 394817 -25744 394903 -25688
rect 394959 -25744 395045 -25688
rect 395101 -25744 395187 -25688
rect 395243 -25744 395329 -25688
rect 395385 -25744 395471 -25688
rect 395527 -25744 395613 -25688
rect 395669 -25744 395755 -25688
rect 395811 -25744 395897 -25688
rect 395953 -25744 396039 -25688
rect 396095 -25744 396181 -25688
rect 396237 -25744 396323 -25688
rect 396379 -25744 396465 -25688
rect 396521 -25744 396607 -25688
rect 396663 -25744 396749 -25688
rect 396805 -25744 396891 -25688
rect 396947 -25744 397033 -25688
rect 397089 -25744 397175 -25688
rect 397231 -25744 397317 -25688
rect 397373 -25744 397459 -25688
rect 397515 -25744 397601 -25688
rect 397657 -25744 397743 -25688
rect 397799 -25744 397885 -25688
rect 397941 -25744 398027 -25688
rect 398083 -25744 398169 -25688
rect 398225 -25744 398311 -25688
rect 398367 -25744 398453 -25688
rect 398509 -25744 398595 -25688
rect 398651 -25744 398737 -25688
rect 398793 -25744 398879 -25688
rect 398935 -25744 399021 -25688
rect 399077 -25744 399163 -25688
rect 399219 -25744 399305 -25688
rect 399361 -25744 399447 -25688
rect 399503 -25744 399589 -25688
rect 399645 -25744 399731 -25688
rect 399787 -25744 399873 -25688
rect 399929 -25744 400015 -25688
rect 400071 -25744 400157 -25688
rect 400213 -25744 400299 -25688
rect 400355 -25744 400441 -25688
rect 400497 -25744 400583 -25688
rect 400639 -25716 400766 -25688
rect 400822 -25716 400890 -25660
rect 400946 -25716 401014 -25660
rect 401070 -25716 401138 -25660
rect 401194 -25716 401262 -25660
rect 401318 -25716 401440 -25660
rect 400639 -25744 401440 -25716
rect 387840 -25784 401440 -25744
rect 387840 -25840 387954 -25784
rect 388010 -25840 388078 -25784
rect 388134 -25840 388202 -25784
rect 388258 -25840 388326 -25784
rect 388382 -25840 388450 -25784
rect 388506 -25830 400766 -25784
rect 388506 -25840 388655 -25830
rect 387840 -25886 388655 -25840
rect 388711 -25886 388797 -25830
rect 388853 -25886 388939 -25830
rect 388995 -25886 389081 -25830
rect 389137 -25886 389223 -25830
rect 389279 -25886 389365 -25830
rect 389421 -25886 389507 -25830
rect 389563 -25886 389649 -25830
rect 389705 -25886 389791 -25830
rect 389847 -25886 389933 -25830
rect 389989 -25886 390075 -25830
rect 390131 -25886 390217 -25830
rect 390273 -25886 390359 -25830
rect 390415 -25886 390501 -25830
rect 390557 -25886 390643 -25830
rect 390699 -25886 390785 -25830
rect 390841 -25886 390927 -25830
rect 390983 -25886 391069 -25830
rect 391125 -25886 391211 -25830
rect 391267 -25886 391353 -25830
rect 391409 -25886 391495 -25830
rect 391551 -25886 391637 -25830
rect 391693 -25886 391779 -25830
rect 391835 -25886 391921 -25830
rect 391977 -25886 392063 -25830
rect 392119 -25886 392205 -25830
rect 392261 -25886 392347 -25830
rect 392403 -25886 392489 -25830
rect 392545 -25886 392631 -25830
rect 392687 -25886 392773 -25830
rect 392829 -25886 392915 -25830
rect 392971 -25886 393057 -25830
rect 393113 -25886 393199 -25830
rect 393255 -25886 393341 -25830
rect 393397 -25886 393483 -25830
rect 393539 -25886 393625 -25830
rect 393681 -25886 393767 -25830
rect 393823 -25886 393909 -25830
rect 393965 -25886 394051 -25830
rect 394107 -25886 394193 -25830
rect 394249 -25886 394335 -25830
rect 394391 -25886 394477 -25830
rect 394533 -25886 394619 -25830
rect 394675 -25886 394761 -25830
rect 394817 -25886 394903 -25830
rect 394959 -25886 395045 -25830
rect 395101 -25886 395187 -25830
rect 395243 -25886 395329 -25830
rect 395385 -25886 395471 -25830
rect 395527 -25886 395613 -25830
rect 395669 -25886 395755 -25830
rect 395811 -25886 395897 -25830
rect 395953 -25886 396039 -25830
rect 396095 -25886 396181 -25830
rect 396237 -25886 396323 -25830
rect 396379 -25886 396465 -25830
rect 396521 -25886 396607 -25830
rect 396663 -25886 396749 -25830
rect 396805 -25886 396891 -25830
rect 396947 -25886 397033 -25830
rect 397089 -25886 397175 -25830
rect 397231 -25886 397317 -25830
rect 397373 -25886 397459 -25830
rect 397515 -25886 397601 -25830
rect 397657 -25886 397743 -25830
rect 397799 -25886 397885 -25830
rect 397941 -25886 398027 -25830
rect 398083 -25886 398169 -25830
rect 398225 -25886 398311 -25830
rect 398367 -25886 398453 -25830
rect 398509 -25886 398595 -25830
rect 398651 -25886 398737 -25830
rect 398793 -25886 398879 -25830
rect 398935 -25886 399021 -25830
rect 399077 -25886 399163 -25830
rect 399219 -25886 399305 -25830
rect 399361 -25886 399447 -25830
rect 399503 -25886 399589 -25830
rect 399645 -25886 399731 -25830
rect 399787 -25886 399873 -25830
rect 399929 -25886 400015 -25830
rect 400071 -25886 400157 -25830
rect 400213 -25886 400299 -25830
rect 400355 -25886 400441 -25830
rect 400497 -25886 400583 -25830
rect 400639 -25840 400766 -25830
rect 400822 -25840 400890 -25784
rect 400946 -25840 401014 -25784
rect 401070 -25840 401138 -25784
rect 401194 -25840 401262 -25784
rect 401318 -25840 401440 -25784
rect 400639 -25886 401440 -25840
rect 387840 -25990 401440 -25886
<< via3 >>
rect 387986 -13097 388042 -13041
rect 388110 -13097 388166 -13041
rect 388234 -13097 388290 -13041
rect 388358 -13097 388414 -13041
rect 388482 -13097 388538 -13041
rect 388606 -13097 388662 -13041
rect 388730 -13097 388786 -13041
rect 388854 -13097 388910 -13041
rect 388978 -13097 389034 -13041
rect 389102 -13097 389158 -13041
rect 389226 -13097 389282 -13041
rect 389350 -13097 389406 -13041
rect 389474 -13097 389530 -13041
rect 389598 -13097 389654 -13041
rect 389722 -13097 389778 -13041
rect 389846 -13097 389902 -13041
rect 389970 -13097 390026 -13041
rect 390094 -13097 390150 -13041
rect 390218 -13097 390274 -13041
rect 390342 -13097 390398 -13041
rect 390466 -13097 390522 -13041
rect 390590 -13097 390646 -13041
rect 390714 -13097 390770 -13041
rect 390838 -13097 390894 -13041
rect 390962 -13097 391018 -13041
rect 391086 -13097 391142 -13041
rect 391210 -13097 391266 -13041
rect 391334 -13097 391390 -13041
rect 391458 -13097 391514 -13041
rect 391582 -13097 391638 -13041
rect 391706 -13097 391762 -13041
rect 391830 -13097 391886 -13041
rect 391954 -13097 392010 -13041
rect 392078 -13097 392134 -13041
rect 392202 -13097 392258 -13041
rect 392326 -13097 392382 -13041
rect 392450 -13097 392506 -13041
rect 392574 -13097 392630 -13041
rect 392698 -13097 392754 -13041
rect 392822 -13097 392878 -13041
rect 392946 -13097 393002 -13041
rect 393070 -13097 393126 -13041
rect 393194 -13097 393250 -13041
rect 393318 -13097 393374 -13041
rect 393442 -13097 393498 -13041
rect 393566 -13097 393622 -13041
rect 393690 -13097 393746 -13041
rect 393814 -13097 393870 -13041
rect 393938 -13097 393994 -13041
rect 394062 -13097 394118 -13041
rect 394186 -13097 394242 -13041
rect 394310 -13097 394366 -13041
rect 394434 -13097 394490 -13041
rect 394558 -13097 394614 -13041
rect 394682 -13097 394738 -13041
rect 394806 -13097 394862 -13041
rect 394930 -13097 394986 -13041
rect 395054 -13097 395110 -13041
rect 395178 -13097 395234 -13041
rect 395302 -13097 395358 -13041
rect 395426 -13097 395482 -13041
rect 395550 -13097 395606 -13041
rect 395674 -13097 395730 -13041
rect 395798 -13097 395854 -13041
rect 395922 -13097 395978 -13041
rect 396046 -13097 396102 -13041
rect 396170 -13097 396226 -13041
rect 396294 -13097 396350 -13041
rect 396418 -13097 396474 -13041
rect 396542 -13097 396598 -13041
rect 396666 -13097 396722 -13041
rect 396790 -13097 396846 -13041
rect 396914 -13097 396970 -13041
rect 397038 -13097 397094 -13041
rect 397162 -13097 397218 -13041
rect 397286 -13097 397342 -13041
rect 397410 -13097 397466 -13041
rect 397534 -13097 397590 -13041
rect 397658 -13097 397714 -13041
rect 397782 -13097 397838 -13041
rect 397906 -13097 397962 -13041
rect 398030 -13097 398086 -13041
rect 398154 -13097 398210 -13041
rect 398278 -13097 398334 -13041
rect 398402 -13097 398458 -13041
rect 398526 -13097 398582 -13041
rect 398650 -13097 398706 -13041
rect 398774 -13097 398830 -13041
rect 398898 -13097 398954 -13041
rect 399022 -13097 399078 -13041
rect 399146 -13097 399202 -13041
rect 399270 -13097 399326 -13041
rect 399394 -13097 399450 -13041
rect 399518 -13097 399574 -13041
rect 399642 -13097 399698 -13041
rect 399766 -13097 399822 -13041
rect 399890 -13097 399946 -13041
rect 400014 -13097 400070 -13041
rect 400138 -13097 400194 -13041
rect 400262 -13097 400318 -13041
rect 400386 -13097 400442 -13041
rect 400510 -13097 400566 -13041
rect 400634 -13097 400690 -13041
rect 400758 -13097 400814 -13041
rect 400882 -13097 400938 -13041
rect 401006 -13097 401062 -13041
rect 401130 -13097 401186 -13041
rect 401254 -13097 401310 -13041
rect 387986 -13221 388042 -13165
rect 388110 -13221 388166 -13165
rect 388234 -13221 388290 -13165
rect 388358 -13221 388414 -13165
rect 388482 -13221 388538 -13165
rect 388606 -13221 388662 -13165
rect 388730 -13221 388786 -13165
rect 388854 -13221 388910 -13165
rect 388978 -13221 389034 -13165
rect 389102 -13221 389158 -13165
rect 389226 -13221 389282 -13165
rect 389350 -13221 389406 -13165
rect 389474 -13221 389530 -13165
rect 389598 -13221 389654 -13165
rect 389722 -13221 389778 -13165
rect 389846 -13221 389902 -13165
rect 389970 -13221 390026 -13165
rect 390094 -13221 390150 -13165
rect 390218 -13221 390274 -13165
rect 390342 -13221 390398 -13165
rect 390466 -13221 390522 -13165
rect 390590 -13221 390646 -13165
rect 390714 -13221 390770 -13165
rect 390838 -13221 390894 -13165
rect 390962 -13221 391018 -13165
rect 391086 -13221 391142 -13165
rect 391210 -13221 391266 -13165
rect 391334 -13221 391390 -13165
rect 391458 -13221 391514 -13165
rect 391582 -13221 391638 -13165
rect 391706 -13221 391762 -13165
rect 391830 -13221 391886 -13165
rect 391954 -13221 392010 -13165
rect 392078 -13221 392134 -13165
rect 392202 -13221 392258 -13165
rect 392326 -13221 392382 -13165
rect 392450 -13221 392506 -13165
rect 392574 -13221 392630 -13165
rect 392698 -13221 392754 -13165
rect 392822 -13221 392878 -13165
rect 392946 -13221 393002 -13165
rect 393070 -13221 393126 -13165
rect 393194 -13221 393250 -13165
rect 393318 -13221 393374 -13165
rect 393442 -13221 393498 -13165
rect 393566 -13221 393622 -13165
rect 393690 -13221 393746 -13165
rect 393814 -13221 393870 -13165
rect 393938 -13221 393994 -13165
rect 394062 -13221 394118 -13165
rect 394186 -13221 394242 -13165
rect 394310 -13221 394366 -13165
rect 394434 -13221 394490 -13165
rect 394558 -13221 394614 -13165
rect 394682 -13221 394738 -13165
rect 394806 -13221 394862 -13165
rect 394930 -13221 394986 -13165
rect 395054 -13221 395110 -13165
rect 395178 -13221 395234 -13165
rect 395302 -13221 395358 -13165
rect 395426 -13221 395482 -13165
rect 395550 -13221 395606 -13165
rect 395674 -13221 395730 -13165
rect 395798 -13221 395854 -13165
rect 395922 -13221 395978 -13165
rect 396046 -13221 396102 -13165
rect 396170 -13221 396226 -13165
rect 396294 -13221 396350 -13165
rect 396418 -13221 396474 -13165
rect 396542 -13221 396598 -13165
rect 396666 -13221 396722 -13165
rect 396790 -13221 396846 -13165
rect 396914 -13221 396970 -13165
rect 397038 -13221 397094 -13165
rect 397162 -13221 397218 -13165
rect 397286 -13221 397342 -13165
rect 397410 -13221 397466 -13165
rect 397534 -13221 397590 -13165
rect 397658 -13221 397714 -13165
rect 397782 -13221 397838 -13165
rect 397906 -13221 397962 -13165
rect 398030 -13221 398086 -13165
rect 398154 -13221 398210 -13165
rect 398278 -13221 398334 -13165
rect 398402 -13221 398458 -13165
rect 398526 -13221 398582 -13165
rect 398650 -13221 398706 -13165
rect 398774 -13221 398830 -13165
rect 398898 -13221 398954 -13165
rect 399022 -13221 399078 -13165
rect 399146 -13221 399202 -13165
rect 399270 -13221 399326 -13165
rect 399394 -13221 399450 -13165
rect 399518 -13221 399574 -13165
rect 399642 -13221 399698 -13165
rect 399766 -13221 399822 -13165
rect 399890 -13221 399946 -13165
rect 400014 -13221 400070 -13165
rect 400138 -13221 400194 -13165
rect 400262 -13221 400318 -13165
rect 400386 -13221 400442 -13165
rect 400510 -13221 400566 -13165
rect 400634 -13221 400690 -13165
rect 400758 -13221 400814 -13165
rect 400882 -13221 400938 -13165
rect 401006 -13221 401062 -13165
rect 401130 -13221 401186 -13165
rect 401254 -13221 401310 -13165
rect 387986 -13345 388042 -13289
rect 388110 -13345 388166 -13289
rect 388234 -13345 388290 -13289
rect 388358 -13345 388414 -13289
rect 388482 -13345 388538 -13289
rect 388606 -13345 388662 -13289
rect 388730 -13345 388786 -13289
rect 388854 -13345 388910 -13289
rect 388978 -13345 389034 -13289
rect 389102 -13345 389158 -13289
rect 389226 -13345 389282 -13289
rect 389350 -13345 389406 -13289
rect 389474 -13345 389530 -13289
rect 389598 -13345 389654 -13289
rect 389722 -13345 389778 -13289
rect 389846 -13345 389902 -13289
rect 389970 -13345 390026 -13289
rect 390094 -13345 390150 -13289
rect 390218 -13345 390274 -13289
rect 390342 -13345 390398 -13289
rect 390466 -13345 390522 -13289
rect 390590 -13345 390646 -13289
rect 390714 -13345 390770 -13289
rect 390838 -13345 390894 -13289
rect 390962 -13345 391018 -13289
rect 391086 -13345 391142 -13289
rect 391210 -13345 391266 -13289
rect 391334 -13345 391390 -13289
rect 391458 -13345 391514 -13289
rect 391582 -13345 391638 -13289
rect 391706 -13345 391762 -13289
rect 391830 -13345 391886 -13289
rect 391954 -13345 392010 -13289
rect 392078 -13345 392134 -13289
rect 392202 -13345 392258 -13289
rect 392326 -13345 392382 -13289
rect 392450 -13345 392506 -13289
rect 392574 -13345 392630 -13289
rect 392698 -13345 392754 -13289
rect 392822 -13345 392878 -13289
rect 392946 -13345 393002 -13289
rect 393070 -13345 393126 -13289
rect 393194 -13345 393250 -13289
rect 393318 -13345 393374 -13289
rect 393442 -13345 393498 -13289
rect 393566 -13345 393622 -13289
rect 393690 -13345 393746 -13289
rect 393814 -13345 393870 -13289
rect 393938 -13345 393994 -13289
rect 394062 -13345 394118 -13289
rect 394186 -13345 394242 -13289
rect 394310 -13345 394366 -13289
rect 394434 -13345 394490 -13289
rect 394558 -13345 394614 -13289
rect 394682 -13345 394738 -13289
rect 394806 -13345 394862 -13289
rect 394930 -13345 394986 -13289
rect 395054 -13345 395110 -13289
rect 395178 -13345 395234 -13289
rect 395302 -13345 395358 -13289
rect 395426 -13345 395482 -13289
rect 395550 -13345 395606 -13289
rect 395674 -13345 395730 -13289
rect 395798 -13345 395854 -13289
rect 395922 -13345 395978 -13289
rect 396046 -13345 396102 -13289
rect 396170 -13345 396226 -13289
rect 396294 -13345 396350 -13289
rect 396418 -13345 396474 -13289
rect 396542 -13345 396598 -13289
rect 396666 -13345 396722 -13289
rect 396790 -13345 396846 -13289
rect 396914 -13345 396970 -13289
rect 397038 -13345 397094 -13289
rect 397162 -13345 397218 -13289
rect 397286 -13345 397342 -13289
rect 397410 -13345 397466 -13289
rect 397534 -13345 397590 -13289
rect 397658 -13345 397714 -13289
rect 397782 -13345 397838 -13289
rect 397906 -13345 397962 -13289
rect 398030 -13345 398086 -13289
rect 398154 -13345 398210 -13289
rect 398278 -13345 398334 -13289
rect 398402 -13345 398458 -13289
rect 398526 -13345 398582 -13289
rect 398650 -13345 398706 -13289
rect 398774 -13345 398830 -13289
rect 398898 -13345 398954 -13289
rect 399022 -13345 399078 -13289
rect 399146 -13345 399202 -13289
rect 399270 -13345 399326 -13289
rect 399394 -13345 399450 -13289
rect 399518 -13345 399574 -13289
rect 399642 -13345 399698 -13289
rect 399766 -13345 399822 -13289
rect 399890 -13345 399946 -13289
rect 400014 -13345 400070 -13289
rect 400138 -13345 400194 -13289
rect 400262 -13345 400318 -13289
rect 400386 -13345 400442 -13289
rect 400510 -13345 400566 -13289
rect 400634 -13345 400690 -13289
rect 400758 -13345 400814 -13289
rect 400882 -13345 400938 -13289
rect 401006 -13345 401062 -13289
rect 401130 -13345 401186 -13289
rect 401254 -13345 401310 -13289
rect 387986 -13469 388042 -13413
rect 388110 -13469 388166 -13413
rect 388234 -13469 388290 -13413
rect 388358 -13469 388414 -13413
rect 388482 -13469 388538 -13413
rect 388606 -13469 388662 -13413
rect 388730 -13469 388786 -13413
rect 388854 -13469 388910 -13413
rect 388978 -13469 389034 -13413
rect 389102 -13469 389158 -13413
rect 389226 -13469 389282 -13413
rect 389350 -13469 389406 -13413
rect 389474 -13469 389530 -13413
rect 389598 -13469 389654 -13413
rect 389722 -13469 389778 -13413
rect 389846 -13469 389902 -13413
rect 389970 -13469 390026 -13413
rect 390094 -13469 390150 -13413
rect 390218 -13469 390274 -13413
rect 390342 -13469 390398 -13413
rect 390466 -13469 390522 -13413
rect 390590 -13469 390646 -13413
rect 390714 -13469 390770 -13413
rect 390838 -13469 390894 -13413
rect 390962 -13469 391018 -13413
rect 391086 -13469 391142 -13413
rect 391210 -13469 391266 -13413
rect 391334 -13469 391390 -13413
rect 391458 -13469 391514 -13413
rect 391582 -13469 391638 -13413
rect 391706 -13469 391762 -13413
rect 391830 -13469 391886 -13413
rect 391954 -13469 392010 -13413
rect 392078 -13469 392134 -13413
rect 392202 -13469 392258 -13413
rect 392326 -13469 392382 -13413
rect 392450 -13469 392506 -13413
rect 392574 -13469 392630 -13413
rect 392698 -13469 392754 -13413
rect 392822 -13469 392878 -13413
rect 392946 -13469 393002 -13413
rect 393070 -13469 393126 -13413
rect 393194 -13469 393250 -13413
rect 393318 -13469 393374 -13413
rect 393442 -13469 393498 -13413
rect 393566 -13469 393622 -13413
rect 393690 -13469 393746 -13413
rect 393814 -13469 393870 -13413
rect 393938 -13469 393994 -13413
rect 394062 -13469 394118 -13413
rect 394186 -13469 394242 -13413
rect 394310 -13469 394366 -13413
rect 394434 -13469 394490 -13413
rect 394558 -13469 394614 -13413
rect 394682 -13469 394738 -13413
rect 394806 -13469 394862 -13413
rect 394930 -13469 394986 -13413
rect 395054 -13469 395110 -13413
rect 395178 -13469 395234 -13413
rect 395302 -13469 395358 -13413
rect 395426 -13469 395482 -13413
rect 395550 -13469 395606 -13413
rect 395674 -13469 395730 -13413
rect 395798 -13469 395854 -13413
rect 395922 -13469 395978 -13413
rect 396046 -13469 396102 -13413
rect 396170 -13469 396226 -13413
rect 396294 -13469 396350 -13413
rect 396418 -13469 396474 -13413
rect 396542 -13469 396598 -13413
rect 396666 -13469 396722 -13413
rect 396790 -13469 396846 -13413
rect 396914 -13469 396970 -13413
rect 397038 -13469 397094 -13413
rect 397162 -13469 397218 -13413
rect 397286 -13469 397342 -13413
rect 397410 -13469 397466 -13413
rect 397534 -13469 397590 -13413
rect 397658 -13469 397714 -13413
rect 397782 -13469 397838 -13413
rect 397906 -13469 397962 -13413
rect 398030 -13469 398086 -13413
rect 398154 -13469 398210 -13413
rect 398278 -13469 398334 -13413
rect 398402 -13469 398458 -13413
rect 398526 -13469 398582 -13413
rect 398650 -13469 398706 -13413
rect 398774 -13469 398830 -13413
rect 398898 -13469 398954 -13413
rect 399022 -13469 399078 -13413
rect 399146 -13469 399202 -13413
rect 399270 -13469 399326 -13413
rect 399394 -13469 399450 -13413
rect 399518 -13469 399574 -13413
rect 399642 -13469 399698 -13413
rect 399766 -13469 399822 -13413
rect 399890 -13469 399946 -13413
rect 400014 -13469 400070 -13413
rect 400138 -13469 400194 -13413
rect 400262 -13469 400318 -13413
rect 400386 -13469 400442 -13413
rect 400510 -13469 400566 -13413
rect 400634 -13469 400690 -13413
rect 400758 -13469 400814 -13413
rect 400882 -13469 400938 -13413
rect 401006 -13469 401062 -13413
rect 401130 -13469 401186 -13413
rect 401254 -13469 401310 -13413
rect 387954 -13688 388010 -13632
rect 388078 -13688 388134 -13632
rect 388202 -13688 388258 -13632
rect 388326 -13688 388382 -13632
rect 388450 -13688 388506 -13632
rect 387954 -13812 388010 -13756
rect 388078 -13812 388134 -13756
rect 388202 -13812 388258 -13756
rect 388326 -13812 388382 -13756
rect 388450 -13812 388506 -13756
rect 387954 -13936 388010 -13880
rect 388078 -13936 388134 -13880
rect 388202 -13936 388258 -13880
rect 388326 -13936 388382 -13880
rect 388450 -13936 388506 -13880
rect 387954 -14060 388010 -14004
rect 388078 -14060 388134 -14004
rect 388202 -14060 388258 -14004
rect 388326 -14060 388382 -14004
rect 388450 -14060 388506 -14004
rect 387954 -14184 388010 -14128
rect 388078 -14184 388134 -14128
rect 388202 -14184 388258 -14128
rect 388326 -14184 388382 -14128
rect 388450 -14184 388506 -14128
rect 387954 -14308 388010 -14252
rect 388078 -14308 388134 -14252
rect 388202 -14308 388258 -14252
rect 388326 -14308 388382 -14252
rect 388450 -14308 388506 -14252
rect 387954 -14432 388010 -14376
rect 388078 -14432 388134 -14376
rect 388202 -14432 388258 -14376
rect 388326 -14432 388382 -14376
rect 388450 -14432 388506 -14376
rect 387954 -14556 388010 -14500
rect 388078 -14556 388134 -14500
rect 388202 -14556 388258 -14500
rect 388326 -14556 388382 -14500
rect 388450 -14556 388506 -14500
rect 387954 -14680 388010 -14624
rect 388078 -14680 388134 -14624
rect 388202 -14680 388258 -14624
rect 388326 -14680 388382 -14624
rect 388450 -14680 388506 -14624
rect 387954 -14804 388010 -14748
rect 388078 -14804 388134 -14748
rect 388202 -14804 388258 -14748
rect 388326 -14804 388382 -14748
rect 388450 -14804 388506 -14748
rect 387954 -14928 388010 -14872
rect 388078 -14928 388134 -14872
rect 388202 -14928 388258 -14872
rect 388326 -14928 388382 -14872
rect 388450 -14928 388506 -14872
rect 387954 -15052 388010 -14996
rect 388078 -15052 388134 -14996
rect 388202 -15052 388258 -14996
rect 388326 -15052 388382 -14996
rect 388450 -15052 388506 -14996
rect 387954 -15176 388010 -15120
rect 388078 -15176 388134 -15120
rect 388202 -15176 388258 -15120
rect 388326 -15176 388382 -15120
rect 388450 -15176 388506 -15120
rect 387954 -15300 388010 -15244
rect 388078 -15300 388134 -15244
rect 388202 -15300 388258 -15244
rect 388326 -15300 388382 -15244
rect 388450 -15300 388506 -15244
rect 387954 -15424 388010 -15368
rect 388078 -15424 388134 -15368
rect 388202 -15424 388258 -15368
rect 388326 -15424 388382 -15368
rect 388450 -15424 388506 -15368
rect 387954 -15548 388010 -15492
rect 388078 -15548 388134 -15492
rect 388202 -15548 388258 -15492
rect 388326 -15548 388382 -15492
rect 388450 -15548 388506 -15492
rect 387954 -15672 388010 -15616
rect 388078 -15672 388134 -15616
rect 388202 -15672 388258 -15616
rect 388326 -15672 388382 -15616
rect 388450 -15672 388506 -15616
rect 387954 -15796 388010 -15740
rect 388078 -15796 388134 -15740
rect 388202 -15796 388258 -15740
rect 388326 -15796 388382 -15740
rect 388450 -15796 388506 -15740
rect 387954 -15920 388010 -15864
rect 388078 -15920 388134 -15864
rect 388202 -15920 388258 -15864
rect 388326 -15920 388382 -15864
rect 388450 -15920 388506 -15864
rect 387954 -16044 388010 -15988
rect 388078 -16044 388134 -15988
rect 388202 -16044 388258 -15988
rect 388326 -16044 388382 -15988
rect 388450 -16044 388506 -15988
rect 387954 -16168 388010 -16112
rect 388078 -16168 388134 -16112
rect 388202 -16168 388258 -16112
rect 388326 -16168 388382 -16112
rect 388450 -16168 388506 -16112
rect 387954 -16292 388010 -16236
rect 388078 -16292 388134 -16236
rect 388202 -16292 388258 -16236
rect 388326 -16292 388382 -16236
rect 388450 -16292 388506 -16236
rect 387954 -16416 388010 -16360
rect 388078 -16416 388134 -16360
rect 388202 -16416 388258 -16360
rect 388326 -16416 388382 -16360
rect 388450 -16416 388506 -16360
rect 387954 -16540 388010 -16484
rect 388078 -16540 388134 -16484
rect 388202 -16540 388258 -16484
rect 388326 -16540 388382 -16484
rect 388450 -16540 388506 -16484
rect 387954 -16664 388010 -16608
rect 388078 -16664 388134 -16608
rect 388202 -16664 388258 -16608
rect 388326 -16664 388382 -16608
rect 388450 -16664 388506 -16608
rect 387954 -16788 388010 -16732
rect 388078 -16788 388134 -16732
rect 388202 -16788 388258 -16732
rect 388326 -16788 388382 -16732
rect 388450 -16788 388506 -16732
rect 387954 -16912 388010 -16856
rect 388078 -16912 388134 -16856
rect 388202 -16912 388258 -16856
rect 388326 -16912 388382 -16856
rect 388450 -16912 388506 -16856
rect 387954 -17036 388010 -16980
rect 388078 -17036 388134 -16980
rect 388202 -17036 388258 -16980
rect 388326 -17036 388382 -16980
rect 388450 -17036 388506 -16980
rect 387954 -17160 388010 -17104
rect 388078 -17160 388134 -17104
rect 388202 -17160 388258 -17104
rect 388326 -17160 388382 -17104
rect 388450 -17160 388506 -17104
rect 387954 -17284 388010 -17228
rect 388078 -17284 388134 -17228
rect 388202 -17284 388258 -17228
rect 388326 -17284 388382 -17228
rect 388450 -17284 388506 -17228
rect 387954 -17408 388010 -17352
rect 388078 -17408 388134 -17352
rect 388202 -17408 388258 -17352
rect 388326 -17408 388382 -17352
rect 388450 -17408 388506 -17352
rect 387954 -17532 388010 -17476
rect 388078 -17532 388134 -17476
rect 388202 -17532 388258 -17476
rect 388326 -17532 388382 -17476
rect 388450 -17532 388506 -17476
rect 387954 -17656 388010 -17600
rect 388078 -17656 388134 -17600
rect 388202 -17656 388258 -17600
rect 388326 -17656 388382 -17600
rect 388450 -17656 388506 -17600
rect 387954 -17780 388010 -17724
rect 388078 -17780 388134 -17724
rect 388202 -17780 388258 -17724
rect 388326 -17780 388382 -17724
rect 388450 -17780 388506 -17724
rect 387954 -17904 388010 -17848
rect 388078 -17904 388134 -17848
rect 388202 -17904 388258 -17848
rect 388326 -17904 388382 -17848
rect 388450 -17904 388506 -17848
rect 387954 -18028 388010 -17972
rect 388078 -18028 388134 -17972
rect 388202 -18028 388258 -17972
rect 388326 -18028 388382 -17972
rect 388450 -18028 388506 -17972
rect 387954 -18152 388010 -18096
rect 388078 -18152 388134 -18096
rect 388202 -18152 388258 -18096
rect 388326 -18152 388382 -18096
rect 388450 -18152 388506 -18096
rect 387954 -18276 388010 -18220
rect 388078 -18276 388134 -18220
rect 388202 -18276 388258 -18220
rect 388326 -18276 388382 -18220
rect 388450 -18276 388506 -18220
rect 387954 -18400 388010 -18344
rect 388078 -18400 388134 -18344
rect 388202 -18400 388258 -18344
rect 388326 -18400 388382 -18344
rect 388450 -18400 388506 -18344
rect 387954 -18524 388010 -18468
rect 388078 -18524 388134 -18468
rect 388202 -18524 388258 -18468
rect 388326 -18524 388382 -18468
rect 388450 -18524 388506 -18468
rect 387954 -18648 388010 -18592
rect 388078 -18648 388134 -18592
rect 388202 -18648 388258 -18592
rect 388326 -18648 388382 -18592
rect 388450 -18648 388506 -18592
rect 387954 -18772 388010 -18716
rect 388078 -18772 388134 -18716
rect 388202 -18772 388258 -18716
rect 388326 -18772 388382 -18716
rect 388450 -18772 388506 -18716
rect 387954 -18896 388010 -18840
rect 388078 -18896 388134 -18840
rect 388202 -18896 388258 -18840
rect 388326 -18896 388382 -18840
rect 388450 -18896 388506 -18840
rect 387954 -19020 388010 -18964
rect 388078 -19020 388134 -18964
rect 388202 -19020 388258 -18964
rect 388326 -19020 388382 -18964
rect 388450 -19020 388506 -18964
rect 387954 -19144 388010 -19088
rect 388078 -19144 388134 -19088
rect 388202 -19144 388258 -19088
rect 388326 -19144 388382 -19088
rect 388450 -19144 388506 -19088
rect 387954 -19268 388010 -19212
rect 388078 -19268 388134 -19212
rect 388202 -19268 388258 -19212
rect 388326 -19268 388382 -19212
rect 388450 -19268 388506 -19212
rect 387954 -19392 388010 -19336
rect 388078 -19392 388134 -19336
rect 388202 -19392 388258 -19336
rect 388326 -19392 388382 -19336
rect 388450 -19392 388506 -19336
rect 387954 -19516 388010 -19460
rect 388078 -19516 388134 -19460
rect 388202 -19516 388258 -19460
rect 388326 -19516 388382 -19460
rect 388450 -19516 388506 -19460
rect 387954 -19640 388010 -19584
rect 388078 -19640 388134 -19584
rect 388202 -19640 388258 -19584
rect 388326 -19640 388382 -19584
rect 388450 -19640 388506 -19584
rect 387954 -19764 388010 -19708
rect 388078 -19764 388134 -19708
rect 388202 -19764 388258 -19708
rect 388326 -19764 388382 -19708
rect 388450 -19764 388506 -19708
rect 387954 -19888 388010 -19832
rect 388078 -19888 388134 -19832
rect 388202 -19888 388258 -19832
rect 388326 -19888 388382 -19832
rect 388450 -19888 388506 -19832
rect 387954 -20012 388010 -19956
rect 388078 -20012 388134 -19956
rect 388202 -20012 388258 -19956
rect 388326 -20012 388382 -19956
rect 388450 -20012 388506 -19956
rect 387954 -20136 388010 -20080
rect 388078 -20136 388134 -20080
rect 388202 -20136 388258 -20080
rect 388326 -20136 388382 -20080
rect 388450 -20136 388506 -20080
rect 387954 -20260 388010 -20204
rect 388078 -20260 388134 -20204
rect 388202 -20260 388258 -20204
rect 388326 -20260 388382 -20204
rect 388450 -20260 388506 -20204
rect 387954 -20384 388010 -20328
rect 388078 -20384 388134 -20328
rect 388202 -20384 388258 -20328
rect 388326 -20384 388382 -20328
rect 388450 -20384 388506 -20328
rect 387954 -20508 388010 -20452
rect 388078 -20508 388134 -20452
rect 388202 -20508 388258 -20452
rect 388326 -20508 388382 -20452
rect 388450 -20508 388506 -20452
rect 387954 -20632 388010 -20576
rect 388078 -20632 388134 -20576
rect 388202 -20632 388258 -20576
rect 388326 -20632 388382 -20576
rect 388450 -20632 388506 -20576
rect 387954 -20756 388010 -20700
rect 388078 -20756 388134 -20700
rect 388202 -20756 388258 -20700
rect 388326 -20756 388382 -20700
rect 388450 -20756 388506 -20700
rect 387954 -20880 388010 -20824
rect 388078 -20880 388134 -20824
rect 388202 -20880 388258 -20824
rect 388326 -20880 388382 -20824
rect 388450 -20880 388506 -20824
rect 387954 -21004 388010 -20948
rect 388078 -21004 388134 -20948
rect 388202 -21004 388258 -20948
rect 388326 -21004 388382 -20948
rect 388450 -21004 388506 -20948
rect 387954 -21128 388010 -21072
rect 388078 -21128 388134 -21072
rect 388202 -21128 388258 -21072
rect 388326 -21128 388382 -21072
rect 388450 -21128 388506 -21072
rect 387954 -21252 388010 -21196
rect 388078 -21252 388134 -21196
rect 388202 -21252 388258 -21196
rect 388326 -21252 388382 -21196
rect 388450 -21252 388506 -21196
rect 387954 -21376 388010 -21320
rect 388078 -21376 388134 -21320
rect 388202 -21376 388258 -21320
rect 388326 -21376 388382 -21320
rect 388450 -21376 388506 -21320
rect 387954 -21500 388010 -21444
rect 388078 -21500 388134 -21444
rect 388202 -21500 388258 -21444
rect 388326 -21500 388382 -21444
rect 388450 -21500 388506 -21444
rect 387954 -21624 388010 -21568
rect 388078 -21624 388134 -21568
rect 388202 -21624 388258 -21568
rect 388326 -21624 388382 -21568
rect 388450 -21624 388506 -21568
rect 387954 -21748 388010 -21692
rect 388078 -21748 388134 -21692
rect 388202 -21748 388258 -21692
rect 388326 -21748 388382 -21692
rect 388450 -21748 388506 -21692
rect 387954 -21872 388010 -21816
rect 388078 -21872 388134 -21816
rect 388202 -21872 388258 -21816
rect 388326 -21872 388382 -21816
rect 388450 -21872 388506 -21816
rect 387954 -21996 388010 -21940
rect 388078 -21996 388134 -21940
rect 388202 -21996 388258 -21940
rect 388326 -21996 388382 -21940
rect 388450 -21996 388506 -21940
rect 387954 -22120 388010 -22064
rect 388078 -22120 388134 -22064
rect 388202 -22120 388258 -22064
rect 388326 -22120 388382 -22064
rect 388450 -22120 388506 -22064
rect 387954 -22244 388010 -22188
rect 388078 -22244 388134 -22188
rect 388202 -22244 388258 -22188
rect 388326 -22244 388382 -22188
rect 388450 -22244 388506 -22188
rect 387954 -22368 388010 -22312
rect 388078 -22368 388134 -22312
rect 388202 -22368 388258 -22312
rect 388326 -22368 388382 -22312
rect 388450 -22368 388506 -22312
rect 387954 -22492 388010 -22436
rect 388078 -22492 388134 -22436
rect 388202 -22492 388258 -22436
rect 388326 -22492 388382 -22436
rect 388450 -22492 388506 -22436
rect 387954 -22616 388010 -22560
rect 388078 -22616 388134 -22560
rect 388202 -22616 388258 -22560
rect 388326 -22616 388382 -22560
rect 388450 -22616 388506 -22560
rect 387954 -22740 388010 -22684
rect 388078 -22740 388134 -22684
rect 388202 -22740 388258 -22684
rect 388326 -22740 388382 -22684
rect 388450 -22740 388506 -22684
rect 387954 -22864 388010 -22808
rect 388078 -22864 388134 -22808
rect 388202 -22864 388258 -22808
rect 388326 -22864 388382 -22808
rect 388450 -22864 388506 -22808
rect 387954 -22988 388010 -22932
rect 388078 -22988 388134 -22932
rect 388202 -22988 388258 -22932
rect 388326 -22988 388382 -22932
rect 388450 -22988 388506 -22932
rect 387954 -23112 388010 -23056
rect 388078 -23112 388134 -23056
rect 388202 -23112 388258 -23056
rect 388326 -23112 388382 -23056
rect 388450 -23112 388506 -23056
rect 387954 -23236 388010 -23180
rect 388078 -23236 388134 -23180
rect 388202 -23236 388258 -23180
rect 388326 -23236 388382 -23180
rect 388450 -23236 388506 -23180
rect 387954 -23360 388010 -23304
rect 388078 -23360 388134 -23304
rect 388202 -23360 388258 -23304
rect 388326 -23360 388382 -23304
rect 388450 -23360 388506 -23304
rect 387954 -23484 388010 -23428
rect 388078 -23484 388134 -23428
rect 388202 -23484 388258 -23428
rect 388326 -23484 388382 -23428
rect 388450 -23484 388506 -23428
rect 387954 -23608 388010 -23552
rect 388078 -23608 388134 -23552
rect 388202 -23608 388258 -23552
rect 388326 -23608 388382 -23552
rect 388450 -23608 388506 -23552
rect 387954 -23732 388010 -23676
rect 388078 -23732 388134 -23676
rect 388202 -23732 388258 -23676
rect 388326 -23732 388382 -23676
rect 388450 -23732 388506 -23676
rect 387954 -23856 388010 -23800
rect 388078 -23856 388134 -23800
rect 388202 -23856 388258 -23800
rect 388326 -23856 388382 -23800
rect 388450 -23856 388506 -23800
rect 387954 -23980 388010 -23924
rect 388078 -23980 388134 -23924
rect 388202 -23980 388258 -23924
rect 388326 -23980 388382 -23924
rect 388450 -23980 388506 -23924
rect 387954 -24104 388010 -24048
rect 388078 -24104 388134 -24048
rect 388202 -24104 388258 -24048
rect 388326 -24104 388382 -24048
rect 388450 -24104 388506 -24048
rect 387954 -24228 388010 -24172
rect 388078 -24228 388134 -24172
rect 388202 -24228 388258 -24172
rect 388326 -24228 388382 -24172
rect 388450 -24228 388506 -24172
rect 387954 -24352 388010 -24296
rect 388078 -24352 388134 -24296
rect 388202 -24352 388258 -24296
rect 388326 -24352 388382 -24296
rect 388450 -24352 388506 -24296
rect 387954 -24476 388010 -24420
rect 388078 -24476 388134 -24420
rect 388202 -24476 388258 -24420
rect 388326 -24476 388382 -24420
rect 388450 -24476 388506 -24420
rect 387954 -24600 388010 -24544
rect 388078 -24600 388134 -24544
rect 388202 -24600 388258 -24544
rect 388326 -24600 388382 -24544
rect 388450 -24600 388506 -24544
rect 387954 -24724 388010 -24668
rect 388078 -24724 388134 -24668
rect 388202 -24724 388258 -24668
rect 388326 -24724 388382 -24668
rect 388450 -24724 388506 -24668
rect 387954 -24848 388010 -24792
rect 388078 -24848 388134 -24792
rect 388202 -24848 388258 -24792
rect 388326 -24848 388382 -24792
rect 388450 -24848 388506 -24792
rect 387954 -24972 388010 -24916
rect 388078 -24972 388134 -24916
rect 388202 -24972 388258 -24916
rect 388326 -24972 388382 -24916
rect 388450 -24972 388506 -24916
rect 387954 -25096 388010 -25040
rect 388078 -25096 388134 -25040
rect 388202 -25096 388258 -25040
rect 388326 -25096 388382 -25040
rect 388450 -25096 388506 -25040
rect 387954 -25220 388010 -25164
rect 388078 -25220 388134 -25164
rect 388202 -25220 388258 -25164
rect 388326 -25220 388382 -25164
rect 388450 -25220 388506 -25164
rect 387954 -25344 388010 -25288
rect 388078 -25344 388134 -25288
rect 388202 -25344 388258 -25288
rect 388326 -25344 388382 -25288
rect 388450 -25344 388506 -25288
rect 387954 -25468 388010 -25412
rect 388078 -25468 388134 -25412
rect 388202 -25468 388258 -25412
rect 388326 -25468 388382 -25412
rect 388450 -25468 388506 -25412
rect 388981 -13736 389037 -13680
rect 389123 -13736 389179 -13680
rect 388981 -13878 389037 -13822
rect 389123 -13878 389179 -13822
rect 388981 -14020 389037 -13964
rect 389123 -14020 389179 -13964
rect 388981 -14162 389037 -14106
rect 389123 -14162 389179 -14106
rect 388981 -14304 389037 -14248
rect 389123 -14304 389179 -14248
rect 388981 -14446 389037 -14390
rect 389123 -14446 389179 -14390
rect 388981 -14588 389037 -14532
rect 389123 -14588 389179 -14532
rect 388981 -14730 389037 -14674
rect 389123 -14730 389179 -14674
rect 388981 -14872 389037 -14816
rect 389123 -14872 389179 -14816
rect 388981 -15014 389037 -14958
rect 389123 -15014 389179 -14958
rect 388981 -15156 389037 -15100
rect 389123 -15156 389179 -15100
rect 388981 -15298 389037 -15242
rect 389123 -15298 389179 -15242
rect 388981 -15440 389037 -15384
rect 389123 -15440 389179 -15384
rect 388981 -15582 389037 -15526
rect 389123 -15582 389179 -15526
rect 388981 -15724 389037 -15668
rect 389123 -15724 389179 -15668
rect 388981 -15866 389037 -15810
rect 389123 -15866 389179 -15810
rect 388981 -16008 389037 -15952
rect 389123 -16008 389179 -15952
rect 388981 -16150 389037 -16094
rect 389123 -16150 389179 -16094
rect 388981 -16292 389037 -16236
rect 389123 -16292 389179 -16236
rect 388981 -16434 389037 -16378
rect 389123 -16434 389179 -16378
rect 388981 -16576 389037 -16520
rect 389123 -16576 389179 -16520
rect 388981 -16718 389037 -16662
rect 389123 -16718 389179 -16662
rect 388981 -16860 389037 -16804
rect 389123 -16860 389179 -16804
rect 388981 -17002 389037 -16946
rect 389123 -17002 389179 -16946
rect 388981 -17144 389037 -17088
rect 389123 -17144 389179 -17088
rect 388981 -17286 389037 -17230
rect 389123 -17286 389179 -17230
rect 388981 -17428 389037 -17372
rect 389123 -17428 389179 -17372
rect 388981 -17570 389037 -17514
rect 389123 -17570 389179 -17514
rect 388981 -17712 389037 -17656
rect 389123 -17712 389179 -17656
rect 388981 -17854 389037 -17798
rect 389123 -17854 389179 -17798
rect 388981 -17996 389037 -17940
rect 389123 -17996 389179 -17940
rect 388981 -18138 389037 -18082
rect 389123 -18138 389179 -18082
rect 388981 -18280 389037 -18224
rect 389123 -18280 389179 -18224
rect 388981 -18422 389037 -18366
rect 389123 -18422 389179 -18366
rect 388981 -18564 389037 -18508
rect 389123 -18564 389179 -18508
rect 388981 -18706 389037 -18650
rect 389123 -18706 389179 -18650
rect 388981 -18848 389037 -18792
rect 389123 -18848 389179 -18792
rect 388981 -18990 389037 -18934
rect 389123 -18990 389179 -18934
rect 388981 -19132 389037 -19076
rect 389123 -19132 389179 -19076
rect 388981 -19274 389037 -19218
rect 389123 -19274 389179 -19218
rect 388981 -19416 389037 -19360
rect 389123 -19416 389179 -19360
rect 388981 -19558 389037 -19502
rect 389123 -19558 389179 -19502
rect 388981 -19700 389037 -19644
rect 389123 -19700 389179 -19644
rect 388981 -19842 389037 -19786
rect 389123 -19842 389179 -19786
rect 388981 -19984 389037 -19928
rect 389123 -19984 389179 -19928
rect 388981 -20126 389037 -20070
rect 389123 -20126 389179 -20070
rect 388981 -20268 389037 -20212
rect 389123 -20268 389179 -20212
rect 388981 -20410 389037 -20354
rect 389123 -20410 389179 -20354
rect 388981 -20552 389037 -20496
rect 389123 -20552 389179 -20496
rect 388981 -20694 389037 -20638
rect 389123 -20694 389179 -20638
rect 388981 -20836 389037 -20780
rect 389123 -20836 389179 -20780
rect 388981 -20978 389037 -20922
rect 389123 -20978 389179 -20922
rect 388981 -21120 389037 -21064
rect 389123 -21120 389179 -21064
rect 388981 -21262 389037 -21206
rect 389123 -21262 389179 -21206
rect 388981 -21404 389037 -21348
rect 389123 -21404 389179 -21348
rect 388981 -21546 389037 -21490
rect 389123 -21546 389179 -21490
rect 388981 -21688 389037 -21632
rect 389123 -21688 389179 -21632
rect 388981 -21830 389037 -21774
rect 389123 -21830 389179 -21774
rect 388981 -21972 389037 -21916
rect 389123 -21972 389179 -21916
rect 388981 -22114 389037 -22058
rect 389123 -22114 389179 -22058
rect 388981 -22256 389037 -22200
rect 389123 -22256 389179 -22200
rect 388981 -22398 389037 -22342
rect 389123 -22398 389179 -22342
rect 388981 -22540 389037 -22484
rect 389123 -22540 389179 -22484
rect 388981 -22682 389037 -22626
rect 389123 -22682 389179 -22626
rect 388981 -22824 389037 -22768
rect 389123 -22824 389179 -22768
rect 388981 -22966 389037 -22910
rect 389123 -22966 389179 -22910
rect 388981 -23108 389037 -23052
rect 389123 -23108 389179 -23052
rect 388981 -23250 389037 -23194
rect 389123 -23250 389179 -23194
rect 388981 -23392 389037 -23336
rect 389123 -23392 389179 -23336
rect 388981 -23534 389037 -23478
rect 389123 -23534 389179 -23478
rect 388981 -23676 389037 -23620
rect 389123 -23676 389179 -23620
rect 388981 -23818 389037 -23762
rect 389123 -23818 389179 -23762
rect 388981 -23960 389037 -23904
rect 389123 -23960 389179 -23904
rect 388981 -24102 389037 -24046
rect 389123 -24102 389179 -24046
rect 388981 -24244 389037 -24188
rect 389123 -24244 389179 -24188
rect 388981 -24386 389037 -24330
rect 389123 -24386 389179 -24330
rect 388981 -24528 389037 -24472
rect 389123 -24528 389179 -24472
rect 388981 -24670 389037 -24614
rect 389123 -24670 389179 -24614
rect 388981 -24812 389037 -24756
rect 389123 -24812 389179 -24756
rect 388981 -24954 389037 -24898
rect 389123 -24954 389179 -24898
rect 388981 -25096 389037 -25040
rect 389123 -25096 389179 -25040
rect 388981 -25238 389037 -25182
rect 389123 -25238 389179 -25182
rect 388981 -25380 389037 -25324
rect 389123 -25380 389179 -25324
rect 388981 -25522 389037 -25466
rect 389123 -25522 389179 -25466
rect 389382 -13736 389438 -13680
rect 389524 -13736 389580 -13680
rect 389382 -13878 389438 -13822
rect 389524 -13878 389580 -13822
rect 389382 -14020 389438 -13964
rect 389524 -14020 389580 -13964
rect 389382 -14162 389438 -14106
rect 389524 -14162 389580 -14106
rect 389382 -14304 389438 -14248
rect 389524 -14304 389580 -14248
rect 389382 -14446 389438 -14390
rect 389524 -14446 389580 -14390
rect 389382 -14588 389438 -14532
rect 389524 -14588 389580 -14532
rect 389382 -14730 389438 -14674
rect 389524 -14730 389580 -14674
rect 389382 -14872 389438 -14816
rect 389524 -14872 389580 -14816
rect 389382 -15014 389438 -14958
rect 389524 -15014 389580 -14958
rect 389382 -15156 389438 -15100
rect 389524 -15156 389580 -15100
rect 389382 -15298 389438 -15242
rect 389524 -15298 389580 -15242
rect 389382 -15440 389438 -15384
rect 389524 -15440 389580 -15384
rect 389382 -15582 389438 -15526
rect 389524 -15582 389580 -15526
rect 389382 -15724 389438 -15668
rect 389524 -15724 389580 -15668
rect 389382 -15866 389438 -15810
rect 389524 -15866 389580 -15810
rect 389382 -16008 389438 -15952
rect 389524 -16008 389580 -15952
rect 389382 -16150 389438 -16094
rect 389524 -16150 389580 -16094
rect 389382 -16292 389438 -16236
rect 389524 -16292 389580 -16236
rect 389382 -16434 389438 -16378
rect 389524 -16434 389580 -16378
rect 389382 -16576 389438 -16520
rect 389524 -16576 389580 -16520
rect 389382 -16718 389438 -16662
rect 389524 -16718 389580 -16662
rect 389382 -16860 389438 -16804
rect 389524 -16860 389580 -16804
rect 389382 -17002 389438 -16946
rect 389524 -17002 389580 -16946
rect 389382 -17144 389438 -17088
rect 389524 -17144 389580 -17088
rect 389382 -17286 389438 -17230
rect 389524 -17286 389580 -17230
rect 389382 -17428 389438 -17372
rect 389524 -17428 389580 -17372
rect 389382 -17570 389438 -17514
rect 389524 -17570 389580 -17514
rect 389382 -17712 389438 -17656
rect 389524 -17712 389580 -17656
rect 389382 -17854 389438 -17798
rect 389524 -17854 389580 -17798
rect 389382 -17996 389438 -17940
rect 389524 -17996 389580 -17940
rect 389382 -18138 389438 -18082
rect 389524 -18138 389580 -18082
rect 389382 -18280 389438 -18224
rect 389524 -18280 389580 -18224
rect 389382 -18422 389438 -18366
rect 389524 -18422 389580 -18366
rect 389382 -18564 389438 -18508
rect 389524 -18564 389580 -18508
rect 389382 -18706 389438 -18650
rect 389524 -18706 389580 -18650
rect 389382 -18848 389438 -18792
rect 389524 -18848 389580 -18792
rect 389382 -18990 389438 -18934
rect 389524 -18990 389580 -18934
rect 389382 -19132 389438 -19076
rect 389524 -19132 389580 -19076
rect 389382 -19274 389438 -19218
rect 389524 -19274 389580 -19218
rect 389382 -19416 389438 -19360
rect 389524 -19416 389580 -19360
rect 389382 -19558 389438 -19502
rect 389524 -19558 389580 -19502
rect 389382 -19700 389438 -19644
rect 389524 -19700 389580 -19644
rect 389382 -19842 389438 -19786
rect 389524 -19842 389580 -19786
rect 389382 -19984 389438 -19928
rect 389524 -19984 389580 -19928
rect 389382 -20126 389438 -20070
rect 389524 -20126 389580 -20070
rect 389382 -20268 389438 -20212
rect 389524 -20268 389580 -20212
rect 389382 -20410 389438 -20354
rect 389524 -20410 389580 -20354
rect 389382 -20552 389438 -20496
rect 389524 -20552 389580 -20496
rect 389382 -20694 389438 -20638
rect 389524 -20694 389580 -20638
rect 389382 -20836 389438 -20780
rect 389524 -20836 389580 -20780
rect 389382 -20978 389438 -20922
rect 389524 -20978 389580 -20922
rect 389382 -21120 389438 -21064
rect 389524 -21120 389580 -21064
rect 389382 -21262 389438 -21206
rect 389524 -21262 389580 -21206
rect 389382 -21404 389438 -21348
rect 389524 -21404 389580 -21348
rect 389382 -21546 389438 -21490
rect 389524 -21546 389580 -21490
rect 389382 -21688 389438 -21632
rect 389524 -21688 389580 -21632
rect 389382 -21830 389438 -21774
rect 389524 -21830 389580 -21774
rect 389382 -21972 389438 -21916
rect 389524 -21972 389580 -21916
rect 389382 -22114 389438 -22058
rect 389524 -22114 389580 -22058
rect 389382 -22256 389438 -22200
rect 389524 -22256 389580 -22200
rect 389382 -22398 389438 -22342
rect 389524 -22398 389580 -22342
rect 389382 -22540 389438 -22484
rect 389524 -22540 389580 -22484
rect 389382 -22682 389438 -22626
rect 389524 -22682 389580 -22626
rect 389382 -22824 389438 -22768
rect 389524 -22824 389580 -22768
rect 389382 -22966 389438 -22910
rect 389524 -22966 389580 -22910
rect 389382 -23108 389438 -23052
rect 389524 -23108 389580 -23052
rect 389382 -23250 389438 -23194
rect 389524 -23250 389580 -23194
rect 389382 -23392 389438 -23336
rect 389524 -23392 389580 -23336
rect 389382 -23534 389438 -23478
rect 389524 -23534 389580 -23478
rect 389382 -23676 389438 -23620
rect 389524 -23676 389580 -23620
rect 389382 -23818 389438 -23762
rect 389524 -23818 389580 -23762
rect 389382 -23960 389438 -23904
rect 389524 -23960 389580 -23904
rect 389382 -24102 389438 -24046
rect 389524 -24102 389580 -24046
rect 389382 -24244 389438 -24188
rect 389524 -24244 389580 -24188
rect 389382 -24386 389438 -24330
rect 389524 -24386 389580 -24330
rect 389382 -24528 389438 -24472
rect 389524 -24528 389580 -24472
rect 389382 -24670 389438 -24614
rect 389524 -24670 389580 -24614
rect 389382 -24812 389438 -24756
rect 389524 -24812 389580 -24756
rect 389382 -24954 389438 -24898
rect 389524 -24954 389580 -24898
rect 389382 -25096 389438 -25040
rect 389524 -25096 389580 -25040
rect 389382 -25238 389438 -25182
rect 389524 -25238 389580 -25182
rect 389382 -25380 389438 -25324
rect 389524 -25380 389580 -25324
rect 389382 -25522 389438 -25466
rect 389524 -25522 389580 -25466
rect 389782 -13736 389838 -13680
rect 389924 -13736 389980 -13680
rect 389782 -13878 389838 -13822
rect 389924 -13878 389980 -13822
rect 389782 -14020 389838 -13964
rect 389924 -14020 389980 -13964
rect 389782 -14162 389838 -14106
rect 389924 -14162 389980 -14106
rect 389782 -14304 389838 -14248
rect 389924 -14304 389980 -14248
rect 389782 -14446 389838 -14390
rect 389924 -14446 389980 -14390
rect 389782 -14588 389838 -14532
rect 389924 -14588 389980 -14532
rect 389782 -14730 389838 -14674
rect 389924 -14730 389980 -14674
rect 389782 -14872 389838 -14816
rect 389924 -14872 389980 -14816
rect 389782 -15014 389838 -14958
rect 389924 -15014 389980 -14958
rect 389782 -15156 389838 -15100
rect 389924 -15156 389980 -15100
rect 389782 -15298 389838 -15242
rect 389924 -15298 389980 -15242
rect 389782 -15440 389838 -15384
rect 389924 -15440 389980 -15384
rect 389782 -15582 389838 -15526
rect 389924 -15582 389980 -15526
rect 389782 -15724 389838 -15668
rect 389924 -15724 389980 -15668
rect 389782 -15866 389838 -15810
rect 389924 -15866 389980 -15810
rect 389782 -16008 389838 -15952
rect 389924 -16008 389980 -15952
rect 389782 -16150 389838 -16094
rect 389924 -16150 389980 -16094
rect 389782 -16292 389838 -16236
rect 389924 -16292 389980 -16236
rect 389782 -16434 389838 -16378
rect 389924 -16434 389980 -16378
rect 389782 -16576 389838 -16520
rect 389924 -16576 389980 -16520
rect 389782 -16718 389838 -16662
rect 389924 -16718 389980 -16662
rect 389782 -16860 389838 -16804
rect 389924 -16860 389980 -16804
rect 389782 -17002 389838 -16946
rect 389924 -17002 389980 -16946
rect 389782 -17144 389838 -17088
rect 389924 -17144 389980 -17088
rect 389782 -17286 389838 -17230
rect 389924 -17286 389980 -17230
rect 389782 -17428 389838 -17372
rect 389924 -17428 389980 -17372
rect 389782 -17570 389838 -17514
rect 389924 -17570 389980 -17514
rect 389782 -17712 389838 -17656
rect 389924 -17712 389980 -17656
rect 389782 -17854 389838 -17798
rect 389924 -17854 389980 -17798
rect 389782 -17996 389838 -17940
rect 389924 -17996 389980 -17940
rect 389782 -18138 389838 -18082
rect 389924 -18138 389980 -18082
rect 389782 -18280 389838 -18224
rect 389924 -18280 389980 -18224
rect 389782 -18422 389838 -18366
rect 389924 -18422 389980 -18366
rect 389782 -18564 389838 -18508
rect 389924 -18564 389980 -18508
rect 389782 -18706 389838 -18650
rect 389924 -18706 389980 -18650
rect 389782 -18848 389838 -18792
rect 389924 -18848 389980 -18792
rect 389782 -18990 389838 -18934
rect 389924 -18990 389980 -18934
rect 389782 -19132 389838 -19076
rect 389924 -19132 389980 -19076
rect 389782 -19274 389838 -19218
rect 389924 -19274 389980 -19218
rect 389782 -19416 389838 -19360
rect 389924 -19416 389980 -19360
rect 389782 -19558 389838 -19502
rect 389924 -19558 389980 -19502
rect 389782 -19700 389838 -19644
rect 389924 -19700 389980 -19644
rect 389782 -19842 389838 -19786
rect 389924 -19842 389980 -19786
rect 389782 -19984 389838 -19928
rect 389924 -19984 389980 -19928
rect 389782 -20126 389838 -20070
rect 389924 -20126 389980 -20070
rect 389782 -20268 389838 -20212
rect 389924 -20268 389980 -20212
rect 389782 -20410 389838 -20354
rect 389924 -20410 389980 -20354
rect 389782 -20552 389838 -20496
rect 389924 -20552 389980 -20496
rect 389782 -20694 389838 -20638
rect 389924 -20694 389980 -20638
rect 389782 -20836 389838 -20780
rect 389924 -20836 389980 -20780
rect 389782 -20978 389838 -20922
rect 389924 -20978 389980 -20922
rect 389782 -21120 389838 -21064
rect 389924 -21120 389980 -21064
rect 389782 -21262 389838 -21206
rect 389924 -21262 389980 -21206
rect 389782 -21404 389838 -21348
rect 389924 -21404 389980 -21348
rect 389782 -21546 389838 -21490
rect 389924 -21546 389980 -21490
rect 389782 -21688 389838 -21632
rect 389924 -21688 389980 -21632
rect 389782 -21830 389838 -21774
rect 389924 -21830 389980 -21774
rect 389782 -21972 389838 -21916
rect 389924 -21972 389980 -21916
rect 389782 -22114 389838 -22058
rect 389924 -22114 389980 -22058
rect 389782 -22256 389838 -22200
rect 389924 -22256 389980 -22200
rect 389782 -22398 389838 -22342
rect 389924 -22398 389980 -22342
rect 389782 -22540 389838 -22484
rect 389924 -22540 389980 -22484
rect 389782 -22682 389838 -22626
rect 389924 -22682 389980 -22626
rect 389782 -22824 389838 -22768
rect 389924 -22824 389980 -22768
rect 389782 -22966 389838 -22910
rect 389924 -22966 389980 -22910
rect 389782 -23108 389838 -23052
rect 389924 -23108 389980 -23052
rect 389782 -23250 389838 -23194
rect 389924 -23250 389980 -23194
rect 389782 -23392 389838 -23336
rect 389924 -23392 389980 -23336
rect 389782 -23534 389838 -23478
rect 389924 -23534 389980 -23478
rect 389782 -23676 389838 -23620
rect 389924 -23676 389980 -23620
rect 389782 -23818 389838 -23762
rect 389924 -23818 389980 -23762
rect 389782 -23960 389838 -23904
rect 389924 -23960 389980 -23904
rect 389782 -24102 389838 -24046
rect 389924 -24102 389980 -24046
rect 389782 -24244 389838 -24188
rect 389924 -24244 389980 -24188
rect 389782 -24386 389838 -24330
rect 389924 -24386 389980 -24330
rect 389782 -24528 389838 -24472
rect 389924 -24528 389980 -24472
rect 389782 -24670 389838 -24614
rect 389924 -24670 389980 -24614
rect 389782 -24812 389838 -24756
rect 389924 -24812 389980 -24756
rect 389782 -24954 389838 -24898
rect 389924 -24954 389980 -24898
rect 389782 -25096 389838 -25040
rect 389924 -25096 389980 -25040
rect 389782 -25238 389838 -25182
rect 389924 -25238 389980 -25182
rect 389782 -25380 389838 -25324
rect 389924 -25380 389980 -25324
rect 389782 -25522 389838 -25466
rect 389924 -25522 389980 -25466
rect 390179 -13736 390235 -13680
rect 390321 -13736 390377 -13680
rect 390179 -13878 390235 -13822
rect 390321 -13878 390377 -13822
rect 390179 -14020 390235 -13964
rect 390321 -14020 390377 -13964
rect 390179 -14162 390235 -14106
rect 390321 -14162 390377 -14106
rect 390179 -14304 390235 -14248
rect 390321 -14304 390377 -14248
rect 390179 -14446 390235 -14390
rect 390321 -14446 390377 -14390
rect 390179 -14588 390235 -14532
rect 390321 -14588 390377 -14532
rect 390179 -14730 390235 -14674
rect 390321 -14730 390377 -14674
rect 390179 -14872 390235 -14816
rect 390321 -14872 390377 -14816
rect 390179 -15014 390235 -14958
rect 390321 -15014 390377 -14958
rect 390179 -15156 390235 -15100
rect 390321 -15156 390377 -15100
rect 390179 -15298 390235 -15242
rect 390321 -15298 390377 -15242
rect 390179 -15440 390235 -15384
rect 390321 -15440 390377 -15384
rect 390179 -15582 390235 -15526
rect 390321 -15582 390377 -15526
rect 390179 -15724 390235 -15668
rect 390321 -15724 390377 -15668
rect 390179 -15866 390235 -15810
rect 390321 -15866 390377 -15810
rect 390179 -16008 390235 -15952
rect 390321 -16008 390377 -15952
rect 390179 -16150 390235 -16094
rect 390321 -16150 390377 -16094
rect 390179 -16292 390235 -16236
rect 390321 -16292 390377 -16236
rect 390179 -16434 390235 -16378
rect 390321 -16434 390377 -16378
rect 390179 -16576 390235 -16520
rect 390321 -16576 390377 -16520
rect 390179 -16718 390235 -16662
rect 390321 -16718 390377 -16662
rect 390179 -16860 390235 -16804
rect 390321 -16860 390377 -16804
rect 390179 -17002 390235 -16946
rect 390321 -17002 390377 -16946
rect 390179 -17144 390235 -17088
rect 390321 -17144 390377 -17088
rect 390179 -17286 390235 -17230
rect 390321 -17286 390377 -17230
rect 390179 -17428 390235 -17372
rect 390321 -17428 390377 -17372
rect 390179 -17570 390235 -17514
rect 390321 -17570 390377 -17514
rect 390179 -17712 390235 -17656
rect 390321 -17712 390377 -17656
rect 390179 -17854 390235 -17798
rect 390321 -17854 390377 -17798
rect 390179 -17996 390235 -17940
rect 390321 -17996 390377 -17940
rect 390179 -18138 390235 -18082
rect 390321 -18138 390377 -18082
rect 390179 -18280 390235 -18224
rect 390321 -18280 390377 -18224
rect 390179 -18422 390235 -18366
rect 390321 -18422 390377 -18366
rect 390179 -18564 390235 -18508
rect 390321 -18564 390377 -18508
rect 390179 -18706 390235 -18650
rect 390321 -18706 390377 -18650
rect 390179 -18848 390235 -18792
rect 390321 -18848 390377 -18792
rect 390179 -18990 390235 -18934
rect 390321 -18990 390377 -18934
rect 390179 -19132 390235 -19076
rect 390321 -19132 390377 -19076
rect 390179 -19274 390235 -19218
rect 390321 -19274 390377 -19218
rect 390179 -19416 390235 -19360
rect 390321 -19416 390377 -19360
rect 390179 -19558 390235 -19502
rect 390321 -19558 390377 -19502
rect 390179 -19700 390235 -19644
rect 390321 -19700 390377 -19644
rect 390179 -19842 390235 -19786
rect 390321 -19842 390377 -19786
rect 390179 -19984 390235 -19928
rect 390321 -19984 390377 -19928
rect 390179 -20126 390235 -20070
rect 390321 -20126 390377 -20070
rect 390179 -20268 390235 -20212
rect 390321 -20268 390377 -20212
rect 390179 -20410 390235 -20354
rect 390321 -20410 390377 -20354
rect 390179 -20552 390235 -20496
rect 390321 -20552 390377 -20496
rect 390179 -20694 390235 -20638
rect 390321 -20694 390377 -20638
rect 390179 -20836 390235 -20780
rect 390321 -20836 390377 -20780
rect 390179 -20978 390235 -20922
rect 390321 -20978 390377 -20922
rect 390179 -21120 390235 -21064
rect 390321 -21120 390377 -21064
rect 390179 -21262 390235 -21206
rect 390321 -21262 390377 -21206
rect 390179 -21404 390235 -21348
rect 390321 -21404 390377 -21348
rect 390179 -21546 390235 -21490
rect 390321 -21546 390377 -21490
rect 390179 -21688 390235 -21632
rect 390321 -21688 390377 -21632
rect 390179 -21830 390235 -21774
rect 390321 -21830 390377 -21774
rect 390179 -21972 390235 -21916
rect 390321 -21972 390377 -21916
rect 390179 -22114 390235 -22058
rect 390321 -22114 390377 -22058
rect 390179 -22256 390235 -22200
rect 390321 -22256 390377 -22200
rect 390179 -22398 390235 -22342
rect 390321 -22398 390377 -22342
rect 390179 -22540 390235 -22484
rect 390321 -22540 390377 -22484
rect 390179 -22682 390235 -22626
rect 390321 -22682 390377 -22626
rect 390179 -22824 390235 -22768
rect 390321 -22824 390377 -22768
rect 390179 -22966 390235 -22910
rect 390321 -22966 390377 -22910
rect 390179 -23108 390235 -23052
rect 390321 -23108 390377 -23052
rect 390179 -23250 390235 -23194
rect 390321 -23250 390377 -23194
rect 390179 -23392 390235 -23336
rect 390321 -23392 390377 -23336
rect 390179 -23534 390235 -23478
rect 390321 -23534 390377 -23478
rect 390179 -23676 390235 -23620
rect 390321 -23676 390377 -23620
rect 390179 -23818 390235 -23762
rect 390321 -23818 390377 -23762
rect 390179 -23960 390235 -23904
rect 390321 -23960 390377 -23904
rect 390179 -24102 390235 -24046
rect 390321 -24102 390377 -24046
rect 390179 -24244 390235 -24188
rect 390321 -24244 390377 -24188
rect 390179 -24386 390235 -24330
rect 390321 -24386 390377 -24330
rect 390179 -24528 390235 -24472
rect 390321 -24528 390377 -24472
rect 390179 -24670 390235 -24614
rect 390321 -24670 390377 -24614
rect 390179 -24812 390235 -24756
rect 390321 -24812 390377 -24756
rect 390179 -24954 390235 -24898
rect 390321 -24954 390377 -24898
rect 390179 -25096 390235 -25040
rect 390321 -25096 390377 -25040
rect 390179 -25238 390235 -25182
rect 390321 -25238 390377 -25182
rect 390179 -25380 390235 -25324
rect 390321 -25380 390377 -25324
rect 390179 -25522 390235 -25466
rect 390321 -25522 390377 -25466
rect 390576 -13736 390632 -13680
rect 390718 -13736 390774 -13680
rect 390576 -13878 390632 -13822
rect 390718 -13878 390774 -13822
rect 390576 -14020 390632 -13964
rect 390718 -14020 390774 -13964
rect 390576 -14162 390632 -14106
rect 390718 -14162 390774 -14106
rect 390576 -14304 390632 -14248
rect 390718 -14304 390774 -14248
rect 390576 -14446 390632 -14390
rect 390718 -14446 390774 -14390
rect 390576 -14588 390632 -14532
rect 390718 -14588 390774 -14532
rect 390576 -14730 390632 -14674
rect 390718 -14730 390774 -14674
rect 390576 -14872 390632 -14816
rect 390718 -14872 390774 -14816
rect 390576 -15014 390632 -14958
rect 390718 -15014 390774 -14958
rect 390576 -15156 390632 -15100
rect 390718 -15156 390774 -15100
rect 390576 -15298 390632 -15242
rect 390718 -15298 390774 -15242
rect 390576 -15440 390632 -15384
rect 390718 -15440 390774 -15384
rect 390576 -15582 390632 -15526
rect 390718 -15582 390774 -15526
rect 390576 -15724 390632 -15668
rect 390718 -15724 390774 -15668
rect 390576 -15866 390632 -15810
rect 390718 -15866 390774 -15810
rect 390576 -16008 390632 -15952
rect 390718 -16008 390774 -15952
rect 390576 -16150 390632 -16094
rect 390718 -16150 390774 -16094
rect 390576 -16292 390632 -16236
rect 390718 -16292 390774 -16236
rect 390576 -16434 390632 -16378
rect 390718 -16434 390774 -16378
rect 390576 -16576 390632 -16520
rect 390718 -16576 390774 -16520
rect 390576 -16718 390632 -16662
rect 390718 -16718 390774 -16662
rect 390576 -16860 390632 -16804
rect 390718 -16860 390774 -16804
rect 390576 -17002 390632 -16946
rect 390718 -17002 390774 -16946
rect 390576 -17144 390632 -17088
rect 390718 -17144 390774 -17088
rect 390576 -17286 390632 -17230
rect 390718 -17286 390774 -17230
rect 390576 -17428 390632 -17372
rect 390718 -17428 390774 -17372
rect 390576 -17570 390632 -17514
rect 390718 -17570 390774 -17514
rect 390576 -17712 390632 -17656
rect 390718 -17712 390774 -17656
rect 390576 -17854 390632 -17798
rect 390718 -17854 390774 -17798
rect 390576 -17996 390632 -17940
rect 390718 -17996 390774 -17940
rect 390576 -18138 390632 -18082
rect 390718 -18138 390774 -18082
rect 390576 -18280 390632 -18224
rect 390718 -18280 390774 -18224
rect 390576 -18422 390632 -18366
rect 390718 -18422 390774 -18366
rect 390576 -18564 390632 -18508
rect 390718 -18564 390774 -18508
rect 390576 -18706 390632 -18650
rect 390718 -18706 390774 -18650
rect 390576 -18848 390632 -18792
rect 390718 -18848 390774 -18792
rect 390576 -18990 390632 -18934
rect 390718 -18990 390774 -18934
rect 390576 -19132 390632 -19076
rect 390718 -19132 390774 -19076
rect 390576 -19274 390632 -19218
rect 390718 -19274 390774 -19218
rect 390576 -19416 390632 -19360
rect 390718 -19416 390774 -19360
rect 390576 -19558 390632 -19502
rect 390718 -19558 390774 -19502
rect 390576 -19700 390632 -19644
rect 390718 -19700 390774 -19644
rect 390576 -19842 390632 -19786
rect 390718 -19842 390774 -19786
rect 390576 -19984 390632 -19928
rect 390718 -19984 390774 -19928
rect 390576 -20126 390632 -20070
rect 390718 -20126 390774 -20070
rect 390576 -20268 390632 -20212
rect 390718 -20268 390774 -20212
rect 390576 -20410 390632 -20354
rect 390718 -20410 390774 -20354
rect 390576 -20552 390632 -20496
rect 390718 -20552 390774 -20496
rect 390576 -20694 390632 -20638
rect 390718 -20694 390774 -20638
rect 390576 -20836 390632 -20780
rect 390718 -20836 390774 -20780
rect 390576 -20978 390632 -20922
rect 390718 -20978 390774 -20922
rect 390576 -21120 390632 -21064
rect 390718 -21120 390774 -21064
rect 390576 -21262 390632 -21206
rect 390718 -21262 390774 -21206
rect 390576 -21404 390632 -21348
rect 390718 -21404 390774 -21348
rect 390576 -21546 390632 -21490
rect 390718 -21546 390774 -21490
rect 390576 -21688 390632 -21632
rect 390718 -21688 390774 -21632
rect 390576 -21830 390632 -21774
rect 390718 -21830 390774 -21774
rect 390576 -21972 390632 -21916
rect 390718 -21972 390774 -21916
rect 390576 -22114 390632 -22058
rect 390718 -22114 390774 -22058
rect 390576 -22256 390632 -22200
rect 390718 -22256 390774 -22200
rect 390576 -22398 390632 -22342
rect 390718 -22398 390774 -22342
rect 390576 -22540 390632 -22484
rect 390718 -22540 390774 -22484
rect 390576 -22682 390632 -22626
rect 390718 -22682 390774 -22626
rect 390576 -22824 390632 -22768
rect 390718 -22824 390774 -22768
rect 390576 -22966 390632 -22910
rect 390718 -22966 390774 -22910
rect 390576 -23108 390632 -23052
rect 390718 -23108 390774 -23052
rect 390576 -23250 390632 -23194
rect 390718 -23250 390774 -23194
rect 390576 -23392 390632 -23336
rect 390718 -23392 390774 -23336
rect 390576 -23534 390632 -23478
rect 390718 -23534 390774 -23478
rect 390576 -23676 390632 -23620
rect 390718 -23676 390774 -23620
rect 390576 -23818 390632 -23762
rect 390718 -23818 390774 -23762
rect 390576 -23960 390632 -23904
rect 390718 -23960 390774 -23904
rect 390576 -24102 390632 -24046
rect 390718 -24102 390774 -24046
rect 390576 -24244 390632 -24188
rect 390718 -24244 390774 -24188
rect 390576 -24386 390632 -24330
rect 390718 -24386 390774 -24330
rect 390576 -24528 390632 -24472
rect 390718 -24528 390774 -24472
rect 390576 -24670 390632 -24614
rect 390718 -24670 390774 -24614
rect 390576 -24812 390632 -24756
rect 390718 -24812 390774 -24756
rect 390576 -24954 390632 -24898
rect 390718 -24954 390774 -24898
rect 390576 -25096 390632 -25040
rect 390718 -25096 390774 -25040
rect 390576 -25238 390632 -25182
rect 390718 -25238 390774 -25182
rect 390576 -25380 390632 -25324
rect 390718 -25380 390774 -25324
rect 390576 -25522 390632 -25466
rect 390718 -25522 390774 -25466
rect 390980 -13736 391036 -13680
rect 391122 -13736 391178 -13680
rect 390980 -13878 391036 -13822
rect 391122 -13878 391178 -13822
rect 390980 -14020 391036 -13964
rect 391122 -14020 391178 -13964
rect 390980 -14162 391036 -14106
rect 391122 -14162 391178 -14106
rect 390980 -14304 391036 -14248
rect 391122 -14304 391178 -14248
rect 390980 -14446 391036 -14390
rect 391122 -14446 391178 -14390
rect 390980 -14588 391036 -14532
rect 391122 -14588 391178 -14532
rect 390980 -14730 391036 -14674
rect 391122 -14730 391178 -14674
rect 390980 -14872 391036 -14816
rect 391122 -14872 391178 -14816
rect 390980 -15014 391036 -14958
rect 391122 -15014 391178 -14958
rect 390980 -15156 391036 -15100
rect 391122 -15156 391178 -15100
rect 390980 -15298 391036 -15242
rect 391122 -15298 391178 -15242
rect 390980 -15440 391036 -15384
rect 391122 -15440 391178 -15384
rect 390980 -15582 391036 -15526
rect 391122 -15582 391178 -15526
rect 390980 -15724 391036 -15668
rect 391122 -15724 391178 -15668
rect 390980 -15866 391036 -15810
rect 391122 -15866 391178 -15810
rect 390980 -16008 391036 -15952
rect 391122 -16008 391178 -15952
rect 390980 -16150 391036 -16094
rect 391122 -16150 391178 -16094
rect 390980 -16292 391036 -16236
rect 391122 -16292 391178 -16236
rect 390980 -16434 391036 -16378
rect 391122 -16434 391178 -16378
rect 390980 -16576 391036 -16520
rect 391122 -16576 391178 -16520
rect 390980 -16718 391036 -16662
rect 391122 -16718 391178 -16662
rect 390980 -16860 391036 -16804
rect 391122 -16860 391178 -16804
rect 390980 -17002 391036 -16946
rect 391122 -17002 391178 -16946
rect 390980 -17144 391036 -17088
rect 391122 -17144 391178 -17088
rect 390980 -17286 391036 -17230
rect 391122 -17286 391178 -17230
rect 390980 -17428 391036 -17372
rect 391122 -17428 391178 -17372
rect 390980 -17570 391036 -17514
rect 391122 -17570 391178 -17514
rect 390980 -17712 391036 -17656
rect 391122 -17712 391178 -17656
rect 390980 -17854 391036 -17798
rect 391122 -17854 391178 -17798
rect 390980 -17996 391036 -17940
rect 391122 -17996 391178 -17940
rect 390980 -18138 391036 -18082
rect 391122 -18138 391178 -18082
rect 390980 -18280 391036 -18224
rect 391122 -18280 391178 -18224
rect 390980 -18422 391036 -18366
rect 391122 -18422 391178 -18366
rect 390980 -18564 391036 -18508
rect 391122 -18564 391178 -18508
rect 390980 -18706 391036 -18650
rect 391122 -18706 391178 -18650
rect 390980 -18848 391036 -18792
rect 391122 -18848 391178 -18792
rect 390980 -18990 391036 -18934
rect 391122 -18990 391178 -18934
rect 390980 -19132 391036 -19076
rect 391122 -19132 391178 -19076
rect 390980 -19274 391036 -19218
rect 391122 -19274 391178 -19218
rect 390980 -19416 391036 -19360
rect 391122 -19416 391178 -19360
rect 390980 -19558 391036 -19502
rect 391122 -19558 391178 -19502
rect 390980 -19700 391036 -19644
rect 391122 -19700 391178 -19644
rect 390980 -19842 391036 -19786
rect 391122 -19842 391178 -19786
rect 390980 -19984 391036 -19928
rect 391122 -19984 391178 -19928
rect 390980 -20126 391036 -20070
rect 391122 -20126 391178 -20070
rect 390980 -20268 391036 -20212
rect 391122 -20268 391178 -20212
rect 390980 -20410 391036 -20354
rect 391122 -20410 391178 -20354
rect 390980 -20552 391036 -20496
rect 391122 -20552 391178 -20496
rect 390980 -20694 391036 -20638
rect 391122 -20694 391178 -20638
rect 390980 -20836 391036 -20780
rect 391122 -20836 391178 -20780
rect 390980 -20978 391036 -20922
rect 391122 -20978 391178 -20922
rect 390980 -21120 391036 -21064
rect 391122 -21120 391178 -21064
rect 390980 -21262 391036 -21206
rect 391122 -21262 391178 -21206
rect 390980 -21404 391036 -21348
rect 391122 -21404 391178 -21348
rect 390980 -21546 391036 -21490
rect 391122 -21546 391178 -21490
rect 390980 -21688 391036 -21632
rect 391122 -21688 391178 -21632
rect 390980 -21830 391036 -21774
rect 391122 -21830 391178 -21774
rect 390980 -21972 391036 -21916
rect 391122 -21972 391178 -21916
rect 390980 -22114 391036 -22058
rect 391122 -22114 391178 -22058
rect 390980 -22256 391036 -22200
rect 391122 -22256 391178 -22200
rect 390980 -22398 391036 -22342
rect 391122 -22398 391178 -22342
rect 390980 -22540 391036 -22484
rect 391122 -22540 391178 -22484
rect 390980 -22682 391036 -22626
rect 391122 -22682 391178 -22626
rect 390980 -22824 391036 -22768
rect 391122 -22824 391178 -22768
rect 390980 -22966 391036 -22910
rect 391122 -22966 391178 -22910
rect 390980 -23108 391036 -23052
rect 391122 -23108 391178 -23052
rect 390980 -23250 391036 -23194
rect 391122 -23250 391178 -23194
rect 390980 -23392 391036 -23336
rect 391122 -23392 391178 -23336
rect 390980 -23534 391036 -23478
rect 391122 -23534 391178 -23478
rect 390980 -23676 391036 -23620
rect 391122 -23676 391178 -23620
rect 390980 -23818 391036 -23762
rect 391122 -23818 391178 -23762
rect 390980 -23960 391036 -23904
rect 391122 -23960 391178 -23904
rect 390980 -24102 391036 -24046
rect 391122 -24102 391178 -24046
rect 390980 -24244 391036 -24188
rect 391122 -24244 391178 -24188
rect 390980 -24386 391036 -24330
rect 391122 -24386 391178 -24330
rect 390980 -24528 391036 -24472
rect 391122 -24528 391178 -24472
rect 390980 -24670 391036 -24614
rect 391122 -24670 391178 -24614
rect 390980 -24812 391036 -24756
rect 391122 -24812 391178 -24756
rect 390980 -24954 391036 -24898
rect 391122 -24954 391178 -24898
rect 390980 -25096 391036 -25040
rect 391122 -25096 391178 -25040
rect 390980 -25238 391036 -25182
rect 391122 -25238 391178 -25182
rect 390980 -25380 391036 -25324
rect 391122 -25380 391178 -25324
rect 390980 -25522 391036 -25466
rect 391122 -25522 391178 -25466
rect 391376 -13736 391432 -13680
rect 391518 -13736 391574 -13680
rect 391376 -13878 391432 -13822
rect 391518 -13878 391574 -13822
rect 391376 -14020 391432 -13964
rect 391518 -14020 391574 -13964
rect 391376 -14162 391432 -14106
rect 391518 -14162 391574 -14106
rect 391376 -14304 391432 -14248
rect 391518 -14304 391574 -14248
rect 391376 -14446 391432 -14390
rect 391518 -14446 391574 -14390
rect 391376 -14588 391432 -14532
rect 391518 -14588 391574 -14532
rect 391376 -14730 391432 -14674
rect 391518 -14730 391574 -14674
rect 391376 -14872 391432 -14816
rect 391518 -14872 391574 -14816
rect 391376 -15014 391432 -14958
rect 391518 -15014 391574 -14958
rect 391376 -15156 391432 -15100
rect 391518 -15156 391574 -15100
rect 391376 -15298 391432 -15242
rect 391518 -15298 391574 -15242
rect 391376 -15440 391432 -15384
rect 391518 -15440 391574 -15384
rect 391376 -15582 391432 -15526
rect 391518 -15582 391574 -15526
rect 391376 -15724 391432 -15668
rect 391518 -15724 391574 -15668
rect 391376 -15866 391432 -15810
rect 391518 -15866 391574 -15810
rect 391376 -16008 391432 -15952
rect 391518 -16008 391574 -15952
rect 391376 -16150 391432 -16094
rect 391518 -16150 391574 -16094
rect 391376 -16292 391432 -16236
rect 391518 -16292 391574 -16236
rect 391376 -16434 391432 -16378
rect 391518 -16434 391574 -16378
rect 391376 -16576 391432 -16520
rect 391518 -16576 391574 -16520
rect 391376 -16718 391432 -16662
rect 391518 -16718 391574 -16662
rect 391376 -16860 391432 -16804
rect 391518 -16860 391574 -16804
rect 391376 -17002 391432 -16946
rect 391518 -17002 391574 -16946
rect 391376 -17144 391432 -17088
rect 391518 -17144 391574 -17088
rect 391376 -17286 391432 -17230
rect 391518 -17286 391574 -17230
rect 391376 -17428 391432 -17372
rect 391518 -17428 391574 -17372
rect 391376 -17570 391432 -17514
rect 391518 -17570 391574 -17514
rect 391376 -17712 391432 -17656
rect 391518 -17712 391574 -17656
rect 391376 -17854 391432 -17798
rect 391518 -17854 391574 -17798
rect 391376 -17996 391432 -17940
rect 391518 -17996 391574 -17940
rect 391376 -18138 391432 -18082
rect 391518 -18138 391574 -18082
rect 391376 -18280 391432 -18224
rect 391518 -18280 391574 -18224
rect 391376 -18422 391432 -18366
rect 391518 -18422 391574 -18366
rect 391376 -18564 391432 -18508
rect 391518 -18564 391574 -18508
rect 391376 -18706 391432 -18650
rect 391518 -18706 391574 -18650
rect 391376 -18848 391432 -18792
rect 391518 -18848 391574 -18792
rect 391376 -18990 391432 -18934
rect 391518 -18990 391574 -18934
rect 391376 -19132 391432 -19076
rect 391518 -19132 391574 -19076
rect 391376 -19274 391432 -19218
rect 391518 -19274 391574 -19218
rect 391376 -19416 391432 -19360
rect 391518 -19416 391574 -19360
rect 391376 -19558 391432 -19502
rect 391518 -19558 391574 -19502
rect 391376 -19700 391432 -19644
rect 391518 -19700 391574 -19644
rect 391376 -19842 391432 -19786
rect 391518 -19842 391574 -19786
rect 391376 -19984 391432 -19928
rect 391518 -19984 391574 -19928
rect 391376 -20126 391432 -20070
rect 391518 -20126 391574 -20070
rect 391376 -20268 391432 -20212
rect 391518 -20268 391574 -20212
rect 391376 -20410 391432 -20354
rect 391518 -20410 391574 -20354
rect 391376 -20552 391432 -20496
rect 391518 -20552 391574 -20496
rect 391376 -20694 391432 -20638
rect 391518 -20694 391574 -20638
rect 391376 -20836 391432 -20780
rect 391518 -20836 391574 -20780
rect 391376 -20978 391432 -20922
rect 391518 -20978 391574 -20922
rect 391376 -21120 391432 -21064
rect 391518 -21120 391574 -21064
rect 391376 -21262 391432 -21206
rect 391518 -21262 391574 -21206
rect 391376 -21404 391432 -21348
rect 391518 -21404 391574 -21348
rect 391376 -21546 391432 -21490
rect 391518 -21546 391574 -21490
rect 391376 -21688 391432 -21632
rect 391518 -21688 391574 -21632
rect 391376 -21830 391432 -21774
rect 391518 -21830 391574 -21774
rect 391376 -21972 391432 -21916
rect 391518 -21972 391574 -21916
rect 391376 -22114 391432 -22058
rect 391518 -22114 391574 -22058
rect 391376 -22256 391432 -22200
rect 391518 -22256 391574 -22200
rect 391376 -22398 391432 -22342
rect 391518 -22398 391574 -22342
rect 391376 -22540 391432 -22484
rect 391518 -22540 391574 -22484
rect 391376 -22682 391432 -22626
rect 391518 -22682 391574 -22626
rect 391376 -22824 391432 -22768
rect 391518 -22824 391574 -22768
rect 391376 -22966 391432 -22910
rect 391518 -22966 391574 -22910
rect 391376 -23108 391432 -23052
rect 391518 -23108 391574 -23052
rect 391376 -23250 391432 -23194
rect 391518 -23250 391574 -23194
rect 391376 -23392 391432 -23336
rect 391518 -23392 391574 -23336
rect 391376 -23534 391432 -23478
rect 391518 -23534 391574 -23478
rect 391376 -23676 391432 -23620
rect 391518 -23676 391574 -23620
rect 391376 -23818 391432 -23762
rect 391518 -23818 391574 -23762
rect 391376 -23960 391432 -23904
rect 391518 -23960 391574 -23904
rect 391376 -24102 391432 -24046
rect 391518 -24102 391574 -24046
rect 391376 -24244 391432 -24188
rect 391518 -24244 391574 -24188
rect 391376 -24386 391432 -24330
rect 391518 -24386 391574 -24330
rect 391376 -24528 391432 -24472
rect 391518 -24528 391574 -24472
rect 391376 -24670 391432 -24614
rect 391518 -24670 391574 -24614
rect 391376 -24812 391432 -24756
rect 391518 -24812 391574 -24756
rect 391376 -24954 391432 -24898
rect 391518 -24954 391574 -24898
rect 391376 -25096 391432 -25040
rect 391518 -25096 391574 -25040
rect 391376 -25238 391432 -25182
rect 391518 -25238 391574 -25182
rect 391376 -25380 391432 -25324
rect 391518 -25380 391574 -25324
rect 391376 -25522 391432 -25466
rect 391518 -25522 391574 -25466
rect 391776 -13736 391832 -13680
rect 391918 -13736 391974 -13680
rect 391776 -13878 391832 -13822
rect 391918 -13878 391974 -13822
rect 391776 -14020 391832 -13964
rect 391918 -14020 391974 -13964
rect 391776 -14162 391832 -14106
rect 391918 -14162 391974 -14106
rect 391776 -14304 391832 -14248
rect 391918 -14304 391974 -14248
rect 391776 -14446 391832 -14390
rect 391918 -14446 391974 -14390
rect 391776 -14588 391832 -14532
rect 391918 -14588 391974 -14532
rect 391776 -14730 391832 -14674
rect 391918 -14730 391974 -14674
rect 391776 -14872 391832 -14816
rect 391918 -14872 391974 -14816
rect 391776 -15014 391832 -14958
rect 391918 -15014 391974 -14958
rect 391776 -15156 391832 -15100
rect 391918 -15156 391974 -15100
rect 391776 -15298 391832 -15242
rect 391918 -15298 391974 -15242
rect 391776 -15440 391832 -15384
rect 391918 -15440 391974 -15384
rect 391776 -15582 391832 -15526
rect 391918 -15582 391974 -15526
rect 391776 -15724 391832 -15668
rect 391918 -15724 391974 -15668
rect 391776 -15866 391832 -15810
rect 391918 -15866 391974 -15810
rect 391776 -16008 391832 -15952
rect 391918 -16008 391974 -15952
rect 391776 -16150 391832 -16094
rect 391918 -16150 391974 -16094
rect 391776 -16292 391832 -16236
rect 391918 -16292 391974 -16236
rect 391776 -16434 391832 -16378
rect 391918 -16434 391974 -16378
rect 391776 -16576 391832 -16520
rect 391918 -16576 391974 -16520
rect 391776 -16718 391832 -16662
rect 391918 -16718 391974 -16662
rect 391776 -16860 391832 -16804
rect 391918 -16860 391974 -16804
rect 391776 -17002 391832 -16946
rect 391918 -17002 391974 -16946
rect 391776 -17144 391832 -17088
rect 391918 -17144 391974 -17088
rect 391776 -17286 391832 -17230
rect 391918 -17286 391974 -17230
rect 391776 -17428 391832 -17372
rect 391918 -17428 391974 -17372
rect 391776 -17570 391832 -17514
rect 391918 -17570 391974 -17514
rect 391776 -17712 391832 -17656
rect 391918 -17712 391974 -17656
rect 391776 -17854 391832 -17798
rect 391918 -17854 391974 -17798
rect 391776 -17996 391832 -17940
rect 391918 -17996 391974 -17940
rect 391776 -18138 391832 -18082
rect 391918 -18138 391974 -18082
rect 391776 -18280 391832 -18224
rect 391918 -18280 391974 -18224
rect 391776 -18422 391832 -18366
rect 391918 -18422 391974 -18366
rect 391776 -18564 391832 -18508
rect 391918 -18564 391974 -18508
rect 391776 -18706 391832 -18650
rect 391918 -18706 391974 -18650
rect 391776 -18848 391832 -18792
rect 391918 -18848 391974 -18792
rect 391776 -18990 391832 -18934
rect 391918 -18990 391974 -18934
rect 391776 -19132 391832 -19076
rect 391918 -19132 391974 -19076
rect 391776 -19274 391832 -19218
rect 391918 -19274 391974 -19218
rect 391776 -19416 391832 -19360
rect 391918 -19416 391974 -19360
rect 391776 -19558 391832 -19502
rect 391918 -19558 391974 -19502
rect 391776 -19700 391832 -19644
rect 391918 -19700 391974 -19644
rect 391776 -19842 391832 -19786
rect 391918 -19842 391974 -19786
rect 391776 -19984 391832 -19928
rect 391918 -19984 391974 -19928
rect 391776 -20126 391832 -20070
rect 391918 -20126 391974 -20070
rect 391776 -20268 391832 -20212
rect 391918 -20268 391974 -20212
rect 391776 -20410 391832 -20354
rect 391918 -20410 391974 -20354
rect 391776 -20552 391832 -20496
rect 391918 -20552 391974 -20496
rect 391776 -20694 391832 -20638
rect 391918 -20694 391974 -20638
rect 391776 -20836 391832 -20780
rect 391918 -20836 391974 -20780
rect 391776 -20978 391832 -20922
rect 391918 -20978 391974 -20922
rect 391776 -21120 391832 -21064
rect 391918 -21120 391974 -21064
rect 391776 -21262 391832 -21206
rect 391918 -21262 391974 -21206
rect 391776 -21404 391832 -21348
rect 391918 -21404 391974 -21348
rect 391776 -21546 391832 -21490
rect 391918 -21546 391974 -21490
rect 391776 -21688 391832 -21632
rect 391918 -21688 391974 -21632
rect 391776 -21830 391832 -21774
rect 391918 -21830 391974 -21774
rect 391776 -21972 391832 -21916
rect 391918 -21972 391974 -21916
rect 391776 -22114 391832 -22058
rect 391918 -22114 391974 -22058
rect 391776 -22256 391832 -22200
rect 391918 -22256 391974 -22200
rect 391776 -22398 391832 -22342
rect 391918 -22398 391974 -22342
rect 391776 -22540 391832 -22484
rect 391918 -22540 391974 -22484
rect 391776 -22682 391832 -22626
rect 391918 -22682 391974 -22626
rect 391776 -22824 391832 -22768
rect 391918 -22824 391974 -22768
rect 391776 -22966 391832 -22910
rect 391918 -22966 391974 -22910
rect 391776 -23108 391832 -23052
rect 391918 -23108 391974 -23052
rect 391776 -23250 391832 -23194
rect 391918 -23250 391974 -23194
rect 391776 -23392 391832 -23336
rect 391918 -23392 391974 -23336
rect 391776 -23534 391832 -23478
rect 391918 -23534 391974 -23478
rect 391776 -23676 391832 -23620
rect 391918 -23676 391974 -23620
rect 391776 -23818 391832 -23762
rect 391918 -23818 391974 -23762
rect 391776 -23960 391832 -23904
rect 391918 -23960 391974 -23904
rect 391776 -24102 391832 -24046
rect 391918 -24102 391974 -24046
rect 391776 -24244 391832 -24188
rect 391918 -24244 391974 -24188
rect 391776 -24386 391832 -24330
rect 391918 -24386 391974 -24330
rect 391776 -24528 391832 -24472
rect 391918 -24528 391974 -24472
rect 391776 -24670 391832 -24614
rect 391918 -24670 391974 -24614
rect 391776 -24812 391832 -24756
rect 391918 -24812 391974 -24756
rect 391776 -24954 391832 -24898
rect 391918 -24954 391974 -24898
rect 391776 -25096 391832 -25040
rect 391918 -25096 391974 -25040
rect 391776 -25238 391832 -25182
rect 391918 -25238 391974 -25182
rect 391776 -25380 391832 -25324
rect 391918 -25380 391974 -25324
rect 391776 -25522 391832 -25466
rect 391918 -25522 391974 -25466
rect 392173 -13736 392229 -13680
rect 392315 -13736 392371 -13680
rect 392173 -13878 392229 -13822
rect 392315 -13878 392371 -13822
rect 392173 -14020 392229 -13964
rect 392315 -14020 392371 -13964
rect 392173 -14162 392229 -14106
rect 392315 -14162 392371 -14106
rect 392173 -14304 392229 -14248
rect 392315 -14304 392371 -14248
rect 392173 -14446 392229 -14390
rect 392315 -14446 392371 -14390
rect 392173 -14588 392229 -14532
rect 392315 -14588 392371 -14532
rect 392173 -14730 392229 -14674
rect 392315 -14730 392371 -14674
rect 392173 -14872 392229 -14816
rect 392315 -14872 392371 -14816
rect 392173 -15014 392229 -14958
rect 392315 -15014 392371 -14958
rect 392173 -15156 392229 -15100
rect 392315 -15156 392371 -15100
rect 392173 -15298 392229 -15242
rect 392315 -15298 392371 -15242
rect 392173 -15440 392229 -15384
rect 392315 -15440 392371 -15384
rect 392173 -15582 392229 -15526
rect 392315 -15582 392371 -15526
rect 392173 -15724 392229 -15668
rect 392315 -15724 392371 -15668
rect 392173 -15866 392229 -15810
rect 392315 -15866 392371 -15810
rect 392173 -16008 392229 -15952
rect 392315 -16008 392371 -15952
rect 392173 -16150 392229 -16094
rect 392315 -16150 392371 -16094
rect 392173 -16292 392229 -16236
rect 392315 -16292 392371 -16236
rect 392173 -16434 392229 -16378
rect 392315 -16434 392371 -16378
rect 392173 -16576 392229 -16520
rect 392315 -16576 392371 -16520
rect 392173 -16718 392229 -16662
rect 392315 -16718 392371 -16662
rect 392173 -16860 392229 -16804
rect 392315 -16860 392371 -16804
rect 392173 -17002 392229 -16946
rect 392315 -17002 392371 -16946
rect 392173 -17144 392229 -17088
rect 392315 -17144 392371 -17088
rect 392173 -17286 392229 -17230
rect 392315 -17286 392371 -17230
rect 392173 -17428 392229 -17372
rect 392315 -17428 392371 -17372
rect 392173 -17570 392229 -17514
rect 392315 -17570 392371 -17514
rect 392173 -17712 392229 -17656
rect 392315 -17712 392371 -17656
rect 392173 -17854 392229 -17798
rect 392315 -17854 392371 -17798
rect 392173 -17996 392229 -17940
rect 392315 -17996 392371 -17940
rect 392173 -18138 392229 -18082
rect 392315 -18138 392371 -18082
rect 392173 -18280 392229 -18224
rect 392315 -18280 392371 -18224
rect 392173 -18422 392229 -18366
rect 392315 -18422 392371 -18366
rect 392173 -18564 392229 -18508
rect 392315 -18564 392371 -18508
rect 392173 -18706 392229 -18650
rect 392315 -18706 392371 -18650
rect 392173 -18848 392229 -18792
rect 392315 -18848 392371 -18792
rect 392173 -18990 392229 -18934
rect 392315 -18990 392371 -18934
rect 392173 -19132 392229 -19076
rect 392315 -19132 392371 -19076
rect 392173 -19274 392229 -19218
rect 392315 -19274 392371 -19218
rect 392173 -19416 392229 -19360
rect 392315 -19416 392371 -19360
rect 392173 -19558 392229 -19502
rect 392315 -19558 392371 -19502
rect 392173 -19700 392229 -19644
rect 392315 -19700 392371 -19644
rect 392173 -19842 392229 -19786
rect 392315 -19842 392371 -19786
rect 392173 -19984 392229 -19928
rect 392315 -19984 392371 -19928
rect 392173 -20126 392229 -20070
rect 392315 -20126 392371 -20070
rect 392173 -20268 392229 -20212
rect 392315 -20268 392371 -20212
rect 392173 -20410 392229 -20354
rect 392315 -20410 392371 -20354
rect 392173 -20552 392229 -20496
rect 392315 -20552 392371 -20496
rect 392173 -20694 392229 -20638
rect 392315 -20694 392371 -20638
rect 392173 -20836 392229 -20780
rect 392315 -20836 392371 -20780
rect 392173 -20978 392229 -20922
rect 392315 -20978 392371 -20922
rect 392173 -21120 392229 -21064
rect 392315 -21120 392371 -21064
rect 392173 -21262 392229 -21206
rect 392315 -21262 392371 -21206
rect 392173 -21404 392229 -21348
rect 392315 -21404 392371 -21348
rect 392173 -21546 392229 -21490
rect 392315 -21546 392371 -21490
rect 392173 -21688 392229 -21632
rect 392315 -21688 392371 -21632
rect 392173 -21830 392229 -21774
rect 392315 -21830 392371 -21774
rect 392173 -21972 392229 -21916
rect 392315 -21972 392371 -21916
rect 392173 -22114 392229 -22058
rect 392315 -22114 392371 -22058
rect 392173 -22256 392229 -22200
rect 392315 -22256 392371 -22200
rect 392173 -22398 392229 -22342
rect 392315 -22398 392371 -22342
rect 392173 -22540 392229 -22484
rect 392315 -22540 392371 -22484
rect 392173 -22682 392229 -22626
rect 392315 -22682 392371 -22626
rect 392173 -22824 392229 -22768
rect 392315 -22824 392371 -22768
rect 392173 -22966 392229 -22910
rect 392315 -22966 392371 -22910
rect 392173 -23108 392229 -23052
rect 392315 -23108 392371 -23052
rect 392173 -23250 392229 -23194
rect 392315 -23250 392371 -23194
rect 392173 -23392 392229 -23336
rect 392315 -23392 392371 -23336
rect 392173 -23534 392229 -23478
rect 392315 -23534 392371 -23478
rect 392173 -23676 392229 -23620
rect 392315 -23676 392371 -23620
rect 392173 -23818 392229 -23762
rect 392315 -23818 392371 -23762
rect 392173 -23960 392229 -23904
rect 392315 -23960 392371 -23904
rect 392173 -24102 392229 -24046
rect 392315 -24102 392371 -24046
rect 392173 -24244 392229 -24188
rect 392315 -24244 392371 -24188
rect 392173 -24386 392229 -24330
rect 392315 -24386 392371 -24330
rect 392173 -24528 392229 -24472
rect 392315 -24528 392371 -24472
rect 392173 -24670 392229 -24614
rect 392315 -24670 392371 -24614
rect 392173 -24812 392229 -24756
rect 392315 -24812 392371 -24756
rect 392173 -24954 392229 -24898
rect 392315 -24954 392371 -24898
rect 392173 -25096 392229 -25040
rect 392315 -25096 392371 -25040
rect 392173 -25238 392229 -25182
rect 392315 -25238 392371 -25182
rect 392173 -25380 392229 -25324
rect 392315 -25380 392371 -25324
rect 392173 -25522 392229 -25466
rect 392315 -25522 392371 -25466
rect 392578 -13736 392634 -13680
rect 392720 -13736 392776 -13680
rect 392578 -13878 392634 -13822
rect 392720 -13878 392776 -13822
rect 392578 -14020 392634 -13964
rect 392720 -14020 392776 -13964
rect 392578 -14162 392634 -14106
rect 392720 -14162 392776 -14106
rect 392578 -14304 392634 -14248
rect 392720 -14304 392776 -14248
rect 392578 -14446 392634 -14390
rect 392720 -14446 392776 -14390
rect 392578 -14588 392634 -14532
rect 392720 -14588 392776 -14532
rect 392578 -14730 392634 -14674
rect 392720 -14730 392776 -14674
rect 392578 -14872 392634 -14816
rect 392720 -14872 392776 -14816
rect 392578 -15014 392634 -14958
rect 392720 -15014 392776 -14958
rect 392578 -15156 392634 -15100
rect 392720 -15156 392776 -15100
rect 392578 -15298 392634 -15242
rect 392720 -15298 392776 -15242
rect 392578 -15440 392634 -15384
rect 392720 -15440 392776 -15384
rect 392578 -15582 392634 -15526
rect 392720 -15582 392776 -15526
rect 392578 -15724 392634 -15668
rect 392720 -15724 392776 -15668
rect 392578 -15866 392634 -15810
rect 392720 -15866 392776 -15810
rect 392578 -16008 392634 -15952
rect 392720 -16008 392776 -15952
rect 392578 -16150 392634 -16094
rect 392720 -16150 392776 -16094
rect 392578 -16292 392634 -16236
rect 392720 -16292 392776 -16236
rect 392578 -16434 392634 -16378
rect 392720 -16434 392776 -16378
rect 392578 -16576 392634 -16520
rect 392720 -16576 392776 -16520
rect 392578 -16718 392634 -16662
rect 392720 -16718 392776 -16662
rect 392578 -16860 392634 -16804
rect 392720 -16860 392776 -16804
rect 392578 -17002 392634 -16946
rect 392720 -17002 392776 -16946
rect 392578 -17144 392634 -17088
rect 392720 -17144 392776 -17088
rect 392578 -17286 392634 -17230
rect 392720 -17286 392776 -17230
rect 392578 -17428 392634 -17372
rect 392720 -17428 392776 -17372
rect 392578 -17570 392634 -17514
rect 392720 -17570 392776 -17514
rect 392578 -17712 392634 -17656
rect 392720 -17712 392776 -17656
rect 392578 -17854 392634 -17798
rect 392720 -17854 392776 -17798
rect 392578 -17996 392634 -17940
rect 392720 -17996 392776 -17940
rect 392578 -18138 392634 -18082
rect 392720 -18138 392776 -18082
rect 392578 -18280 392634 -18224
rect 392720 -18280 392776 -18224
rect 392578 -18422 392634 -18366
rect 392720 -18422 392776 -18366
rect 392578 -18564 392634 -18508
rect 392720 -18564 392776 -18508
rect 392578 -18706 392634 -18650
rect 392720 -18706 392776 -18650
rect 392578 -18848 392634 -18792
rect 392720 -18848 392776 -18792
rect 392578 -18990 392634 -18934
rect 392720 -18990 392776 -18934
rect 392578 -19132 392634 -19076
rect 392720 -19132 392776 -19076
rect 392578 -19274 392634 -19218
rect 392720 -19274 392776 -19218
rect 392578 -19416 392634 -19360
rect 392720 -19416 392776 -19360
rect 392578 -19558 392634 -19502
rect 392720 -19558 392776 -19502
rect 392578 -19700 392634 -19644
rect 392720 -19700 392776 -19644
rect 392578 -19842 392634 -19786
rect 392720 -19842 392776 -19786
rect 392578 -19984 392634 -19928
rect 392720 -19984 392776 -19928
rect 392578 -20126 392634 -20070
rect 392720 -20126 392776 -20070
rect 392578 -20268 392634 -20212
rect 392720 -20268 392776 -20212
rect 392578 -20410 392634 -20354
rect 392720 -20410 392776 -20354
rect 392578 -20552 392634 -20496
rect 392720 -20552 392776 -20496
rect 392578 -20694 392634 -20638
rect 392720 -20694 392776 -20638
rect 392578 -20836 392634 -20780
rect 392720 -20836 392776 -20780
rect 392578 -20978 392634 -20922
rect 392720 -20978 392776 -20922
rect 392578 -21120 392634 -21064
rect 392720 -21120 392776 -21064
rect 392578 -21262 392634 -21206
rect 392720 -21262 392776 -21206
rect 392578 -21404 392634 -21348
rect 392720 -21404 392776 -21348
rect 392578 -21546 392634 -21490
rect 392720 -21546 392776 -21490
rect 392578 -21688 392634 -21632
rect 392720 -21688 392776 -21632
rect 392578 -21830 392634 -21774
rect 392720 -21830 392776 -21774
rect 392578 -21972 392634 -21916
rect 392720 -21972 392776 -21916
rect 392578 -22114 392634 -22058
rect 392720 -22114 392776 -22058
rect 392578 -22256 392634 -22200
rect 392720 -22256 392776 -22200
rect 392578 -22398 392634 -22342
rect 392720 -22398 392776 -22342
rect 392578 -22540 392634 -22484
rect 392720 -22540 392776 -22484
rect 392578 -22682 392634 -22626
rect 392720 -22682 392776 -22626
rect 392578 -22824 392634 -22768
rect 392720 -22824 392776 -22768
rect 392578 -22966 392634 -22910
rect 392720 -22966 392776 -22910
rect 392578 -23108 392634 -23052
rect 392720 -23108 392776 -23052
rect 392578 -23250 392634 -23194
rect 392720 -23250 392776 -23194
rect 392578 -23392 392634 -23336
rect 392720 -23392 392776 -23336
rect 392578 -23534 392634 -23478
rect 392720 -23534 392776 -23478
rect 392578 -23676 392634 -23620
rect 392720 -23676 392776 -23620
rect 392578 -23818 392634 -23762
rect 392720 -23818 392776 -23762
rect 392578 -23960 392634 -23904
rect 392720 -23960 392776 -23904
rect 392578 -24102 392634 -24046
rect 392720 -24102 392776 -24046
rect 392578 -24244 392634 -24188
rect 392720 -24244 392776 -24188
rect 392578 -24386 392634 -24330
rect 392720 -24386 392776 -24330
rect 392578 -24528 392634 -24472
rect 392720 -24528 392776 -24472
rect 392578 -24670 392634 -24614
rect 392720 -24670 392776 -24614
rect 392578 -24812 392634 -24756
rect 392720 -24812 392776 -24756
rect 392578 -24954 392634 -24898
rect 392720 -24954 392776 -24898
rect 392578 -25096 392634 -25040
rect 392720 -25096 392776 -25040
rect 392578 -25238 392634 -25182
rect 392720 -25238 392776 -25182
rect 392578 -25380 392634 -25324
rect 392720 -25380 392776 -25324
rect 392578 -25522 392634 -25466
rect 392720 -25522 392776 -25466
rect 392978 -13736 393034 -13680
rect 393120 -13736 393176 -13680
rect 392978 -13878 393034 -13822
rect 393120 -13878 393176 -13822
rect 392978 -14020 393034 -13964
rect 393120 -14020 393176 -13964
rect 392978 -14162 393034 -14106
rect 393120 -14162 393176 -14106
rect 392978 -14304 393034 -14248
rect 393120 -14304 393176 -14248
rect 392978 -14446 393034 -14390
rect 393120 -14446 393176 -14390
rect 392978 -14588 393034 -14532
rect 393120 -14588 393176 -14532
rect 392978 -14730 393034 -14674
rect 393120 -14730 393176 -14674
rect 392978 -14872 393034 -14816
rect 393120 -14872 393176 -14816
rect 392978 -15014 393034 -14958
rect 393120 -15014 393176 -14958
rect 392978 -15156 393034 -15100
rect 393120 -15156 393176 -15100
rect 392978 -15298 393034 -15242
rect 393120 -15298 393176 -15242
rect 392978 -15440 393034 -15384
rect 393120 -15440 393176 -15384
rect 392978 -15582 393034 -15526
rect 393120 -15582 393176 -15526
rect 392978 -15724 393034 -15668
rect 393120 -15724 393176 -15668
rect 392978 -15866 393034 -15810
rect 393120 -15866 393176 -15810
rect 392978 -16008 393034 -15952
rect 393120 -16008 393176 -15952
rect 392978 -16150 393034 -16094
rect 393120 -16150 393176 -16094
rect 392978 -16292 393034 -16236
rect 393120 -16292 393176 -16236
rect 392978 -16434 393034 -16378
rect 393120 -16434 393176 -16378
rect 392978 -16576 393034 -16520
rect 393120 -16576 393176 -16520
rect 392978 -16718 393034 -16662
rect 393120 -16718 393176 -16662
rect 392978 -16860 393034 -16804
rect 393120 -16860 393176 -16804
rect 392978 -17002 393034 -16946
rect 393120 -17002 393176 -16946
rect 392978 -17144 393034 -17088
rect 393120 -17144 393176 -17088
rect 392978 -17286 393034 -17230
rect 393120 -17286 393176 -17230
rect 392978 -17428 393034 -17372
rect 393120 -17428 393176 -17372
rect 392978 -17570 393034 -17514
rect 393120 -17570 393176 -17514
rect 392978 -17712 393034 -17656
rect 393120 -17712 393176 -17656
rect 392978 -17854 393034 -17798
rect 393120 -17854 393176 -17798
rect 392978 -17996 393034 -17940
rect 393120 -17996 393176 -17940
rect 392978 -18138 393034 -18082
rect 393120 -18138 393176 -18082
rect 392978 -18280 393034 -18224
rect 393120 -18280 393176 -18224
rect 392978 -18422 393034 -18366
rect 393120 -18422 393176 -18366
rect 392978 -18564 393034 -18508
rect 393120 -18564 393176 -18508
rect 392978 -18706 393034 -18650
rect 393120 -18706 393176 -18650
rect 392978 -18848 393034 -18792
rect 393120 -18848 393176 -18792
rect 392978 -18990 393034 -18934
rect 393120 -18990 393176 -18934
rect 392978 -19132 393034 -19076
rect 393120 -19132 393176 -19076
rect 392978 -19274 393034 -19218
rect 393120 -19274 393176 -19218
rect 392978 -19416 393034 -19360
rect 393120 -19416 393176 -19360
rect 392978 -19558 393034 -19502
rect 393120 -19558 393176 -19502
rect 392978 -19700 393034 -19644
rect 393120 -19700 393176 -19644
rect 392978 -19842 393034 -19786
rect 393120 -19842 393176 -19786
rect 392978 -19984 393034 -19928
rect 393120 -19984 393176 -19928
rect 392978 -20126 393034 -20070
rect 393120 -20126 393176 -20070
rect 392978 -20268 393034 -20212
rect 393120 -20268 393176 -20212
rect 392978 -20410 393034 -20354
rect 393120 -20410 393176 -20354
rect 392978 -20552 393034 -20496
rect 393120 -20552 393176 -20496
rect 392978 -20694 393034 -20638
rect 393120 -20694 393176 -20638
rect 392978 -20836 393034 -20780
rect 393120 -20836 393176 -20780
rect 392978 -20978 393034 -20922
rect 393120 -20978 393176 -20922
rect 392978 -21120 393034 -21064
rect 393120 -21120 393176 -21064
rect 392978 -21262 393034 -21206
rect 393120 -21262 393176 -21206
rect 392978 -21404 393034 -21348
rect 393120 -21404 393176 -21348
rect 392978 -21546 393034 -21490
rect 393120 -21546 393176 -21490
rect 392978 -21688 393034 -21632
rect 393120 -21688 393176 -21632
rect 392978 -21830 393034 -21774
rect 393120 -21830 393176 -21774
rect 392978 -21972 393034 -21916
rect 393120 -21972 393176 -21916
rect 392978 -22114 393034 -22058
rect 393120 -22114 393176 -22058
rect 392978 -22256 393034 -22200
rect 393120 -22256 393176 -22200
rect 392978 -22398 393034 -22342
rect 393120 -22398 393176 -22342
rect 392978 -22540 393034 -22484
rect 393120 -22540 393176 -22484
rect 392978 -22682 393034 -22626
rect 393120 -22682 393176 -22626
rect 392978 -22824 393034 -22768
rect 393120 -22824 393176 -22768
rect 392978 -22966 393034 -22910
rect 393120 -22966 393176 -22910
rect 392978 -23108 393034 -23052
rect 393120 -23108 393176 -23052
rect 392978 -23250 393034 -23194
rect 393120 -23250 393176 -23194
rect 392978 -23392 393034 -23336
rect 393120 -23392 393176 -23336
rect 392978 -23534 393034 -23478
rect 393120 -23534 393176 -23478
rect 392978 -23676 393034 -23620
rect 393120 -23676 393176 -23620
rect 392978 -23818 393034 -23762
rect 393120 -23818 393176 -23762
rect 392978 -23960 393034 -23904
rect 393120 -23960 393176 -23904
rect 392978 -24102 393034 -24046
rect 393120 -24102 393176 -24046
rect 392978 -24244 393034 -24188
rect 393120 -24244 393176 -24188
rect 392978 -24386 393034 -24330
rect 393120 -24386 393176 -24330
rect 392978 -24528 393034 -24472
rect 393120 -24528 393176 -24472
rect 392978 -24670 393034 -24614
rect 393120 -24670 393176 -24614
rect 392978 -24812 393034 -24756
rect 393120 -24812 393176 -24756
rect 392978 -24954 393034 -24898
rect 393120 -24954 393176 -24898
rect 392978 -25096 393034 -25040
rect 393120 -25096 393176 -25040
rect 392978 -25238 393034 -25182
rect 393120 -25238 393176 -25182
rect 392978 -25380 393034 -25324
rect 393120 -25380 393176 -25324
rect 392978 -25522 393034 -25466
rect 393120 -25522 393176 -25466
rect 393383 -13736 393439 -13680
rect 393525 -13736 393581 -13680
rect 393383 -13878 393439 -13822
rect 393525 -13878 393581 -13822
rect 393383 -14020 393439 -13964
rect 393525 -14020 393581 -13964
rect 393383 -14162 393439 -14106
rect 393525 -14162 393581 -14106
rect 393383 -14304 393439 -14248
rect 393525 -14304 393581 -14248
rect 393383 -14446 393439 -14390
rect 393525 -14446 393581 -14390
rect 393383 -14588 393439 -14532
rect 393525 -14588 393581 -14532
rect 393383 -14730 393439 -14674
rect 393525 -14730 393581 -14674
rect 393383 -14872 393439 -14816
rect 393525 -14872 393581 -14816
rect 393383 -15014 393439 -14958
rect 393525 -15014 393581 -14958
rect 393383 -15156 393439 -15100
rect 393525 -15156 393581 -15100
rect 393383 -15298 393439 -15242
rect 393525 -15298 393581 -15242
rect 393383 -15440 393439 -15384
rect 393525 -15440 393581 -15384
rect 393383 -15582 393439 -15526
rect 393525 -15582 393581 -15526
rect 393383 -15724 393439 -15668
rect 393525 -15724 393581 -15668
rect 393383 -15866 393439 -15810
rect 393525 -15866 393581 -15810
rect 393383 -16008 393439 -15952
rect 393525 -16008 393581 -15952
rect 393383 -16150 393439 -16094
rect 393525 -16150 393581 -16094
rect 393383 -16292 393439 -16236
rect 393525 -16292 393581 -16236
rect 393383 -16434 393439 -16378
rect 393525 -16434 393581 -16378
rect 393383 -16576 393439 -16520
rect 393525 -16576 393581 -16520
rect 393383 -16718 393439 -16662
rect 393525 -16718 393581 -16662
rect 393383 -16860 393439 -16804
rect 393525 -16860 393581 -16804
rect 393383 -17002 393439 -16946
rect 393525 -17002 393581 -16946
rect 393383 -17144 393439 -17088
rect 393525 -17144 393581 -17088
rect 393383 -17286 393439 -17230
rect 393525 -17286 393581 -17230
rect 393383 -17428 393439 -17372
rect 393525 -17428 393581 -17372
rect 393383 -17570 393439 -17514
rect 393525 -17570 393581 -17514
rect 393383 -17712 393439 -17656
rect 393525 -17712 393581 -17656
rect 393383 -17854 393439 -17798
rect 393525 -17854 393581 -17798
rect 393383 -17996 393439 -17940
rect 393525 -17996 393581 -17940
rect 393383 -18138 393439 -18082
rect 393525 -18138 393581 -18082
rect 393383 -18280 393439 -18224
rect 393525 -18280 393581 -18224
rect 393383 -18422 393439 -18366
rect 393525 -18422 393581 -18366
rect 393383 -18564 393439 -18508
rect 393525 -18564 393581 -18508
rect 393383 -18706 393439 -18650
rect 393525 -18706 393581 -18650
rect 393383 -18848 393439 -18792
rect 393525 -18848 393581 -18792
rect 393383 -18990 393439 -18934
rect 393525 -18990 393581 -18934
rect 393383 -19132 393439 -19076
rect 393525 -19132 393581 -19076
rect 393383 -19274 393439 -19218
rect 393525 -19274 393581 -19218
rect 393383 -19416 393439 -19360
rect 393525 -19416 393581 -19360
rect 393383 -19558 393439 -19502
rect 393525 -19558 393581 -19502
rect 393383 -19700 393439 -19644
rect 393525 -19700 393581 -19644
rect 393383 -19842 393439 -19786
rect 393525 -19842 393581 -19786
rect 393383 -19984 393439 -19928
rect 393525 -19984 393581 -19928
rect 393383 -20126 393439 -20070
rect 393525 -20126 393581 -20070
rect 393383 -20268 393439 -20212
rect 393525 -20268 393581 -20212
rect 393383 -20410 393439 -20354
rect 393525 -20410 393581 -20354
rect 393383 -20552 393439 -20496
rect 393525 -20552 393581 -20496
rect 393383 -20694 393439 -20638
rect 393525 -20694 393581 -20638
rect 393383 -20836 393439 -20780
rect 393525 -20836 393581 -20780
rect 393383 -20978 393439 -20922
rect 393525 -20978 393581 -20922
rect 393383 -21120 393439 -21064
rect 393525 -21120 393581 -21064
rect 393383 -21262 393439 -21206
rect 393525 -21262 393581 -21206
rect 393383 -21404 393439 -21348
rect 393525 -21404 393581 -21348
rect 393383 -21546 393439 -21490
rect 393525 -21546 393581 -21490
rect 393383 -21688 393439 -21632
rect 393525 -21688 393581 -21632
rect 393383 -21830 393439 -21774
rect 393525 -21830 393581 -21774
rect 393383 -21972 393439 -21916
rect 393525 -21972 393581 -21916
rect 393383 -22114 393439 -22058
rect 393525 -22114 393581 -22058
rect 393383 -22256 393439 -22200
rect 393525 -22256 393581 -22200
rect 393383 -22398 393439 -22342
rect 393525 -22398 393581 -22342
rect 393383 -22540 393439 -22484
rect 393525 -22540 393581 -22484
rect 393383 -22682 393439 -22626
rect 393525 -22682 393581 -22626
rect 393383 -22824 393439 -22768
rect 393525 -22824 393581 -22768
rect 393383 -22966 393439 -22910
rect 393525 -22966 393581 -22910
rect 393383 -23108 393439 -23052
rect 393525 -23108 393581 -23052
rect 393383 -23250 393439 -23194
rect 393525 -23250 393581 -23194
rect 393383 -23392 393439 -23336
rect 393525 -23392 393581 -23336
rect 393383 -23534 393439 -23478
rect 393525 -23534 393581 -23478
rect 393383 -23676 393439 -23620
rect 393525 -23676 393581 -23620
rect 393383 -23818 393439 -23762
rect 393525 -23818 393581 -23762
rect 393383 -23960 393439 -23904
rect 393525 -23960 393581 -23904
rect 393383 -24102 393439 -24046
rect 393525 -24102 393581 -24046
rect 393383 -24244 393439 -24188
rect 393525 -24244 393581 -24188
rect 393383 -24386 393439 -24330
rect 393525 -24386 393581 -24330
rect 393383 -24528 393439 -24472
rect 393525 -24528 393581 -24472
rect 393383 -24670 393439 -24614
rect 393525 -24670 393581 -24614
rect 393383 -24812 393439 -24756
rect 393525 -24812 393581 -24756
rect 393383 -24954 393439 -24898
rect 393525 -24954 393581 -24898
rect 393383 -25096 393439 -25040
rect 393525 -25096 393581 -25040
rect 393383 -25238 393439 -25182
rect 393525 -25238 393581 -25182
rect 393383 -25380 393439 -25324
rect 393525 -25380 393581 -25324
rect 393383 -25522 393439 -25466
rect 393525 -25522 393581 -25466
rect 393780 -13736 393836 -13680
rect 393922 -13736 393978 -13680
rect 393780 -13878 393836 -13822
rect 393922 -13878 393978 -13822
rect 393780 -14020 393836 -13964
rect 393922 -14020 393978 -13964
rect 393780 -14162 393836 -14106
rect 393922 -14162 393978 -14106
rect 393780 -14304 393836 -14248
rect 393922 -14304 393978 -14248
rect 393780 -14446 393836 -14390
rect 393922 -14446 393978 -14390
rect 393780 -14588 393836 -14532
rect 393922 -14588 393978 -14532
rect 393780 -14730 393836 -14674
rect 393922 -14730 393978 -14674
rect 393780 -14872 393836 -14816
rect 393922 -14872 393978 -14816
rect 393780 -15014 393836 -14958
rect 393922 -15014 393978 -14958
rect 393780 -15156 393836 -15100
rect 393922 -15156 393978 -15100
rect 393780 -15298 393836 -15242
rect 393922 -15298 393978 -15242
rect 393780 -15440 393836 -15384
rect 393922 -15440 393978 -15384
rect 393780 -15582 393836 -15526
rect 393922 -15582 393978 -15526
rect 393780 -15724 393836 -15668
rect 393922 -15724 393978 -15668
rect 393780 -15866 393836 -15810
rect 393922 -15866 393978 -15810
rect 393780 -16008 393836 -15952
rect 393922 -16008 393978 -15952
rect 393780 -16150 393836 -16094
rect 393922 -16150 393978 -16094
rect 393780 -16292 393836 -16236
rect 393922 -16292 393978 -16236
rect 393780 -16434 393836 -16378
rect 393922 -16434 393978 -16378
rect 393780 -16576 393836 -16520
rect 393922 -16576 393978 -16520
rect 393780 -16718 393836 -16662
rect 393922 -16718 393978 -16662
rect 393780 -16860 393836 -16804
rect 393922 -16860 393978 -16804
rect 393780 -17002 393836 -16946
rect 393922 -17002 393978 -16946
rect 393780 -17144 393836 -17088
rect 393922 -17144 393978 -17088
rect 393780 -17286 393836 -17230
rect 393922 -17286 393978 -17230
rect 393780 -17428 393836 -17372
rect 393922 -17428 393978 -17372
rect 393780 -17570 393836 -17514
rect 393922 -17570 393978 -17514
rect 393780 -17712 393836 -17656
rect 393922 -17712 393978 -17656
rect 393780 -17854 393836 -17798
rect 393922 -17854 393978 -17798
rect 393780 -17996 393836 -17940
rect 393922 -17996 393978 -17940
rect 393780 -18138 393836 -18082
rect 393922 -18138 393978 -18082
rect 393780 -18280 393836 -18224
rect 393922 -18280 393978 -18224
rect 393780 -18422 393836 -18366
rect 393922 -18422 393978 -18366
rect 393780 -18564 393836 -18508
rect 393922 -18564 393978 -18508
rect 393780 -18706 393836 -18650
rect 393922 -18706 393978 -18650
rect 393780 -18848 393836 -18792
rect 393922 -18848 393978 -18792
rect 393780 -18990 393836 -18934
rect 393922 -18990 393978 -18934
rect 393780 -19132 393836 -19076
rect 393922 -19132 393978 -19076
rect 393780 -19274 393836 -19218
rect 393922 -19274 393978 -19218
rect 393780 -19416 393836 -19360
rect 393922 -19416 393978 -19360
rect 393780 -19558 393836 -19502
rect 393922 -19558 393978 -19502
rect 393780 -19700 393836 -19644
rect 393922 -19700 393978 -19644
rect 393780 -19842 393836 -19786
rect 393922 -19842 393978 -19786
rect 393780 -19984 393836 -19928
rect 393922 -19984 393978 -19928
rect 393780 -20126 393836 -20070
rect 393922 -20126 393978 -20070
rect 393780 -20268 393836 -20212
rect 393922 -20268 393978 -20212
rect 393780 -20410 393836 -20354
rect 393922 -20410 393978 -20354
rect 393780 -20552 393836 -20496
rect 393922 -20552 393978 -20496
rect 393780 -20694 393836 -20638
rect 393922 -20694 393978 -20638
rect 393780 -20836 393836 -20780
rect 393922 -20836 393978 -20780
rect 393780 -20978 393836 -20922
rect 393922 -20978 393978 -20922
rect 393780 -21120 393836 -21064
rect 393922 -21120 393978 -21064
rect 393780 -21262 393836 -21206
rect 393922 -21262 393978 -21206
rect 393780 -21404 393836 -21348
rect 393922 -21404 393978 -21348
rect 393780 -21546 393836 -21490
rect 393922 -21546 393978 -21490
rect 393780 -21688 393836 -21632
rect 393922 -21688 393978 -21632
rect 393780 -21830 393836 -21774
rect 393922 -21830 393978 -21774
rect 393780 -21972 393836 -21916
rect 393922 -21972 393978 -21916
rect 393780 -22114 393836 -22058
rect 393922 -22114 393978 -22058
rect 393780 -22256 393836 -22200
rect 393922 -22256 393978 -22200
rect 393780 -22398 393836 -22342
rect 393922 -22398 393978 -22342
rect 393780 -22540 393836 -22484
rect 393922 -22540 393978 -22484
rect 393780 -22682 393836 -22626
rect 393922 -22682 393978 -22626
rect 393780 -22824 393836 -22768
rect 393922 -22824 393978 -22768
rect 393780 -22966 393836 -22910
rect 393922 -22966 393978 -22910
rect 393780 -23108 393836 -23052
rect 393922 -23108 393978 -23052
rect 393780 -23250 393836 -23194
rect 393922 -23250 393978 -23194
rect 393780 -23392 393836 -23336
rect 393922 -23392 393978 -23336
rect 393780 -23534 393836 -23478
rect 393922 -23534 393978 -23478
rect 393780 -23676 393836 -23620
rect 393922 -23676 393978 -23620
rect 393780 -23818 393836 -23762
rect 393922 -23818 393978 -23762
rect 393780 -23960 393836 -23904
rect 393922 -23960 393978 -23904
rect 393780 -24102 393836 -24046
rect 393922 -24102 393978 -24046
rect 393780 -24244 393836 -24188
rect 393922 -24244 393978 -24188
rect 393780 -24386 393836 -24330
rect 393922 -24386 393978 -24330
rect 393780 -24528 393836 -24472
rect 393922 -24528 393978 -24472
rect 393780 -24670 393836 -24614
rect 393922 -24670 393978 -24614
rect 393780 -24812 393836 -24756
rect 393922 -24812 393978 -24756
rect 393780 -24954 393836 -24898
rect 393922 -24954 393978 -24898
rect 393780 -25096 393836 -25040
rect 393922 -25096 393978 -25040
rect 393780 -25238 393836 -25182
rect 393922 -25238 393978 -25182
rect 393780 -25380 393836 -25324
rect 393922 -25380 393978 -25324
rect 393780 -25522 393836 -25466
rect 393922 -25522 393978 -25466
rect 394177 -13736 394233 -13680
rect 394319 -13736 394375 -13680
rect 394177 -13878 394233 -13822
rect 394319 -13878 394375 -13822
rect 394177 -14020 394233 -13964
rect 394319 -14020 394375 -13964
rect 394177 -14162 394233 -14106
rect 394319 -14162 394375 -14106
rect 394177 -14304 394233 -14248
rect 394319 -14304 394375 -14248
rect 394177 -14446 394233 -14390
rect 394319 -14446 394375 -14390
rect 394177 -14588 394233 -14532
rect 394319 -14588 394375 -14532
rect 394177 -14730 394233 -14674
rect 394319 -14730 394375 -14674
rect 394177 -14872 394233 -14816
rect 394319 -14872 394375 -14816
rect 394177 -15014 394233 -14958
rect 394319 -15014 394375 -14958
rect 394177 -15156 394233 -15100
rect 394319 -15156 394375 -15100
rect 394177 -15298 394233 -15242
rect 394319 -15298 394375 -15242
rect 394177 -15440 394233 -15384
rect 394319 -15440 394375 -15384
rect 394177 -15582 394233 -15526
rect 394319 -15582 394375 -15526
rect 394177 -15724 394233 -15668
rect 394319 -15724 394375 -15668
rect 394177 -15866 394233 -15810
rect 394319 -15866 394375 -15810
rect 394177 -16008 394233 -15952
rect 394319 -16008 394375 -15952
rect 394177 -16150 394233 -16094
rect 394319 -16150 394375 -16094
rect 394177 -16292 394233 -16236
rect 394319 -16292 394375 -16236
rect 394177 -16434 394233 -16378
rect 394319 -16434 394375 -16378
rect 394177 -16576 394233 -16520
rect 394319 -16576 394375 -16520
rect 394177 -16718 394233 -16662
rect 394319 -16718 394375 -16662
rect 394177 -16860 394233 -16804
rect 394319 -16860 394375 -16804
rect 394177 -17002 394233 -16946
rect 394319 -17002 394375 -16946
rect 394177 -17144 394233 -17088
rect 394319 -17144 394375 -17088
rect 394177 -17286 394233 -17230
rect 394319 -17286 394375 -17230
rect 394177 -17428 394233 -17372
rect 394319 -17428 394375 -17372
rect 394177 -17570 394233 -17514
rect 394319 -17570 394375 -17514
rect 394177 -17712 394233 -17656
rect 394319 -17712 394375 -17656
rect 394177 -17854 394233 -17798
rect 394319 -17854 394375 -17798
rect 394177 -17996 394233 -17940
rect 394319 -17996 394375 -17940
rect 394177 -18138 394233 -18082
rect 394319 -18138 394375 -18082
rect 394177 -18280 394233 -18224
rect 394319 -18280 394375 -18224
rect 394177 -18422 394233 -18366
rect 394319 -18422 394375 -18366
rect 394177 -18564 394233 -18508
rect 394319 -18564 394375 -18508
rect 394177 -18706 394233 -18650
rect 394319 -18706 394375 -18650
rect 394177 -18848 394233 -18792
rect 394319 -18848 394375 -18792
rect 394177 -18990 394233 -18934
rect 394319 -18990 394375 -18934
rect 394177 -19132 394233 -19076
rect 394319 -19132 394375 -19076
rect 394177 -19274 394233 -19218
rect 394319 -19274 394375 -19218
rect 394177 -19416 394233 -19360
rect 394319 -19416 394375 -19360
rect 394177 -19558 394233 -19502
rect 394319 -19558 394375 -19502
rect 394177 -19700 394233 -19644
rect 394319 -19700 394375 -19644
rect 394177 -19842 394233 -19786
rect 394319 -19842 394375 -19786
rect 394177 -19984 394233 -19928
rect 394319 -19984 394375 -19928
rect 394177 -20126 394233 -20070
rect 394319 -20126 394375 -20070
rect 394177 -20268 394233 -20212
rect 394319 -20268 394375 -20212
rect 394177 -20410 394233 -20354
rect 394319 -20410 394375 -20354
rect 394177 -20552 394233 -20496
rect 394319 -20552 394375 -20496
rect 394177 -20694 394233 -20638
rect 394319 -20694 394375 -20638
rect 394177 -20836 394233 -20780
rect 394319 -20836 394375 -20780
rect 394177 -20978 394233 -20922
rect 394319 -20978 394375 -20922
rect 394177 -21120 394233 -21064
rect 394319 -21120 394375 -21064
rect 394177 -21262 394233 -21206
rect 394319 -21262 394375 -21206
rect 394177 -21404 394233 -21348
rect 394319 -21404 394375 -21348
rect 394177 -21546 394233 -21490
rect 394319 -21546 394375 -21490
rect 394177 -21688 394233 -21632
rect 394319 -21688 394375 -21632
rect 394177 -21830 394233 -21774
rect 394319 -21830 394375 -21774
rect 394177 -21972 394233 -21916
rect 394319 -21972 394375 -21916
rect 394177 -22114 394233 -22058
rect 394319 -22114 394375 -22058
rect 394177 -22256 394233 -22200
rect 394319 -22256 394375 -22200
rect 394177 -22398 394233 -22342
rect 394319 -22398 394375 -22342
rect 394177 -22540 394233 -22484
rect 394319 -22540 394375 -22484
rect 394177 -22682 394233 -22626
rect 394319 -22682 394375 -22626
rect 394177 -22824 394233 -22768
rect 394319 -22824 394375 -22768
rect 394177 -22966 394233 -22910
rect 394319 -22966 394375 -22910
rect 394177 -23108 394233 -23052
rect 394319 -23108 394375 -23052
rect 394177 -23250 394233 -23194
rect 394319 -23250 394375 -23194
rect 394177 -23392 394233 -23336
rect 394319 -23392 394375 -23336
rect 394177 -23534 394233 -23478
rect 394319 -23534 394375 -23478
rect 394177 -23676 394233 -23620
rect 394319 -23676 394375 -23620
rect 394177 -23818 394233 -23762
rect 394319 -23818 394375 -23762
rect 394177 -23960 394233 -23904
rect 394319 -23960 394375 -23904
rect 394177 -24102 394233 -24046
rect 394319 -24102 394375 -24046
rect 394177 -24244 394233 -24188
rect 394319 -24244 394375 -24188
rect 394177 -24386 394233 -24330
rect 394319 -24386 394375 -24330
rect 394177 -24528 394233 -24472
rect 394319 -24528 394375 -24472
rect 394177 -24670 394233 -24614
rect 394319 -24670 394375 -24614
rect 394177 -24812 394233 -24756
rect 394319 -24812 394375 -24756
rect 394177 -24954 394233 -24898
rect 394319 -24954 394375 -24898
rect 394177 -25096 394233 -25040
rect 394319 -25096 394375 -25040
rect 394177 -25238 394233 -25182
rect 394319 -25238 394375 -25182
rect 394177 -25380 394233 -25324
rect 394319 -25380 394375 -25324
rect 394177 -25522 394233 -25466
rect 394319 -25522 394375 -25466
rect 394580 -13736 394636 -13680
rect 394722 -13736 394778 -13680
rect 394580 -13878 394636 -13822
rect 394722 -13878 394778 -13822
rect 394580 -14020 394636 -13964
rect 394722 -14020 394778 -13964
rect 394580 -14162 394636 -14106
rect 394722 -14162 394778 -14106
rect 394580 -14304 394636 -14248
rect 394722 -14304 394778 -14248
rect 394580 -14446 394636 -14390
rect 394722 -14446 394778 -14390
rect 394580 -14588 394636 -14532
rect 394722 -14588 394778 -14532
rect 394580 -14730 394636 -14674
rect 394722 -14730 394778 -14674
rect 394580 -14872 394636 -14816
rect 394722 -14872 394778 -14816
rect 394580 -15014 394636 -14958
rect 394722 -15014 394778 -14958
rect 394580 -15156 394636 -15100
rect 394722 -15156 394778 -15100
rect 394580 -15298 394636 -15242
rect 394722 -15298 394778 -15242
rect 394580 -15440 394636 -15384
rect 394722 -15440 394778 -15384
rect 394580 -15582 394636 -15526
rect 394722 -15582 394778 -15526
rect 394580 -15724 394636 -15668
rect 394722 -15724 394778 -15668
rect 394580 -15866 394636 -15810
rect 394722 -15866 394778 -15810
rect 394580 -16008 394636 -15952
rect 394722 -16008 394778 -15952
rect 394580 -16150 394636 -16094
rect 394722 -16150 394778 -16094
rect 394580 -16292 394636 -16236
rect 394722 -16292 394778 -16236
rect 394580 -16434 394636 -16378
rect 394722 -16434 394778 -16378
rect 394580 -16576 394636 -16520
rect 394722 -16576 394778 -16520
rect 394580 -16718 394636 -16662
rect 394722 -16718 394778 -16662
rect 394580 -16860 394636 -16804
rect 394722 -16860 394778 -16804
rect 394580 -17002 394636 -16946
rect 394722 -17002 394778 -16946
rect 394580 -17144 394636 -17088
rect 394722 -17144 394778 -17088
rect 394580 -17286 394636 -17230
rect 394722 -17286 394778 -17230
rect 394580 -17428 394636 -17372
rect 394722 -17428 394778 -17372
rect 394580 -17570 394636 -17514
rect 394722 -17570 394778 -17514
rect 394580 -17712 394636 -17656
rect 394722 -17712 394778 -17656
rect 394580 -17854 394636 -17798
rect 394722 -17854 394778 -17798
rect 394580 -17996 394636 -17940
rect 394722 -17996 394778 -17940
rect 394580 -18138 394636 -18082
rect 394722 -18138 394778 -18082
rect 394580 -18280 394636 -18224
rect 394722 -18280 394778 -18224
rect 394580 -18422 394636 -18366
rect 394722 -18422 394778 -18366
rect 394580 -18564 394636 -18508
rect 394722 -18564 394778 -18508
rect 394580 -18706 394636 -18650
rect 394722 -18706 394778 -18650
rect 394580 -18848 394636 -18792
rect 394722 -18848 394778 -18792
rect 394580 -18990 394636 -18934
rect 394722 -18990 394778 -18934
rect 394580 -19132 394636 -19076
rect 394722 -19132 394778 -19076
rect 394580 -19274 394636 -19218
rect 394722 -19274 394778 -19218
rect 394580 -19416 394636 -19360
rect 394722 -19416 394778 -19360
rect 394580 -19558 394636 -19502
rect 394722 -19558 394778 -19502
rect 394580 -19700 394636 -19644
rect 394722 -19700 394778 -19644
rect 394580 -19842 394636 -19786
rect 394722 -19842 394778 -19786
rect 394580 -19984 394636 -19928
rect 394722 -19984 394778 -19928
rect 394580 -20126 394636 -20070
rect 394722 -20126 394778 -20070
rect 394580 -20268 394636 -20212
rect 394722 -20268 394778 -20212
rect 394580 -20410 394636 -20354
rect 394722 -20410 394778 -20354
rect 394580 -20552 394636 -20496
rect 394722 -20552 394778 -20496
rect 394580 -20694 394636 -20638
rect 394722 -20694 394778 -20638
rect 394580 -20836 394636 -20780
rect 394722 -20836 394778 -20780
rect 394580 -20978 394636 -20922
rect 394722 -20978 394778 -20922
rect 394580 -21120 394636 -21064
rect 394722 -21120 394778 -21064
rect 394580 -21262 394636 -21206
rect 394722 -21262 394778 -21206
rect 394580 -21404 394636 -21348
rect 394722 -21404 394778 -21348
rect 394580 -21546 394636 -21490
rect 394722 -21546 394778 -21490
rect 394580 -21688 394636 -21632
rect 394722 -21688 394778 -21632
rect 394580 -21830 394636 -21774
rect 394722 -21830 394778 -21774
rect 394580 -21972 394636 -21916
rect 394722 -21972 394778 -21916
rect 394580 -22114 394636 -22058
rect 394722 -22114 394778 -22058
rect 394580 -22256 394636 -22200
rect 394722 -22256 394778 -22200
rect 394580 -22398 394636 -22342
rect 394722 -22398 394778 -22342
rect 394580 -22540 394636 -22484
rect 394722 -22540 394778 -22484
rect 394580 -22682 394636 -22626
rect 394722 -22682 394778 -22626
rect 394580 -22824 394636 -22768
rect 394722 -22824 394778 -22768
rect 394580 -22966 394636 -22910
rect 394722 -22966 394778 -22910
rect 394580 -23108 394636 -23052
rect 394722 -23108 394778 -23052
rect 394580 -23250 394636 -23194
rect 394722 -23250 394778 -23194
rect 394580 -23392 394636 -23336
rect 394722 -23392 394778 -23336
rect 394580 -23534 394636 -23478
rect 394722 -23534 394778 -23478
rect 394580 -23676 394636 -23620
rect 394722 -23676 394778 -23620
rect 394580 -23818 394636 -23762
rect 394722 -23818 394778 -23762
rect 394580 -23960 394636 -23904
rect 394722 -23960 394778 -23904
rect 394580 -24102 394636 -24046
rect 394722 -24102 394778 -24046
rect 394580 -24244 394636 -24188
rect 394722 -24244 394778 -24188
rect 394580 -24386 394636 -24330
rect 394722 -24386 394778 -24330
rect 394580 -24528 394636 -24472
rect 394722 -24528 394778 -24472
rect 394580 -24670 394636 -24614
rect 394722 -24670 394778 -24614
rect 394580 -24812 394636 -24756
rect 394722 -24812 394778 -24756
rect 394580 -24954 394636 -24898
rect 394722 -24954 394778 -24898
rect 394580 -25096 394636 -25040
rect 394722 -25096 394778 -25040
rect 394580 -25238 394636 -25182
rect 394722 -25238 394778 -25182
rect 394580 -25380 394636 -25324
rect 394722 -25380 394778 -25324
rect 394580 -25522 394636 -25466
rect 394722 -25522 394778 -25466
rect 394982 -13736 395038 -13680
rect 395124 -13736 395180 -13680
rect 394982 -13878 395038 -13822
rect 395124 -13878 395180 -13822
rect 394982 -14020 395038 -13964
rect 395124 -14020 395180 -13964
rect 394982 -14162 395038 -14106
rect 395124 -14162 395180 -14106
rect 394982 -14304 395038 -14248
rect 395124 -14304 395180 -14248
rect 394982 -14446 395038 -14390
rect 395124 -14446 395180 -14390
rect 394982 -14588 395038 -14532
rect 395124 -14588 395180 -14532
rect 394982 -14730 395038 -14674
rect 395124 -14730 395180 -14674
rect 394982 -14872 395038 -14816
rect 395124 -14872 395180 -14816
rect 394982 -15014 395038 -14958
rect 395124 -15014 395180 -14958
rect 394982 -15156 395038 -15100
rect 395124 -15156 395180 -15100
rect 394982 -15298 395038 -15242
rect 395124 -15298 395180 -15242
rect 394982 -15440 395038 -15384
rect 395124 -15440 395180 -15384
rect 394982 -15582 395038 -15526
rect 395124 -15582 395180 -15526
rect 394982 -15724 395038 -15668
rect 395124 -15724 395180 -15668
rect 394982 -15866 395038 -15810
rect 395124 -15866 395180 -15810
rect 394982 -16008 395038 -15952
rect 395124 -16008 395180 -15952
rect 394982 -16150 395038 -16094
rect 395124 -16150 395180 -16094
rect 394982 -16292 395038 -16236
rect 395124 -16292 395180 -16236
rect 394982 -16434 395038 -16378
rect 395124 -16434 395180 -16378
rect 394982 -16576 395038 -16520
rect 395124 -16576 395180 -16520
rect 394982 -16718 395038 -16662
rect 395124 -16718 395180 -16662
rect 394982 -16860 395038 -16804
rect 395124 -16860 395180 -16804
rect 394982 -17002 395038 -16946
rect 395124 -17002 395180 -16946
rect 394982 -17144 395038 -17088
rect 395124 -17144 395180 -17088
rect 394982 -17286 395038 -17230
rect 395124 -17286 395180 -17230
rect 394982 -17428 395038 -17372
rect 395124 -17428 395180 -17372
rect 394982 -17570 395038 -17514
rect 395124 -17570 395180 -17514
rect 394982 -17712 395038 -17656
rect 395124 -17712 395180 -17656
rect 394982 -17854 395038 -17798
rect 395124 -17854 395180 -17798
rect 394982 -17996 395038 -17940
rect 395124 -17996 395180 -17940
rect 394982 -18138 395038 -18082
rect 395124 -18138 395180 -18082
rect 394982 -18280 395038 -18224
rect 395124 -18280 395180 -18224
rect 394982 -18422 395038 -18366
rect 395124 -18422 395180 -18366
rect 394982 -18564 395038 -18508
rect 395124 -18564 395180 -18508
rect 394982 -18706 395038 -18650
rect 395124 -18706 395180 -18650
rect 394982 -18848 395038 -18792
rect 395124 -18848 395180 -18792
rect 394982 -18990 395038 -18934
rect 395124 -18990 395180 -18934
rect 394982 -19132 395038 -19076
rect 395124 -19132 395180 -19076
rect 394982 -19274 395038 -19218
rect 395124 -19274 395180 -19218
rect 394982 -19416 395038 -19360
rect 395124 -19416 395180 -19360
rect 394982 -19558 395038 -19502
rect 395124 -19558 395180 -19502
rect 394982 -19700 395038 -19644
rect 395124 -19700 395180 -19644
rect 394982 -19842 395038 -19786
rect 395124 -19842 395180 -19786
rect 394982 -19984 395038 -19928
rect 395124 -19984 395180 -19928
rect 394982 -20126 395038 -20070
rect 395124 -20126 395180 -20070
rect 394982 -20268 395038 -20212
rect 395124 -20268 395180 -20212
rect 394982 -20410 395038 -20354
rect 395124 -20410 395180 -20354
rect 394982 -20552 395038 -20496
rect 395124 -20552 395180 -20496
rect 394982 -20694 395038 -20638
rect 395124 -20694 395180 -20638
rect 394982 -20836 395038 -20780
rect 395124 -20836 395180 -20780
rect 394982 -20978 395038 -20922
rect 395124 -20978 395180 -20922
rect 394982 -21120 395038 -21064
rect 395124 -21120 395180 -21064
rect 394982 -21262 395038 -21206
rect 395124 -21262 395180 -21206
rect 394982 -21404 395038 -21348
rect 395124 -21404 395180 -21348
rect 394982 -21546 395038 -21490
rect 395124 -21546 395180 -21490
rect 394982 -21688 395038 -21632
rect 395124 -21688 395180 -21632
rect 394982 -21830 395038 -21774
rect 395124 -21830 395180 -21774
rect 394982 -21972 395038 -21916
rect 395124 -21972 395180 -21916
rect 394982 -22114 395038 -22058
rect 395124 -22114 395180 -22058
rect 394982 -22256 395038 -22200
rect 395124 -22256 395180 -22200
rect 394982 -22398 395038 -22342
rect 395124 -22398 395180 -22342
rect 394982 -22540 395038 -22484
rect 395124 -22540 395180 -22484
rect 394982 -22682 395038 -22626
rect 395124 -22682 395180 -22626
rect 394982 -22824 395038 -22768
rect 395124 -22824 395180 -22768
rect 394982 -22966 395038 -22910
rect 395124 -22966 395180 -22910
rect 394982 -23108 395038 -23052
rect 395124 -23108 395180 -23052
rect 394982 -23250 395038 -23194
rect 395124 -23250 395180 -23194
rect 394982 -23392 395038 -23336
rect 395124 -23392 395180 -23336
rect 394982 -23534 395038 -23478
rect 395124 -23534 395180 -23478
rect 394982 -23676 395038 -23620
rect 395124 -23676 395180 -23620
rect 394982 -23818 395038 -23762
rect 395124 -23818 395180 -23762
rect 394982 -23960 395038 -23904
rect 395124 -23960 395180 -23904
rect 394982 -24102 395038 -24046
rect 395124 -24102 395180 -24046
rect 394982 -24244 395038 -24188
rect 395124 -24244 395180 -24188
rect 394982 -24386 395038 -24330
rect 395124 -24386 395180 -24330
rect 394982 -24528 395038 -24472
rect 395124 -24528 395180 -24472
rect 394982 -24670 395038 -24614
rect 395124 -24670 395180 -24614
rect 394982 -24812 395038 -24756
rect 395124 -24812 395180 -24756
rect 394982 -24954 395038 -24898
rect 395124 -24954 395180 -24898
rect 394982 -25096 395038 -25040
rect 395124 -25096 395180 -25040
rect 394982 -25238 395038 -25182
rect 395124 -25238 395180 -25182
rect 394982 -25380 395038 -25324
rect 395124 -25380 395180 -25324
rect 394982 -25522 395038 -25466
rect 395124 -25522 395180 -25466
rect 395385 -13736 395441 -13680
rect 395527 -13736 395583 -13680
rect 395385 -13878 395441 -13822
rect 395527 -13878 395583 -13822
rect 395385 -14020 395441 -13964
rect 395527 -14020 395583 -13964
rect 395385 -14162 395441 -14106
rect 395527 -14162 395583 -14106
rect 395385 -14304 395441 -14248
rect 395527 -14304 395583 -14248
rect 395385 -14446 395441 -14390
rect 395527 -14446 395583 -14390
rect 395385 -14588 395441 -14532
rect 395527 -14588 395583 -14532
rect 395385 -14730 395441 -14674
rect 395527 -14730 395583 -14674
rect 395385 -14872 395441 -14816
rect 395527 -14872 395583 -14816
rect 395385 -15014 395441 -14958
rect 395527 -15014 395583 -14958
rect 395385 -15156 395441 -15100
rect 395527 -15156 395583 -15100
rect 395385 -15298 395441 -15242
rect 395527 -15298 395583 -15242
rect 395385 -15440 395441 -15384
rect 395527 -15440 395583 -15384
rect 395385 -15582 395441 -15526
rect 395527 -15582 395583 -15526
rect 395385 -15724 395441 -15668
rect 395527 -15724 395583 -15668
rect 395385 -15866 395441 -15810
rect 395527 -15866 395583 -15810
rect 395385 -16008 395441 -15952
rect 395527 -16008 395583 -15952
rect 395385 -16150 395441 -16094
rect 395527 -16150 395583 -16094
rect 395385 -16292 395441 -16236
rect 395527 -16292 395583 -16236
rect 395385 -16434 395441 -16378
rect 395527 -16434 395583 -16378
rect 395385 -16576 395441 -16520
rect 395527 -16576 395583 -16520
rect 395385 -16718 395441 -16662
rect 395527 -16718 395583 -16662
rect 395385 -16860 395441 -16804
rect 395527 -16860 395583 -16804
rect 395385 -17002 395441 -16946
rect 395527 -17002 395583 -16946
rect 395385 -17144 395441 -17088
rect 395527 -17144 395583 -17088
rect 395385 -17286 395441 -17230
rect 395527 -17286 395583 -17230
rect 395385 -17428 395441 -17372
rect 395527 -17428 395583 -17372
rect 395385 -17570 395441 -17514
rect 395527 -17570 395583 -17514
rect 395385 -17712 395441 -17656
rect 395527 -17712 395583 -17656
rect 395385 -17854 395441 -17798
rect 395527 -17854 395583 -17798
rect 395385 -17996 395441 -17940
rect 395527 -17996 395583 -17940
rect 395385 -18138 395441 -18082
rect 395527 -18138 395583 -18082
rect 395385 -18280 395441 -18224
rect 395527 -18280 395583 -18224
rect 395385 -18422 395441 -18366
rect 395527 -18422 395583 -18366
rect 395385 -18564 395441 -18508
rect 395527 -18564 395583 -18508
rect 395385 -18706 395441 -18650
rect 395527 -18706 395583 -18650
rect 395385 -18848 395441 -18792
rect 395527 -18848 395583 -18792
rect 395385 -18990 395441 -18934
rect 395527 -18990 395583 -18934
rect 395385 -19132 395441 -19076
rect 395527 -19132 395583 -19076
rect 395385 -19274 395441 -19218
rect 395527 -19274 395583 -19218
rect 395385 -19416 395441 -19360
rect 395527 -19416 395583 -19360
rect 395385 -19558 395441 -19502
rect 395527 -19558 395583 -19502
rect 395385 -19700 395441 -19644
rect 395527 -19700 395583 -19644
rect 395385 -19842 395441 -19786
rect 395527 -19842 395583 -19786
rect 395385 -19984 395441 -19928
rect 395527 -19984 395583 -19928
rect 395385 -20126 395441 -20070
rect 395527 -20126 395583 -20070
rect 395385 -20268 395441 -20212
rect 395527 -20268 395583 -20212
rect 395385 -20410 395441 -20354
rect 395527 -20410 395583 -20354
rect 395385 -20552 395441 -20496
rect 395527 -20552 395583 -20496
rect 395385 -20694 395441 -20638
rect 395527 -20694 395583 -20638
rect 395385 -20836 395441 -20780
rect 395527 -20836 395583 -20780
rect 395385 -20978 395441 -20922
rect 395527 -20978 395583 -20922
rect 395385 -21120 395441 -21064
rect 395527 -21120 395583 -21064
rect 395385 -21262 395441 -21206
rect 395527 -21262 395583 -21206
rect 395385 -21404 395441 -21348
rect 395527 -21404 395583 -21348
rect 395385 -21546 395441 -21490
rect 395527 -21546 395583 -21490
rect 395385 -21688 395441 -21632
rect 395527 -21688 395583 -21632
rect 395385 -21830 395441 -21774
rect 395527 -21830 395583 -21774
rect 395385 -21972 395441 -21916
rect 395527 -21972 395583 -21916
rect 395385 -22114 395441 -22058
rect 395527 -22114 395583 -22058
rect 395385 -22256 395441 -22200
rect 395527 -22256 395583 -22200
rect 395385 -22398 395441 -22342
rect 395527 -22398 395583 -22342
rect 395385 -22540 395441 -22484
rect 395527 -22540 395583 -22484
rect 395385 -22682 395441 -22626
rect 395527 -22682 395583 -22626
rect 395385 -22824 395441 -22768
rect 395527 -22824 395583 -22768
rect 395385 -22966 395441 -22910
rect 395527 -22966 395583 -22910
rect 395385 -23108 395441 -23052
rect 395527 -23108 395583 -23052
rect 395385 -23250 395441 -23194
rect 395527 -23250 395583 -23194
rect 395385 -23392 395441 -23336
rect 395527 -23392 395583 -23336
rect 395385 -23534 395441 -23478
rect 395527 -23534 395583 -23478
rect 395385 -23676 395441 -23620
rect 395527 -23676 395583 -23620
rect 395385 -23818 395441 -23762
rect 395527 -23818 395583 -23762
rect 395385 -23960 395441 -23904
rect 395527 -23960 395583 -23904
rect 395385 -24102 395441 -24046
rect 395527 -24102 395583 -24046
rect 395385 -24244 395441 -24188
rect 395527 -24244 395583 -24188
rect 395385 -24386 395441 -24330
rect 395527 -24386 395583 -24330
rect 395385 -24528 395441 -24472
rect 395527 -24528 395583 -24472
rect 395385 -24670 395441 -24614
rect 395527 -24670 395583 -24614
rect 395385 -24812 395441 -24756
rect 395527 -24812 395583 -24756
rect 395385 -24954 395441 -24898
rect 395527 -24954 395583 -24898
rect 395385 -25096 395441 -25040
rect 395527 -25096 395583 -25040
rect 395385 -25238 395441 -25182
rect 395527 -25238 395583 -25182
rect 395385 -25380 395441 -25324
rect 395527 -25380 395583 -25324
rect 395385 -25522 395441 -25466
rect 395527 -25522 395583 -25466
rect 395779 -13736 395835 -13680
rect 395921 -13736 395977 -13680
rect 395779 -13878 395835 -13822
rect 395921 -13878 395977 -13822
rect 395779 -14020 395835 -13964
rect 395921 -14020 395977 -13964
rect 395779 -14162 395835 -14106
rect 395921 -14162 395977 -14106
rect 395779 -14304 395835 -14248
rect 395921 -14304 395977 -14248
rect 395779 -14446 395835 -14390
rect 395921 -14446 395977 -14390
rect 395779 -14588 395835 -14532
rect 395921 -14588 395977 -14532
rect 395779 -14730 395835 -14674
rect 395921 -14730 395977 -14674
rect 395779 -14872 395835 -14816
rect 395921 -14872 395977 -14816
rect 395779 -15014 395835 -14958
rect 395921 -15014 395977 -14958
rect 395779 -15156 395835 -15100
rect 395921 -15156 395977 -15100
rect 395779 -15298 395835 -15242
rect 395921 -15298 395977 -15242
rect 395779 -15440 395835 -15384
rect 395921 -15440 395977 -15384
rect 395779 -15582 395835 -15526
rect 395921 -15582 395977 -15526
rect 395779 -15724 395835 -15668
rect 395921 -15724 395977 -15668
rect 395779 -15866 395835 -15810
rect 395921 -15866 395977 -15810
rect 395779 -16008 395835 -15952
rect 395921 -16008 395977 -15952
rect 395779 -16150 395835 -16094
rect 395921 -16150 395977 -16094
rect 395779 -16292 395835 -16236
rect 395921 -16292 395977 -16236
rect 395779 -16434 395835 -16378
rect 395921 -16434 395977 -16378
rect 395779 -16576 395835 -16520
rect 395921 -16576 395977 -16520
rect 395779 -16718 395835 -16662
rect 395921 -16718 395977 -16662
rect 395779 -16860 395835 -16804
rect 395921 -16860 395977 -16804
rect 395779 -17002 395835 -16946
rect 395921 -17002 395977 -16946
rect 395779 -17144 395835 -17088
rect 395921 -17144 395977 -17088
rect 395779 -17286 395835 -17230
rect 395921 -17286 395977 -17230
rect 395779 -17428 395835 -17372
rect 395921 -17428 395977 -17372
rect 395779 -17570 395835 -17514
rect 395921 -17570 395977 -17514
rect 395779 -17712 395835 -17656
rect 395921 -17712 395977 -17656
rect 395779 -17854 395835 -17798
rect 395921 -17854 395977 -17798
rect 395779 -17996 395835 -17940
rect 395921 -17996 395977 -17940
rect 395779 -18138 395835 -18082
rect 395921 -18138 395977 -18082
rect 395779 -18280 395835 -18224
rect 395921 -18280 395977 -18224
rect 395779 -18422 395835 -18366
rect 395921 -18422 395977 -18366
rect 395779 -18564 395835 -18508
rect 395921 -18564 395977 -18508
rect 395779 -18706 395835 -18650
rect 395921 -18706 395977 -18650
rect 395779 -18848 395835 -18792
rect 395921 -18848 395977 -18792
rect 395779 -18990 395835 -18934
rect 395921 -18990 395977 -18934
rect 395779 -19132 395835 -19076
rect 395921 -19132 395977 -19076
rect 395779 -19274 395835 -19218
rect 395921 -19274 395977 -19218
rect 395779 -19416 395835 -19360
rect 395921 -19416 395977 -19360
rect 395779 -19558 395835 -19502
rect 395921 -19558 395977 -19502
rect 395779 -19700 395835 -19644
rect 395921 -19700 395977 -19644
rect 395779 -19842 395835 -19786
rect 395921 -19842 395977 -19786
rect 395779 -19984 395835 -19928
rect 395921 -19984 395977 -19928
rect 395779 -20126 395835 -20070
rect 395921 -20126 395977 -20070
rect 395779 -20268 395835 -20212
rect 395921 -20268 395977 -20212
rect 395779 -20410 395835 -20354
rect 395921 -20410 395977 -20354
rect 395779 -20552 395835 -20496
rect 395921 -20552 395977 -20496
rect 395779 -20694 395835 -20638
rect 395921 -20694 395977 -20638
rect 395779 -20836 395835 -20780
rect 395921 -20836 395977 -20780
rect 395779 -20978 395835 -20922
rect 395921 -20978 395977 -20922
rect 395779 -21120 395835 -21064
rect 395921 -21120 395977 -21064
rect 395779 -21262 395835 -21206
rect 395921 -21262 395977 -21206
rect 395779 -21404 395835 -21348
rect 395921 -21404 395977 -21348
rect 395779 -21546 395835 -21490
rect 395921 -21546 395977 -21490
rect 395779 -21688 395835 -21632
rect 395921 -21688 395977 -21632
rect 395779 -21830 395835 -21774
rect 395921 -21830 395977 -21774
rect 395779 -21972 395835 -21916
rect 395921 -21972 395977 -21916
rect 395779 -22114 395835 -22058
rect 395921 -22114 395977 -22058
rect 395779 -22256 395835 -22200
rect 395921 -22256 395977 -22200
rect 395779 -22398 395835 -22342
rect 395921 -22398 395977 -22342
rect 395779 -22540 395835 -22484
rect 395921 -22540 395977 -22484
rect 395779 -22682 395835 -22626
rect 395921 -22682 395977 -22626
rect 395779 -22824 395835 -22768
rect 395921 -22824 395977 -22768
rect 395779 -22966 395835 -22910
rect 395921 -22966 395977 -22910
rect 395779 -23108 395835 -23052
rect 395921 -23108 395977 -23052
rect 395779 -23250 395835 -23194
rect 395921 -23250 395977 -23194
rect 395779 -23392 395835 -23336
rect 395921 -23392 395977 -23336
rect 395779 -23534 395835 -23478
rect 395921 -23534 395977 -23478
rect 395779 -23676 395835 -23620
rect 395921 -23676 395977 -23620
rect 395779 -23818 395835 -23762
rect 395921 -23818 395977 -23762
rect 395779 -23960 395835 -23904
rect 395921 -23960 395977 -23904
rect 395779 -24102 395835 -24046
rect 395921 -24102 395977 -24046
rect 395779 -24244 395835 -24188
rect 395921 -24244 395977 -24188
rect 395779 -24386 395835 -24330
rect 395921 -24386 395977 -24330
rect 395779 -24528 395835 -24472
rect 395921 -24528 395977 -24472
rect 395779 -24670 395835 -24614
rect 395921 -24670 395977 -24614
rect 395779 -24812 395835 -24756
rect 395921 -24812 395977 -24756
rect 395779 -24954 395835 -24898
rect 395921 -24954 395977 -24898
rect 395779 -25096 395835 -25040
rect 395921 -25096 395977 -25040
rect 395779 -25238 395835 -25182
rect 395921 -25238 395977 -25182
rect 395779 -25380 395835 -25324
rect 395921 -25380 395977 -25324
rect 395779 -25522 395835 -25466
rect 395921 -25522 395977 -25466
rect 396180 -13736 396236 -13680
rect 396322 -13736 396378 -13680
rect 396180 -13878 396236 -13822
rect 396322 -13878 396378 -13822
rect 396180 -14020 396236 -13964
rect 396322 -14020 396378 -13964
rect 396180 -14162 396236 -14106
rect 396322 -14162 396378 -14106
rect 396180 -14304 396236 -14248
rect 396322 -14304 396378 -14248
rect 396180 -14446 396236 -14390
rect 396322 -14446 396378 -14390
rect 396180 -14588 396236 -14532
rect 396322 -14588 396378 -14532
rect 396180 -14730 396236 -14674
rect 396322 -14730 396378 -14674
rect 396180 -14872 396236 -14816
rect 396322 -14872 396378 -14816
rect 396180 -15014 396236 -14958
rect 396322 -15014 396378 -14958
rect 396180 -15156 396236 -15100
rect 396322 -15156 396378 -15100
rect 396180 -15298 396236 -15242
rect 396322 -15298 396378 -15242
rect 396180 -15440 396236 -15384
rect 396322 -15440 396378 -15384
rect 396180 -15582 396236 -15526
rect 396322 -15582 396378 -15526
rect 396180 -15724 396236 -15668
rect 396322 -15724 396378 -15668
rect 396180 -15866 396236 -15810
rect 396322 -15866 396378 -15810
rect 396180 -16008 396236 -15952
rect 396322 -16008 396378 -15952
rect 396180 -16150 396236 -16094
rect 396322 -16150 396378 -16094
rect 396180 -16292 396236 -16236
rect 396322 -16292 396378 -16236
rect 396180 -16434 396236 -16378
rect 396322 -16434 396378 -16378
rect 396180 -16576 396236 -16520
rect 396322 -16576 396378 -16520
rect 396180 -16718 396236 -16662
rect 396322 -16718 396378 -16662
rect 396180 -16860 396236 -16804
rect 396322 -16860 396378 -16804
rect 396180 -17002 396236 -16946
rect 396322 -17002 396378 -16946
rect 396180 -17144 396236 -17088
rect 396322 -17144 396378 -17088
rect 396180 -17286 396236 -17230
rect 396322 -17286 396378 -17230
rect 396180 -17428 396236 -17372
rect 396322 -17428 396378 -17372
rect 396180 -17570 396236 -17514
rect 396322 -17570 396378 -17514
rect 396180 -17712 396236 -17656
rect 396322 -17712 396378 -17656
rect 396180 -17854 396236 -17798
rect 396322 -17854 396378 -17798
rect 396180 -17996 396236 -17940
rect 396322 -17996 396378 -17940
rect 396180 -18138 396236 -18082
rect 396322 -18138 396378 -18082
rect 396180 -18280 396236 -18224
rect 396322 -18280 396378 -18224
rect 396180 -18422 396236 -18366
rect 396322 -18422 396378 -18366
rect 396180 -18564 396236 -18508
rect 396322 -18564 396378 -18508
rect 396180 -18706 396236 -18650
rect 396322 -18706 396378 -18650
rect 396180 -18848 396236 -18792
rect 396322 -18848 396378 -18792
rect 396180 -18990 396236 -18934
rect 396322 -18990 396378 -18934
rect 396180 -19132 396236 -19076
rect 396322 -19132 396378 -19076
rect 396180 -19274 396236 -19218
rect 396322 -19274 396378 -19218
rect 396180 -19416 396236 -19360
rect 396322 -19416 396378 -19360
rect 396180 -19558 396236 -19502
rect 396322 -19558 396378 -19502
rect 396180 -19700 396236 -19644
rect 396322 -19700 396378 -19644
rect 396180 -19842 396236 -19786
rect 396322 -19842 396378 -19786
rect 396180 -19984 396236 -19928
rect 396322 -19984 396378 -19928
rect 396180 -20126 396236 -20070
rect 396322 -20126 396378 -20070
rect 396180 -20268 396236 -20212
rect 396322 -20268 396378 -20212
rect 396180 -20410 396236 -20354
rect 396322 -20410 396378 -20354
rect 396180 -20552 396236 -20496
rect 396322 -20552 396378 -20496
rect 396180 -20694 396236 -20638
rect 396322 -20694 396378 -20638
rect 396180 -20836 396236 -20780
rect 396322 -20836 396378 -20780
rect 396180 -20978 396236 -20922
rect 396322 -20978 396378 -20922
rect 396180 -21120 396236 -21064
rect 396322 -21120 396378 -21064
rect 396180 -21262 396236 -21206
rect 396322 -21262 396378 -21206
rect 396180 -21404 396236 -21348
rect 396322 -21404 396378 -21348
rect 396180 -21546 396236 -21490
rect 396322 -21546 396378 -21490
rect 396180 -21688 396236 -21632
rect 396322 -21688 396378 -21632
rect 396180 -21830 396236 -21774
rect 396322 -21830 396378 -21774
rect 396180 -21972 396236 -21916
rect 396322 -21972 396378 -21916
rect 396180 -22114 396236 -22058
rect 396322 -22114 396378 -22058
rect 396180 -22256 396236 -22200
rect 396322 -22256 396378 -22200
rect 396180 -22398 396236 -22342
rect 396322 -22398 396378 -22342
rect 396180 -22540 396236 -22484
rect 396322 -22540 396378 -22484
rect 396180 -22682 396236 -22626
rect 396322 -22682 396378 -22626
rect 396180 -22824 396236 -22768
rect 396322 -22824 396378 -22768
rect 396180 -22966 396236 -22910
rect 396322 -22966 396378 -22910
rect 396180 -23108 396236 -23052
rect 396322 -23108 396378 -23052
rect 396180 -23250 396236 -23194
rect 396322 -23250 396378 -23194
rect 396180 -23392 396236 -23336
rect 396322 -23392 396378 -23336
rect 396180 -23534 396236 -23478
rect 396322 -23534 396378 -23478
rect 396180 -23676 396236 -23620
rect 396322 -23676 396378 -23620
rect 396180 -23818 396236 -23762
rect 396322 -23818 396378 -23762
rect 396180 -23960 396236 -23904
rect 396322 -23960 396378 -23904
rect 396180 -24102 396236 -24046
rect 396322 -24102 396378 -24046
rect 396180 -24244 396236 -24188
rect 396322 -24244 396378 -24188
rect 396180 -24386 396236 -24330
rect 396322 -24386 396378 -24330
rect 396180 -24528 396236 -24472
rect 396322 -24528 396378 -24472
rect 396180 -24670 396236 -24614
rect 396322 -24670 396378 -24614
rect 396180 -24812 396236 -24756
rect 396322 -24812 396378 -24756
rect 396180 -24954 396236 -24898
rect 396322 -24954 396378 -24898
rect 396180 -25096 396236 -25040
rect 396322 -25096 396378 -25040
rect 396180 -25238 396236 -25182
rect 396322 -25238 396378 -25182
rect 396180 -25380 396236 -25324
rect 396322 -25380 396378 -25324
rect 396180 -25522 396236 -25466
rect 396322 -25522 396378 -25466
rect 396580 -13736 396636 -13680
rect 396722 -13736 396778 -13680
rect 396580 -13878 396636 -13822
rect 396722 -13878 396778 -13822
rect 396580 -14020 396636 -13964
rect 396722 -14020 396778 -13964
rect 396580 -14162 396636 -14106
rect 396722 -14162 396778 -14106
rect 396580 -14304 396636 -14248
rect 396722 -14304 396778 -14248
rect 396580 -14446 396636 -14390
rect 396722 -14446 396778 -14390
rect 396580 -14588 396636 -14532
rect 396722 -14588 396778 -14532
rect 396580 -14730 396636 -14674
rect 396722 -14730 396778 -14674
rect 396580 -14872 396636 -14816
rect 396722 -14872 396778 -14816
rect 396580 -15014 396636 -14958
rect 396722 -15014 396778 -14958
rect 396580 -15156 396636 -15100
rect 396722 -15156 396778 -15100
rect 396580 -15298 396636 -15242
rect 396722 -15298 396778 -15242
rect 396580 -15440 396636 -15384
rect 396722 -15440 396778 -15384
rect 396580 -15582 396636 -15526
rect 396722 -15582 396778 -15526
rect 396580 -15724 396636 -15668
rect 396722 -15724 396778 -15668
rect 396580 -15866 396636 -15810
rect 396722 -15866 396778 -15810
rect 396580 -16008 396636 -15952
rect 396722 -16008 396778 -15952
rect 396580 -16150 396636 -16094
rect 396722 -16150 396778 -16094
rect 396580 -16292 396636 -16236
rect 396722 -16292 396778 -16236
rect 396580 -16434 396636 -16378
rect 396722 -16434 396778 -16378
rect 396580 -16576 396636 -16520
rect 396722 -16576 396778 -16520
rect 396580 -16718 396636 -16662
rect 396722 -16718 396778 -16662
rect 396580 -16860 396636 -16804
rect 396722 -16860 396778 -16804
rect 396580 -17002 396636 -16946
rect 396722 -17002 396778 -16946
rect 396580 -17144 396636 -17088
rect 396722 -17144 396778 -17088
rect 396580 -17286 396636 -17230
rect 396722 -17286 396778 -17230
rect 396580 -17428 396636 -17372
rect 396722 -17428 396778 -17372
rect 396580 -17570 396636 -17514
rect 396722 -17570 396778 -17514
rect 396580 -17712 396636 -17656
rect 396722 -17712 396778 -17656
rect 396580 -17854 396636 -17798
rect 396722 -17854 396778 -17798
rect 396580 -17996 396636 -17940
rect 396722 -17996 396778 -17940
rect 396580 -18138 396636 -18082
rect 396722 -18138 396778 -18082
rect 396580 -18280 396636 -18224
rect 396722 -18280 396778 -18224
rect 396580 -18422 396636 -18366
rect 396722 -18422 396778 -18366
rect 396580 -18564 396636 -18508
rect 396722 -18564 396778 -18508
rect 396580 -18706 396636 -18650
rect 396722 -18706 396778 -18650
rect 396580 -18848 396636 -18792
rect 396722 -18848 396778 -18792
rect 396580 -18990 396636 -18934
rect 396722 -18990 396778 -18934
rect 396580 -19132 396636 -19076
rect 396722 -19132 396778 -19076
rect 396580 -19274 396636 -19218
rect 396722 -19274 396778 -19218
rect 396580 -19416 396636 -19360
rect 396722 -19416 396778 -19360
rect 396580 -19558 396636 -19502
rect 396722 -19558 396778 -19502
rect 396580 -19700 396636 -19644
rect 396722 -19700 396778 -19644
rect 396580 -19842 396636 -19786
rect 396722 -19842 396778 -19786
rect 396580 -19984 396636 -19928
rect 396722 -19984 396778 -19928
rect 396580 -20126 396636 -20070
rect 396722 -20126 396778 -20070
rect 396580 -20268 396636 -20212
rect 396722 -20268 396778 -20212
rect 396580 -20410 396636 -20354
rect 396722 -20410 396778 -20354
rect 396580 -20552 396636 -20496
rect 396722 -20552 396778 -20496
rect 396580 -20694 396636 -20638
rect 396722 -20694 396778 -20638
rect 396580 -20836 396636 -20780
rect 396722 -20836 396778 -20780
rect 396580 -20978 396636 -20922
rect 396722 -20978 396778 -20922
rect 396580 -21120 396636 -21064
rect 396722 -21120 396778 -21064
rect 396580 -21262 396636 -21206
rect 396722 -21262 396778 -21206
rect 396580 -21404 396636 -21348
rect 396722 -21404 396778 -21348
rect 396580 -21546 396636 -21490
rect 396722 -21546 396778 -21490
rect 396580 -21688 396636 -21632
rect 396722 -21688 396778 -21632
rect 396580 -21830 396636 -21774
rect 396722 -21830 396778 -21774
rect 396580 -21972 396636 -21916
rect 396722 -21972 396778 -21916
rect 396580 -22114 396636 -22058
rect 396722 -22114 396778 -22058
rect 396580 -22256 396636 -22200
rect 396722 -22256 396778 -22200
rect 396580 -22398 396636 -22342
rect 396722 -22398 396778 -22342
rect 396580 -22540 396636 -22484
rect 396722 -22540 396778 -22484
rect 396580 -22682 396636 -22626
rect 396722 -22682 396778 -22626
rect 396580 -22824 396636 -22768
rect 396722 -22824 396778 -22768
rect 396580 -22966 396636 -22910
rect 396722 -22966 396778 -22910
rect 396580 -23108 396636 -23052
rect 396722 -23108 396778 -23052
rect 396580 -23250 396636 -23194
rect 396722 -23250 396778 -23194
rect 396580 -23392 396636 -23336
rect 396722 -23392 396778 -23336
rect 396580 -23534 396636 -23478
rect 396722 -23534 396778 -23478
rect 396580 -23676 396636 -23620
rect 396722 -23676 396778 -23620
rect 396580 -23818 396636 -23762
rect 396722 -23818 396778 -23762
rect 396580 -23960 396636 -23904
rect 396722 -23960 396778 -23904
rect 396580 -24102 396636 -24046
rect 396722 -24102 396778 -24046
rect 396580 -24244 396636 -24188
rect 396722 -24244 396778 -24188
rect 396580 -24386 396636 -24330
rect 396722 -24386 396778 -24330
rect 396580 -24528 396636 -24472
rect 396722 -24528 396778 -24472
rect 396580 -24670 396636 -24614
rect 396722 -24670 396778 -24614
rect 396580 -24812 396636 -24756
rect 396722 -24812 396778 -24756
rect 396580 -24954 396636 -24898
rect 396722 -24954 396778 -24898
rect 396580 -25096 396636 -25040
rect 396722 -25096 396778 -25040
rect 396580 -25238 396636 -25182
rect 396722 -25238 396778 -25182
rect 396580 -25380 396636 -25324
rect 396722 -25380 396778 -25324
rect 396580 -25522 396636 -25466
rect 396722 -25522 396778 -25466
rect 396977 -13736 397033 -13680
rect 397119 -13736 397175 -13680
rect 396977 -13878 397033 -13822
rect 397119 -13878 397175 -13822
rect 396977 -14020 397033 -13964
rect 397119 -14020 397175 -13964
rect 396977 -14162 397033 -14106
rect 397119 -14162 397175 -14106
rect 396977 -14304 397033 -14248
rect 397119 -14304 397175 -14248
rect 396977 -14446 397033 -14390
rect 397119 -14446 397175 -14390
rect 396977 -14588 397033 -14532
rect 397119 -14588 397175 -14532
rect 396977 -14730 397033 -14674
rect 397119 -14730 397175 -14674
rect 396977 -14872 397033 -14816
rect 397119 -14872 397175 -14816
rect 396977 -15014 397033 -14958
rect 397119 -15014 397175 -14958
rect 396977 -15156 397033 -15100
rect 397119 -15156 397175 -15100
rect 396977 -15298 397033 -15242
rect 397119 -15298 397175 -15242
rect 396977 -15440 397033 -15384
rect 397119 -15440 397175 -15384
rect 396977 -15582 397033 -15526
rect 397119 -15582 397175 -15526
rect 396977 -15724 397033 -15668
rect 397119 -15724 397175 -15668
rect 396977 -15866 397033 -15810
rect 397119 -15866 397175 -15810
rect 396977 -16008 397033 -15952
rect 397119 -16008 397175 -15952
rect 396977 -16150 397033 -16094
rect 397119 -16150 397175 -16094
rect 396977 -16292 397033 -16236
rect 397119 -16292 397175 -16236
rect 396977 -16434 397033 -16378
rect 397119 -16434 397175 -16378
rect 396977 -16576 397033 -16520
rect 397119 -16576 397175 -16520
rect 396977 -16718 397033 -16662
rect 397119 -16718 397175 -16662
rect 396977 -16860 397033 -16804
rect 397119 -16860 397175 -16804
rect 396977 -17002 397033 -16946
rect 397119 -17002 397175 -16946
rect 396977 -17144 397033 -17088
rect 397119 -17144 397175 -17088
rect 396977 -17286 397033 -17230
rect 397119 -17286 397175 -17230
rect 396977 -17428 397033 -17372
rect 397119 -17428 397175 -17372
rect 396977 -17570 397033 -17514
rect 397119 -17570 397175 -17514
rect 396977 -17712 397033 -17656
rect 397119 -17712 397175 -17656
rect 396977 -17854 397033 -17798
rect 397119 -17854 397175 -17798
rect 396977 -17996 397033 -17940
rect 397119 -17996 397175 -17940
rect 396977 -18138 397033 -18082
rect 397119 -18138 397175 -18082
rect 396977 -18280 397033 -18224
rect 397119 -18280 397175 -18224
rect 396977 -18422 397033 -18366
rect 397119 -18422 397175 -18366
rect 396977 -18564 397033 -18508
rect 397119 -18564 397175 -18508
rect 396977 -18706 397033 -18650
rect 397119 -18706 397175 -18650
rect 396977 -18848 397033 -18792
rect 397119 -18848 397175 -18792
rect 396977 -18990 397033 -18934
rect 397119 -18990 397175 -18934
rect 396977 -19132 397033 -19076
rect 397119 -19132 397175 -19076
rect 396977 -19274 397033 -19218
rect 397119 -19274 397175 -19218
rect 396977 -19416 397033 -19360
rect 397119 -19416 397175 -19360
rect 396977 -19558 397033 -19502
rect 397119 -19558 397175 -19502
rect 396977 -19700 397033 -19644
rect 397119 -19700 397175 -19644
rect 396977 -19842 397033 -19786
rect 397119 -19842 397175 -19786
rect 396977 -19984 397033 -19928
rect 397119 -19984 397175 -19928
rect 396977 -20126 397033 -20070
rect 397119 -20126 397175 -20070
rect 396977 -20268 397033 -20212
rect 397119 -20268 397175 -20212
rect 396977 -20410 397033 -20354
rect 397119 -20410 397175 -20354
rect 396977 -20552 397033 -20496
rect 397119 -20552 397175 -20496
rect 396977 -20694 397033 -20638
rect 397119 -20694 397175 -20638
rect 396977 -20836 397033 -20780
rect 397119 -20836 397175 -20780
rect 396977 -20978 397033 -20922
rect 397119 -20978 397175 -20922
rect 396977 -21120 397033 -21064
rect 397119 -21120 397175 -21064
rect 396977 -21262 397033 -21206
rect 397119 -21262 397175 -21206
rect 396977 -21404 397033 -21348
rect 397119 -21404 397175 -21348
rect 396977 -21546 397033 -21490
rect 397119 -21546 397175 -21490
rect 396977 -21688 397033 -21632
rect 397119 -21688 397175 -21632
rect 396977 -21830 397033 -21774
rect 397119 -21830 397175 -21774
rect 396977 -21972 397033 -21916
rect 397119 -21972 397175 -21916
rect 396977 -22114 397033 -22058
rect 397119 -22114 397175 -22058
rect 396977 -22256 397033 -22200
rect 397119 -22256 397175 -22200
rect 396977 -22398 397033 -22342
rect 397119 -22398 397175 -22342
rect 396977 -22540 397033 -22484
rect 397119 -22540 397175 -22484
rect 396977 -22682 397033 -22626
rect 397119 -22682 397175 -22626
rect 396977 -22824 397033 -22768
rect 397119 -22824 397175 -22768
rect 396977 -22966 397033 -22910
rect 397119 -22966 397175 -22910
rect 396977 -23108 397033 -23052
rect 397119 -23108 397175 -23052
rect 396977 -23250 397033 -23194
rect 397119 -23250 397175 -23194
rect 396977 -23392 397033 -23336
rect 397119 -23392 397175 -23336
rect 396977 -23534 397033 -23478
rect 397119 -23534 397175 -23478
rect 396977 -23676 397033 -23620
rect 397119 -23676 397175 -23620
rect 396977 -23818 397033 -23762
rect 397119 -23818 397175 -23762
rect 396977 -23960 397033 -23904
rect 397119 -23960 397175 -23904
rect 396977 -24102 397033 -24046
rect 397119 -24102 397175 -24046
rect 396977 -24244 397033 -24188
rect 397119 -24244 397175 -24188
rect 396977 -24386 397033 -24330
rect 397119 -24386 397175 -24330
rect 396977 -24528 397033 -24472
rect 397119 -24528 397175 -24472
rect 396977 -24670 397033 -24614
rect 397119 -24670 397175 -24614
rect 396977 -24812 397033 -24756
rect 397119 -24812 397175 -24756
rect 396977 -24954 397033 -24898
rect 397119 -24954 397175 -24898
rect 396977 -25096 397033 -25040
rect 397119 -25096 397175 -25040
rect 396977 -25238 397033 -25182
rect 397119 -25238 397175 -25182
rect 396977 -25380 397033 -25324
rect 397119 -25380 397175 -25324
rect 396977 -25522 397033 -25466
rect 397119 -25522 397175 -25466
rect 397374 -13736 397430 -13680
rect 397516 -13736 397572 -13680
rect 397374 -13878 397430 -13822
rect 397516 -13878 397572 -13822
rect 397374 -14020 397430 -13964
rect 397516 -14020 397572 -13964
rect 397374 -14162 397430 -14106
rect 397516 -14162 397572 -14106
rect 397374 -14304 397430 -14248
rect 397516 -14304 397572 -14248
rect 397374 -14446 397430 -14390
rect 397516 -14446 397572 -14390
rect 397374 -14588 397430 -14532
rect 397516 -14588 397572 -14532
rect 397374 -14730 397430 -14674
rect 397516 -14730 397572 -14674
rect 397374 -14872 397430 -14816
rect 397516 -14872 397572 -14816
rect 397374 -15014 397430 -14958
rect 397516 -15014 397572 -14958
rect 397374 -15156 397430 -15100
rect 397516 -15156 397572 -15100
rect 397374 -15298 397430 -15242
rect 397516 -15298 397572 -15242
rect 397374 -15440 397430 -15384
rect 397516 -15440 397572 -15384
rect 397374 -15582 397430 -15526
rect 397516 -15582 397572 -15526
rect 397374 -15724 397430 -15668
rect 397516 -15724 397572 -15668
rect 397374 -15866 397430 -15810
rect 397516 -15866 397572 -15810
rect 397374 -16008 397430 -15952
rect 397516 -16008 397572 -15952
rect 397374 -16150 397430 -16094
rect 397516 -16150 397572 -16094
rect 397374 -16292 397430 -16236
rect 397516 -16292 397572 -16236
rect 397374 -16434 397430 -16378
rect 397516 -16434 397572 -16378
rect 397374 -16576 397430 -16520
rect 397516 -16576 397572 -16520
rect 397374 -16718 397430 -16662
rect 397516 -16718 397572 -16662
rect 397374 -16860 397430 -16804
rect 397516 -16860 397572 -16804
rect 397374 -17002 397430 -16946
rect 397516 -17002 397572 -16946
rect 397374 -17144 397430 -17088
rect 397516 -17144 397572 -17088
rect 397374 -17286 397430 -17230
rect 397516 -17286 397572 -17230
rect 397374 -17428 397430 -17372
rect 397516 -17428 397572 -17372
rect 397374 -17570 397430 -17514
rect 397516 -17570 397572 -17514
rect 397374 -17712 397430 -17656
rect 397516 -17712 397572 -17656
rect 397374 -17854 397430 -17798
rect 397516 -17854 397572 -17798
rect 397374 -17996 397430 -17940
rect 397516 -17996 397572 -17940
rect 397374 -18138 397430 -18082
rect 397516 -18138 397572 -18082
rect 397374 -18280 397430 -18224
rect 397516 -18280 397572 -18224
rect 397374 -18422 397430 -18366
rect 397516 -18422 397572 -18366
rect 397374 -18564 397430 -18508
rect 397516 -18564 397572 -18508
rect 397374 -18706 397430 -18650
rect 397516 -18706 397572 -18650
rect 397374 -18848 397430 -18792
rect 397516 -18848 397572 -18792
rect 397374 -18990 397430 -18934
rect 397516 -18990 397572 -18934
rect 397374 -19132 397430 -19076
rect 397516 -19132 397572 -19076
rect 397374 -19274 397430 -19218
rect 397516 -19274 397572 -19218
rect 397374 -19416 397430 -19360
rect 397516 -19416 397572 -19360
rect 397374 -19558 397430 -19502
rect 397516 -19558 397572 -19502
rect 397374 -19700 397430 -19644
rect 397516 -19700 397572 -19644
rect 397374 -19842 397430 -19786
rect 397516 -19842 397572 -19786
rect 397374 -19984 397430 -19928
rect 397516 -19984 397572 -19928
rect 397374 -20126 397430 -20070
rect 397516 -20126 397572 -20070
rect 397374 -20268 397430 -20212
rect 397516 -20268 397572 -20212
rect 397374 -20410 397430 -20354
rect 397516 -20410 397572 -20354
rect 397374 -20552 397430 -20496
rect 397516 -20552 397572 -20496
rect 397374 -20694 397430 -20638
rect 397516 -20694 397572 -20638
rect 397374 -20836 397430 -20780
rect 397516 -20836 397572 -20780
rect 397374 -20978 397430 -20922
rect 397516 -20978 397572 -20922
rect 397374 -21120 397430 -21064
rect 397516 -21120 397572 -21064
rect 397374 -21262 397430 -21206
rect 397516 -21262 397572 -21206
rect 397374 -21404 397430 -21348
rect 397516 -21404 397572 -21348
rect 397374 -21546 397430 -21490
rect 397516 -21546 397572 -21490
rect 397374 -21688 397430 -21632
rect 397516 -21688 397572 -21632
rect 397374 -21830 397430 -21774
rect 397516 -21830 397572 -21774
rect 397374 -21972 397430 -21916
rect 397516 -21972 397572 -21916
rect 397374 -22114 397430 -22058
rect 397516 -22114 397572 -22058
rect 397374 -22256 397430 -22200
rect 397516 -22256 397572 -22200
rect 397374 -22398 397430 -22342
rect 397516 -22398 397572 -22342
rect 397374 -22540 397430 -22484
rect 397516 -22540 397572 -22484
rect 397374 -22682 397430 -22626
rect 397516 -22682 397572 -22626
rect 397374 -22824 397430 -22768
rect 397516 -22824 397572 -22768
rect 397374 -22966 397430 -22910
rect 397516 -22966 397572 -22910
rect 397374 -23108 397430 -23052
rect 397516 -23108 397572 -23052
rect 397374 -23250 397430 -23194
rect 397516 -23250 397572 -23194
rect 397374 -23392 397430 -23336
rect 397516 -23392 397572 -23336
rect 397374 -23534 397430 -23478
rect 397516 -23534 397572 -23478
rect 397374 -23676 397430 -23620
rect 397516 -23676 397572 -23620
rect 397374 -23818 397430 -23762
rect 397516 -23818 397572 -23762
rect 397374 -23960 397430 -23904
rect 397516 -23960 397572 -23904
rect 397374 -24102 397430 -24046
rect 397516 -24102 397572 -24046
rect 397374 -24244 397430 -24188
rect 397516 -24244 397572 -24188
rect 397374 -24386 397430 -24330
rect 397516 -24386 397572 -24330
rect 397374 -24528 397430 -24472
rect 397516 -24528 397572 -24472
rect 397374 -24670 397430 -24614
rect 397516 -24670 397572 -24614
rect 397374 -24812 397430 -24756
rect 397516 -24812 397572 -24756
rect 397374 -24954 397430 -24898
rect 397516 -24954 397572 -24898
rect 397374 -25096 397430 -25040
rect 397516 -25096 397572 -25040
rect 397374 -25238 397430 -25182
rect 397516 -25238 397572 -25182
rect 397374 -25380 397430 -25324
rect 397516 -25380 397572 -25324
rect 397374 -25522 397430 -25466
rect 397516 -25522 397572 -25466
rect 397778 -13736 397834 -13680
rect 397920 -13736 397976 -13680
rect 397778 -13878 397834 -13822
rect 397920 -13878 397976 -13822
rect 397778 -14020 397834 -13964
rect 397920 -14020 397976 -13964
rect 397778 -14162 397834 -14106
rect 397920 -14162 397976 -14106
rect 397778 -14304 397834 -14248
rect 397920 -14304 397976 -14248
rect 397778 -14446 397834 -14390
rect 397920 -14446 397976 -14390
rect 397778 -14588 397834 -14532
rect 397920 -14588 397976 -14532
rect 397778 -14730 397834 -14674
rect 397920 -14730 397976 -14674
rect 397778 -14872 397834 -14816
rect 397920 -14872 397976 -14816
rect 397778 -15014 397834 -14958
rect 397920 -15014 397976 -14958
rect 397778 -15156 397834 -15100
rect 397920 -15156 397976 -15100
rect 397778 -15298 397834 -15242
rect 397920 -15298 397976 -15242
rect 397778 -15440 397834 -15384
rect 397920 -15440 397976 -15384
rect 397778 -15582 397834 -15526
rect 397920 -15582 397976 -15526
rect 397778 -15724 397834 -15668
rect 397920 -15724 397976 -15668
rect 397778 -15866 397834 -15810
rect 397920 -15866 397976 -15810
rect 397778 -16008 397834 -15952
rect 397920 -16008 397976 -15952
rect 397778 -16150 397834 -16094
rect 397920 -16150 397976 -16094
rect 397778 -16292 397834 -16236
rect 397920 -16292 397976 -16236
rect 397778 -16434 397834 -16378
rect 397920 -16434 397976 -16378
rect 397778 -16576 397834 -16520
rect 397920 -16576 397976 -16520
rect 397778 -16718 397834 -16662
rect 397920 -16718 397976 -16662
rect 397778 -16860 397834 -16804
rect 397920 -16860 397976 -16804
rect 397778 -17002 397834 -16946
rect 397920 -17002 397976 -16946
rect 397778 -17144 397834 -17088
rect 397920 -17144 397976 -17088
rect 397778 -17286 397834 -17230
rect 397920 -17286 397976 -17230
rect 397778 -17428 397834 -17372
rect 397920 -17428 397976 -17372
rect 397778 -17570 397834 -17514
rect 397920 -17570 397976 -17514
rect 397778 -17712 397834 -17656
rect 397920 -17712 397976 -17656
rect 397778 -17854 397834 -17798
rect 397920 -17854 397976 -17798
rect 397778 -17996 397834 -17940
rect 397920 -17996 397976 -17940
rect 397778 -18138 397834 -18082
rect 397920 -18138 397976 -18082
rect 397778 -18280 397834 -18224
rect 397920 -18280 397976 -18224
rect 397778 -18422 397834 -18366
rect 397920 -18422 397976 -18366
rect 397778 -18564 397834 -18508
rect 397920 -18564 397976 -18508
rect 397778 -18706 397834 -18650
rect 397920 -18706 397976 -18650
rect 397778 -18848 397834 -18792
rect 397920 -18848 397976 -18792
rect 397778 -18990 397834 -18934
rect 397920 -18990 397976 -18934
rect 397778 -19132 397834 -19076
rect 397920 -19132 397976 -19076
rect 397778 -19274 397834 -19218
rect 397920 -19274 397976 -19218
rect 397778 -19416 397834 -19360
rect 397920 -19416 397976 -19360
rect 397778 -19558 397834 -19502
rect 397920 -19558 397976 -19502
rect 397778 -19700 397834 -19644
rect 397920 -19700 397976 -19644
rect 397778 -19842 397834 -19786
rect 397920 -19842 397976 -19786
rect 397778 -19984 397834 -19928
rect 397920 -19984 397976 -19928
rect 397778 -20126 397834 -20070
rect 397920 -20126 397976 -20070
rect 397778 -20268 397834 -20212
rect 397920 -20268 397976 -20212
rect 397778 -20410 397834 -20354
rect 397920 -20410 397976 -20354
rect 397778 -20552 397834 -20496
rect 397920 -20552 397976 -20496
rect 397778 -20694 397834 -20638
rect 397920 -20694 397976 -20638
rect 397778 -20836 397834 -20780
rect 397920 -20836 397976 -20780
rect 397778 -20978 397834 -20922
rect 397920 -20978 397976 -20922
rect 397778 -21120 397834 -21064
rect 397920 -21120 397976 -21064
rect 397778 -21262 397834 -21206
rect 397920 -21262 397976 -21206
rect 397778 -21404 397834 -21348
rect 397920 -21404 397976 -21348
rect 397778 -21546 397834 -21490
rect 397920 -21546 397976 -21490
rect 397778 -21688 397834 -21632
rect 397920 -21688 397976 -21632
rect 397778 -21830 397834 -21774
rect 397920 -21830 397976 -21774
rect 397778 -21972 397834 -21916
rect 397920 -21972 397976 -21916
rect 397778 -22114 397834 -22058
rect 397920 -22114 397976 -22058
rect 397778 -22256 397834 -22200
rect 397920 -22256 397976 -22200
rect 397778 -22398 397834 -22342
rect 397920 -22398 397976 -22342
rect 397778 -22540 397834 -22484
rect 397920 -22540 397976 -22484
rect 397778 -22682 397834 -22626
rect 397920 -22682 397976 -22626
rect 397778 -22824 397834 -22768
rect 397920 -22824 397976 -22768
rect 397778 -22966 397834 -22910
rect 397920 -22966 397976 -22910
rect 397778 -23108 397834 -23052
rect 397920 -23108 397976 -23052
rect 397778 -23250 397834 -23194
rect 397920 -23250 397976 -23194
rect 397778 -23392 397834 -23336
rect 397920 -23392 397976 -23336
rect 397778 -23534 397834 -23478
rect 397920 -23534 397976 -23478
rect 397778 -23676 397834 -23620
rect 397920 -23676 397976 -23620
rect 397778 -23818 397834 -23762
rect 397920 -23818 397976 -23762
rect 397778 -23960 397834 -23904
rect 397920 -23960 397976 -23904
rect 397778 -24102 397834 -24046
rect 397920 -24102 397976 -24046
rect 397778 -24244 397834 -24188
rect 397920 -24244 397976 -24188
rect 397778 -24386 397834 -24330
rect 397920 -24386 397976 -24330
rect 397778 -24528 397834 -24472
rect 397920 -24528 397976 -24472
rect 397778 -24670 397834 -24614
rect 397920 -24670 397976 -24614
rect 397778 -24812 397834 -24756
rect 397920 -24812 397976 -24756
rect 397778 -24954 397834 -24898
rect 397920 -24954 397976 -24898
rect 397778 -25096 397834 -25040
rect 397920 -25096 397976 -25040
rect 397778 -25238 397834 -25182
rect 397920 -25238 397976 -25182
rect 397778 -25380 397834 -25324
rect 397920 -25380 397976 -25324
rect 397778 -25522 397834 -25466
rect 397920 -25522 397976 -25466
rect 398174 -13736 398230 -13680
rect 398316 -13736 398372 -13680
rect 398174 -13878 398230 -13822
rect 398316 -13878 398372 -13822
rect 398174 -14020 398230 -13964
rect 398316 -14020 398372 -13964
rect 398174 -14162 398230 -14106
rect 398316 -14162 398372 -14106
rect 398174 -14304 398230 -14248
rect 398316 -14304 398372 -14248
rect 398174 -14446 398230 -14390
rect 398316 -14446 398372 -14390
rect 398174 -14588 398230 -14532
rect 398316 -14588 398372 -14532
rect 398174 -14730 398230 -14674
rect 398316 -14730 398372 -14674
rect 398174 -14872 398230 -14816
rect 398316 -14872 398372 -14816
rect 398174 -15014 398230 -14958
rect 398316 -15014 398372 -14958
rect 398174 -15156 398230 -15100
rect 398316 -15156 398372 -15100
rect 398174 -15298 398230 -15242
rect 398316 -15298 398372 -15242
rect 398174 -15440 398230 -15384
rect 398316 -15440 398372 -15384
rect 398174 -15582 398230 -15526
rect 398316 -15582 398372 -15526
rect 398174 -15724 398230 -15668
rect 398316 -15724 398372 -15668
rect 398174 -15866 398230 -15810
rect 398316 -15866 398372 -15810
rect 398174 -16008 398230 -15952
rect 398316 -16008 398372 -15952
rect 398174 -16150 398230 -16094
rect 398316 -16150 398372 -16094
rect 398174 -16292 398230 -16236
rect 398316 -16292 398372 -16236
rect 398174 -16434 398230 -16378
rect 398316 -16434 398372 -16378
rect 398174 -16576 398230 -16520
rect 398316 -16576 398372 -16520
rect 398174 -16718 398230 -16662
rect 398316 -16718 398372 -16662
rect 398174 -16860 398230 -16804
rect 398316 -16860 398372 -16804
rect 398174 -17002 398230 -16946
rect 398316 -17002 398372 -16946
rect 398174 -17144 398230 -17088
rect 398316 -17144 398372 -17088
rect 398174 -17286 398230 -17230
rect 398316 -17286 398372 -17230
rect 398174 -17428 398230 -17372
rect 398316 -17428 398372 -17372
rect 398174 -17570 398230 -17514
rect 398316 -17570 398372 -17514
rect 398174 -17712 398230 -17656
rect 398316 -17712 398372 -17656
rect 398174 -17854 398230 -17798
rect 398316 -17854 398372 -17798
rect 398174 -17996 398230 -17940
rect 398316 -17996 398372 -17940
rect 398174 -18138 398230 -18082
rect 398316 -18138 398372 -18082
rect 398174 -18280 398230 -18224
rect 398316 -18280 398372 -18224
rect 398174 -18422 398230 -18366
rect 398316 -18422 398372 -18366
rect 398174 -18564 398230 -18508
rect 398316 -18564 398372 -18508
rect 398174 -18706 398230 -18650
rect 398316 -18706 398372 -18650
rect 398174 -18848 398230 -18792
rect 398316 -18848 398372 -18792
rect 398174 -18990 398230 -18934
rect 398316 -18990 398372 -18934
rect 398174 -19132 398230 -19076
rect 398316 -19132 398372 -19076
rect 398174 -19274 398230 -19218
rect 398316 -19274 398372 -19218
rect 398174 -19416 398230 -19360
rect 398316 -19416 398372 -19360
rect 398174 -19558 398230 -19502
rect 398316 -19558 398372 -19502
rect 398174 -19700 398230 -19644
rect 398316 -19700 398372 -19644
rect 398174 -19842 398230 -19786
rect 398316 -19842 398372 -19786
rect 398174 -19984 398230 -19928
rect 398316 -19984 398372 -19928
rect 398174 -20126 398230 -20070
rect 398316 -20126 398372 -20070
rect 398174 -20268 398230 -20212
rect 398316 -20268 398372 -20212
rect 398174 -20410 398230 -20354
rect 398316 -20410 398372 -20354
rect 398174 -20552 398230 -20496
rect 398316 -20552 398372 -20496
rect 398174 -20694 398230 -20638
rect 398316 -20694 398372 -20638
rect 398174 -20836 398230 -20780
rect 398316 -20836 398372 -20780
rect 398174 -20978 398230 -20922
rect 398316 -20978 398372 -20922
rect 398174 -21120 398230 -21064
rect 398316 -21120 398372 -21064
rect 398174 -21262 398230 -21206
rect 398316 -21262 398372 -21206
rect 398174 -21404 398230 -21348
rect 398316 -21404 398372 -21348
rect 398174 -21546 398230 -21490
rect 398316 -21546 398372 -21490
rect 398174 -21688 398230 -21632
rect 398316 -21688 398372 -21632
rect 398174 -21830 398230 -21774
rect 398316 -21830 398372 -21774
rect 398174 -21972 398230 -21916
rect 398316 -21972 398372 -21916
rect 398174 -22114 398230 -22058
rect 398316 -22114 398372 -22058
rect 398174 -22256 398230 -22200
rect 398316 -22256 398372 -22200
rect 398174 -22398 398230 -22342
rect 398316 -22398 398372 -22342
rect 398174 -22540 398230 -22484
rect 398316 -22540 398372 -22484
rect 398174 -22682 398230 -22626
rect 398316 -22682 398372 -22626
rect 398174 -22824 398230 -22768
rect 398316 -22824 398372 -22768
rect 398174 -22966 398230 -22910
rect 398316 -22966 398372 -22910
rect 398174 -23108 398230 -23052
rect 398316 -23108 398372 -23052
rect 398174 -23250 398230 -23194
rect 398316 -23250 398372 -23194
rect 398174 -23392 398230 -23336
rect 398316 -23392 398372 -23336
rect 398174 -23534 398230 -23478
rect 398316 -23534 398372 -23478
rect 398174 -23676 398230 -23620
rect 398316 -23676 398372 -23620
rect 398174 -23818 398230 -23762
rect 398316 -23818 398372 -23762
rect 398174 -23960 398230 -23904
rect 398316 -23960 398372 -23904
rect 398174 -24102 398230 -24046
rect 398316 -24102 398372 -24046
rect 398174 -24244 398230 -24188
rect 398316 -24244 398372 -24188
rect 398174 -24386 398230 -24330
rect 398316 -24386 398372 -24330
rect 398174 -24528 398230 -24472
rect 398316 -24528 398372 -24472
rect 398174 -24670 398230 -24614
rect 398316 -24670 398372 -24614
rect 398174 -24812 398230 -24756
rect 398316 -24812 398372 -24756
rect 398174 -24954 398230 -24898
rect 398316 -24954 398372 -24898
rect 398174 -25096 398230 -25040
rect 398316 -25096 398372 -25040
rect 398174 -25238 398230 -25182
rect 398316 -25238 398372 -25182
rect 398174 -25380 398230 -25324
rect 398316 -25380 398372 -25324
rect 398174 -25522 398230 -25466
rect 398316 -25522 398372 -25466
rect 398574 -13736 398630 -13680
rect 398716 -13736 398772 -13680
rect 398574 -13878 398630 -13822
rect 398716 -13878 398772 -13822
rect 398574 -14020 398630 -13964
rect 398716 -14020 398772 -13964
rect 398574 -14162 398630 -14106
rect 398716 -14162 398772 -14106
rect 398574 -14304 398630 -14248
rect 398716 -14304 398772 -14248
rect 398574 -14446 398630 -14390
rect 398716 -14446 398772 -14390
rect 398574 -14588 398630 -14532
rect 398716 -14588 398772 -14532
rect 398574 -14730 398630 -14674
rect 398716 -14730 398772 -14674
rect 398574 -14872 398630 -14816
rect 398716 -14872 398772 -14816
rect 398574 -15014 398630 -14958
rect 398716 -15014 398772 -14958
rect 398574 -15156 398630 -15100
rect 398716 -15156 398772 -15100
rect 398574 -15298 398630 -15242
rect 398716 -15298 398772 -15242
rect 398574 -15440 398630 -15384
rect 398716 -15440 398772 -15384
rect 398574 -15582 398630 -15526
rect 398716 -15582 398772 -15526
rect 398574 -15724 398630 -15668
rect 398716 -15724 398772 -15668
rect 398574 -15866 398630 -15810
rect 398716 -15866 398772 -15810
rect 398574 -16008 398630 -15952
rect 398716 -16008 398772 -15952
rect 398574 -16150 398630 -16094
rect 398716 -16150 398772 -16094
rect 398574 -16292 398630 -16236
rect 398716 -16292 398772 -16236
rect 398574 -16434 398630 -16378
rect 398716 -16434 398772 -16378
rect 398574 -16576 398630 -16520
rect 398716 -16576 398772 -16520
rect 398574 -16718 398630 -16662
rect 398716 -16718 398772 -16662
rect 398574 -16860 398630 -16804
rect 398716 -16860 398772 -16804
rect 398574 -17002 398630 -16946
rect 398716 -17002 398772 -16946
rect 398574 -17144 398630 -17088
rect 398716 -17144 398772 -17088
rect 398574 -17286 398630 -17230
rect 398716 -17286 398772 -17230
rect 398574 -17428 398630 -17372
rect 398716 -17428 398772 -17372
rect 398574 -17570 398630 -17514
rect 398716 -17570 398772 -17514
rect 398574 -17712 398630 -17656
rect 398716 -17712 398772 -17656
rect 398574 -17854 398630 -17798
rect 398716 -17854 398772 -17798
rect 398574 -17996 398630 -17940
rect 398716 -17996 398772 -17940
rect 398574 -18138 398630 -18082
rect 398716 -18138 398772 -18082
rect 398574 -18280 398630 -18224
rect 398716 -18280 398772 -18224
rect 398574 -18422 398630 -18366
rect 398716 -18422 398772 -18366
rect 398574 -18564 398630 -18508
rect 398716 -18564 398772 -18508
rect 398574 -18706 398630 -18650
rect 398716 -18706 398772 -18650
rect 398574 -18848 398630 -18792
rect 398716 -18848 398772 -18792
rect 398574 -18990 398630 -18934
rect 398716 -18990 398772 -18934
rect 398574 -19132 398630 -19076
rect 398716 -19132 398772 -19076
rect 398574 -19274 398630 -19218
rect 398716 -19274 398772 -19218
rect 398574 -19416 398630 -19360
rect 398716 -19416 398772 -19360
rect 398574 -19558 398630 -19502
rect 398716 -19558 398772 -19502
rect 398574 -19700 398630 -19644
rect 398716 -19700 398772 -19644
rect 398574 -19842 398630 -19786
rect 398716 -19842 398772 -19786
rect 398574 -19984 398630 -19928
rect 398716 -19984 398772 -19928
rect 398574 -20126 398630 -20070
rect 398716 -20126 398772 -20070
rect 398574 -20268 398630 -20212
rect 398716 -20268 398772 -20212
rect 398574 -20410 398630 -20354
rect 398716 -20410 398772 -20354
rect 398574 -20552 398630 -20496
rect 398716 -20552 398772 -20496
rect 398574 -20694 398630 -20638
rect 398716 -20694 398772 -20638
rect 398574 -20836 398630 -20780
rect 398716 -20836 398772 -20780
rect 398574 -20978 398630 -20922
rect 398716 -20978 398772 -20922
rect 398574 -21120 398630 -21064
rect 398716 -21120 398772 -21064
rect 398574 -21262 398630 -21206
rect 398716 -21262 398772 -21206
rect 398574 -21404 398630 -21348
rect 398716 -21404 398772 -21348
rect 398574 -21546 398630 -21490
rect 398716 -21546 398772 -21490
rect 398574 -21688 398630 -21632
rect 398716 -21688 398772 -21632
rect 398574 -21830 398630 -21774
rect 398716 -21830 398772 -21774
rect 398574 -21972 398630 -21916
rect 398716 -21972 398772 -21916
rect 398574 -22114 398630 -22058
rect 398716 -22114 398772 -22058
rect 398574 -22256 398630 -22200
rect 398716 -22256 398772 -22200
rect 398574 -22398 398630 -22342
rect 398716 -22398 398772 -22342
rect 398574 -22540 398630 -22484
rect 398716 -22540 398772 -22484
rect 398574 -22682 398630 -22626
rect 398716 -22682 398772 -22626
rect 398574 -22824 398630 -22768
rect 398716 -22824 398772 -22768
rect 398574 -22966 398630 -22910
rect 398716 -22966 398772 -22910
rect 398574 -23108 398630 -23052
rect 398716 -23108 398772 -23052
rect 398574 -23250 398630 -23194
rect 398716 -23250 398772 -23194
rect 398574 -23392 398630 -23336
rect 398716 -23392 398772 -23336
rect 398574 -23534 398630 -23478
rect 398716 -23534 398772 -23478
rect 398574 -23676 398630 -23620
rect 398716 -23676 398772 -23620
rect 398574 -23818 398630 -23762
rect 398716 -23818 398772 -23762
rect 398574 -23960 398630 -23904
rect 398716 -23960 398772 -23904
rect 398574 -24102 398630 -24046
rect 398716 -24102 398772 -24046
rect 398574 -24244 398630 -24188
rect 398716 -24244 398772 -24188
rect 398574 -24386 398630 -24330
rect 398716 -24386 398772 -24330
rect 398574 -24528 398630 -24472
rect 398716 -24528 398772 -24472
rect 398574 -24670 398630 -24614
rect 398716 -24670 398772 -24614
rect 398574 -24812 398630 -24756
rect 398716 -24812 398772 -24756
rect 398574 -24954 398630 -24898
rect 398716 -24954 398772 -24898
rect 398574 -25096 398630 -25040
rect 398716 -25096 398772 -25040
rect 398574 -25238 398630 -25182
rect 398716 -25238 398772 -25182
rect 398574 -25380 398630 -25324
rect 398716 -25380 398772 -25324
rect 398574 -25522 398630 -25466
rect 398716 -25522 398772 -25466
rect 398971 -13736 399027 -13680
rect 399113 -13736 399169 -13680
rect 398971 -13878 399027 -13822
rect 399113 -13878 399169 -13822
rect 398971 -14020 399027 -13964
rect 399113 -14020 399169 -13964
rect 398971 -14162 399027 -14106
rect 399113 -14162 399169 -14106
rect 398971 -14304 399027 -14248
rect 399113 -14304 399169 -14248
rect 398971 -14446 399027 -14390
rect 399113 -14446 399169 -14390
rect 398971 -14588 399027 -14532
rect 399113 -14588 399169 -14532
rect 398971 -14730 399027 -14674
rect 399113 -14730 399169 -14674
rect 398971 -14872 399027 -14816
rect 399113 -14872 399169 -14816
rect 398971 -15014 399027 -14958
rect 399113 -15014 399169 -14958
rect 398971 -15156 399027 -15100
rect 399113 -15156 399169 -15100
rect 398971 -15298 399027 -15242
rect 399113 -15298 399169 -15242
rect 398971 -15440 399027 -15384
rect 399113 -15440 399169 -15384
rect 398971 -15582 399027 -15526
rect 399113 -15582 399169 -15526
rect 398971 -15724 399027 -15668
rect 399113 -15724 399169 -15668
rect 398971 -15866 399027 -15810
rect 399113 -15866 399169 -15810
rect 398971 -16008 399027 -15952
rect 399113 -16008 399169 -15952
rect 398971 -16150 399027 -16094
rect 399113 -16150 399169 -16094
rect 398971 -16292 399027 -16236
rect 399113 -16292 399169 -16236
rect 398971 -16434 399027 -16378
rect 399113 -16434 399169 -16378
rect 398971 -16576 399027 -16520
rect 399113 -16576 399169 -16520
rect 398971 -16718 399027 -16662
rect 399113 -16718 399169 -16662
rect 398971 -16860 399027 -16804
rect 399113 -16860 399169 -16804
rect 398971 -17002 399027 -16946
rect 399113 -17002 399169 -16946
rect 398971 -17144 399027 -17088
rect 399113 -17144 399169 -17088
rect 398971 -17286 399027 -17230
rect 399113 -17286 399169 -17230
rect 398971 -17428 399027 -17372
rect 399113 -17428 399169 -17372
rect 398971 -17570 399027 -17514
rect 399113 -17570 399169 -17514
rect 398971 -17712 399027 -17656
rect 399113 -17712 399169 -17656
rect 398971 -17854 399027 -17798
rect 399113 -17854 399169 -17798
rect 398971 -17996 399027 -17940
rect 399113 -17996 399169 -17940
rect 398971 -18138 399027 -18082
rect 399113 -18138 399169 -18082
rect 398971 -18280 399027 -18224
rect 399113 -18280 399169 -18224
rect 398971 -18422 399027 -18366
rect 399113 -18422 399169 -18366
rect 398971 -18564 399027 -18508
rect 399113 -18564 399169 -18508
rect 398971 -18706 399027 -18650
rect 399113 -18706 399169 -18650
rect 398971 -18848 399027 -18792
rect 399113 -18848 399169 -18792
rect 398971 -18990 399027 -18934
rect 399113 -18990 399169 -18934
rect 398971 -19132 399027 -19076
rect 399113 -19132 399169 -19076
rect 398971 -19274 399027 -19218
rect 399113 -19274 399169 -19218
rect 398971 -19416 399027 -19360
rect 399113 -19416 399169 -19360
rect 398971 -19558 399027 -19502
rect 399113 -19558 399169 -19502
rect 398971 -19700 399027 -19644
rect 399113 -19700 399169 -19644
rect 398971 -19842 399027 -19786
rect 399113 -19842 399169 -19786
rect 398971 -19984 399027 -19928
rect 399113 -19984 399169 -19928
rect 398971 -20126 399027 -20070
rect 399113 -20126 399169 -20070
rect 398971 -20268 399027 -20212
rect 399113 -20268 399169 -20212
rect 398971 -20410 399027 -20354
rect 399113 -20410 399169 -20354
rect 398971 -20552 399027 -20496
rect 399113 -20552 399169 -20496
rect 398971 -20694 399027 -20638
rect 399113 -20694 399169 -20638
rect 398971 -20836 399027 -20780
rect 399113 -20836 399169 -20780
rect 398971 -20978 399027 -20922
rect 399113 -20978 399169 -20922
rect 398971 -21120 399027 -21064
rect 399113 -21120 399169 -21064
rect 398971 -21262 399027 -21206
rect 399113 -21262 399169 -21206
rect 398971 -21404 399027 -21348
rect 399113 -21404 399169 -21348
rect 398971 -21546 399027 -21490
rect 399113 -21546 399169 -21490
rect 398971 -21688 399027 -21632
rect 399113 -21688 399169 -21632
rect 398971 -21830 399027 -21774
rect 399113 -21830 399169 -21774
rect 398971 -21972 399027 -21916
rect 399113 -21972 399169 -21916
rect 398971 -22114 399027 -22058
rect 399113 -22114 399169 -22058
rect 398971 -22256 399027 -22200
rect 399113 -22256 399169 -22200
rect 398971 -22398 399027 -22342
rect 399113 -22398 399169 -22342
rect 398971 -22540 399027 -22484
rect 399113 -22540 399169 -22484
rect 398971 -22682 399027 -22626
rect 399113 -22682 399169 -22626
rect 398971 -22824 399027 -22768
rect 399113 -22824 399169 -22768
rect 398971 -22966 399027 -22910
rect 399113 -22966 399169 -22910
rect 398971 -23108 399027 -23052
rect 399113 -23108 399169 -23052
rect 398971 -23250 399027 -23194
rect 399113 -23250 399169 -23194
rect 398971 -23392 399027 -23336
rect 399113 -23392 399169 -23336
rect 398971 -23534 399027 -23478
rect 399113 -23534 399169 -23478
rect 398971 -23676 399027 -23620
rect 399113 -23676 399169 -23620
rect 398971 -23818 399027 -23762
rect 399113 -23818 399169 -23762
rect 398971 -23960 399027 -23904
rect 399113 -23960 399169 -23904
rect 398971 -24102 399027 -24046
rect 399113 -24102 399169 -24046
rect 398971 -24244 399027 -24188
rect 399113 -24244 399169 -24188
rect 398971 -24386 399027 -24330
rect 399113 -24386 399169 -24330
rect 398971 -24528 399027 -24472
rect 399113 -24528 399169 -24472
rect 398971 -24670 399027 -24614
rect 399113 -24670 399169 -24614
rect 398971 -24812 399027 -24756
rect 399113 -24812 399169 -24756
rect 398971 -24954 399027 -24898
rect 399113 -24954 399169 -24898
rect 398971 -25096 399027 -25040
rect 399113 -25096 399169 -25040
rect 398971 -25238 399027 -25182
rect 399113 -25238 399169 -25182
rect 398971 -25380 399027 -25324
rect 399113 -25380 399169 -25324
rect 398971 -25522 399027 -25466
rect 399113 -25522 399169 -25466
rect 399376 -13736 399432 -13680
rect 399518 -13736 399574 -13680
rect 399376 -13878 399432 -13822
rect 399518 -13878 399574 -13822
rect 399376 -14020 399432 -13964
rect 399518 -14020 399574 -13964
rect 399376 -14162 399432 -14106
rect 399518 -14162 399574 -14106
rect 399376 -14304 399432 -14248
rect 399518 -14304 399574 -14248
rect 399376 -14446 399432 -14390
rect 399518 -14446 399574 -14390
rect 399376 -14588 399432 -14532
rect 399518 -14588 399574 -14532
rect 399376 -14730 399432 -14674
rect 399518 -14730 399574 -14674
rect 399376 -14872 399432 -14816
rect 399518 -14872 399574 -14816
rect 399376 -15014 399432 -14958
rect 399518 -15014 399574 -14958
rect 399376 -15156 399432 -15100
rect 399518 -15156 399574 -15100
rect 399376 -15298 399432 -15242
rect 399518 -15298 399574 -15242
rect 399376 -15440 399432 -15384
rect 399518 -15440 399574 -15384
rect 399376 -15582 399432 -15526
rect 399518 -15582 399574 -15526
rect 399376 -15724 399432 -15668
rect 399518 -15724 399574 -15668
rect 399376 -15866 399432 -15810
rect 399518 -15866 399574 -15810
rect 399376 -16008 399432 -15952
rect 399518 -16008 399574 -15952
rect 399376 -16150 399432 -16094
rect 399518 -16150 399574 -16094
rect 399376 -16292 399432 -16236
rect 399518 -16292 399574 -16236
rect 399376 -16434 399432 -16378
rect 399518 -16434 399574 -16378
rect 399376 -16576 399432 -16520
rect 399518 -16576 399574 -16520
rect 399376 -16718 399432 -16662
rect 399518 -16718 399574 -16662
rect 399376 -16860 399432 -16804
rect 399518 -16860 399574 -16804
rect 399376 -17002 399432 -16946
rect 399518 -17002 399574 -16946
rect 399376 -17144 399432 -17088
rect 399518 -17144 399574 -17088
rect 399376 -17286 399432 -17230
rect 399518 -17286 399574 -17230
rect 399376 -17428 399432 -17372
rect 399518 -17428 399574 -17372
rect 399376 -17570 399432 -17514
rect 399518 -17570 399574 -17514
rect 399376 -17712 399432 -17656
rect 399518 -17712 399574 -17656
rect 399376 -17854 399432 -17798
rect 399518 -17854 399574 -17798
rect 399376 -17996 399432 -17940
rect 399518 -17996 399574 -17940
rect 399376 -18138 399432 -18082
rect 399518 -18138 399574 -18082
rect 399376 -18280 399432 -18224
rect 399518 -18280 399574 -18224
rect 399376 -18422 399432 -18366
rect 399518 -18422 399574 -18366
rect 399376 -18564 399432 -18508
rect 399518 -18564 399574 -18508
rect 399376 -18706 399432 -18650
rect 399518 -18706 399574 -18650
rect 399376 -18848 399432 -18792
rect 399518 -18848 399574 -18792
rect 399376 -18990 399432 -18934
rect 399518 -18990 399574 -18934
rect 399376 -19132 399432 -19076
rect 399518 -19132 399574 -19076
rect 399376 -19274 399432 -19218
rect 399518 -19274 399574 -19218
rect 399376 -19416 399432 -19360
rect 399518 -19416 399574 -19360
rect 399376 -19558 399432 -19502
rect 399518 -19558 399574 -19502
rect 399376 -19700 399432 -19644
rect 399518 -19700 399574 -19644
rect 399376 -19842 399432 -19786
rect 399518 -19842 399574 -19786
rect 399376 -19984 399432 -19928
rect 399518 -19984 399574 -19928
rect 399376 -20126 399432 -20070
rect 399518 -20126 399574 -20070
rect 399376 -20268 399432 -20212
rect 399518 -20268 399574 -20212
rect 399376 -20410 399432 -20354
rect 399518 -20410 399574 -20354
rect 399376 -20552 399432 -20496
rect 399518 -20552 399574 -20496
rect 399376 -20694 399432 -20638
rect 399518 -20694 399574 -20638
rect 399376 -20836 399432 -20780
rect 399518 -20836 399574 -20780
rect 399376 -20978 399432 -20922
rect 399518 -20978 399574 -20922
rect 399376 -21120 399432 -21064
rect 399518 -21120 399574 -21064
rect 399376 -21262 399432 -21206
rect 399518 -21262 399574 -21206
rect 399376 -21404 399432 -21348
rect 399518 -21404 399574 -21348
rect 399376 -21546 399432 -21490
rect 399518 -21546 399574 -21490
rect 399376 -21688 399432 -21632
rect 399518 -21688 399574 -21632
rect 399376 -21830 399432 -21774
rect 399518 -21830 399574 -21774
rect 399376 -21972 399432 -21916
rect 399518 -21972 399574 -21916
rect 399376 -22114 399432 -22058
rect 399518 -22114 399574 -22058
rect 399376 -22256 399432 -22200
rect 399518 -22256 399574 -22200
rect 399376 -22398 399432 -22342
rect 399518 -22398 399574 -22342
rect 399376 -22540 399432 -22484
rect 399518 -22540 399574 -22484
rect 399376 -22682 399432 -22626
rect 399518 -22682 399574 -22626
rect 399376 -22824 399432 -22768
rect 399518 -22824 399574 -22768
rect 399376 -22966 399432 -22910
rect 399518 -22966 399574 -22910
rect 399376 -23108 399432 -23052
rect 399518 -23108 399574 -23052
rect 399376 -23250 399432 -23194
rect 399518 -23250 399574 -23194
rect 399376 -23392 399432 -23336
rect 399518 -23392 399574 -23336
rect 399376 -23534 399432 -23478
rect 399518 -23534 399574 -23478
rect 399376 -23676 399432 -23620
rect 399518 -23676 399574 -23620
rect 399376 -23818 399432 -23762
rect 399518 -23818 399574 -23762
rect 399376 -23960 399432 -23904
rect 399518 -23960 399574 -23904
rect 399376 -24102 399432 -24046
rect 399518 -24102 399574 -24046
rect 399376 -24244 399432 -24188
rect 399518 -24244 399574 -24188
rect 399376 -24386 399432 -24330
rect 399518 -24386 399574 -24330
rect 399376 -24528 399432 -24472
rect 399518 -24528 399574 -24472
rect 399376 -24670 399432 -24614
rect 399518 -24670 399574 -24614
rect 399376 -24812 399432 -24756
rect 399518 -24812 399574 -24756
rect 399376 -24954 399432 -24898
rect 399518 -24954 399574 -24898
rect 399376 -25096 399432 -25040
rect 399518 -25096 399574 -25040
rect 399376 -25238 399432 -25182
rect 399518 -25238 399574 -25182
rect 399376 -25380 399432 -25324
rect 399518 -25380 399574 -25324
rect 399376 -25522 399432 -25466
rect 399518 -25522 399574 -25466
rect 399776 -13736 399832 -13680
rect 399918 -13736 399974 -13680
rect 399776 -13878 399832 -13822
rect 399918 -13878 399974 -13822
rect 399776 -14020 399832 -13964
rect 399918 -14020 399974 -13964
rect 399776 -14162 399832 -14106
rect 399918 -14162 399974 -14106
rect 399776 -14304 399832 -14248
rect 399918 -14304 399974 -14248
rect 399776 -14446 399832 -14390
rect 399918 -14446 399974 -14390
rect 399776 -14588 399832 -14532
rect 399918 -14588 399974 -14532
rect 399776 -14730 399832 -14674
rect 399918 -14730 399974 -14674
rect 399776 -14872 399832 -14816
rect 399918 -14872 399974 -14816
rect 399776 -15014 399832 -14958
rect 399918 -15014 399974 -14958
rect 399776 -15156 399832 -15100
rect 399918 -15156 399974 -15100
rect 399776 -15298 399832 -15242
rect 399918 -15298 399974 -15242
rect 399776 -15440 399832 -15384
rect 399918 -15440 399974 -15384
rect 399776 -15582 399832 -15526
rect 399918 -15582 399974 -15526
rect 399776 -15724 399832 -15668
rect 399918 -15724 399974 -15668
rect 399776 -15866 399832 -15810
rect 399918 -15866 399974 -15810
rect 399776 -16008 399832 -15952
rect 399918 -16008 399974 -15952
rect 399776 -16150 399832 -16094
rect 399918 -16150 399974 -16094
rect 399776 -16292 399832 -16236
rect 399918 -16292 399974 -16236
rect 399776 -16434 399832 -16378
rect 399918 -16434 399974 -16378
rect 399776 -16576 399832 -16520
rect 399918 -16576 399974 -16520
rect 399776 -16718 399832 -16662
rect 399918 -16718 399974 -16662
rect 399776 -16860 399832 -16804
rect 399918 -16860 399974 -16804
rect 399776 -17002 399832 -16946
rect 399918 -17002 399974 -16946
rect 399776 -17144 399832 -17088
rect 399918 -17144 399974 -17088
rect 399776 -17286 399832 -17230
rect 399918 -17286 399974 -17230
rect 399776 -17428 399832 -17372
rect 399918 -17428 399974 -17372
rect 399776 -17570 399832 -17514
rect 399918 -17570 399974 -17514
rect 399776 -17712 399832 -17656
rect 399918 -17712 399974 -17656
rect 399776 -17854 399832 -17798
rect 399918 -17854 399974 -17798
rect 399776 -17996 399832 -17940
rect 399918 -17996 399974 -17940
rect 399776 -18138 399832 -18082
rect 399918 -18138 399974 -18082
rect 399776 -18280 399832 -18224
rect 399918 -18280 399974 -18224
rect 399776 -18422 399832 -18366
rect 399918 -18422 399974 -18366
rect 399776 -18564 399832 -18508
rect 399918 -18564 399974 -18508
rect 399776 -18706 399832 -18650
rect 399918 -18706 399974 -18650
rect 399776 -18848 399832 -18792
rect 399918 -18848 399974 -18792
rect 399776 -18990 399832 -18934
rect 399918 -18990 399974 -18934
rect 399776 -19132 399832 -19076
rect 399918 -19132 399974 -19076
rect 399776 -19274 399832 -19218
rect 399918 -19274 399974 -19218
rect 399776 -19416 399832 -19360
rect 399918 -19416 399974 -19360
rect 399776 -19558 399832 -19502
rect 399918 -19558 399974 -19502
rect 399776 -19700 399832 -19644
rect 399918 -19700 399974 -19644
rect 399776 -19842 399832 -19786
rect 399918 -19842 399974 -19786
rect 399776 -19984 399832 -19928
rect 399918 -19984 399974 -19928
rect 399776 -20126 399832 -20070
rect 399918 -20126 399974 -20070
rect 399776 -20268 399832 -20212
rect 399918 -20268 399974 -20212
rect 399776 -20410 399832 -20354
rect 399918 -20410 399974 -20354
rect 399776 -20552 399832 -20496
rect 399918 -20552 399974 -20496
rect 399776 -20694 399832 -20638
rect 399918 -20694 399974 -20638
rect 399776 -20836 399832 -20780
rect 399918 -20836 399974 -20780
rect 399776 -20978 399832 -20922
rect 399918 -20978 399974 -20922
rect 399776 -21120 399832 -21064
rect 399918 -21120 399974 -21064
rect 399776 -21262 399832 -21206
rect 399918 -21262 399974 -21206
rect 399776 -21404 399832 -21348
rect 399918 -21404 399974 -21348
rect 399776 -21546 399832 -21490
rect 399918 -21546 399974 -21490
rect 399776 -21688 399832 -21632
rect 399918 -21688 399974 -21632
rect 399776 -21830 399832 -21774
rect 399918 -21830 399974 -21774
rect 399776 -21972 399832 -21916
rect 399918 -21972 399974 -21916
rect 399776 -22114 399832 -22058
rect 399918 -22114 399974 -22058
rect 399776 -22256 399832 -22200
rect 399918 -22256 399974 -22200
rect 399776 -22398 399832 -22342
rect 399918 -22398 399974 -22342
rect 399776 -22540 399832 -22484
rect 399918 -22540 399974 -22484
rect 399776 -22682 399832 -22626
rect 399918 -22682 399974 -22626
rect 399776 -22824 399832 -22768
rect 399918 -22824 399974 -22768
rect 399776 -22966 399832 -22910
rect 399918 -22966 399974 -22910
rect 399776 -23108 399832 -23052
rect 399918 -23108 399974 -23052
rect 399776 -23250 399832 -23194
rect 399918 -23250 399974 -23194
rect 399776 -23392 399832 -23336
rect 399918 -23392 399974 -23336
rect 399776 -23534 399832 -23478
rect 399918 -23534 399974 -23478
rect 399776 -23676 399832 -23620
rect 399918 -23676 399974 -23620
rect 399776 -23818 399832 -23762
rect 399918 -23818 399974 -23762
rect 399776 -23960 399832 -23904
rect 399918 -23960 399974 -23904
rect 399776 -24102 399832 -24046
rect 399918 -24102 399974 -24046
rect 399776 -24244 399832 -24188
rect 399918 -24244 399974 -24188
rect 399776 -24386 399832 -24330
rect 399918 -24386 399974 -24330
rect 399776 -24528 399832 -24472
rect 399918 -24528 399974 -24472
rect 399776 -24670 399832 -24614
rect 399918 -24670 399974 -24614
rect 399776 -24812 399832 -24756
rect 399918 -24812 399974 -24756
rect 399776 -24954 399832 -24898
rect 399918 -24954 399974 -24898
rect 399776 -25096 399832 -25040
rect 399918 -25096 399974 -25040
rect 399776 -25238 399832 -25182
rect 399918 -25238 399974 -25182
rect 399776 -25380 399832 -25324
rect 399918 -25380 399974 -25324
rect 399776 -25522 399832 -25466
rect 399918 -25522 399974 -25466
rect 400181 -13736 400237 -13680
rect 400323 -13736 400379 -13680
rect 400181 -13878 400237 -13822
rect 400323 -13878 400379 -13822
rect 400181 -14020 400237 -13964
rect 400323 -14020 400379 -13964
rect 400181 -14162 400237 -14106
rect 400323 -14162 400379 -14106
rect 400181 -14304 400237 -14248
rect 400323 -14304 400379 -14248
rect 400181 -14446 400237 -14390
rect 400323 -14446 400379 -14390
rect 400181 -14588 400237 -14532
rect 400323 -14588 400379 -14532
rect 400181 -14730 400237 -14674
rect 400323 -14730 400379 -14674
rect 400181 -14872 400237 -14816
rect 400323 -14872 400379 -14816
rect 400181 -15014 400237 -14958
rect 400323 -15014 400379 -14958
rect 400181 -15156 400237 -15100
rect 400323 -15156 400379 -15100
rect 400181 -15298 400237 -15242
rect 400323 -15298 400379 -15242
rect 400181 -15440 400237 -15384
rect 400323 -15440 400379 -15384
rect 400181 -15582 400237 -15526
rect 400323 -15582 400379 -15526
rect 400181 -15724 400237 -15668
rect 400323 -15724 400379 -15668
rect 400181 -15866 400237 -15810
rect 400323 -15866 400379 -15810
rect 400181 -16008 400237 -15952
rect 400323 -16008 400379 -15952
rect 400181 -16150 400237 -16094
rect 400323 -16150 400379 -16094
rect 400181 -16292 400237 -16236
rect 400323 -16292 400379 -16236
rect 400181 -16434 400237 -16378
rect 400323 -16434 400379 -16378
rect 400181 -16576 400237 -16520
rect 400323 -16576 400379 -16520
rect 400181 -16718 400237 -16662
rect 400323 -16718 400379 -16662
rect 400181 -16860 400237 -16804
rect 400323 -16860 400379 -16804
rect 400181 -17002 400237 -16946
rect 400323 -17002 400379 -16946
rect 400181 -17144 400237 -17088
rect 400323 -17144 400379 -17088
rect 400181 -17286 400237 -17230
rect 400323 -17286 400379 -17230
rect 400181 -17428 400237 -17372
rect 400323 -17428 400379 -17372
rect 400181 -17570 400237 -17514
rect 400323 -17570 400379 -17514
rect 400181 -17712 400237 -17656
rect 400323 -17712 400379 -17656
rect 400181 -17854 400237 -17798
rect 400323 -17854 400379 -17798
rect 400181 -17996 400237 -17940
rect 400323 -17996 400379 -17940
rect 400181 -18138 400237 -18082
rect 400323 -18138 400379 -18082
rect 400181 -18280 400237 -18224
rect 400323 -18280 400379 -18224
rect 400181 -18422 400237 -18366
rect 400323 -18422 400379 -18366
rect 400181 -18564 400237 -18508
rect 400323 -18564 400379 -18508
rect 400181 -18706 400237 -18650
rect 400323 -18706 400379 -18650
rect 400181 -18848 400237 -18792
rect 400323 -18848 400379 -18792
rect 400181 -18990 400237 -18934
rect 400323 -18990 400379 -18934
rect 400181 -19132 400237 -19076
rect 400323 -19132 400379 -19076
rect 400181 -19274 400237 -19218
rect 400323 -19274 400379 -19218
rect 400181 -19416 400237 -19360
rect 400323 -19416 400379 -19360
rect 400181 -19558 400237 -19502
rect 400323 -19558 400379 -19502
rect 400181 -19700 400237 -19644
rect 400323 -19700 400379 -19644
rect 400181 -19842 400237 -19786
rect 400323 -19842 400379 -19786
rect 400181 -19984 400237 -19928
rect 400323 -19984 400379 -19928
rect 400181 -20126 400237 -20070
rect 400323 -20126 400379 -20070
rect 400181 -20268 400237 -20212
rect 400323 -20268 400379 -20212
rect 400181 -20410 400237 -20354
rect 400323 -20410 400379 -20354
rect 400181 -20552 400237 -20496
rect 400323 -20552 400379 -20496
rect 400181 -20694 400237 -20638
rect 400323 -20694 400379 -20638
rect 400181 -20836 400237 -20780
rect 400323 -20836 400379 -20780
rect 400181 -20978 400237 -20922
rect 400323 -20978 400379 -20922
rect 400181 -21120 400237 -21064
rect 400323 -21120 400379 -21064
rect 400181 -21262 400237 -21206
rect 400323 -21262 400379 -21206
rect 400181 -21404 400237 -21348
rect 400323 -21404 400379 -21348
rect 400181 -21546 400237 -21490
rect 400323 -21546 400379 -21490
rect 400181 -21688 400237 -21632
rect 400323 -21688 400379 -21632
rect 400181 -21830 400237 -21774
rect 400323 -21830 400379 -21774
rect 400181 -21972 400237 -21916
rect 400323 -21972 400379 -21916
rect 400181 -22114 400237 -22058
rect 400323 -22114 400379 -22058
rect 400181 -22256 400237 -22200
rect 400323 -22256 400379 -22200
rect 400181 -22398 400237 -22342
rect 400323 -22398 400379 -22342
rect 400181 -22540 400237 -22484
rect 400323 -22540 400379 -22484
rect 400181 -22682 400237 -22626
rect 400323 -22682 400379 -22626
rect 400181 -22824 400237 -22768
rect 400323 -22824 400379 -22768
rect 400181 -22966 400237 -22910
rect 400323 -22966 400379 -22910
rect 400181 -23108 400237 -23052
rect 400323 -23108 400379 -23052
rect 400181 -23250 400237 -23194
rect 400323 -23250 400379 -23194
rect 400181 -23392 400237 -23336
rect 400323 -23392 400379 -23336
rect 400181 -23534 400237 -23478
rect 400323 -23534 400379 -23478
rect 400181 -23676 400237 -23620
rect 400323 -23676 400379 -23620
rect 400181 -23818 400237 -23762
rect 400323 -23818 400379 -23762
rect 400181 -23960 400237 -23904
rect 400323 -23960 400379 -23904
rect 400181 -24102 400237 -24046
rect 400323 -24102 400379 -24046
rect 400181 -24244 400237 -24188
rect 400323 -24244 400379 -24188
rect 400181 -24386 400237 -24330
rect 400323 -24386 400379 -24330
rect 400181 -24528 400237 -24472
rect 400323 -24528 400379 -24472
rect 400181 -24670 400237 -24614
rect 400323 -24670 400379 -24614
rect 400181 -24812 400237 -24756
rect 400323 -24812 400379 -24756
rect 400181 -24954 400237 -24898
rect 400323 -24954 400379 -24898
rect 400181 -25096 400237 -25040
rect 400323 -25096 400379 -25040
rect 400181 -25238 400237 -25182
rect 400323 -25238 400379 -25182
rect 400181 -25380 400237 -25324
rect 400323 -25380 400379 -25324
rect 400181 -25522 400237 -25466
rect 400323 -25522 400379 -25466
rect 400766 -13688 400822 -13632
rect 400890 -13688 400946 -13632
rect 401014 -13688 401070 -13632
rect 401138 -13688 401194 -13632
rect 401262 -13688 401318 -13632
rect 400766 -13812 400822 -13756
rect 400890 -13812 400946 -13756
rect 401014 -13812 401070 -13756
rect 401138 -13812 401194 -13756
rect 401262 -13812 401318 -13756
rect 400766 -13936 400822 -13880
rect 400890 -13936 400946 -13880
rect 401014 -13936 401070 -13880
rect 401138 -13936 401194 -13880
rect 401262 -13936 401318 -13880
rect 400766 -14060 400822 -14004
rect 400890 -14060 400946 -14004
rect 401014 -14060 401070 -14004
rect 401138 -14060 401194 -14004
rect 401262 -14060 401318 -14004
rect 400766 -14184 400822 -14128
rect 400890 -14184 400946 -14128
rect 401014 -14184 401070 -14128
rect 401138 -14184 401194 -14128
rect 401262 -14184 401318 -14128
rect 400766 -14308 400822 -14252
rect 400890 -14308 400946 -14252
rect 401014 -14308 401070 -14252
rect 401138 -14308 401194 -14252
rect 401262 -14308 401318 -14252
rect 400766 -14432 400822 -14376
rect 400890 -14432 400946 -14376
rect 401014 -14432 401070 -14376
rect 401138 -14432 401194 -14376
rect 401262 -14432 401318 -14376
rect 400766 -14556 400822 -14500
rect 400890 -14556 400946 -14500
rect 401014 -14556 401070 -14500
rect 401138 -14556 401194 -14500
rect 401262 -14556 401318 -14500
rect 400766 -14680 400822 -14624
rect 400890 -14680 400946 -14624
rect 401014 -14680 401070 -14624
rect 401138 -14680 401194 -14624
rect 401262 -14680 401318 -14624
rect 400766 -14804 400822 -14748
rect 400890 -14804 400946 -14748
rect 401014 -14804 401070 -14748
rect 401138 -14804 401194 -14748
rect 401262 -14804 401318 -14748
rect 400766 -14928 400822 -14872
rect 400890 -14928 400946 -14872
rect 401014 -14928 401070 -14872
rect 401138 -14928 401194 -14872
rect 401262 -14928 401318 -14872
rect 400766 -15052 400822 -14996
rect 400890 -15052 400946 -14996
rect 401014 -15052 401070 -14996
rect 401138 -15052 401194 -14996
rect 401262 -15052 401318 -14996
rect 400766 -15176 400822 -15120
rect 400890 -15176 400946 -15120
rect 401014 -15176 401070 -15120
rect 401138 -15176 401194 -15120
rect 401262 -15176 401318 -15120
rect 400766 -15300 400822 -15244
rect 400890 -15300 400946 -15244
rect 401014 -15300 401070 -15244
rect 401138 -15300 401194 -15244
rect 401262 -15300 401318 -15244
rect 400766 -15424 400822 -15368
rect 400890 -15424 400946 -15368
rect 401014 -15424 401070 -15368
rect 401138 -15424 401194 -15368
rect 401262 -15424 401318 -15368
rect 400766 -15548 400822 -15492
rect 400890 -15548 400946 -15492
rect 401014 -15548 401070 -15492
rect 401138 -15548 401194 -15492
rect 401262 -15548 401318 -15492
rect 400766 -15672 400822 -15616
rect 400890 -15672 400946 -15616
rect 401014 -15672 401070 -15616
rect 401138 -15672 401194 -15616
rect 401262 -15672 401318 -15616
rect 400766 -15796 400822 -15740
rect 400890 -15796 400946 -15740
rect 401014 -15796 401070 -15740
rect 401138 -15796 401194 -15740
rect 401262 -15796 401318 -15740
rect 400766 -15920 400822 -15864
rect 400890 -15920 400946 -15864
rect 401014 -15920 401070 -15864
rect 401138 -15920 401194 -15864
rect 401262 -15920 401318 -15864
rect 400766 -16044 400822 -15988
rect 400890 -16044 400946 -15988
rect 401014 -16044 401070 -15988
rect 401138 -16044 401194 -15988
rect 401262 -16044 401318 -15988
rect 400766 -16168 400822 -16112
rect 400890 -16168 400946 -16112
rect 401014 -16168 401070 -16112
rect 401138 -16168 401194 -16112
rect 401262 -16168 401318 -16112
rect 400766 -16292 400822 -16236
rect 400890 -16292 400946 -16236
rect 401014 -16292 401070 -16236
rect 401138 -16292 401194 -16236
rect 401262 -16292 401318 -16236
rect 400766 -16416 400822 -16360
rect 400890 -16416 400946 -16360
rect 401014 -16416 401070 -16360
rect 401138 -16416 401194 -16360
rect 401262 -16416 401318 -16360
rect 400766 -16540 400822 -16484
rect 400890 -16540 400946 -16484
rect 401014 -16540 401070 -16484
rect 401138 -16540 401194 -16484
rect 401262 -16540 401318 -16484
rect 400766 -16664 400822 -16608
rect 400890 -16664 400946 -16608
rect 401014 -16664 401070 -16608
rect 401138 -16664 401194 -16608
rect 401262 -16664 401318 -16608
rect 400766 -16788 400822 -16732
rect 400890 -16788 400946 -16732
rect 401014 -16788 401070 -16732
rect 401138 -16788 401194 -16732
rect 401262 -16788 401318 -16732
rect 400766 -16912 400822 -16856
rect 400890 -16912 400946 -16856
rect 401014 -16912 401070 -16856
rect 401138 -16912 401194 -16856
rect 401262 -16912 401318 -16856
rect 400766 -17036 400822 -16980
rect 400890 -17036 400946 -16980
rect 401014 -17036 401070 -16980
rect 401138 -17036 401194 -16980
rect 401262 -17036 401318 -16980
rect 400766 -17160 400822 -17104
rect 400890 -17160 400946 -17104
rect 401014 -17160 401070 -17104
rect 401138 -17160 401194 -17104
rect 401262 -17160 401318 -17104
rect 400766 -17284 400822 -17228
rect 400890 -17284 400946 -17228
rect 401014 -17284 401070 -17228
rect 401138 -17284 401194 -17228
rect 401262 -17284 401318 -17228
rect 400766 -17408 400822 -17352
rect 400890 -17408 400946 -17352
rect 401014 -17408 401070 -17352
rect 401138 -17408 401194 -17352
rect 401262 -17408 401318 -17352
rect 400766 -17532 400822 -17476
rect 400890 -17532 400946 -17476
rect 401014 -17532 401070 -17476
rect 401138 -17532 401194 -17476
rect 401262 -17532 401318 -17476
rect 400766 -17656 400822 -17600
rect 400890 -17656 400946 -17600
rect 401014 -17656 401070 -17600
rect 401138 -17656 401194 -17600
rect 401262 -17656 401318 -17600
rect 400766 -17780 400822 -17724
rect 400890 -17780 400946 -17724
rect 401014 -17780 401070 -17724
rect 401138 -17780 401194 -17724
rect 401262 -17780 401318 -17724
rect 400766 -17904 400822 -17848
rect 400890 -17904 400946 -17848
rect 401014 -17904 401070 -17848
rect 401138 -17904 401194 -17848
rect 401262 -17904 401318 -17848
rect 400766 -18028 400822 -17972
rect 400890 -18028 400946 -17972
rect 401014 -18028 401070 -17972
rect 401138 -18028 401194 -17972
rect 401262 -18028 401318 -17972
rect 400766 -18152 400822 -18096
rect 400890 -18152 400946 -18096
rect 401014 -18152 401070 -18096
rect 401138 -18152 401194 -18096
rect 401262 -18152 401318 -18096
rect 400766 -18276 400822 -18220
rect 400890 -18276 400946 -18220
rect 401014 -18276 401070 -18220
rect 401138 -18276 401194 -18220
rect 401262 -18276 401318 -18220
rect 400766 -18400 400822 -18344
rect 400890 -18400 400946 -18344
rect 401014 -18400 401070 -18344
rect 401138 -18400 401194 -18344
rect 401262 -18400 401318 -18344
rect 400766 -18524 400822 -18468
rect 400890 -18524 400946 -18468
rect 401014 -18524 401070 -18468
rect 401138 -18524 401194 -18468
rect 401262 -18524 401318 -18468
rect 400766 -18648 400822 -18592
rect 400890 -18648 400946 -18592
rect 401014 -18648 401070 -18592
rect 401138 -18648 401194 -18592
rect 401262 -18648 401318 -18592
rect 400766 -18772 400822 -18716
rect 400890 -18772 400946 -18716
rect 401014 -18772 401070 -18716
rect 401138 -18772 401194 -18716
rect 401262 -18772 401318 -18716
rect 400766 -18896 400822 -18840
rect 400890 -18896 400946 -18840
rect 401014 -18896 401070 -18840
rect 401138 -18896 401194 -18840
rect 401262 -18896 401318 -18840
rect 400766 -19020 400822 -18964
rect 400890 -19020 400946 -18964
rect 401014 -19020 401070 -18964
rect 401138 -19020 401194 -18964
rect 401262 -19020 401318 -18964
rect 400766 -19144 400822 -19088
rect 400890 -19144 400946 -19088
rect 401014 -19144 401070 -19088
rect 401138 -19144 401194 -19088
rect 401262 -19144 401318 -19088
rect 400766 -19268 400822 -19212
rect 400890 -19268 400946 -19212
rect 401014 -19268 401070 -19212
rect 401138 -19268 401194 -19212
rect 401262 -19268 401318 -19212
rect 400766 -19392 400822 -19336
rect 400890 -19392 400946 -19336
rect 401014 -19392 401070 -19336
rect 401138 -19392 401194 -19336
rect 401262 -19392 401318 -19336
rect 400766 -19516 400822 -19460
rect 400890 -19516 400946 -19460
rect 401014 -19516 401070 -19460
rect 401138 -19516 401194 -19460
rect 401262 -19516 401318 -19460
rect 400766 -19640 400822 -19584
rect 400890 -19640 400946 -19584
rect 401014 -19640 401070 -19584
rect 401138 -19640 401194 -19584
rect 401262 -19640 401318 -19584
rect 400766 -19764 400822 -19708
rect 400890 -19764 400946 -19708
rect 401014 -19764 401070 -19708
rect 401138 -19764 401194 -19708
rect 401262 -19764 401318 -19708
rect 400766 -19888 400822 -19832
rect 400890 -19888 400946 -19832
rect 401014 -19888 401070 -19832
rect 401138 -19888 401194 -19832
rect 401262 -19888 401318 -19832
rect 400766 -20012 400822 -19956
rect 400890 -20012 400946 -19956
rect 401014 -20012 401070 -19956
rect 401138 -20012 401194 -19956
rect 401262 -20012 401318 -19956
rect 400766 -20136 400822 -20080
rect 400890 -20136 400946 -20080
rect 401014 -20136 401070 -20080
rect 401138 -20136 401194 -20080
rect 401262 -20136 401318 -20080
rect 400766 -20260 400822 -20204
rect 400890 -20260 400946 -20204
rect 401014 -20260 401070 -20204
rect 401138 -20260 401194 -20204
rect 401262 -20260 401318 -20204
rect 400766 -20384 400822 -20328
rect 400890 -20384 400946 -20328
rect 401014 -20384 401070 -20328
rect 401138 -20384 401194 -20328
rect 401262 -20384 401318 -20328
rect 400766 -20508 400822 -20452
rect 400890 -20508 400946 -20452
rect 401014 -20508 401070 -20452
rect 401138 -20508 401194 -20452
rect 401262 -20508 401318 -20452
rect 400766 -20632 400822 -20576
rect 400890 -20632 400946 -20576
rect 401014 -20632 401070 -20576
rect 401138 -20632 401194 -20576
rect 401262 -20632 401318 -20576
rect 400766 -20756 400822 -20700
rect 400890 -20756 400946 -20700
rect 401014 -20756 401070 -20700
rect 401138 -20756 401194 -20700
rect 401262 -20756 401318 -20700
rect 400766 -20880 400822 -20824
rect 400890 -20880 400946 -20824
rect 401014 -20880 401070 -20824
rect 401138 -20880 401194 -20824
rect 401262 -20880 401318 -20824
rect 400766 -21004 400822 -20948
rect 400890 -21004 400946 -20948
rect 401014 -21004 401070 -20948
rect 401138 -21004 401194 -20948
rect 401262 -21004 401318 -20948
rect 400766 -21128 400822 -21072
rect 400890 -21128 400946 -21072
rect 401014 -21128 401070 -21072
rect 401138 -21128 401194 -21072
rect 401262 -21128 401318 -21072
rect 400766 -21252 400822 -21196
rect 400890 -21252 400946 -21196
rect 401014 -21252 401070 -21196
rect 401138 -21252 401194 -21196
rect 401262 -21252 401318 -21196
rect 400766 -21376 400822 -21320
rect 400890 -21376 400946 -21320
rect 401014 -21376 401070 -21320
rect 401138 -21376 401194 -21320
rect 401262 -21376 401318 -21320
rect 400766 -21500 400822 -21444
rect 400890 -21500 400946 -21444
rect 401014 -21500 401070 -21444
rect 401138 -21500 401194 -21444
rect 401262 -21500 401318 -21444
rect 400766 -21624 400822 -21568
rect 400890 -21624 400946 -21568
rect 401014 -21624 401070 -21568
rect 401138 -21624 401194 -21568
rect 401262 -21624 401318 -21568
rect 400766 -21748 400822 -21692
rect 400890 -21748 400946 -21692
rect 401014 -21748 401070 -21692
rect 401138 -21748 401194 -21692
rect 401262 -21748 401318 -21692
rect 400766 -21872 400822 -21816
rect 400890 -21872 400946 -21816
rect 401014 -21872 401070 -21816
rect 401138 -21872 401194 -21816
rect 401262 -21872 401318 -21816
rect 400766 -21996 400822 -21940
rect 400890 -21996 400946 -21940
rect 401014 -21996 401070 -21940
rect 401138 -21996 401194 -21940
rect 401262 -21996 401318 -21940
rect 400766 -22120 400822 -22064
rect 400890 -22120 400946 -22064
rect 401014 -22120 401070 -22064
rect 401138 -22120 401194 -22064
rect 401262 -22120 401318 -22064
rect 400766 -22244 400822 -22188
rect 400890 -22244 400946 -22188
rect 401014 -22244 401070 -22188
rect 401138 -22244 401194 -22188
rect 401262 -22244 401318 -22188
rect 400766 -22368 400822 -22312
rect 400890 -22368 400946 -22312
rect 401014 -22368 401070 -22312
rect 401138 -22368 401194 -22312
rect 401262 -22368 401318 -22312
rect 400766 -22492 400822 -22436
rect 400890 -22492 400946 -22436
rect 401014 -22492 401070 -22436
rect 401138 -22492 401194 -22436
rect 401262 -22492 401318 -22436
rect 400766 -22616 400822 -22560
rect 400890 -22616 400946 -22560
rect 401014 -22616 401070 -22560
rect 401138 -22616 401194 -22560
rect 401262 -22616 401318 -22560
rect 400766 -22740 400822 -22684
rect 400890 -22740 400946 -22684
rect 401014 -22740 401070 -22684
rect 401138 -22740 401194 -22684
rect 401262 -22740 401318 -22684
rect 400766 -22864 400822 -22808
rect 400890 -22864 400946 -22808
rect 401014 -22864 401070 -22808
rect 401138 -22864 401194 -22808
rect 401262 -22864 401318 -22808
rect 400766 -22988 400822 -22932
rect 400890 -22988 400946 -22932
rect 401014 -22988 401070 -22932
rect 401138 -22988 401194 -22932
rect 401262 -22988 401318 -22932
rect 400766 -23112 400822 -23056
rect 400890 -23112 400946 -23056
rect 401014 -23112 401070 -23056
rect 401138 -23112 401194 -23056
rect 401262 -23112 401318 -23056
rect 400766 -23236 400822 -23180
rect 400890 -23236 400946 -23180
rect 401014 -23236 401070 -23180
rect 401138 -23236 401194 -23180
rect 401262 -23236 401318 -23180
rect 400766 -23360 400822 -23304
rect 400890 -23360 400946 -23304
rect 401014 -23360 401070 -23304
rect 401138 -23360 401194 -23304
rect 401262 -23360 401318 -23304
rect 400766 -23484 400822 -23428
rect 400890 -23484 400946 -23428
rect 401014 -23484 401070 -23428
rect 401138 -23484 401194 -23428
rect 401262 -23484 401318 -23428
rect 400766 -23608 400822 -23552
rect 400890 -23608 400946 -23552
rect 401014 -23608 401070 -23552
rect 401138 -23608 401194 -23552
rect 401262 -23608 401318 -23552
rect 400766 -23732 400822 -23676
rect 400890 -23732 400946 -23676
rect 401014 -23732 401070 -23676
rect 401138 -23732 401194 -23676
rect 401262 -23732 401318 -23676
rect 400766 -23856 400822 -23800
rect 400890 -23856 400946 -23800
rect 401014 -23856 401070 -23800
rect 401138 -23856 401194 -23800
rect 401262 -23856 401318 -23800
rect 400766 -23980 400822 -23924
rect 400890 -23980 400946 -23924
rect 401014 -23980 401070 -23924
rect 401138 -23980 401194 -23924
rect 401262 -23980 401318 -23924
rect 400766 -24104 400822 -24048
rect 400890 -24104 400946 -24048
rect 401014 -24104 401070 -24048
rect 401138 -24104 401194 -24048
rect 401262 -24104 401318 -24048
rect 400766 -24228 400822 -24172
rect 400890 -24228 400946 -24172
rect 401014 -24228 401070 -24172
rect 401138 -24228 401194 -24172
rect 401262 -24228 401318 -24172
rect 400766 -24352 400822 -24296
rect 400890 -24352 400946 -24296
rect 401014 -24352 401070 -24296
rect 401138 -24352 401194 -24296
rect 401262 -24352 401318 -24296
rect 400766 -24476 400822 -24420
rect 400890 -24476 400946 -24420
rect 401014 -24476 401070 -24420
rect 401138 -24476 401194 -24420
rect 401262 -24476 401318 -24420
rect 400766 -24600 400822 -24544
rect 400890 -24600 400946 -24544
rect 401014 -24600 401070 -24544
rect 401138 -24600 401194 -24544
rect 401262 -24600 401318 -24544
rect 400766 -24724 400822 -24668
rect 400890 -24724 400946 -24668
rect 401014 -24724 401070 -24668
rect 401138 -24724 401194 -24668
rect 401262 -24724 401318 -24668
rect 400766 -24848 400822 -24792
rect 400890 -24848 400946 -24792
rect 401014 -24848 401070 -24792
rect 401138 -24848 401194 -24792
rect 401262 -24848 401318 -24792
rect 400766 -24972 400822 -24916
rect 400890 -24972 400946 -24916
rect 401014 -24972 401070 -24916
rect 401138 -24972 401194 -24916
rect 401262 -24972 401318 -24916
rect 400766 -25096 400822 -25040
rect 400890 -25096 400946 -25040
rect 401014 -25096 401070 -25040
rect 401138 -25096 401194 -25040
rect 401262 -25096 401318 -25040
rect 400766 -25220 400822 -25164
rect 400890 -25220 400946 -25164
rect 401014 -25220 401070 -25164
rect 401138 -25220 401194 -25164
rect 401262 -25220 401318 -25164
rect 400766 -25344 400822 -25288
rect 400890 -25344 400946 -25288
rect 401014 -25344 401070 -25288
rect 401138 -25344 401194 -25288
rect 401262 -25344 401318 -25288
rect 400766 -25468 400822 -25412
rect 400890 -25468 400946 -25412
rect 401014 -25468 401070 -25412
rect 401138 -25468 401194 -25412
rect 401262 -25468 401318 -25412
rect 387954 -25592 388010 -25536
rect 388078 -25592 388134 -25536
rect 388202 -25592 388258 -25536
rect 388326 -25592 388382 -25536
rect 388450 -25592 388506 -25536
rect 400766 -25592 400822 -25536
rect 400890 -25592 400946 -25536
rect 401014 -25592 401070 -25536
rect 401138 -25592 401194 -25536
rect 401262 -25592 401318 -25536
rect 387954 -25716 388010 -25660
rect 388078 -25716 388134 -25660
rect 388202 -25716 388258 -25660
rect 388326 -25716 388382 -25660
rect 388450 -25716 388506 -25660
rect 388655 -25744 388711 -25688
rect 388797 -25744 388853 -25688
rect 388939 -25744 388995 -25688
rect 389081 -25744 389137 -25688
rect 389223 -25744 389279 -25688
rect 389365 -25744 389421 -25688
rect 389507 -25744 389563 -25688
rect 389649 -25744 389705 -25688
rect 389791 -25744 389847 -25688
rect 389933 -25744 389989 -25688
rect 390075 -25744 390131 -25688
rect 390217 -25744 390273 -25688
rect 390359 -25744 390415 -25688
rect 390501 -25744 390557 -25688
rect 390643 -25744 390699 -25688
rect 390785 -25744 390841 -25688
rect 390927 -25744 390983 -25688
rect 391069 -25744 391125 -25688
rect 391211 -25744 391267 -25688
rect 391353 -25744 391409 -25688
rect 391495 -25744 391551 -25688
rect 391637 -25744 391693 -25688
rect 391779 -25744 391835 -25688
rect 391921 -25744 391977 -25688
rect 392063 -25744 392119 -25688
rect 392205 -25744 392261 -25688
rect 392347 -25744 392403 -25688
rect 392489 -25744 392545 -25688
rect 392631 -25744 392687 -25688
rect 392773 -25744 392829 -25688
rect 392915 -25744 392971 -25688
rect 393057 -25744 393113 -25688
rect 393199 -25744 393255 -25688
rect 393341 -25744 393397 -25688
rect 393483 -25744 393539 -25688
rect 393625 -25744 393681 -25688
rect 393767 -25744 393823 -25688
rect 393909 -25744 393965 -25688
rect 394051 -25744 394107 -25688
rect 394193 -25744 394249 -25688
rect 394335 -25744 394391 -25688
rect 394477 -25744 394533 -25688
rect 394619 -25744 394675 -25688
rect 394761 -25744 394817 -25688
rect 394903 -25744 394959 -25688
rect 395045 -25744 395101 -25688
rect 395187 -25744 395243 -25688
rect 395329 -25744 395385 -25688
rect 395471 -25744 395527 -25688
rect 395613 -25744 395669 -25688
rect 395755 -25744 395811 -25688
rect 395897 -25744 395953 -25688
rect 396039 -25744 396095 -25688
rect 396181 -25744 396237 -25688
rect 396323 -25744 396379 -25688
rect 396465 -25744 396521 -25688
rect 396607 -25744 396663 -25688
rect 396749 -25744 396805 -25688
rect 396891 -25744 396947 -25688
rect 397033 -25744 397089 -25688
rect 397175 -25744 397231 -25688
rect 397317 -25744 397373 -25688
rect 397459 -25744 397515 -25688
rect 397601 -25744 397657 -25688
rect 397743 -25744 397799 -25688
rect 397885 -25744 397941 -25688
rect 398027 -25744 398083 -25688
rect 398169 -25744 398225 -25688
rect 398311 -25744 398367 -25688
rect 398453 -25744 398509 -25688
rect 398595 -25744 398651 -25688
rect 398737 -25744 398793 -25688
rect 398879 -25744 398935 -25688
rect 399021 -25744 399077 -25688
rect 399163 -25744 399219 -25688
rect 399305 -25744 399361 -25688
rect 399447 -25744 399503 -25688
rect 399589 -25744 399645 -25688
rect 399731 -25744 399787 -25688
rect 399873 -25744 399929 -25688
rect 400015 -25744 400071 -25688
rect 400157 -25744 400213 -25688
rect 400299 -25744 400355 -25688
rect 400441 -25744 400497 -25688
rect 400583 -25744 400639 -25688
rect 400766 -25716 400822 -25660
rect 400890 -25716 400946 -25660
rect 401014 -25716 401070 -25660
rect 401138 -25716 401194 -25660
rect 401262 -25716 401318 -25660
rect 387954 -25840 388010 -25784
rect 388078 -25840 388134 -25784
rect 388202 -25840 388258 -25784
rect 388326 -25840 388382 -25784
rect 388450 -25840 388506 -25784
rect 388655 -25886 388711 -25830
rect 388797 -25886 388853 -25830
rect 388939 -25886 388995 -25830
rect 389081 -25886 389137 -25830
rect 389223 -25886 389279 -25830
rect 389365 -25886 389421 -25830
rect 389507 -25886 389563 -25830
rect 389649 -25886 389705 -25830
rect 389791 -25886 389847 -25830
rect 389933 -25886 389989 -25830
rect 390075 -25886 390131 -25830
rect 390217 -25886 390273 -25830
rect 390359 -25886 390415 -25830
rect 390501 -25886 390557 -25830
rect 390643 -25886 390699 -25830
rect 390785 -25886 390841 -25830
rect 390927 -25886 390983 -25830
rect 391069 -25886 391125 -25830
rect 391211 -25886 391267 -25830
rect 391353 -25886 391409 -25830
rect 391495 -25886 391551 -25830
rect 391637 -25886 391693 -25830
rect 391779 -25886 391835 -25830
rect 391921 -25886 391977 -25830
rect 392063 -25886 392119 -25830
rect 392205 -25886 392261 -25830
rect 392347 -25886 392403 -25830
rect 392489 -25886 392545 -25830
rect 392631 -25886 392687 -25830
rect 392773 -25886 392829 -25830
rect 392915 -25886 392971 -25830
rect 393057 -25886 393113 -25830
rect 393199 -25886 393255 -25830
rect 393341 -25886 393397 -25830
rect 393483 -25886 393539 -25830
rect 393625 -25886 393681 -25830
rect 393767 -25886 393823 -25830
rect 393909 -25886 393965 -25830
rect 394051 -25886 394107 -25830
rect 394193 -25886 394249 -25830
rect 394335 -25886 394391 -25830
rect 394477 -25886 394533 -25830
rect 394619 -25886 394675 -25830
rect 394761 -25886 394817 -25830
rect 394903 -25886 394959 -25830
rect 395045 -25886 395101 -25830
rect 395187 -25886 395243 -25830
rect 395329 -25886 395385 -25830
rect 395471 -25886 395527 -25830
rect 395613 -25886 395669 -25830
rect 395755 -25886 395811 -25830
rect 395897 -25886 395953 -25830
rect 396039 -25886 396095 -25830
rect 396181 -25886 396237 -25830
rect 396323 -25886 396379 -25830
rect 396465 -25886 396521 -25830
rect 396607 -25886 396663 -25830
rect 396749 -25886 396805 -25830
rect 396891 -25886 396947 -25830
rect 397033 -25886 397089 -25830
rect 397175 -25886 397231 -25830
rect 397317 -25886 397373 -25830
rect 397459 -25886 397515 -25830
rect 397601 -25886 397657 -25830
rect 397743 -25886 397799 -25830
rect 397885 -25886 397941 -25830
rect 398027 -25886 398083 -25830
rect 398169 -25886 398225 -25830
rect 398311 -25886 398367 -25830
rect 398453 -25886 398509 -25830
rect 398595 -25886 398651 -25830
rect 398737 -25886 398793 -25830
rect 398879 -25886 398935 -25830
rect 399021 -25886 399077 -25830
rect 399163 -25886 399219 -25830
rect 399305 -25886 399361 -25830
rect 399447 -25886 399503 -25830
rect 399589 -25886 399645 -25830
rect 399731 -25886 399787 -25830
rect 399873 -25886 399929 -25830
rect 400015 -25886 400071 -25830
rect 400157 -25886 400213 -25830
rect 400299 -25886 400355 -25830
rect 400441 -25886 400497 -25830
rect 400583 -25886 400639 -25830
rect 400766 -25840 400822 -25784
rect 400890 -25840 400946 -25784
rect 401014 -25840 401070 -25784
rect 401138 -25840 401194 -25784
rect 401262 -25840 401318 -25784
<< metal4 >>
rect 387840 -13041 401440 -12925
rect 387840 -13097 387986 -13041
rect 388042 -13097 388110 -13041
rect 388166 -13097 388234 -13041
rect 388290 -13097 388358 -13041
rect 388414 -13097 388482 -13041
rect 388538 -13097 388606 -13041
rect 388662 -13097 388730 -13041
rect 388786 -13097 388854 -13041
rect 388910 -13097 388978 -13041
rect 389034 -13097 389102 -13041
rect 389158 -13097 389226 -13041
rect 389282 -13097 389350 -13041
rect 389406 -13097 389474 -13041
rect 389530 -13097 389598 -13041
rect 389654 -13097 389722 -13041
rect 389778 -13097 389846 -13041
rect 389902 -13097 389970 -13041
rect 390026 -13097 390094 -13041
rect 390150 -13097 390218 -13041
rect 390274 -13097 390342 -13041
rect 390398 -13097 390466 -13041
rect 390522 -13097 390590 -13041
rect 390646 -13097 390714 -13041
rect 390770 -13097 390838 -13041
rect 390894 -13097 390962 -13041
rect 391018 -13097 391086 -13041
rect 391142 -13097 391210 -13041
rect 391266 -13097 391334 -13041
rect 391390 -13097 391458 -13041
rect 391514 -13097 391582 -13041
rect 391638 -13097 391706 -13041
rect 391762 -13097 391830 -13041
rect 391886 -13097 391954 -13041
rect 392010 -13097 392078 -13041
rect 392134 -13097 392202 -13041
rect 392258 -13097 392326 -13041
rect 392382 -13097 392450 -13041
rect 392506 -13097 392574 -13041
rect 392630 -13097 392698 -13041
rect 392754 -13097 392822 -13041
rect 392878 -13097 392946 -13041
rect 393002 -13097 393070 -13041
rect 393126 -13097 393194 -13041
rect 393250 -13097 393318 -13041
rect 393374 -13097 393442 -13041
rect 393498 -13097 393566 -13041
rect 393622 -13097 393690 -13041
rect 393746 -13097 393814 -13041
rect 393870 -13097 393938 -13041
rect 393994 -13097 394062 -13041
rect 394118 -13097 394186 -13041
rect 394242 -13097 394310 -13041
rect 394366 -13097 394434 -13041
rect 394490 -13097 394558 -13041
rect 394614 -13097 394682 -13041
rect 394738 -13097 394806 -13041
rect 394862 -13097 394930 -13041
rect 394986 -13097 395054 -13041
rect 395110 -13097 395178 -13041
rect 395234 -13097 395302 -13041
rect 395358 -13097 395426 -13041
rect 395482 -13097 395550 -13041
rect 395606 -13097 395674 -13041
rect 395730 -13097 395798 -13041
rect 395854 -13097 395922 -13041
rect 395978 -13097 396046 -13041
rect 396102 -13097 396170 -13041
rect 396226 -13097 396294 -13041
rect 396350 -13097 396418 -13041
rect 396474 -13097 396542 -13041
rect 396598 -13097 396666 -13041
rect 396722 -13097 396790 -13041
rect 396846 -13097 396914 -13041
rect 396970 -13097 397038 -13041
rect 397094 -13097 397162 -13041
rect 397218 -13097 397286 -13041
rect 397342 -13097 397410 -13041
rect 397466 -13097 397534 -13041
rect 397590 -13097 397658 -13041
rect 397714 -13097 397782 -13041
rect 397838 -13097 397906 -13041
rect 397962 -13097 398030 -13041
rect 398086 -13097 398154 -13041
rect 398210 -13097 398278 -13041
rect 398334 -13097 398402 -13041
rect 398458 -13097 398526 -13041
rect 398582 -13097 398650 -13041
rect 398706 -13097 398774 -13041
rect 398830 -13097 398898 -13041
rect 398954 -13097 399022 -13041
rect 399078 -13097 399146 -13041
rect 399202 -13097 399270 -13041
rect 399326 -13097 399394 -13041
rect 399450 -13097 399518 -13041
rect 399574 -13097 399642 -13041
rect 399698 -13097 399766 -13041
rect 399822 -13097 399890 -13041
rect 399946 -13097 400014 -13041
rect 400070 -13097 400138 -13041
rect 400194 -13097 400262 -13041
rect 400318 -13097 400386 -13041
rect 400442 -13097 400510 -13041
rect 400566 -13097 400634 -13041
rect 400690 -13097 400758 -13041
rect 400814 -13097 400882 -13041
rect 400938 -13097 401006 -13041
rect 401062 -13097 401130 -13041
rect 401186 -13097 401254 -13041
rect 401310 -13097 401440 -13041
rect 387840 -13165 401440 -13097
rect 387840 -13221 387986 -13165
rect 388042 -13221 388110 -13165
rect 388166 -13221 388234 -13165
rect 388290 -13221 388358 -13165
rect 388414 -13221 388482 -13165
rect 388538 -13221 388606 -13165
rect 388662 -13221 388730 -13165
rect 388786 -13221 388854 -13165
rect 388910 -13221 388978 -13165
rect 389034 -13221 389102 -13165
rect 389158 -13221 389226 -13165
rect 389282 -13221 389350 -13165
rect 389406 -13221 389474 -13165
rect 389530 -13221 389598 -13165
rect 389654 -13221 389722 -13165
rect 389778 -13221 389846 -13165
rect 389902 -13221 389970 -13165
rect 390026 -13221 390094 -13165
rect 390150 -13221 390218 -13165
rect 390274 -13221 390342 -13165
rect 390398 -13221 390466 -13165
rect 390522 -13221 390590 -13165
rect 390646 -13221 390714 -13165
rect 390770 -13221 390838 -13165
rect 390894 -13221 390962 -13165
rect 391018 -13221 391086 -13165
rect 391142 -13221 391210 -13165
rect 391266 -13221 391334 -13165
rect 391390 -13221 391458 -13165
rect 391514 -13221 391582 -13165
rect 391638 -13221 391706 -13165
rect 391762 -13221 391830 -13165
rect 391886 -13221 391954 -13165
rect 392010 -13221 392078 -13165
rect 392134 -13221 392202 -13165
rect 392258 -13221 392326 -13165
rect 392382 -13221 392450 -13165
rect 392506 -13221 392574 -13165
rect 392630 -13221 392698 -13165
rect 392754 -13221 392822 -13165
rect 392878 -13221 392946 -13165
rect 393002 -13221 393070 -13165
rect 393126 -13221 393194 -13165
rect 393250 -13221 393318 -13165
rect 393374 -13221 393442 -13165
rect 393498 -13221 393566 -13165
rect 393622 -13221 393690 -13165
rect 393746 -13221 393814 -13165
rect 393870 -13221 393938 -13165
rect 393994 -13221 394062 -13165
rect 394118 -13221 394186 -13165
rect 394242 -13221 394310 -13165
rect 394366 -13221 394434 -13165
rect 394490 -13221 394558 -13165
rect 394614 -13221 394682 -13165
rect 394738 -13221 394806 -13165
rect 394862 -13221 394930 -13165
rect 394986 -13221 395054 -13165
rect 395110 -13221 395178 -13165
rect 395234 -13221 395302 -13165
rect 395358 -13221 395426 -13165
rect 395482 -13221 395550 -13165
rect 395606 -13221 395674 -13165
rect 395730 -13221 395798 -13165
rect 395854 -13221 395922 -13165
rect 395978 -13221 396046 -13165
rect 396102 -13221 396170 -13165
rect 396226 -13221 396294 -13165
rect 396350 -13221 396418 -13165
rect 396474 -13221 396542 -13165
rect 396598 -13221 396666 -13165
rect 396722 -13221 396790 -13165
rect 396846 -13221 396914 -13165
rect 396970 -13221 397038 -13165
rect 397094 -13221 397162 -13165
rect 397218 -13221 397286 -13165
rect 397342 -13221 397410 -13165
rect 397466 -13221 397534 -13165
rect 397590 -13221 397658 -13165
rect 397714 -13221 397782 -13165
rect 397838 -13221 397906 -13165
rect 397962 -13221 398030 -13165
rect 398086 -13221 398154 -13165
rect 398210 -13221 398278 -13165
rect 398334 -13221 398402 -13165
rect 398458 -13221 398526 -13165
rect 398582 -13221 398650 -13165
rect 398706 -13221 398774 -13165
rect 398830 -13221 398898 -13165
rect 398954 -13221 399022 -13165
rect 399078 -13221 399146 -13165
rect 399202 -13221 399270 -13165
rect 399326 -13221 399394 -13165
rect 399450 -13221 399518 -13165
rect 399574 -13221 399642 -13165
rect 399698 -13221 399766 -13165
rect 399822 -13221 399890 -13165
rect 399946 -13221 400014 -13165
rect 400070 -13221 400138 -13165
rect 400194 -13221 400262 -13165
rect 400318 -13221 400386 -13165
rect 400442 -13221 400510 -13165
rect 400566 -13221 400634 -13165
rect 400690 -13221 400758 -13165
rect 400814 -13221 400882 -13165
rect 400938 -13221 401006 -13165
rect 401062 -13221 401130 -13165
rect 401186 -13221 401254 -13165
rect 401310 -13221 401440 -13165
rect 387840 -13289 401440 -13221
rect 387840 -13345 387986 -13289
rect 388042 -13345 388110 -13289
rect 388166 -13345 388234 -13289
rect 388290 -13345 388358 -13289
rect 388414 -13345 388482 -13289
rect 388538 -13345 388606 -13289
rect 388662 -13345 388730 -13289
rect 388786 -13345 388854 -13289
rect 388910 -13345 388978 -13289
rect 389034 -13345 389102 -13289
rect 389158 -13345 389226 -13289
rect 389282 -13345 389350 -13289
rect 389406 -13345 389474 -13289
rect 389530 -13345 389598 -13289
rect 389654 -13345 389722 -13289
rect 389778 -13345 389846 -13289
rect 389902 -13345 389970 -13289
rect 390026 -13345 390094 -13289
rect 390150 -13345 390218 -13289
rect 390274 -13345 390342 -13289
rect 390398 -13345 390466 -13289
rect 390522 -13345 390590 -13289
rect 390646 -13345 390714 -13289
rect 390770 -13345 390838 -13289
rect 390894 -13345 390962 -13289
rect 391018 -13345 391086 -13289
rect 391142 -13345 391210 -13289
rect 391266 -13345 391334 -13289
rect 391390 -13345 391458 -13289
rect 391514 -13345 391582 -13289
rect 391638 -13345 391706 -13289
rect 391762 -13345 391830 -13289
rect 391886 -13345 391954 -13289
rect 392010 -13345 392078 -13289
rect 392134 -13345 392202 -13289
rect 392258 -13345 392326 -13289
rect 392382 -13345 392450 -13289
rect 392506 -13345 392574 -13289
rect 392630 -13345 392698 -13289
rect 392754 -13345 392822 -13289
rect 392878 -13345 392946 -13289
rect 393002 -13345 393070 -13289
rect 393126 -13345 393194 -13289
rect 393250 -13345 393318 -13289
rect 393374 -13345 393442 -13289
rect 393498 -13345 393566 -13289
rect 393622 -13345 393690 -13289
rect 393746 -13345 393814 -13289
rect 393870 -13345 393938 -13289
rect 393994 -13345 394062 -13289
rect 394118 -13345 394186 -13289
rect 394242 -13345 394310 -13289
rect 394366 -13345 394434 -13289
rect 394490 -13345 394558 -13289
rect 394614 -13345 394682 -13289
rect 394738 -13345 394806 -13289
rect 394862 -13345 394930 -13289
rect 394986 -13345 395054 -13289
rect 395110 -13345 395178 -13289
rect 395234 -13345 395302 -13289
rect 395358 -13345 395426 -13289
rect 395482 -13345 395550 -13289
rect 395606 -13345 395674 -13289
rect 395730 -13345 395798 -13289
rect 395854 -13345 395922 -13289
rect 395978 -13345 396046 -13289
rect 396102 -13345 396170 -13289
rect 396226 -13345 396294 -13289
rect 396350 -13345 396418 -13289
rect 396474 -13345 396542 -13289
rect 396598 -13345 396666 -13289
rect 396722 -13345 396790 -13289
rect 396846 -13345 396914 -13289
rect 396970 -13345 397038 -13289
rect 397094 -13345 397162 -13289
rect 397218 -13345 397286 -13289
rect 397342 -13345 397410 -13289
rect 397466 -13345 397534 -13289
rect 397590 -13345 397658 -13289
rect 397714 -13345 397782 -13289
rect 397838 -13345 397906 -13289
rect 397962 -13345 398030 -13289
rect 398086 -13345 398154 -13289
rect 398210 -13345 398278 -13289
rect 398334 -13345 398402 -13289
rect 398458 -13345 398526 -13289
rect 398582 -13345 398650 -13289
rect 398706 -13345 398774 -13289
rect 398830 -13345 398898 -13289
rect 398954 -13345 399022 -13289
rect 399078 -13345 399146 -13289
rect 399202 -13345 399270 -13289
rect 399326 -13345 399394 -13289
rect 399450 -13345 399518 -13289
rect 399574 -13345 399642 -13289
rect 399698 -13345 399766 -13289
rect 399822 -13345 399890 -13289
rect 399946 -13345 400014 -13289
rect 400070 -13345 400138 -13289
rect 400194 -13345 400262 -13289
rect 400318 -13345 400386 -13289
rect 400442 -13345 400510 -13289
rect 400566 -13345 400634 -13289
rect 400690 -13345 400758 -13289
rect 400814 -13345 400882 -13289
rect 400938 -13345 401006 -13289
rect 401062 -13345 401130 -13289
rect 401186 -13345 401254 -13289
rect 401310 -13345 401440 -13289
rect 387840 -13413 401440 -13345
rect 387840 -13469 387986 -13413
rect 388042 -13469 388110 -13413
rect 388166 -13469 388234 -13413
rect 388290 -13469 388358 -13413
rect 388414 -13469 388482 -13413
rect 388538 -13469 388606 -13413
rect 388662 -13469 388730 -13413
rect 388786 -13469 388854 -13413
rect 388910 -13469 388978 -13413
rect 389034 -13469 389102 -13413
rect 389158 -13469 389226 -13413
rect 389282 -13469 389350 -13413
rect 389406 -13469 389474 -13413
rect 389530 -13469 389598 -13413
rect 389654 -13469 389722 -13413
rect 389778 -13469 389846 -13413
rect 389902 -13469 389970 -13413
rect 390026 -13469 390094 -13413
rect 390150 -13469 390218 -13413
rect 390274 -13469 390342 -13413
rect 390398 -13469 390466 -13413
rect 390522 -13469 390590 -13413
rect 390646 -13469 390714 -13413
rect 390770 -13469 390838 -13413
rect 390894 -13469 390962 -13413
rect 391018 -13469 391086 -13413
rect 391142 -13469 391210 -13413
rect 391266 -13469 391334 -13413
rect 391390 -13469 391458 -13413
rect 391514 -13469 391582 -13413
rect 391638 -13469 391706 -13413
rect 391762 -13469 391830 -13413
rect 391886 -13469 391954 -13413
rect 392010 -13469 392078 -13413
rect 392134 -13469 392202 -13413
rect 392258 -13469 392326 -13413
rect 392382 -13469 392450 -13413
rect 392506 -13469 392574 -13413
rect 392630 -13469 392698 -13413
rect 392754 -13469 392822 -13413
rect 392878 -13469 392946 -13413
rect 393002 -13469 393070 -13413
rect 393126 -13469 393194 -13413
rect 393250 -13469 393318 -13413
rect 393374 -13469 393442 -13413
rect 393498 -13469 393566 -13413
rect 393622 -13469 393690 -13413
rect 393746 -13469 393814 -13413
rect 393870 -13469 393938 -13413
rect 393994 -13469 394062 -13413
rect 394118 -13469 394186 -13413
rect 394242 -13469 394310 -13413
rect 394366 -13469 394434 -13413
rect 394490 -13469 394558 -13413
rect 394614 -13469 394682 -13413
rect 394738 -13469 394806 -13413
rect 394862 -13469 394930 -13413
rect 394986 -13469 395054 -13413
rect 395110 -13469 395178 -13413
rect 395234 -13469 395302 -13413
rect 395358 -13469 395426 -13413
rect 395482 -13469 395550 -13413
rect 395606 -13469 395674 -13413
rect 395730 -13469 395798 -13413
rect 395854 -13469 395922 -13413
rect 395978 -13469 396046 -13413
rect 396102 -13469 396170 -13413
rect 396226 -13469 396294 -13413
rect 396350 -13469 396418 -13413
rect 396474 -13469 396542 -13413
rect 396598 -13469 396666 -13413
rect 396722 -13469 396790 -13413
rect 396846 -13469 396914 -13413
rect 396970 -13469 397038 -13413
rect 397094 -13469 397162 -13413
rect 397218 -13469 397286 -13413
rect 397342 -13469 397410 -13413
rect 397466 -13469 397534 -13413
rect 397590 -13469 397658 -13413
rect 397714 -13469 397782 -13413
rect 397838 -13469 397906 -13413
rect 397962 -13469 398030 -13413
rect 398086 -13469 398154 -13413
rect 398210 -13469 398278 -13413
rect 398334 -13469 398402 -13413
rect 398458 -13469 398526 -13413
rect 398582 -13469 398650 -13413
rect 398706 -13469 398774 -13413
rect 398830 -13469 398898 -13413
rect 398954 -13469 399022 -13413
rect 399078 -13469 399146 -13413
rect 399202 -13469 399270 -13413
rect 399326 -13469 399394 -13413
rect 399450 -13469 399518 -13413
rect 399574 -13469 399642 -13413
rect 399698 -13469 399766 -13413
rect 399822 -13469 399890 -13413
rect 399946 -13469 400014 -13413
rect 400070 -13469 400138 -13413
rect 400194 -13469 400262 -13413
rect 400318 -13469 400386 -13413
rect 400442 -13469 400510 -13413
rect 400566 -13469 400634 -13413
rect 400690 -13469 400758 -13413
rect 400814 -13469 400882 -13413
rect 400938 -13469 401006 -13413
rect 401062 -13469 401130 -13413
rect 401186 -13469 401254 -13413
rect 401310 -13469 401440 -13413
rect 387840 -13632 401440 -13469
rect 387840 -13688 387954 -13632
rect 388010 -13688 388078 -13632
rect 388134 -13688 388202 -13632
rect 388258 -13688 388326 -13632
rect 388382 -13688 388450 -13632
rect 388506 -13670 400766 -13632
rect 388506 -13688 388640 -13670
rect 387840 -13756 388640 -13688
rect 387840 -13812 387954 -13756
rect 388010 -13812 388078 -13756
rect 388134 -13812 388202 -13756
rect 388258 -13812 388326 -13756
rect 388382 -13812 388450 -13756
rect 388506 -13812 388640 -13756
rect 387840 -13880 388640 -13812
rect 387840 -13936 387954 -13880
rect 388010 -13936 388078 -13880
rect 388134 -13936 388202 -13880
rect 388258 -13936 388326 -13880
rect 388382 -13936 388450 -13880
rect 388506 -13936 388640 -13880
rect 387840 -14004 388640 -13936
rect 387840 -14060 387954 -14004
rect 388010 -14060 388078 -14004
rect 388134 -14060 388202 -14004
rect 388258 -14060 388326 -14004
rect 388382 -14060 388450 -14004
rect 388506 -14060 388640 -14004
rect 387840 -14128 388640 -14060
rect 387840 -14184 387954 -14128
rect 388010 -14184 388078 -14128
rect 388134 -14184 388202 -14128
rect 388258 -14184 388326 -14128
rect 388382 -14184 388450 -14128
rect 388506 -14184 388640 -14128
rect 387840 -14252 388640 -14184
rect 387840 -14308 387954 -14252
rect 388010 -14308 388078 -14252
rect 388134 -14308 388202 -14252
rect 388258 -14308 388326 -14252
rect 388382 -14308 388450 -14252
rect 388506 -14308 388640 -14252
rect 387840 -14376 388640 -14308
rect 387840 -14432 387954 -14376
rect 388010 -14432 388078 -14376
rect 388134 -14432 388202 -14376
rect 388258 -14432 388326 -14376
rect 388382 -14432 388450 -14376
rect 388506 -14432 388640 -14376
rect 387840 -14500 388640 -14432
rect 387840 -14556 387954 -14500
rect 388010 -14556 388078 -14500
rect 388134 -14556 388202 -14500
rect 388258 -14556 388326 -14500
rect 388382 -14556 388450 -14500
rect 388506 -14556 388640 -14500
rect 387840 -14624 388640 -14556
rect 387840 -14680 387954 -14624
rect 388010 -14680 388078 -14624
rect 388134 -14680 388202 -14624
rect 388258 -14680 388326 -14624
rect 388382 -14680 388450 -14624
rect 388506 -14680 388640 -14624
rect 387840 -14748 388640 -14680
rect 387840 -14804 387954 -14748
rect 388010 -14804 388078 -14748
rect 388134 -14804 388202 -14748
rect 388258 -14804 388326 -14748
rect 388382 -14804 388450 -14748
rect 388506 -14804 388640 -14748
rect 387840 -14872 388640 -14804
rect 387840 -14928 387954 -14872
rect 388010 -14928 388078 -14872
rect 388134 -14928 388202 -14872
rect 388258 -14928 388326 -14872
rect 388382 -14928 388450 -14872
rect 388506 -14928 388640 -14872
rect 387840 -14996 388640 -14928
rect 387840 -15052 387954 -14996
rect 388010 -15052 388078 -14996
rect 388134 -15052 388202 -14996
rect 388258 -15052 388326 -14996
rect 388382 -15052 388450 -14996
rect 388506 -15052 388640 -14996
rect 387840 -15120 388640 -15052
rect 387840 -15176 387954 -15120
rect 388010 -15176 388078 -15120
rect 388134 -15176 388202 -15120
rect 388258 -15176 388326 -15120
rect 388382 -15176 388450 -15120
rect 388506 -15176 388640 -15120
rect 387840 -15244 388640 -15176
rect 387840 -15300 387954 -15244
rect 388010 -15300 388078 -15244
rect 388134 -15300 388202 -15244
rect 388258 -15300 388326 -15244
rect 388382 -15300 388450 -15244
rect 388506 -15300 388640 -15244
rect 387840 -15368 388640 -15300
rect 387840 -15424 387954 -15368
rect 388010 -15424 388078 -15368
rect 388134 -15424 388202 -15368
rect 388258 -15424 388326 -15368
rect 388382 -15424 388450 -15368
rect 388506 -15424 388640 -15368
rect 387840 -15492 388640 -15424
rect 387840 -15548 387954 -15492
rect 388010 -15548 388078 -15492
rect 388134 -15548 388202 -15492
rect 388258 -15548 388326 -15492
rect 388382 -15548 388450 -15492
rect 388506 -15548 388640 -15492
rect 387840 -15616 388640 -15548
rect 387840 -15672 387954 -15616
rect 388010 -15672 388078 -15616
rect 388134 -15672 388202 -15616
rect 388258 -15672 388326 -15616
rect 388382 -15672 388450 -15616
rect 388506 -15672 388640 -15616
rect 387840 -15740 388640 -15672
rect 387840 -15796 387954 -15740
rect 388010 -15796 388078 -15740
rect 388134 -15796 388202 -15740
rect 388258 -15796 388326 -15740
rect 388382 -15796 388450 -15740
rect 388506 -15796 388640 -15740
rect 387840 -15864 388640 -15796
rect 387840 -15920 387954 -15864
rect 388010 -15920 388078 -15864
rect 388134 -15920 388202 -15864
rect 388258 -15920 388326 -15864
rect 388382 -15920 388450 -15864
rect 388506 -15920 388640 -15864
rect 387840 -15988 388640 -15920
rect 387840 -16044 387954 -15988
rect 388010 -16044 388078 -15988
rect 388134 -16044 388202 -15988
rect 388258 -16044 388326 -15988
rect 388382 -16044 388450 -15988
rect 388506 -16044 388640 -15988
rect 387840 -16112 388640 -16044
rect 387840 -16168 387954 -16112
rect 388010 -16168 388078 -16112
rect 388134 -16168 388202 -16112
rect 388258 -16168 388326 -16112
rect 388382 -16168 388450 -16112
rect 388506 -16168 388640 -16112
rect 387840 -16236 388640 -16168
rect 387840 -16292 387954 -16236
rect 388010 -16292 388078 -16236
rect 388134 -16292 388202 -16236
rect 388258 -16292 388326 -16236
rect 388382 -16292 388450 -16236
rect 388506 -16292 388640 -16236
rect 387840 -16360 388640 -16292
rect 387840 -16416 387954 -16360
rect 388010 -16416 388078 -16360
rect 388134 -16416 388202 -16360
rect 388258 -16416 388326 -16360
rect 388382 -16416 388450 -16360
rect 388506 -16416 388640 -16360
rect 387840 -16484 388640 -16416
rect 387840 -16540 387954 -16484
rect 388010 -16540 388078 -16484
rect 388134 -16540 388202 -16484
rect 388258 -16540 388326 -16484
rect 388382 -16540 388450 -16484
rect 388506 -16540 388640 -16484
rect 387840 -16608 388640 -16540
rect 387840 -16664 387954 -16608
rect 388010 -16664 388078 -16608
rect 388134 -16664 388202 -16608
rect 388258 -16664 388326 -16608
rect 388382 -16664 388450 -16608
rect 388506 -16664 388640 -16608
rect 387840 -16732 388640 -16664
rect 387840 -16788 387954 -16732
rect 388010 -16788 388078 -16732
rect 388134 -16788 388202 -16732
rect 388258 -16788 388326 -16732
rect 388382 -16788 388450 -16732
rect 388506 -16788 388640 -16732
rect 387840 -16856 388640 -16788
rect 387840 -16912 387954 -16856
rect 388010 -16912 388078 -16856
rect 388134 -16912 388202 -16856
rect 388258 -16912 388326 -16856
rect 388382 -16912 388450 -16856
rect 388506 -16912 388640 -16856
rect 387840 -16980 388640 -16912
rect 387840 -17036 387954 -16980
rect 388010 -17036 388078 -16980
rect 388134 -17036 388202 -16980
rect 388258 -17036 388326 -16980
rect 388382 -17036 388450 -16980
rect 388506 -17036 388640 -16980
rect 387840 -17104 388640 -17036
rect 387840 -17160 387954 -17104
rect 388010 -17160 388078 -17104
rect 388134 -17160 388202 -17104
rect 388258 -17160 388326 -17104
rect 388382 -17160 388450 -17104
rect 388506 -17160 388640 -17104
rect 387840 -17228 388640 -17160
rect 387840 -17284 387954 -17228
rect 388010 -17284 388078 -17228
rect 388134 -17284 388202 -17228
rect 388258 -17284 388326 -17228
rect 388382 -17284 388450 -17228
rect 388506 -17284 388640 -17228
rect 387840 -17352 388640 -17284
rect 387840 -17408 387954 -17352
rect 388010 -17408 388078 -17352
rect 388134 -17408 388202 -17352
rect 388258 -17408 388326 -17352
rect 388382 -17408 388450 -17352
rect 388506 -17408 388640 -17352
rect 387840 -17476 388640 -17408
rect 387840 -17532 387954 -17476
rect 388010 -17532 388078 -17476
rect 388134 -17532 388202 -17476
rect 388258 -17532 388326 -17476
rect 388382 -17532 388450 -17476
rect 388506 -17532 388640 -17476
rect 387840 -17600 388640 -17532
rect 387840 -17656 387954 -17600
rect 388010 -17656 388078 -17600
rect 388134 -17656 388202 -17600
rect 388258 -17656 388326 -17600
rect 388382 -17656 388450 -17600
rect 388506 -17656 388640 -17600
rect 387840 -17724 388640 -17656
rect 387840 -17780 387954 -17724
rect 388010 -17780 388078 -17724
rect 388134 -17780 388202 -17724
rect 388258 -17780 388326 -17724
rect 388382 -17780 388450 -17724
rect 388506 -17780 388640 -17724
rect 387840 -17848 388640 -17780
rect 387840 -17904 387954 -17848
rect 388010 -17904 388078 -17848
rect 388134 -17904 388202 -17848
rect 388258 -17904 388326 -17848
rect 388382 -17904 388450 -17848
rect 388506 -17904 388640 -17848
rect 387840 -17972 388640 -17904
rect 387840 -18028 387954 -17972
rect 388010 -18028 388078 -17972
rect 388134 -18028 388202 -17972
rect 388258 -18028 388326 -17972
rect 388382 -18028 388450 -17972
rect 388506 -18028 388640 -17972
rect 387840 -18096 388640 -18028
rect 387840 -18152 387954 -18096
rect 388010 -18152 388078 -18096
rect 388134 -18152 388202 -18096
rect 388258 -18152 388326 -18096
rect 388382 -18152 388450 -18096
rect 388506 -18152 388640 -18096
rect 387840 -18220 388640 -18152
rect 387840 -18276 387954 -18220
rect 388010 -18276 388078 -18220
rect 388134 -18276 388202 -18220
rect 388258 -18276 388326 -18220
rect 388382 -18276 388450 -18220
rect 388506 -18276 388640 -18220
rect 387840 -18344 388640 -18276
rect 387840 -18400 387954 -18344
rect 388010 -18400 388078 -18344
rect 388134 -18400 388202 -18344
rect 388258 -18400 388326 -18344
rect 388382 -18400 388450 -18344
rect 388506 -18400 388640 -18344
rect 387840 -18468 388640 -18400
rect 387840 -18524 387954 -18468
rect 388010 -18524 388078 -18468
rect 388134 -18524 388202 -18468
rect 388258 -18524 388326 -18468
rect 388382 -18524 388450 -18468
rect 388506 -18524 388640 -18468
rect 387840 -18592 388640 -18524
rect 387840 -18648 387954 -18592
rect 388010 -18648 388078 -18592
rect 388134 -18648 388202 -18592
rect 388258 -18648 388326 -18592
rect 388382 -18648 388450 -18592
rect 388506 -18648 388640 -18592
rect 387840 -18716 388640 -18648
rect 387840 -18772 387954 -18716
rect 388010 -18772 388078 -18716
rect 388134 -18772 388202 -18716
rect 388258 -18772 388326 -18716
rect 388382 -18772 388450 -18716
rect 388506 -18772 388640 -18716
rect 387840 -18840 388640 -18772
rect 387840 -18896 387954 -18840
rect 388010 -18896 388078 -18840
rect 388134 -18896 388202 -18840
rect 388258 -18896 388326 -18840
rect 388382 -18896 388450 -18840
rect 388506 -18896 388640 -18840
rect 387840 -18964 388640 -18896
rect 387840 -19020 387954 -18964
rect 388010 -19020 388078 -18964
rect 388134 -19020 388202 -18964
rect 388258 -19020 388326 -18964
rect 388382 -19020 388450 -18964
rect 388506 -19020 388640 -18964
rect 387840 -19088 388640 -19020
rect 387840 -19144 387954 -19088
rect 388010 -19144 388078 -19088
rect 388134 -19144 388202 -19088
rect 388258 -19144 388326 -19088
rect 388382 -19144 388450 -19088
rect 388506 -19144 388640 -19088
rect 387840 -19212 388640 -19144
rect 387840 -19268 387954 -19212
rect 388010 -19268 388078 -19212
rect 388134 -19268 388202 -19212
rect 388258 -19268 388326 -19212
rect 388382 -19268 388450 -19212
rect 388506 -19268 388640 -19212
rect 387840 -19336 388640 -19268
rect 387840 -19392 387954 -19336
rect 388010 -19392 388078 -19336
rect 388134 -19392 388202 -19336
rect 388258 -19392 388326 -19336
rect 388382 -19392 388450 -19336
rect 388506 -19392 388640 -19336
rect 387840 -19460 388640 -19392
rect 387840 -19516 387954 -19460
rect 388010 -19516 388078 -19460
rect 388134 -19516 388202 -19460
rect 388258 -19516 388326 -19460
rect 388382 -19516 388450 -19460
rect 388506 -19516 388640 -19460
rect 387840 -19584 388640 -19516
rect 387840 -19640 387954 -19584
rect 388010 -19640 388078 -19584
rect 388134 -19640 388202 -19584
rect 388258 -19640 388326 -19584
rect 388382 -19640 388450 -19584
rect 388506 -19640 388640 -19584
rect 387840 -19708 388640 -19640
rect 387840 -19764 387954 -19708
rect 388010 -19764 388078 -19708
rect 388134 -19764 388202 -19708
rect 388258 -19764 388326 -19708
rect 388382 -19764 388450 -19708
rect 388506 -19764 388640 -19708
rect 387840 -19832 388640 -19764
rect 387840 -19888 387954 -19832
rect 388010 -19888 388078 -19832
rect 388134 -19888 388202 -19832
rect 388258 -19888 388326 -19832
rect 388382 -19888 388450 -19832
rect 388506 -19888 388640 -19832
rect 387840 -19956 388640 -19888
rect 387840 -20012 387954 -19956
rect 388010 -20012 388078 -19956
rect 388134 -20012 388202 -19956
rect 388258 -20012 388326 -19956
rect 388382 -20012 388450 -19956
rect 388506 -20012 388640 -19956
rect 387840 -20080 388640 -20012
rect 387840 -20136 387954 -20080
rect 388010 -20136 388078 -20080
rect 388134 -20136 388202 -20080
rect 388258 -20136 388326 -20080
rect 388382 -20136 388450 -20080
rect 388506 -20136 388640 -20080
rect 387840 -20204 388640 -20136
rect 387840 -20260 387954 -20204
rect 388010 -20260 388078 -20204
rect 388134 -20260 388202 -20204
rect 388258 -20260 388326 -20204
rect 388382 -20260 388450 -20204
rect 388506 -20260 388640 -20204
rect 387840 -20328 388640 -20260
rect 387840 -20384 387954 -20328
rect 388010 -20384 388078 -20328
rect 388134 -20384 388202 -20328
rect 388258 -20384 388326 -20328
rect 388382 -20384 388450 -20328
rect 388506 -20384 388640 -20328
rect 387840 -20452 388640 -20384
rect 387840 -20508 387954 -20452
rect 388010 -20508 388078 -20452
rect 388134 -20508 388202 -20452
rect 388258 -20508 388326 -20452
rect 388382 -20508 388450 -20452
rect 388506 -20508 388640 -20452
rect 387840 -20576 388640 -20508
rect 387840 -20632 387954 -20576
rect 388010 -20632 388078 -20576
rect 388134 -20632 388202 -20576
rect 388258 -20632 388326 -20576
rect 388382 -20632 388450 -20576
rect 388506 -20632 388640 -20576
rect 387840 -20700 388640 -20632
rect 387840 -20756 387954 -20700
rect 388010 -20756 388078 -20700
rect 388134 -20756 388202 -20700
rect 388258 -20756 388326 -20700
rect 388382 -20756 388450 -20700
rect 388506 -20756 388640 -20700
rect 387840 -20824 388640 -20756
rect 387840 -20880 387954 -20824
rect 388010 -20880 388078 -20824
rect 388134 -20880 388202 -20824
rect 388258 -20880 388326 -20824
rect 388382 -20880 388450 -20824
rect 388506 -20880 388640 -20824
rect 387840 -20948 388640 -20880
rect 387840 -21004 387954 -20948
rect 388010 -21004 388078 -20948
rect 388134 -21004 388202 -20948
rect 388258 -21004 388326 -20948
rect 388382 -21004 388450 -20948
rect 388506 -21004 388640 -20948
rect 387840 -21072 388640 -21004
rect 387840 -21128 387954 -21072
rect 388010 -21128 388078 -21072
rect 388134 -21128 388202 -21072
rect 388258 -21128 388326 -21072
rect 388382 -21128 388450 -21072
rect 388506 -21128 388640 -21072
rect 387840 -21196 388640 -21128
rect 387840 -21252 387954 -21196
rect 388010 -21252 388078 -21196
rect 388134 -21252 388202 -21196
rect 388258 -21252 388326 -21196
rect 388382 -21252 388450 -21196
rect 388506 -21252 388640 -21196
rect 387840 -21320 388640 -21252
rect 387840 -21376 387954 -21320
rect 388010 -21376 388078 -21320
rect 388134 -21376 388202 -21320
rect 388258 -21376 388326 -21320
rect 388382 -21376 388450 -21320
rect 388506 -21376 388640 -21320
rect 387840 -21444 388640 -21376
rect 387840 -21500 387954 -21444
rect 388010 -21500 388078 -21444
rect 388134 -21500 388202 -21444
rect 388258 -21500 388326 -21444
rect 388382 -21500 388450 -21444
rect 388506 -21500 388640 -21444
rect 387840 -21568 388640 -21500
rect 387840 -21624 387954 -21568
rect 388010 -21624 388078 -21568
rect 388134 -21624 388202 -21568
rect 388258 -21624 388326 -21568
rect 388382 -21624 388450 -21568
rect 388506 -21624 388640 -21568
rect 387840 -21692 388640 -21624
rect 387840 -21748 387954 -21692
rect 388010 -21748 388078 -21692
rect 388134 -21748 388202 -21692
rect 388258 -21748 388326 -21692
rect 388382 -21748 388450 -21692
rect 388506 -21748 388640 -21692
rect 387840 -21816 388640 -21748
rect 387840 -21872 387954 -21816
rect 388010 -21872 388078 -21816
rect 388134 -21872 388202 -21816
rect 388258 -21872 388326 -21816
rect 388382 -21872 388450 -21816
rect 388506 -21872 388640 -21816
rect 387840 -21940 388640 -21872
rect 387840 -21996 387954 -21940
rect 388010 -21996 388078 -21940
rect 388134 -21996 388202 -21940
rect 388258 -21996 388326 -21940
rect 388382 -21996 388450 -21940
rect 388506 -21996 388640 -21940
rect 387840 -22064 388640 -21996
rect 387840 -22120 387954 -22064
rect 388010 -22120 388078 -22064
rect 388134 -22120 388202 -22064
rect 388258 -22120 388326 -22064
rect 388382 -22120 388450 -22064
rect 388506 -22120 388640 -22064
rect 387840 -22188 388640 -22120
rect 387840 -22244 387954 -22188
rect 388010 -22244 388078 -22188
rect 388134 -22244 388202 -22188
rect 388258 -22244 388326 -22188
rect 388382 -22244 388450 -22188
rect 388506 -22244 388640 -22188
rect 387840 -22312 388640 -22244
rect 387840 -22368 387954 -22312
rect 388010 -22368 388078 -22312
rect 388134 -22368 388202 -22312
rect 388258 -22368 388326 -22312
rect 388382 -22368 388450 -22312
rect 388506 -22368 388640 -22312
rect 387840 -22436 388640 -22368
rect 387840 -22492 387954 -22436
rect 388010 -22492 388078 -22436
rect 388134 -22492 388202 -22436
rect 388258 -22492 388326 -22436
rect 388382 -22492 388450 -22436
rect 388506 -22492 388640 -22436
rect 387840 -22560 388640 -22492
rect 387840 -22616 387954 -22560
rect 388010 -22616 388078 -22560
rect 388134 -22616 388202 -22560
rect 388258 -22616 388326 -22560
rect 388382 -22616 388450 -22560
rect 388506 -22616 388640 -22560
rect 387840 -22684 388640 -22616
rect 387840 -22740 387954 -22684
rect 388010 -22740 388078 -22684
rect 388134 -22740 388202 -22684
rect 388258 -22740 388326 -22684
rect 388382 -22740 388450 -22684
rect 388506 -22740 388640 -22684
rect 387840 -22808 388640 -22740
rect 387840 -22864 387954 -22808
rect 388010 -22864 388078 -22808
rect 388134 -22864 388202 -22808
rect 388258 -22864 388326 -22808
rect 388382 -22864 388450 -22808
rect 388506 -22864 388640 -22808
rect 387840 -22932 388640 -22864
rect 387840 -22988 387954 -22932
rect 388010 -22988 388078 -22932
rect 388134 -22988 388202 -22932
rect 388258 -22988 388326 -22932
rect 388382 -22988 388450 -22932
rect 388506 -22988 388640 -22932
rect 387840 -23056 388640 -22988
rect 387840 -23112 387954 -23056
rect 388010 -23112 388078 -23056
rect 388134 -23112 388202 -23056
rect 388258 -23112 388326 -23056
rect 388382 -23112 388450 -23056
rect 388506 -23112 388640 -23056
rect 387840 -23180 388640 -23112
rect 387840 -23236 387954 -23180
rect 388010 -23236 388078 -23180
rect 388134 -23236 388202 -23180
rect 388258 -23236 388326 -23180
rect 388382 -23236 388450 -23180
rect 388506 -23236 388640 -23180
rect 387840 -23304 388640 -23236
rect 387840 -23360 387954 -23304
rect 388010 -23360 388078 -23304
rect 388134 -23360 388202 -23304
rect 388258 -23360 388326 -23304
rect 388382 -23360 388450 -23304
rect 388506 -23360 388640 -23304
rect 387840 -23428 388640 -23360
rect 387840 -23484 387954 -23428
rect 388010 -23484 388078 -23428
rect 388134 -23484 388202 -23428
rect 388258 -23484 388326 -23428
rect 388382 -23484 388450 -23428
rect 388506 -23484 388640 -23428
rect 387840 -23552 388640 -23484
rect 387840 -23608 387954 -23552
rect 388010 -23608 388078 -23552
rect 388134 -23608 388202 -23552
rect 388258 -23608 388326 -23552
rect 388382 -23608 388450 -23552
rect 388506 -23608 388640 -23552
rect 387840 -23676 388640 -23608
rect 387840 -23732 387954 -23676
rect 388010 -23732 388078 -23676
rect 388134 -23732 388202 -23676
rect 388258 -23732 388326 -23676
rect 388382 -23732 388450 -23676
rect 388506 -23732 388640 -23676
rect 387840 -23800 388640 -23732
rect 387840 -23856 387954 -23800
rect 388010 -23856 388078 -23800
rect 388134 -23856 388202 -23800
rect 388258 -23856 388326 -23800
rect 388382 -23856 388450 -23800
rect 388506 -23856 388640 -23800
rect 387840 -23924 388640 -23856
rect 387840 -23980 387954 -23924
rect 388010 -23980 388078 -23924
rect 388134 -23980 388202 -23924
rect 388258 -23980 388326 -23924
rect 388382 -23980 388450 -23924
rect 388506 -23980 388640 -23924
rect 387840 -24048 388640 -23980
rect 387840 -24104 387954 -24048
rect 388010 -24104 388078 -24048
rect 388134 -24104 388202 -24048
rect 388258 -24104 388326 -24048
rect 388382 -24104 388450 -24048
rect 388506 -24104 388640 -24048
rect 387840 -24172 388640 -24104
rect 387840 -24228 387954 -24172
rect 388010 -24228 388078 -24172
rect 388134 -24228 388202 -24172
rect 388258 -24228 388326 -24172
rect 388382 -24228 388450 -24172
rect 388506 -24228 388640 -24172
rect 387840 -24296 388640 -24228
rect 387840 -24352 387954 -24296
rect 388010 -24352 388078 -24296
rect 388134 -24352 388202 -24296
rect 388258 -24352 388326 -24296
rect 388382 -24352 388450 -24296
rect 388506 -24352 388640 -24296
rect 387840 -24420 388640 -24352
rect 387840 -24476 387954 -24420
rect 388010 -24476 388078 -24420
rect 388134 -24476 388202 -24420
rect 388258 -24476 388326 -24420
rect 388382 -24476 388450 -24420
rect 388506 -24476 388640 -24420
rect 387840 -24544 388640 -24476
rect 387840 -24600 387954 -24544
rect 388010 -24600 388078 -24544
rect 388134 -24600 388202 -24544
rect 388258 -24600 388326 -24544
rect 388382 -24600 388450 -24544
rect 388506 -24600 388640 -24544
rect 387840 -24668 388640 -24600
rect 387840 -24724 387954 -24668
rect 388010 -24724 388078 -24668
rect 388134 -24724 388202 -24668
rect 388258 -24724 388326 -24668
rect 388382 -24724 388450 -24668
rect 388506 -24724 388640 -24668
rect 387840 -24792 388640 -24724
rect 387840 -24848 387954 -24792
rect 388010 -24848 388078 -24792
rect 388134 -24848 388202 -24792
rect 388258 -24848 388326 -24792
rect 388382 -24848 388450 -24792
rect 388506 -24848 388640 -24792
rect 387840 -24916 388640 -24848
rect 387840 -24972 387954 -24916
rect 388010 -24972 388078 -24916
rect 388134 -24972 388202 -24916
rect 388258 -24972 388326 -24916
rect 388382 -24972 388450 -24916
rect 388506 -24972 388640 -24916
rect 387840 -25040 388640 -24972
rect 387840 -25096 387954 -25040
rect 388010 -25096 388078 -25040
rect 388134 -25096 388202 -25040
rect 388258 -25096 388326 -25040
rect 388382 -25096 388450 -25040
rect 388506 -25096 388640 -25040
rect 387840 -25164 388640 -25096
rect 387840 -25220 387954 -25164
rect 388010 -25220 388078 -25164
rect 388134 -25220 388202 -25164
rect 388258 -25220 388326 -25164
rect 388382 -25220 388450 -25164
rect 388506 -25220 388640 -25164
rect 387840 -25288 388640 -25220
rect 387840 -25344 387954 -25288
rect 388010 -25344 388078 -25288
rect 388134 -25344 388202 -25288
rect 388258 -25344 388326 -25288
rect 388382 -25344 388450 -25288
rect 388506 -25344 388640 -25288
rect 387840 -25412 388640 -25344
rect 387840 -25468 387954 -25412
rect 388010 -25468 388078 -25412
rect 388134 -25468 388202 -25412
rect 388258 -25468 388326 -25412
rect 388382 -25468 388450 -25412
rect 388506 -25468 388640 -25412
rect 387840 -25532 388640 -25468
rect 388908 -13680 389248 -13670
rect 388908 -13736 388981 -13680
rect 389037 -13736 389123 -13680
rect 389179 -13736 389248 -13680
rect 388908 -13822 389248 -13736
rect 388908 -13878 388981 -13822
rect 389037 -13878 389123 -13822
rect 389179 -13878 389248 -13822
rect 388908 -13964 389248 -13878
rect 388908 -14020 388981 -13964
rect 389037 -14020 389123 -13964
rect 389179 -14020 389248 -13964
rect 388908 -14106 389248 -14020
rect 388908 -14162 388981 -14106
rect 389037 -14162 389123 -14106
rect 389179 -14162 389248 -14106
rect 388908 -14248 389248 -14162
rect 388908 -14304 388981 -14248
rect 389037 -14304 389123 -14248
rect 389179 -14304 389248 -14248
rect 388908 -14390 389248 -14304
rect 388908 -14446 388981 -14390
rect 389037 -14446 389123 -14390
rect 389179 -14446 389248 -14390
rect 388908 -14532 389248 -14446
rect 388908 -14588 388981 -14532
rect 389037 -14588 389123 -14532
rect 389179 -14588 389248 -14532
rect 388908 -14674 389248 -14588
rect 388908 -14730 388981 -14674
rect 389037 -14730 389123 -14674
rect 389179 -14730 389248 -14674
rect 388908 -14816 389248 -14730
rect 388908 -14872 388981 -14816
rect 389037 -14872 389123 -14816
rect 389179 -14872 389248 -14816
rect 388908 -14958 389248 -14872
rect 388908 -15014 388981 -14958
rect 389037 -15014 389123 -14958
rect 389179 -15014 389248 -14958
rect 388908 -15100 389248 -15014
rect 388908 -15156 388981 -15100
rect 389037 -15156 389123 -15100
rect 389179 -15156 389248 -15100
rect 388908 -15242 389248 -15156
rect 388908 -15298 388981 -15242
rect 389037 -15298 389123 -15242
rect 389179 -15298 389248 -15242
rect 388908 -15384 389248 -15298
rect 388908 -15440 388981 -15384
rect 389037 -15440 389123 -15384
rect 389179 -15440 389248 -15384
rect 388908 -15526 389248 -15440
rect 388908 -15582 388981 -15526
rect 389037 -15582 389123 -15526
rect 389179 -15582 389248 -15526
rect 388908 -15668 389248 -15582
rect 388908 -15724 388981 -15668
rect 389037 -15724 389123 -15668
rect 389179 -15724 389248 -15668
rect 388908 -15810 389248 -15724
rect 388908 -15866 388981 -15810
rect 389037 -15866 389123 -15810
rect 389179 -15866 389248 -15810
rect 388908 -15952 389248 -15866
rect 388908 -16008 388981 -15952
rect 389037 -16008 389123 -15952
rect 389179 -16008 389248 -15952
rect 388908 -16094 389248 -16008
rect 388908 -16150 388981 -16094
rect 389037 -16150 389123 -16094
rect 389179 -16150 389248 -16094
rect 388908 -16236 389248 -16150
rect 388908 -16292 388981 -16236
rect 389037 -16292 389123 -16236
rect 389179 -16292 389248 -16236
rect 388908 -16378 389248 -16292
rect 388908 -16434 388981 -16378
rect 389037 -16434 389123 -16378
rect 389179 -16434 389248 -16378
rect 388908 -16520 389248 -16434
rect 388908 -16576 388981 -16520
rect 389037 -16576 389123 -16520
rect 389179 -16576 389248 -16520
rect 388908 -16662 389248 -16576
rect 388908 -16718 388981 -16662
rect 389037 -16718 389123 -16662
rect 389179 -16718 389248 -16662
rect 388908 -16804 389248 -16718
rect 388908 -16860 388981 -16804
rect 389037 -16860 389123 -16804
rect 389179 -16860 389248 -16804
rect 388908 -16946 389248 -16860
rect 388908 -17002 388981 -16946
rect 389037 -17002 389123 -16946
rect 389179 -17002 389248 -16946
rect 388908 -17088 389248 -17002
rect 388908 -17144 388981 -17088
rect 389037 -17144 389123 -17088
rect 389179 -17144 389248 -17088
rect 388908 -17230 389248 -17144
rect 388908 -17286 388981 -17230
rect 389037 -17286 389123 -17230
rect 389179 -17286 389248 -17230
rect 388908 -17372 389248 -17286
rect 388908 -17428 388981 -17372
rect 389037 -17428 389123 -17372
rect 389179 -17428 389248 -17372
rect 388908 -17514 389248 -17428
rect 388908 -17570 388981 -17514
rect 389037 -17570 389123 -17514
rect 389179 -17570 389248 -17514
rect 388908 -17656 389248 -17570
rect 388908 -17712 388981 -17656
rect 389037 -17712 389123 -17656
rect 389179 -17712 389248 -17656
rect 388908 -17798 389248 -17712
rect 388908 -17854 388981 -17798
rect 389037 -17854 389123 -17798
rect 389179 -17854 389248 -17798
rect 388908 -17940 389248 -17854
rect 388908 -17996 388981 -17940
rect 389037 -17996 389123 -17940
rect 389179 -17996 389248 -17940
rect 388908 -18082 389248 -17996
rect 388908 -18138 388981 -18082
rect 389037 -18138 389123 -18082
rect 389179 -18138 389248 -18082
rect 388908 -18224 389248 -18138
rect 388908 -18280 388981 -18224
rect 389037 -18280 389123 -18224
rect 389179 -18280 389248 -18224
rect 388908 -18366 389248 -18280
rect 388908 -18422 388981 -18366
rect 389037 -18422 389123 -18366
rect 389179 -18422 389248 -18366
rect 388908 -18508 389248 -18422
rect 388908 -18564 388981 -18508
rect 389037 -18564 389123 -18508
rect 389179 -18564 389248 -18508
rect 388908 -18650 389248 -18564
rect 388908 -18706 388981 -18650
rect 389037 -18706 389123 -18650
rect 389179 -18706 389248 -18650
rect 388908 -18792 389248 -18706
rect 388908 -18848 388981 -18792
rect 389037 -18848 389123 -18792
rect 389179 -18848 389248 -18792
rect 388908 -18934 389248 -18848
rect 388908 -18990 388981 -18934
rect 389037 -18990 389123 -18934
rect 389179 -18990 389248 -18934
rect 388908 -19076 389248 -18990
rect 388908 -19132 388981 -19076
rect 389037 -19132 389123 -19076
rect 389179 -19132 389248 -19076
rect 388908 -19218 389248 -19132
rect 388908 -19274 388981 -19218
rect 389037 -19274 389123 -19218
rect 389179 -19274 389248 -19218
rect 388908 -19360 389248 -19274
rect 388908 -19416 388981 -19360
rect 389037 -19416 389123 -19360
rect 389179 -19416 389248 -19360
rect 388908 -19502 389248 -19416
rect 388908 -19558 388981 -19502
rect 389037 -19558 389123 -19502
rect 389179 -19558 389248 -19502
rect 388908 -19644 389248 -19558
rect 388908 -19700 388981 -19644
rect 389037 -19700 389123 -19644
rect 389179 -19700 389248 -19644
rect 388908 -19786 389248 -19700
rect 388908 -19842 388981 -19786
rect 389037 -19842 389123 -19786
rect 389179 -19842 389248 -19786
rect 388908 -19928 389248 -19842
rect 388908 -19984 388981 -19928
rect 389037 -19984 389123 -19928
rect 389179 -19984 389248 -19928
rect 388908 -20070 389248 -19984
rect 388908 -20126 388981 -20070
rect 389037 -20126 389123 -20070
rect 389179 -20126 389248 -20070
rect 388908 -20212 389248 -20126
rect 388908 -20268 388981 -20212
rect 389037 -20268 389123 -20212
rect 389179 -20268 389248 -20212
rect 388908 -20354 389248 -20268
rect 388908 -20410 388981 -20354
rect 389037 -20410 389123 -20354
rect 389179 -20410 389248 -20354
rect 388908 -20496 389248 -20410
rect 388908 -20552 388981 -20496
rect 389037 -20552 389123 -20496
rect 389179 -20552 389248 -20496
rect 388908 -20638 389248 -20552
rect 388908 -20694 388981 -20638
rect 389037 -20694 389123 -20638
rect 389179 -20694 389248 -20638
rect 388908 -20780 389248 -20694
rect 388908 -20836 388981 -20780
rect 389037 -20836 389123 -20780
rect 389179 -20836 389248 -20780
rect 388908 -20922 389248 -20836
rect 388908 -20978 388981 -20922
rect 389037 -20978 389123 -20922
rect 389179 -20978 389248 -20922
rect 388908 -21064 389248 -20978
rect 388908 -21120 388981 -21064
rect 389037 -21120 389123 -21064
rect 389179 -21120 389248 -21064
rect 388908 -21206 389248 -21120
rect 388908 -21262 388981 -21206
rect 389037 -21262 389123 -21206
rect 389179 -21262 389248 -21206
rect 388908 -21348 389248 -21262
rect 388908 -21404 388981 -21348
rect 389037 -21404 389123 -21348
rect 389179 -21404 389248 -21348
rect 388908 -21490 389248 -21404
rect 388908 -21546 388981 -21490
rect 389037 -21546 389123 -21490
rect 389179 -21546 389248 -21490
rect 388908 -21632 389248 -21546
rect 388908 -21688 388981 -21632
rect 389037 -21688 389123 -21632
rect 389179 -21688 389248 -21632
rect 388908 -21774 389248 -21688
rect 388908 -21830 388981 -21774
rect 389037 -21830 389123 -21774
rect 389179 -21830 389248 -21774
rect 388908 -21916 389248 -21830
rect 388908 -21972 388981 -21916
rect 389037 -21972 389123 -21916
rect 389179 -21972 389248 -21916
rect 388908 -22058 389248 -21972
rect 388908 -22114 388981 -22058
rect 389037 -22114 389123 -22058
rect 389179 -22114 389248 -22058
rect 388908 -22200 389248 -22114
rect 388908 -22256 388981 -22200
rect 389037 -22256 389123 -22200
rect 389179 -22256 389248 -22200
rect 388908 -22342 389248 -22256
rect 388908 -22398 388981 -22342
rect 389037 -22398 389123 -22342
rect 389179 -22398 389248 -22342
rect 388908 -22484 389248 -22398
rect 388908 -22540 388981 -22484
rect 389037 -22540 389123 -22484
rect 389179 -22540 389248 -22484
rect 388908 -22626 389248 -22540
rect 388908 -22682 388981 -22626
rect 389037 -22682 389123 -22626
rect 389179 -22682 389248 -22626
rect 388908 -22768 389248 -22682
rect 388908 -22824 388981 -22768
rect 389037 -22824 389123 -22768
rect 389179 -22824 389248 -22768
rect 388908 -22910 389248 -22824
rect 388908 -22966 388981 -22910
rect 389037 -22966 389123 -22910
rect 389179 -22966 389248 -22910
rect 388908 -23052 389248 -22966
rect 388908 -23108 388981 -23052
rect 389037 -23108 389123 -23052
rect 389179 -23108 389248 -23052
rect 388908 -23194 389248 -23108
rect 388908 -23250 388981 -23194
rect 389037 -23250 389123 -23194
rect 389179 -23250 389248 -23194
rect 388908 -23336 389248 -23250
rect 388908 -23392 388981 -23336
rect 389037 -23392 389123 -23336
rect 389179 -23392 389248 -23336
rect 388908 -23478 389248 -23392
rect 388908 -23534 388981 -23478
rect 389037 -23534 389123 -23478
rect 389179 -23534 389248 -23478
rect 388908 -23620 389248 -23534
rect 388908 -23676 388981 -23620
rect 389037 -23676 389123 -23620
rect 389179 -23676 389248 -23620
rect 388908 -23762 389248 -23676
rect 388908 -23818 388981 -23762
rect 389037 -23818 389123 -23762
rect 389179 -23818 389248 -23762
rect 388908 -23904 389248 -23818
rect 388908 -23960 388981 -23904
rect 389037 -23960 389123 -23904
rect 389179 -23960 389248 -23904
rect 388908 -24046 389248 -23960
rect 388908 -24102 388981 -24046
rect 389037 -24102 389123 -24046
rect 389179 -24102 389248 -24046
rect 388908 -24188 389248 -24102
rect 388908 -24244 388981 -24188
rect 389037 -24244 389123 -24188
rect 389179 -24244 389248 -24188
rect 388908 -24330 389248 -24244
rect 388908 -24386 388981 -24330
rect 389037 -24386 389123 -24330
rect 389179 -24386 389248 -24330
rect 388908 -24472 389248 -24386
rect 388908 -24528 388981 -24472
rect 389037 -24528 389123 -24472
rect 389179 -24528 389248 -24472
rect 388908 -24614 389248 -24528
rect 388908 -24670 388981 -24614
rect 389037 -24670 389123 -24614
rect 389179 -24670 389248 -24614
rect 388908 -24756 389248 -24670
rect 388908 -24812 388981 -24756
rect 389037 -24812 389123 -24756
rect 389179 -24812 389248 -24756
rect 388908 -24898 389248 -24812
rect 388908 -24954 388981 -24898
rect 389037 -24954 389123 -24898
rect 389179 -24954 389248 -24898
rect 388908 -25040 389248 -24954
rect 388908 -25096 388981 -25040
rect 389037 -25096 389123 -25040
rect 389179 -25096 389248 -25040
rect 388908 -25182 389248 -25096
rect 388908 -25238 388981 -25182
rect 389037 -25238 389123 -25182
rect 389179 -25238 389248 -25182
rect 388908 -25324 389248 -25238
rect 388908 -25380 388981 -25324
rect 389037 -25380 389123 -25324
rect 389179 -25380 389248 -25324
rect 388908 -25466 389248 -25380
rect 388908 -25522 388981 -25466
rect 389037 -25522 389123 -25466
rect 389179 -25522 389248 -25466
rect 388908 -25532 389248 -25522
rect 389308 -13680 389648 -13670
rect 389308 -13736 389382 -13680
rect 389438 -13736 389524 -13680
rect 389580 -13736 389648 -13680
rect 389308 -13822 389648 -13736
rect 389308 -13878 389382 -13822
rect 389438 -13878 389524 -13822
rect 389580 -13878 389648 -13822
rect 389308 -13964 389648 -13878
rect 389308 -14020 389382 -13964
rect 389438 -14020 389524 -13964
rect 389580 -14020 389648 -13964
rect 389308 -14106 389648 -14020
rect 389308 -14162 389382 -14106
rect 389438 -14162 389524 -14106
rect 389580 -14162 389648 -14106
rect 389308 -14248 389648 -14162
rect 389308 -14304 389382 -14248
rect 389438 -14304 389524 -14248
rect 389580 -14304 389648 -14248
rect 389308 -14390 389648 -14304
rect 389308 -14446 389382 -14390
rect 389438 -14446 389524 -14390
rect 389580 -14446 389648 -14390
rect 389308 -14532 389648 -14446
rect 389308 -14588 389382 -14532
rect 389438 -14588 389524 -14532
rect 389580 -14588 389648 -14532
rect 389308 -14674 389648 -14588
rect 389308 -14730 389382 -14674
rect 389438 -14730 389524 -14674
rect 389580 -14730 389648 -14674
rect 389308 -14816 389648 -14730
rect 389308 -14872 389382 -14816
rect 389438 -14872 389524 -14816
rect 389580 -14872 389648 -14816
rect 389308 -14958 389648 -14872
rect 389308 -15014 389382 -14958
rect 389438 -15014 389524 -14958
rect 389580 -15014 389648 -14958
rect 389308 -15100 389648 -15014
rect 389308 -15156 389382 -15100
rect 389438 -15156 389524 -15100
rect 389580 -15156 389648 -15100
rect 389308 -15242 389648 -15156
rect 389308 -15298 389382 -15242
rect 389438 -15298 389524 -15242
rect 389580 -15298 389648 -15242
rect 389308 -15384 389648 -15298
rect 389308 -15440 389382 -15384
rect 389438 -15440 389524 -15384
rect 389580 -15440 389648 -15384
rect 389308 -15526 389648 -15440
rect 389308 -15582 389382 -15526
rect 389438 -15582 389524 -15526
rect 389580 -15582 389648 -15526
rect 389308 -15668 389648 -15582
rect 389308 -15724 389382 -15668
rect 389438 -15724 389524 -15668
rect 389580 -15724 389648 -15668
rect 389308 -15810 389648 -15724
rect 389308 -15866 389382 -15810
rect 389438 -15866 389524 -15810
rect 389580 -15866 389648 -15810
rect 389308 -15952 389648 -15866
rect 389308 -16008 389382 -15952
rect 389438 -16008 389524 -15952
rect 389580 -16008 389648 -15952
rect 389308 -16094 389648 -16008
rect 389308 -16150 389382 -16094
rect 389438 -16150 389524 -16094
rect 389580 -16150 389648 -16094
rect 389308 -16236 389648 -16150
rect 389308 -16292 389382 -16236
rect 389438 -16292 389524 -16236
rect 389580 -16292 389648 -16236
rect 389308 -16378 389648 -16292
rect 389308 -16434 389382 -16378
rect 389438 -16434 389524 -16378
rect 389580 -16434 389648 -16378
rect 389308 -16520 389648 -16434
rect 389308 -16576 389382 -16520
rect 389438 -16576 389524 -16520
rect 389580 -16576 389648 -16520
rect 389308 -16662 389648 -16576
rect 389308 -16718 389382 -16662
rect 389438 -16718 389524 -16662
rect 389580 -16718 389648 -16662
rect 389308 -16804 389648 -16718
rect 389308 -16860 389382 -16804
rect 389438 -16860 389524 -16804
rect 389580 -16860 389648 -16804
rect 389308 -16946 389648 -16860
rect 389308 -17002 389382 -16946
rect 389438 -17002 389524 -16946
rect 389580 -17002 389648 -16946
rect 389308 -17088 389648 -17002
rect 389308 -17144 389382 -17088
rect 389438 -17144 389524 -17088
rect 389580 -17144 389648 -17088
rect 389308 -17230 389648 -17144
rect 389308 -17286 389382 -17230
rect 389438 -17286 389524 -17230
rect 389580 -17286 389648 -17230
rect 389308 -17372 389648 -17286
rect 389308 -17428 389382 -17372
rect 389438 -17428 389524 -17372
rect 389580 -17428 389648 -17372
rect 389308 -17514 389648 -17428
rect 389308 -17570 389382 -17514
rect 389438 -17570 389524 -17514
rect 389580 -17570 389648 -17514
rect 389308 -17656 389648 -17570
rect 389308 -17712 389382 -17656
rect 389438 -17712 389524 -17656
rect 389580 -17712 389648 -17656
rect 389308 -17798 389648 -17712
rect 389308 -17854 389382 -17798
rect 389438 -17854 389524 -17798
rect 389580 -17854 389648 -17798
rect 389308 -17940 389648 -17854
rect 389308 -17996 389382 -17940
rect 389438 -17996 389524 -17940
rect 389580 -17996 389648 -17940
rect 389308 -18082 389648 -17996
rect 389308 -18138 389382 -18082
rect 389438 -18138 389524 -18082
rect 389580 -18138 389648 -18082
rect 389308 -18224 389648 -18138
rect 389308 -18280 389382 -18224
rect 389438 -18280 389524 -18224
rect 389580 -18280 389648 -18224
rect 389308 -18366 389648 -18280
rect 389308 -18422 389382 -18366
rect 389438 -18422 389524 -18366
rect 389580 -18422 389648 -18366
rect 389308 -18508 389648 -18422
rect 389308 -18564 389382 -18508
rect 389438 -18564 389524 -18508
rect 389580 -18564 389648 -18508
rect 389308 -18650 389648 -18564
rect 389308 -18706 389382 -18650
rect 389438 -18706 389524 -18650
rect 389580 -18706 389648 -18650
rect 389308 -18792 389648 -18706
rect 389308 -18848 389382 -18792
rect 389438 -18848 389524 -18792
rect 389580 -18848 389648 -18792
rect 389308 -18934 389648 -18848
rect 389308 -18990 389382 -18934
rect 389438 -18990 389524 -18934
rect 389580 -18990 389648 -18934
rect 389308 -19076 389648 -18990
rect 389308 -19132 389382 -19076
rect 389438 -19132 389524 -19076
rect 389580 -19132 389648 -19076
rect 389308 -19218 389648 -19132
rect 389308 -19274 389382 -19218
rect 389438 -19274 389524 -19218
rect 389580 -19274 389648 -19218
rect 389308 -19360 389648 -19274
rect 389308 -19416 389382 -19360
rect 389438 -19416 389524 -19360
rect 389580 -19416 389648 -19360
rect 389308 -19502 389648 -19416
rect 389308 -19558 389382 -19502
rect 389438 -19558 389524 -19502
rect 389580 -19558 389648 -19502
rect 389308 -19644 389648 -19558
rect 389308 -19700 389382 -19644
rect 389438 -19700 389524 -19644
rect 389580 -19700 389648 -19644
rect 389308 -19786 389648 -19700
rect 389308 -19842 389382 -19786
rect 389438 -19842 389524 -19786
rect 389580 -19842 389648 -19786
rect 389308 -19928 389648 -19842
rect 389308 -19984 389382 -19928
rect 389438 -19984 389524 -19928
rect 389580 -19984 389648 -19928
rect 389308 -20070 389648 -19984
rect 389308 -20126 389382 -20070
rect 389438 -20126 389524 -20070
rect 389580 -20126 389648 -20070
rect 389308 -20212 389648 -20126
rect 389308 -20268 389382 -20212
rect 389438 -20268 389524 -20212
rect 389580 -20268 389648 -20212
rect 389308 -20354 389648 -20268
rect 389308 -20410 389382 -20354
rect 389438 -20410 389524 -20354
rect 389580 -20410 389648 -20354
rect 389308 -20496 389648 -20410
rect 389308 -20552 389382 -20496
rect 389438 -20552 389524 -20496
rect 389580 -20552 389648 -20496
rect 389308 -20638 389648 -20552
rect 389308 -20694 389382 -20638
rect 389438 -20694 389524 -20638
rect 389580 -20694 389648 -20638
rect 389308 -20780 389648 -20694
rect 389308 -20836 389382 -20780
rect 389438 -20836 389524 -20780
rect 389580 -20836 389648 -20780
rect 389308 -20922 389648 -20836
rect 389308 -20978 389382 -20922
rect 389438 -20978 389524 -20922
rect 389580 -20978 389648 -20922
rect 389308 -21064 389648 -20978
rect 389308 -21120 389382 -21064
rect 389438 -21120 389524 -21064
rect 389580 -21120 389648 -21064
rect 389308 -21206 389648 -21120
rect 389308 -21262 389382 -21206
rect 389438 -21262 389524 -21206
rect 389580 -21262 389648 -21206
rect 389308 -21348 389648 -21262
rect 389308 -21404 389382 -21348
rect 389438 -21404 389524 -21348
rect 389580 -21404 389648 -21348
rect 389308 -21490 389648 -21404
rect 389308 -21546 389382 -21490
rect 389438 -21546 389524 -21490
rect 389580 -21546 389648 -21490
rect 389308 -21632 389648 -21546
rect 389308 -21688 389382 -21632
rect 389438 -21688 389524 -21632
rect 389580 -21688 389648 -21632
rect 389308 -21774 389648 -21688
rect 389308 -21830 389382 -21774
rect 389438 -21830 389524 -21774
rect 389580 -21830 389648 -21774
rect 389308 -21916 389648 -21830
rect 389308 -21972 389382 -21916
rect 389438 -21972 389524 -21916
rect 389580 -21972 389648 -21916
rect 389308 -22058 389648 -21972
rect 389308 -22114 389382 -22058
rect 389438 -22114 389524 -22058
rect 389580 -22114 389648 -22058
rect 389308 -22200 389648 -22114
rect 389308 -22256 389382 -22200
rect 389438 -22256 389524 -22200
rect 389580 -22256 389648 -22200
rect 389308 -22342 389648 -22256
rect 389308 -22398 389382 -22342
rect 389438 -22398 389524 -22342
rect 389580 -22398 389648 -22342
rect 389308 -22484 389648 -22398
rect 389308 -22540 389382 -22484
rect 389438 -22540 389524 -22484
rect 389580 -22540 389648 -22484
rect 389308 -22626 389648 -22540
rect 389308 -22682 389382 -22626
rect 389438 -22682 389524 -22626
rect 389580 -22682 389648 -22626
rect 389308 -22768 389648 -22682
rect 389308 -22824 389382 -22768
rect 389438 -22824 389524 -22768
rect 389580 -22824 389648 -22768
rect 389308 -22910 389648 -22824
rect 389308 -22966 389382 -22910
rect 389438 -22966 389524 -22910
rect 389580 -22966 389648 -22910
rect 389308 -23052 389648 -22966
rect 389308 -23108 389382 -23052
rect 389438 -23108 389524 -23052
rect 389580 -23108 389648 -23052
rect 389308 -23194 389648 -23108
rect 389308 -23250 389382 -23194
rect 389438 -23250 389524 -23194
rect 389580 -23250 389648 -23194
rect 389308 -23336 389648 -23250
rect 389308 -23392 389382 -23336
rect 389438 -23392 389524 -23336
rect 389580 -23392 389648 -23336
rect 389308 -23478 389648 -23392
rect 389308 -23534 389382 -23478
rect 389438 -23534 389524 -23478
rect 389580 -23534 389648 -23478
rect 389308 -23620 389648 -23534
rect 389308 -23676 389382 -23620
rect 389438 -23676 389524 -23620
rect 389580 -23676 389648 -23620
rect 389308 -23762 389648 -23676
rect 389308 -23818 389382 -23762
rect 389438 -23818 389524 -23762
rect 389580 -23818 389648 -23762
rect 389308 -23904 389648 -23818
rect 389308 -23960 389382 -23904
rect 389438 -23960 389524 -23904
rect 389580 -23960 389648 -23904
rect 389308 -24046 389648 -23960
rect 389308 -24102 389382 -24046
rect 389438 -24102 389524 -24046
rect 389580 -24102 389648 -24046
rect 389308 -24188 389648 -24102
rect 389308 -24244 389382 -24188
rect 389438 -24244 389524 -24188
rect 389580 -24244 389648 -24188
rect 389308 -24330 389648 -24244
rect 389308 -24386 389382 -24330
rect 389438 -24386 389524 -24330
rect 389580 -24386 389648 -24330
rect 389308 -24472 389648 -24386
rect 389308 -24528 389382 -24472
rect 389438 -24528 389524 -24472
rect 389580 -24528 389648 -24472
rect 389308 -24614 389648 -24528
rect 389308 -24670 389382 -24614
rect 389438 -24670 389524 -24614
rect 389580 -24670 389648 -24614
rect 389308 -24756 389648 -24670
rect 389308 -24812 389382 -24756
rect 389438 -24812 389524 -24756
rect 389580 -24812 389648 -24756
rect 389308 -24898 389648 -24812
rect 389308 -24954 389382 -24898
rect 389438 -24954 389524 -24898
rect 389580 -24954 389648 -24898
rect 389308 -25040 389648 -24954
rect 389308 -25096 389382 -25040
rect 389438 -25096 389524 -25040
rect 389580 -25096 389648 -25040
rect 389308 -25182 389648 -25096
rect 389308 -25238 389382 -25182
rect 389438 -25238 389524 -25182
rect 389580 -25238 389648 -25182
rect 389308 -25324 389648 -25238
rect 389308 -25380 389382 -25324
rect 389438 -25380 389524 -25324
rect 389580 -25380 389648 -25324
rect 389308 -25466 389648 -25380
rect 389308 -25522 389382 -25466
rect 389438 -25522 389524 -25466
rect 389580 -25522 389648 -25466
rect 389308 -25532 389648 -25522
rect 389708 -13680 390048 -13670
rect 389708 -13736 389782 -13680
rect 389838 -13736 389924 -13680
rect 389980 -13736 390048 -13680
rect 389708 -13822 390048 -13736
rect 389708 -13878 389782 -13822
rect 389838 -13878 389924 -13822
rect 389980 -13878 390048 -13822
rect 389708 -13964 390048 -13878
rect 389708 -14020 389782 -13964
rect 389838 -14020 389924 -13964
rect 389980 -14020 390048 -13964
rect 389708 -14106 390048 -14020
rect 389708 -14162 389782 -14106
rect 389838 -14162 389924 -14106
rect 389980 -14162 390048 -14106
rect 389708 -14248 390048 -14162
rect 389708 -14304 389782 -14248
rect 389838 -14304 389924 -14248
rect 389980 -14304 390048 -14248
rect 389708 -14390 390048 -14304
rect 389708 -14446 389782 -14390
rect 389838 -14446 389924 -14390
rect 389980 -14446 390048 -14390
rect 389708 -14532 390048 -14446
rect 389708 -14588 389782 -14532
rect 389838 -14588 389924 -14532
rect 389980 -14588 390048 -14532
rect 389708 -14674 390048 -14588
rect 389708 -14730 389782 -14674
rect 389838 -14730 389924 -14674
rect 389980 -14730 390048 -14674
rect 389708 -14816 390048 -14730
rect 389708 -14872 389782 -14816
rect 389838 -14872 389924 -14816
rect 389980 -14872 390048 -14816
rect 389708 -14958 390048 -14872
rect 389708 -15014 389782 -14958
rect 389838 -15014 389924 -14958
rect 389980 -15014 390048 -14958
rect 389708 -15100 390048 -15014
rect 389708 -15156 389782 -15100
rect 389838 -15156 389924 -15100
rect 389980 -15156 390048 -15100
rect 389708 -15242 390048 -15156
rect 389708 -15298 389782 -15242
rect 389838 -15298 389924 -15242
rect 389980 -15298 390048 -15242
rect 389708 -15384 390048 -15298
rect 389708 -15440 389782 -15384
rect 389838 -15440 389924 -15384
rect 389980 -15440 390048 -15384
rect 389708 -15526 390048 -15440
rect 389708 -15582 389782 -15526
rect 389838 -15582 389924 -15526
rect 389980 -15582 390048 -15526
rect 389708 -15668 390048 -15582
rect 389708 -15724 389782 -15668
rect 389838 -15724 389924 -15668
rect 389980 -15724 390048 -15668
rect 389708 -15810 390048 -15724
rect 389708 -15866 389782 -15810
rect 389838 -15866 389924 -15810
rect 389980 -15866 390048 -15810
rect 389708 -15952 390048 -15866
rect 389708 -16008 389782 -15952
rect 389838 -16008 389924 -15952
rect 389980 -16008 390048 -15952
rect 389708 -16094 390048 -16008
rect 389708 -16150 389782 -16094
rect 389838 -16150 389924 -16094
rect 389980 -16150 390048 -16094
rect 389708 -16236 390048 -16150
rect 389708 -16292 389782 -16236
rect 389838 -16292 389924 -16236
rect 389980 -16292 390048 -16236
rect 389708 -16378 390048 -16292
rect 389708 -16434 389782 -16378
rect 389838 -16434 389924 -16378
rect 389980 -16434 390048 -16378
rect 389708 -16520 390048 -16434
rect 389708 -16576 389782 -16520
rect 389838 -16576 389924 -16520
rect 389980 -16576 390048 -16520
rect 389708 -16662 390048 -16576
rect 389708 -16718 389782 -16662
rect 389838 -16718 389924 -16662
rect 389980 -16718 390048 -16662
rect 389708 -16804 390048 -16718
rect 389708 -16860 389782 -16804
rect 389838 -16860 389924 -16804
rect 389980 -16860 390048 -16804
rect 389708 -16946 390048 -16860
rect 389708 -17002 389782 -16946
rect 389838 -17002 389924 -16946
rect 389980 -17002 390048 -16946
rect 389708 -17088 390048 -17002
rect 389708 -17144 389782 -17088
rect 389838 -17144 389924 -17088
rect 389980 -17144 390048 -17088
rect 389708 -17230 390048 -17144
rect 389708 -17286 389782 -17230
rect 389838 -17286 389924 -17230
rect 389980 -17286 390048 -17230
rect 389708 -17372 390048 -17286
rect 389708 -17428 389782 -17372
rect 389838 -17428 389924 -17372
rect 389980 -17428 390048 -17372
rect 389708 -17514 390048 -17428
rect 389708 -17570 389782 -17514
rect 389838 -17570 389924 -17514
rect 389980 -17570 390048 -17514
rect 389708 -17656 390048 -17570
rect 389708 -17712 389782 -17656
rect 389838 -17712 389924 -17656
rect 389980 -17712 390048 -17656
rect 389708 -17798 390048 -17712
rect 389708 -17854 389782 -17798
rect 389838 -17854 389924 -17798
rect 389980 -17854 390048 -17798
rect 389708 -17940 390048 -17854
rect 389708 -17996 389782 -17940
rect 389838 -17996 389924 -17940
rect 389980 -17996 390048 -17940
rect 389708 -18082 390048 -17996
rect 389708 -18138 389782 -18082
rect 389838 -18138 389924 -18082
rect 389980 -18138 390048 -18082
rect 389708 -18224 390048 -18138
rect 389708 -18280 389782 -18224
rect 389838 -18280 389924 -18224
rect 389980 -18280 390048 -18224
rect 389708 -18366 390048 -18280
rect 389708 -18422 389782 -18366
rect 389838 -18422 389924 -18366
rect 389980 -18422 390048 -18366
rect 389708 -18508 390048 -18422
rect 389708 -18564 389782 -18508
rect 389838 -18564 389924 -18508
rect 389980 -18564 390048 -18508
rect 389708 -18650 390048 -18564
rect 389708 -18706 389782 -18650
rect 389838 -18706 389924 -18650
rect 389980 -18706 390048 -18650
rect 389708 -18792 390048 -18706
rect 389708 -18848 389782 -18792
rect 389838 -18848 389924 -18792
rect 389980 -18848 390048 -18792
rect 389708 -18934 390048 -18848
rect 389708 -18990 389782 -18934
rect 389838 -18990 389924 -18934
rect 389980 -18990 390048 -18934
rect 389708 -19076 390048 -18990
rect 389708 -19132 389782 -19076
rect 389838 -19132 389924 -19076
rect 389980 -19132 390048 -19076
rect 389708 -19218 390048 -19132
rect 389708 -19274 389782 -19218
rect 389838 -19274 389924 -19218
rect 389980 -19274 390048 -19218
rect 389708 -19360 390048 -19274
rect 389708 -19416 389782 -19360
rect 389838 -19416 389924 -19360
rect 389980 -19416 390048 -19360
rect 389708 -19502 390048 -19416
rect 389708 -19558 389782 -19502
rect 389838 -19558 389924 -19502
rect 389980 -19558 390048 -19502
rect 389708 -19644 390048 -19558
rect 389708 -19700 389782 -19644
rect 389838 -19700 389924 -19644
rect 389980 -19700 390048 -19644
rect 389708 -19786 390048 -19700
rect 389708 -19842 389782 -19786
rect 389838 -19842 389924 -19786
rect 389980 -19842 390048 -19786
rect 389708 -19928 390048 -19842
rect 389708 -19984 389782 -19928
rect 389838 -19984 389924 -19928
rect 389980 -19984 390048 -19928
rect 389708 -20070 390048 -19984
rect 389708 -20126 389782 -20070
rect 389838 -20126 389924 -20070
rect 389980 -20126 390048 -20070
rect 389708 -20212 390048 -20126
rect 389708 -20268 389782 -20212
rect 389838 -20268 389924 -20212
rect 389980 -20268 390048 -20212
rect 389708 -20354 390048 -20268
rect 389708 -20410 389782 -20354
rect 389838 -20410 389924 -20354
rect 389980 -20410 390048 -20354
rect 389708 -20496 390048 -20410
rect 389708 -20552 389782 -20496
rect 389838 -20552 389924 -20496
rect 389980 -20552 390048 -20496
rect 389708 -20638 390048 -20552
rect 389708 -20694 389782 -20638
rect 389838 -20694 389924 -20638
rect 389980 -20694 390048 -20638
rect 389708 -20780 390048 -20694
rect 389708 -20836 389782 -20780
rect 389838 -20836 389924 -20780
rect 389980 -20836 390048 -20780
rect 389708 -20922 390048 -20836
rect 389708 -20978 389782 -20922
rect 389838 -20978 389924 -20922
rect 389980 -20978 390048 -20922
rect 389708 -21064 390048 -20978
rect 389708 -21120 389782 -21064
rect 389838 -21120 389924 -21064
rect 389980 -21120 390048 -21064
rect 389708 -21206 390048 -21120
rect 389708 -21262 389782 -21206
rect 389838 -21262 389924 -21206
rect 389980 -21262 390048 -21206
rect 389708 -21348 390048 -21262
rect 389708 -21404 389782 -21348
rect 389838 -21404 389924 -21348
rect 389980 -21404 390048 -21348
rect 389708 -21490 390048 -21404
rect 389708 -21546 389782 -21490
rect 389838 -21546 389924 -21490
rect 389980 -21546 390048 -21490
rect 389708 -21632 390048 -21546
rect 389708 -21688 389782 -21632
rect 389838 -21688 389924 -21632
rect 389980 -21688 390048 -21632
rect 389708 -21774 390048 -21688
rect 389708 -21830 389782 -21774
rect 389838 -21830 389924 -21774
rect 389980 -21830 390048 -21774
rect 389708 -21916 390048 -21830
rect 389708 -21972 389782 -21916
rect 389838 -21972 389924 -21916
rect 389980 -21972 390048 -21916
rect 389708 -22058 390048 -21972
rect 389708 -22114 389782 -22058
rect 389838 -22114 389924 -22058
rect 389980 -22114 390048 -22058
rect 389708 -22200 390048 -22114
rect 389708 -22256 389782 -22200
rect 389838 -22256 389924 -22200
rect 389980 -22256 390048 -22200
rect 389708 -22342 390048 -22256
rect 389708 -22398 389782 -22342
rect 389838 -22398 389924 -22342
rect 389980 -22398 390048 -22342
rect 389708 -22484 390048 -22398
rect 389708 -22540 389782 -22484
rect 389838 -22540 389924 -22484
rect 389980 -22540 390048 -22484
rect 389708 -22626 390048 -22540
rect 389708 -22682 389782 -22626
rect 389838 -22682 389924 -22626
rect 389980 -22682 390048 -22626
rect 389708 -22768 390048 -22682
rect 389708 -22824 389782 -22768
rect 389838 -22824 389924 -22768
rect 389980 -22824 390048 -22768
rect 389708 -22910 390048 -22824
rect 389708 -22966 389782 -22910
rect 389838 -22966 389924 -22910
rect 389980 -22966 390048 -22910
rect 389708 -23052 390048 -22966
rect 389708 -23108 389782 -23052
rect 389838 -23108 389924 -23052
rect 389980 -23108 390048 -23052
rect 389708 -23194 390048 -23108
rect 389708 -23250 389782 -23194
rect 389838 -23250 389924 -23194
rect 389980 -23250 390048 -23194
rect 389708 -23336 390048 -23250
rect 389708 -23392 389782 -23336
rect 389838 -23392 389924 -23336
rect 389980 -23392 390048 -23336
rect 389708 -23478 390048 -23392
rect 389708 -23534 389782 -23478
rect 389838 -23534 389924 -23478
rect 389980 -23534 390048 -23478
rect 389708 -23620 390048 -23534
rect 389708 -23676 389782 -23620
rect 389838 -23676 389924 -23620
rect 389980 -23676 390048 -23620
rect 389708 -23762 390048 -23676
rect 389708 -23818 389782 -23762
rect 389838 -23818 389924 -23762
rect 389980 -23818 390048 -23762
rect 389708 -23904 390048 -23818
rect 389708 -23960 389782 -23904
rect 389838 -23960 389924 -23904
rect 389980 -23960 390048 -23904
rect 389708 -24046 390048 -23960
rect 389708 -24102 389782 -24046
rect 389838 -24102 389924 -24046
rect 389980 -24102 390048 -24046
rect 389708 -24188 390048 -24102
rect 389708 -24244 389782 -24188
rect 389838 -24244 389924 -24188
rect 389980 -24244 390048 -24188
rect 389708 -24330 390048 -24244
rect 389708 -24386 389782 -24330
rect 389838 -24386 389924 -24330
rect 389980 -24386 390048 -24330
rect 389708 -24472 390048 -24386
rect 389708 -24528 389782 -24472
rect 389838 -24528 389924 -24472
rect 389980 -24528 390048 -24472
rect 389708 -24614 390048 -24528
rect 389708 -24670 389782 -24614
rect 389838 -24670 389924 -24614
rect 389980 -24670 390048 -24614
rect 389708 -24756 390048 -24670
rect 389708 -24812 389782 -24756
rect 389838 -24812 389924 -24756
rect 389980 -24812 390048 -24756
rect 389708 -24898 390048 -24812
rect 389708 -24954 389782 -24898
rect 389838 -24954 389924 -24898
rect 389980 -24954 390048 -24898
rect 389708 -25040 390048 -24954
rect 389708 -25096 389782 -25040
rect 389838 -25096 389924 -25040
rect 389980 -25096 390048 -25040
rect 389708 -25182 390048 -25096
rect 389708 -25238 389782 -25182
rect 389838 -25238 389924 -25182
rect 389980 -25238 390048 -25182
rect 389708 -25324 390048 -25238
rect 389708 -25380 389782 -25324
rect 389838 -25380 389924 -25324
rect 389980 -25380 390048 -25324
rect 389708 -25466 390048 -25380
rect 389708 -25522 389782 -25466
rect 389838 -25522 389924 -25466
rect 389980 -25522 390048 -25466
rect 389708 -25532 390048 -25522
rect 390108 -13680 390448 -13670
rect 390108 -13736 390179 -13680
rect 390235 -13736 390321 -13680
rect 390377 -13736 390448 -13680
rect 390108 -13822 390448 -13736
rect 390108 -13878 390179 -13822
rect 390235 -13878 390321 -13822
rect 390377 -13878 390448 -13822
rect 390108 -13964 390448 -13878
rect 390108 -14020 390179 -13964
rect 390235 -14020 390321 -13964
rect 390377 -14020 390448 -13964
rect 390108 -14106 390448 -14020
rect 390108 -14162 390179 -14106
rect 390235 -14162 390321 -14106
rect 390377 -14162 390448 -14106
rect 390108 -14248 390448 -14162
rect 390108 -14304 390179 -14248
rect 390235 -14304 390321 -14248
rect 390377 -14304 390448 -14248
rect 390108 -14390 390448 -14304
rect 390108 -14446 390179 -14390
rect 390235 -14446 390321 -14390
rect 390377 -14446 390448 -14390
rect 390108 -14532 390448 -14446
rect 390108 -14588 390179 -14532
rect 390235 -14588 390321 -14532
rect 390377 -14588 390448 -14532
rect 390108 -14674 390448 -14588
rect 390108 -14730 390179 -14674
rect 390235 -14730 390321 -14674
rect 390377 -14730 390448 -14674
rect 390108 -14816 390448 -14730
rect 390108 -14872 390179 -14816
rect 390235 -14872 390321 -14816
rect 390377 -14872 390448 -14816
rect 390108 -14958 390448 -14872
rect 390108 -15014 390179 -14958
rect 390235 -15014 390321 -14958
rect 390377 -15014 390448 -14958
rect 390108 -15100 390448 -15014
rect 390108 -15156 390179 -15100
rect 390235 -15156 390321 -15100
rect 390377 -15156 390448 -15100
rect 390108 -15242 390448 -15156
rect 390108 -15298 390179 -15242
rect 390235 -15298 390321 -15242
rect 390377 -15298 390448 -15242
rect 390108 -15384 390448 -15298
rect 390108 -15440 390179 -15384
rect 390235 -15440 390321 -15384
rect 390377 -15440 390448 -15384
rect 390108 -15526 390448 -15440
rect 390108 -15582 390179 -15526
rect 390235 -15582 390321 -15526
rect 390377 -15582 390448 -15526
rect 390108 -15668 390448 -15582
rect 390108 -15724 390179 -15668
rect 390235 -15724 390321 -15668
rect 390377 -15724 390448 -15668
rect 390108 -15810 390448 -15724
rect 390108 -15866 390179 -15810
rect 390235 -15866 390321 -15810
rect 390377 -15866 390448 -15810
rect 390108 -15952 390448 -15866
rect 390108 -16008 390179 -15952
rect 390235 -16008 390321 -15952
rect 390377 -16008 390448 -15952
rect 390108 -16094 390448 -16008
rect 390108 -16150 390179 -16094
rect 390235 -16150 390321 -16094
rect 390377 -16150 390448 -16094
rect 390108 -16236 390448 -16150
rect 390108 -16292 390179 -16236
rect 390235 -16292 390321 -16236
rect 390377 -16292 390448 -16236
rect 390108 -16378 390448 -16292
rect 390108 -16434 390179 -16378
rect 390235 -16434 390321 -16378
rect 390377 -16434 390448 -16378
rect 390108 -16520 390448 -16434
rect 390108 -16576 390179 -16520
rect 390235 -16576 390321 -16520
rect 390377 -16576 390448 -16520
rect 390108 -16662 390448 -16576
rect 390108 -16718 390179 -16662
rect 390235 -16718 390321 -16662
rect 390377 -16718 390448 -16662
rect 390108 -16804 390448 -16718
rect 390108 -16860 390179 -16804
rect 390235 -16860 390321 -16804
rect 390377 -16860 390448 -16804
rect 390108 -16946 390448 -16860
rect 390108 -17002 390179 -16946
rect 390235 -17002 390321 -16946
rect 390377 -17002 390448 -16946
rect 390108 -17088 390448 -17002
rect 390108 -17144 390179 -17088
rect 390235 -17144 390321 -17088
rect 390377 -17144 390448 -17088
rect 390108 -17230 390448 -17144
rect 390108 -17286 390179 -17230
rect 390235 -17286 390321 -17230
rect 390377 -17286 390448 -17230
rect 390108 -17372 390448 -17286
rect 390108 -17428 390179 -17372
rect 390235 -17428 390321 -17372
rect 390377 -17428 390448 -17372
rect 390108 -17514 390448 -17428
rect 390108 -17570 390179 -17514
rect 390235 -17570 390321 -17514
rect 390377 -17570 390448 -17514
rect 390108 -17656 390448 -17570
rect 390108 -17712 390179 -17656
rect 390235 -17712 390321 -17656
rect 390377 -17712 390448 -17656
rect 390108 -17798 390448 -17712
rect 390108 -17854 390179 -17798
rect 390235 -17854 390321 -17798
rect 390377 -17854 390448 -17798
rect 390108 -17940 390448 -17854
rect 390108 -17996 390179 -17940
rect 390235 -17996 390321 -17940
rect 390377 -17996 390448 -17940
rect 390108 -18082 390448 -17996
rect 390108 -18138 390179 -18082
rect 390235 -18138 390321 -18082
rect 390377 -18138 390448 -18082
rect 390108 -18224 390448 -18138
rect 390108 -18280 390179 -18224
rect 390235 -18280 390321 -18224
rect 390377 -18280 390448 -18224
rect 390108 -18366 390448 -18280
rect 390108 -18422 390179 -18366
rect 390235 -18422 390321 -18366
rect 390377 -18422 390448 -18366
rect 390108 -18508 390448 -18422
rect 390108 -18564 390179 -18508
rect 390235 -18564 390321 -18508
rect 390377 -18564 390448 -18508
rect 390108 -18650 390448 -18564
rect 390108 -18706 390179 -18650
rect 390235 -18706 390321 -18650
rect 390377 -18706 390448 -18650
rect 390108 -18792 390448 -18706
rect 390108 -18848 390179 -18792
rect 390235 -18848 390321 -18792
rect 390377 -18848 390448 -18792
rect 390108 -18934 390448 -18848
rect 390108 -18990 390179 -18934
rect 390235 -18990 390321 -18934
rect 390377 -18990 390448 -18934
rect 390108 -19076 390448 -18990
rect 390108 -19132 390179 -19076
rect 390235 -19132 390321 -19076
rect 390377 -19132 390448 -19076
rect 390108 -19218 390448 -19132
rect 390108 -19274 390179 -19218
rect 390235 -19274 390321 -19218
rect 390377 -19274 390448 -19218
rect 390108 -19360 390448 -19274
rect 390108 -19416 390179 -19360
rect 390235 -19416 390321 -19360
rect 390377 -19416 390448 -19360
rect 390108 -19502 390448 -19416
rect 390108 -19558 390179 -19502
rect 390235 -19558 390321 -19502
rect 390377 -19558 390448 -19502
rect 390108 -19644 390448 -19558
rect 390108 -19700 390179 -19644
rect 390235 -19700 390321 -19644
rect 390377 -19700 390448 -19644
rect 390108 -19786 390448 -19700
rect 390108 -19842 390179 -19786
rect 390235 -19842 390321 -19786
rect 390377 -19842 390448 -19786
rect 390108 -19928 390448 -19842
rect 390108 -19984 390179 -19928
rect 390235 -19984 390321 -19928
rect 390377 -19984 390448 -19928
rect 390108 -20070 390448 -19984
rect 390108 -20126 390179 -20070
rect 390235 -20126 390321 -20070
rect 390377 -20126 390448 -20070
rect 390108 -20212 390448 -20126
rect 390108 -20268 390179 -20212
rect 390235 -20268 390321 -20212
rect 390377 -20268 390448 -20212
rect 390108 -20354 390448 -20268
rect 390108 -20410 390179 -20354
rect 390235 -20410 390321 -20354
rect 390377 -20410 390448 -20354
rect 390108 -20496 390448 -20410
rect 390108 -20552 390179 -20496
rect 390235 -20552 390321 -20496
rect 390377 -20552 390448 -20496
rect 390108 -20638 390448 -20552
rect 390108 -20694 390179 -20638
rect 390235 -20694 390321 -20638
rect 390377 -20694 390448 -20638
rect 390108 -20780 390448 -20694
rect 390108 -20836 390179 -20780
rect 390235 -20836 390321 -20780
rect 390377 -20836 390448 -20780
rect 390108 -20922 390448 -20836
rect 390108 -20978 390179 -20922
rect 390235 -20978 390321 -20922
rect 390377 -20978 390448 -20922
rect 390108 -21064 390448 -20978
rect 390108 -21120 390179 -21064
rect 390235 -21120 390321 -21064
rect 390377 -21120 390448 -21064
rect 390108 -21206 390448 -21120
rect 390108 -21262 390179 -21206
rect 390235 -21262 390321 -21206
rect 390377 -21262 390448 -21206
rect 390108 -21348 390448 -21262
rect 390108 -21404 390179 -21348
rect 390235 -21404 390321 -21348
rect 390377 -21404 390448 -21348
rect 390108 -21490 390448 -21404
rect 390108 -21546 390179 -21490
rect 390235 -21546 390321 -21490
rect 390377 -21546 390448 -21490
rect 390108 -21632 390448 -21546
rect 390108 -21688 390179 -21632
rect 390235 -21688 390321 -21632
rect 390377 -21688 390448 -21632
rect 390108 -21774 390448 -21688
rect 390108 -21830 390179 -21774
rect 390235 -21830 390321 -21774
rect 390377 -21830 390448 -21774
rect 390108 -21916 390448 -21830
rect 390108 -21972 390179 -21916
rect 390235 -21972 390321 -21916
rect 390377 -21972 390448 -21916
rect 390108 -22058 390448 -21972
rect 390108 -22114 390179 -22058
rect 390235 -22114 390321 -22058
rect 390377 -22114 390448 -22058
rect 390108 -22200 390448 -22114
rect 390108 -22256 390179 -22200
rect 390235 -22256 390321 -22200
rect 390377 -22256 390448 -22200
rect 390108 -22342 390448 -22256
rect 390108 -22398 390179 -22342
rect 390235 -22398 390321 -22342
rect 390377 -22398 390448 -22342
rect 390108 -22484 390448 -22398
rect 390108 -22540 390179 -22484
rect 390235 -22540 390321 -22484
rect 390377 -22540 390448 -22484
rect 390108 -22626 390448 -22540
rect 390108 -22682 390179 -22626
rect 390235 -22682 390321 -22626
rect 390377 -22682 390448 -22626
rect 390108 -22768 390448 -22682
rect 390108 -22824 390179 -22768
rect 390235 -22824 390321 -22768
rect 390377 -22824 390448 -22768
rect 390108 -22910 390448 -22824
rect 390108 -22966 390179 -22910
rect 390235 -22966 390321 -22910
rect 390377 -22966 390448 -22910
rect 390108 -23052 390448 -22966
rect 390108 -23108 390179 -23052
rect 390235 -23108 390321 -23052
rect 390377 -23108 390448 -23052
rect 390108 -23194 390448 -23108
rect 390108 -23250 390179 -23194
rect 390235 -23250 390321 -23194
rect 390377 -23250 390448 -23194
rect 390108 -23336 390448 -23250
rect 390108 -23392 390179 -23336
rect 390235 -23392 390321 -23336
rect 390377 -23392 390448 -23336
rect 390108 -23478 390448 -23392
rect 390108 -23534 390179 -23478
rect 390235 -23534 390321 -23478
rect 390377 -23534 390448 -23478
rect 390108 -23620 390448 -23534
rect 390108 -23676 390179 -23620
rect 390235 -23676 390321 -23620
rect 390377 -23676 390448 -23620
rect 390108 -23762 390448 -23676
rect 390108 -23818 390179 -23762
rect 390235 -23818 390321 -23762
rect 390377 -23818 390448 -23762
rect 390108 -23904 390448 -23818
rect 390108 -23960 390179 -23904
rect 390235 -23960 390321 -23904
rect 390377 -23960 390448 -23904
rect 390108 -24046 390448 -23960
rect 390108 -24102 390179 -24046
rect 390235 -24102 390321 -24046
rect 390377 -24102 390448 -24046
rect 390108 -24188 390448 -24102
rect 390108 -24244 390179 -24188
rect 390235 -24244 390321 -24188
rect 390377 -24244 390448 -24188
rect 390108 -24330 390448 -24244
rect 390108 -24386 390179 -24330
rect 390235 -24386 390321 -24330
rect 390377 -24386 390448 -24330
rect 390108 -24472 390448 -24386
rect 390108 -24528 390179 -24472
rect 390235 -24528 390321 -24472
rect 390377 -24528 390448 -24472
rect 390108 -24614 390448 -24528
rect 390108 -24670 390179 -24614
rect 390235 -24670 390321 -24614
rect 390377 -24670 390448 -24614
rect 390108 -24756 390448 -24670
rect 390108 -24812 390179 -24756
rect 390235 -24812 390321 -24756
rect 390377 -24812 390448 -24756
rect 390108 -24898 390448 -24812
rect 390108 -24954 390179 -24898
rect 390235 -24954 390321 -24898
rect 390377 -24954 390448 -24898
rect 390108 -25040 390448 -24954
rect 390108 -25096 390179 -25040
rect 390235 -25096 390321 -25040
rect 390377 -25096 390448 -25040
rect 390108 -25182 390448 -25096
rect 390108 -25238 390179 -25182
rect 390235 -25238 390321 -25182
rect 390377 -25238 390448 -25182
rect 390108 -25324 390448 -25238
rect 390108 -25380 390179 -25324
rect 390235 -25380 390321 -25324
rect 390377 -25380 390448 -25324
rect 390108 -25466 390448 -25380
rect 390108 -25522 390179 -25466
rect 390235 -25522 390321 -25466
rect 390377 -25522 390448 -25466
rect 390108 -25532 390448 -25522
rect 390508 -13680 390848 -13670
rect 390508 -13736 390576 -13680
rect 390632 -13736 390718 -13680
rect 390774 -13736 390848 -13680
rect 390508 -13822 390848 -13736
rect 390508 -13878 390576 -13822
rect 390632 -13878 390718 -13822
rect 390774 -13878 390848 -13822
rect 390508 -13964 390848 -13878
rect 390508 -14020 390576 -13964
rect 390632 -14020 390718 -13964
rect 390774 -14020 390848 -13964
rect 390508 -14106 390848 -14020
rect 390508 -14162 390576 -14106
rect 390632 -14162 390718 -14106
rect 390774 -14162 390848 -14106
rect 390508 -14248 390848 -14162
rect 390508 -14304 390576 -14248
rect 390632 -14304 390718 -14248
rect 390774 -14304 390848 -14248
rect 390508 -14390 390848 -14304
rect 390508 -14446 390576 -14390
rect 390632 -14446 390718 -14390
rect 390774 -14446 390848 -14390
rect 390508 -14532 390848 -14446
rect 390508 -14588 390576 -14532
rect 390632 -14588 390718 -14532
rect 390774 -14588 390848 -14532
rect 390508 -14674 390848 -14588
rect 390508 -14730 390576 -14674
rect 390632 -14730 390718 -14674
rect 390774 -14730 390848 -14674
rect 390508 -14816 390848 -14730
rect 390508 -14872 390576 -14816
rect 390632 -14872 390718 -14816
rect 390774 -14872 390848 -14816
rect 390508 -14958 390848 -14872
rect 390508 -15014 390576 -14958
rect 390632 -15014 390718 -14958
rect 390774 -15014 390848 -14958
rect 390508 -15100 390848 -15014
rect 390508 -15156 390576 -15100
rect 390632 -15156 390718 -15100
rect 390774 -15156 390848 -15100
rect 390508 -15242 390848 -15156
rect 390508 -15298 390576 -15242
rect 390632 -15298 390718 -15242
rect 390774 -15298 390848 -15242
rect 390508 -15384 390848 -15298
rect 390508 -15440 390576 -15384
rect 390632 -15440 390718 -15384
rect 390774 -15440 390848 -15384
rect 390508 -15526 390848 -15440
rect 390508 -15582 390576 -15526
rect 390632 -15582 390718 -15526
rect 390774 -15582 390848 -15526
rect 390508 -15668 390848 -15582
rect 390508 -15724 390576 -15668
rect 390632 -15724 390718 -15668
rect 390774 -15724 390848 -15668
rect 390508 -15810 390848 -15724
rect 390508 -15866 390576 -15810
rect 390632 -15866 390718 -15810
rect 390774 -15866 390848 -15810
rect 390508 -15952 390848 -15866
rect 390508 -16008 390576 -15952
rect 390632 -16008 390718 -15952
rect 390774 -16008 390848 -15952
rect 390508 -16094 390848 -16008
rect 390508 -16150 390576 -16094
rect 390632 -16150 390718 -16094
rect 390774 -16150 390848 -16094
rect 390508 -16236 390848 -16150
rect 390508 -16292 390576 -16236
rect 390632 -16292 390718 -16236
rect 390774 -16292 390848 -16236
rect 390508 -16378 390848 -16292
rect 390508 -16434 390576 -16378
rect 390632 -16434 390718 -16378
rect 390774 -16434 390848 -16378
rect 390508 -16520 390848 -16434
rect 390508 -16576 390576 -16520
rect 390632 -16576 390718 -16520
rect 390774 -16576 390848 -16520
rect 390508 -16662 390848 -16576
rect 390508 -16718 390576 -16662
rect 390632 -16718 390718 -16662
rect 390774 -16718 390848 -16662
rect 390508 -16804 390848 -16718
rect 390508 -16860 390576 -16804
rect 390632 -16860 390718 -16804
rect 390774 -16860 390848 -16804
rect 390508 -16946 390848 -16860
rect 390508 -17002 390576 -16946
rect 390632 -17002 390718 -16946
rect 390774 -17002 390848 -16946
rect 390508 -17088 390848 -17002
rect 390508 -17144 390576 -17088
rect 390632 -17144 390718 -17088
rect 390774 -17144 390848 -17088
rect 390508 -17230 390848 -17144
rect 390508 -17286 390576 -17230
rect 390632 -17286 390718 -17230
rect 390774 -17286 390848 -17230
rect 390508 -17372 390848 -17286
rect 390508 -17428 390576 -17372
rect 390632 -17428 390718 -17372
rect 390774 -17428 390848 -17372
rect 390508 -17514 390848 -17428
rect 390508 -17570 390576 -17514
rect 390632 -17570 390718 -17514
rect 390774 -17570 390848 -17514
rect 390508 -17656 390848 -17570
rect 390508 -17712 390576 -17656
rect 390632 -17712 390718 -17656
rect 390774 -17712 390848 -17656
rect 390508 -17798 390848 -17712
rect 390508 -17854 390576 -17798
rect 390632 -17854 390718 -17798
rect 390774 -17854 390848 -17798
rect 390508 -17940 390848 -17854
rect 390508 -17996 390576 -17940
rect 390632 -17996 390718 -17940
rect 390774 -17996 390848 -17940
rect 390508 -18082 390848 -17996
rect 390508 -18138 390576 -18082
rect 390632 -18138 390718 -18082
rect 390774 -18138 390848 -18082
rect 390508 -18224 390848 -18138
rect 390508 -18280 390576 -18224
rect 390632 -18280 390718 -18224
rect 390774 -18280 390848 -18224
rect 390508 -18366 390848 -18280
rect 390508 -18422 390576 -18366
rect 390632 -18422 390718 -18366
rect 390774 -18422 390848 -18366
rect 390508 -18508 390848 -18422
rect 390508 -18564 390576 -18508
rect 390632 -18564 390718 -18508
rect 390774 -18564 390848 -18508
rect 390508 -18650 390848 -18564
rect 390508 -18706 390576 -18650
rect 390632 -18706 390718 -18650
rect 390774 -18706 390848 -18650
rect 390508 -18792 390848 -18706
rect 390508 -18848 390576 -18792
rect 390632 -18848 390718 -18792
rect 390774 -18848 390848 -18792
rect 390508 -18934 390848 -18848
rect 390508 -18990 390576 -18934
rect 390632 -18990 390718 -18934
rect 390774 -18990 390848 -18934
rect 390508 -19076 390848 -18990
rect 390508 -19132 390576 -19076
rect 390632 -19132 390718 -19076
rect 390774 -19132 390848 -19076
rect 390508 -19218 390848 -19132
rect 390508 -19274 390576 -19218
rect 390632 -19274 390718 -19218
rect 390774 -19274 390848 -19218
rect 390508 -19360 390848 -19274
rect 390508 -19416 390576 -19360
rect 390632 -19416 390718 -19360
rect 390774 -19416 390848 -19360
rect 390508 -19502 390848 -19416
rect 390508 -19558 390576 -19502
rect 390632 -19558 390718 -19502
rect 390774 -19558 390848 -19502
rect 390508 -19644 390848 -19558
rect 390508 -19700 390576 -19644
rect 390632 -19700 390718 -19644
rect 390774 -19700 390848 -19644
rect 390508 -19786 390848 -19700
rect 390508 -19842 390576 -19786
rect 390632 -19842 390718 -19786
rect 390774 -19842 390848 -19786
rect 390508 -19928 390848 -19842
rect 390508 -19984 390576 -19928
rect 390632 -19984 390718 -19928
rect 390774 -19984 390848 -19928
rect 390508 -20070 390848 -19984
rect 390508 -20126 390576 -20070
rect 390632 -20126 390718 -20070
rect 390774 -20126 390848 -20070
rect 390508 -20212 390848 -20126
rect 390508 -20268 390576 -20212
rect 390632 -20268 390718 -20212
rect 390774 -20268 390848 -20212
rect 390508 -20354 390848 -20268
rect 390508 -20410 390576 -20354
rect 390632 -20410 390718 -20354
rect 390774 -20410 390848 -20354
rect 390508 -20496 390848 -20410
rect 390508 -20552 390576 -20496
rect 390632 -20552 390718 -20496
rect 390774 -20552 390848 -20496
rect 390508 -20638 390848 -20552
rect 390508 -20694 390576 -20638
rect 390632 -20694 390718 -20638
rect 390774 -20694 390848 -20638
rect 390508 -20780 390848 -20694
rect 390508 -20836 390576 -20780
rect 390632 -20836 390718 -20780
rect 390774 -20836 390848 -20780
rect 390508 -20922 390848 -20836
rect 390508 -20978 390576 -20922
rect 390632 -20978 390718 -20922
rect 390774 -20978 390848 -20922
rect 390508 -21064 390848 -20978
rect 390508 -21120 390576 -21064
rect 390632 -21120 390718 -21064
rect 390774 -21120 390848 -21064
rect 390508 -21206 390848 -21120
rect 390508 -21262 390576 -21206
rect 390632 -21262 390718 -21206
rect 390774 -21262 390848 -21206
rect 390508 -21348 390848 -21262
rect 390508 -21404 390576 -21348
rect 390632 -21404 390718 -21348
rect 390774 -21404 390848 -21348
rect 390508 -21490 390848 -21404
rect 390508 -21546 390576 -21490
rect 390632 -21546 390718 -21490
rect 390774 -21546 390848 -21490
rect 390508 -21632 390848 -21546
rect 390508 -21688 390576 -21632
rect 390632 -21688 390718 -21632
rect 390774 -21688 390848 -21632
rect 390508 -21774 390848 -21688
rect 390508 -21830 390576 -21774
rect 390632 -21830 390718 -21774
rect 390774 -21830 390848 -21774
rect 390508 -21916 390848 -21830
rect 390508 -21972 390576 -21916
rect 390632 -21972 390718 -21916
rect 390774 -21972 390848 -21916
rect 390508 -22058 390848 -21972
rect 390508 -22114 390576 -22058
rect 390632 -22114 390718 -22058
rect 390774 -22114 390848 -22058
rect 390508 -22200 390848 -22114
rect 390508 -22256 390576 -22200
rect 390632 -22256 390718 -22200
rect 390774 -22256 390848 -22200
rect 390508 -22342 390848 -22256
rect 390508 -22398 390576 -22342
rect 390632 -22398 390718 -22342
rect 390774 -22398 390848 -22342
rect 390508 -22484 390848 -22398
rect 390508 -22540 390576 -22484
rect 390632 -22540 390718 -22484
rect 390774 -22540 390848 -22484
rect 390508 -22626 390848 -22540
rect 390508 -22682 390576 -22626
rect 390632 -22682 390718 -22626
rect 390774 -22682 390848 -22626
rect 390508 -22768 390848 -22682
rect 390508 -22824 390576 -22768
rect 390632 -22824 390718 -22768
rect 390774 -22824 390848 -22768
rect 390508 -22910 390848 -22824
rect 390508 -22966 390576 -22910
rect 390632 -22966 390718 -22910
rect 390774 -22966 390848 -22910
rect 390508 -23052 390848 -22966
rect 390508 -23108 390576 -23052
rect 390632 -23108 390718 -23052
rect 390774 -23108 390848 -23052
rect 390508 -23194 390848 -23108
rect 390508 -23250 390576 -23194
rect 390632 -23250 390718 -23194
rect 390774 -23250 390848 -23194
rect 390508 -23336 390848 -23250
rect 390508 -23392 390576 -23336
rect 390632 -23392 390718 -23336
rect 390774 -23392 390848 -23336
rect 390508 -23478 390848 -23392
rect 390508 -23534 390576 -23478
rect 390632 -23534 390718 -23478
rect 390774 -23534 390848 -23478
rect 390508 -23620 390848 -23534
rect 390508 -23676 390576 -23620
rect 390632 -23676 390718 -23620
rect 390774 -23676 390848 -23620
rect 390508 -23762 390848 -23676
rect 390508 -23818 390576 -23762
rect 390632 -23818 390718 -23762
rect 390774 -23818 390848 -23762
rect 390508 -23904 390848 -23818
rect 390508 -23960 390576 -23904
rect 390632 -23960 390718 -23904
rect 390774 -23960 390848 -23904
rect 390508 -24046 390848 -23960
rect 390508 -24102 390576 -24046
rect 390632 -24102 390718 -24046
rect 390774 -24102 390848 -24046
rect 390508 -24188 390848 -24102
rect 390508 -24244 390576 -24188
rect 390632 -24244 390718 -24188
rect 390774 -24244 390848 -24188
rect 390508 -24330 390848 -24244
rect 390508 -24386 390576 -24330
rect 390632 -24386 390718 -24330
rect 390774 -24386 390848 -24330
rect 390508 -24472 390848 -24386
rect 390508 -24528 390576 -24472
rect 390632 -24528 390718 -24472
rect 390774 -24528 390848 -24472
rect 390508 -24614 390848 -24528
rect 390508 -24670 390576 -24614
rect 390632 -24670 390718 -24614
rect 390774 -24670 390848 -24614
rect 390508 -24756 390848 -24670
rect 390508 -24812 390576 -24756
rect 390632 -24812 390718 -24756
rect 390774 -24812 390848 -24756
rect 390508 -24898 390848 -24812
rect 390508 -24954 390576 -24898
rect 390632 -24954 390718 -24898
rect 390774 -24954 390848 -24898
rect 390508 -25040 390848 -24954
rect 390508 -25096 390576 -25040
rect 390632 -25096 390718 -25040
rect 390774 -25096 390848 -25040
rect 390508 -25182 390848 -25096
rect 390508 -25238 390576 -25182
rect 390632 -25238 390718 -25182
rect 390774 -25238 390848 -25182
rect 390508 -25324 390848 -25238
rect 390508 -25380 390576 -25324
rect 390632 -25380 390718 -25324
rect 390774 -25380 390848 -25324
rect 390508 -25466 390848 -25380
rect 390508 -25522 390576 -25466
rect 390632 -25522 390718 -25466
rect 390774 -25522 390848 -25466
rect 390508 -25532 390848 -25522
rect 390908 -13680 391248 -13670
rect 390908 -13736 390980 -13680
rect 391036 -13736 391122 -13680
rect 391178 -13736 391248 -13680
rect 390908 -13822 391248 -13736
rect 390908 -13878 390980 -13822
rect 391036 -13878 391122 -13822
rect 391178 -13878 391248 -13822
rect 390908 -13964 391248 -13878
rect 390908 -14020 390980 -13964
rect 391036 -14020 391122 -13964
rect 391178 -14020 391248 -13964
rect 390908 -14106 391248 -14020
rect 390908 -14162 390980 -14106
rect 391036 -14162 391122 -14106
rect 391178 -14162 391248 -14106
rect 390908 -14248 391248 -14162
rect 390908 -14304 390980 -14248
rect 391036 -14304 391122 -14248
rect 391178 -14304 391248 -14248
rect 390908 -14390 391248 -14304
rect 390908 -14446 390980 -14390
rect 391036 -14446 391122 -14390
rect 391178 -14446 391248 -14390
rect 390908 -14532 391248 -14446
rect 390908 -14588 390980 -14532
rect 391036 -14588 391122 -14532
rect 391178 -14588 391248 -14532
rect 390908 -14674 391248 -14588
rect 390908 -14730 390980 -14674
rect 391036 -14730 391122 -14674
rect 391178 -14730 391248 -14674
rect 390908 -14816 391248 -14730
rect 390908 -14872 390980 -14816
rect 391036 -14872 391122 -14816
rect 391178 -14872 391248 -14816
rect 390908 -14958 391248 -14872
rect 390908 -15014 390980 -14958
rect 391036 -15014 391122 -14958
rect 391178 -15014 391248 -14958
rect 390908 -15100 391248 -15014
rect 390908 -15156 390980 -15100
rect 391036 -15156 391122 -15100
rect 391178 -15156 391248 -15100
rect 390908 -15242 391248 -15156
rect 390908 -15298 390980 -15242
rect 391036 -15298 391122 -15242
rect 391178 -15298 391248 -15242
rect 390908 -15384 391248 -15298
rect 390908 -15440 390980 -15384
rect 391036 -15440 391122 -15384
rect 391178 -15440 391248 -15384
rect 390908 -15526 391248 -15440
rect 390908 -15582 390980 -15526
rect 391036 -15582 391122 -15526
rect 391178 -15582 391248 -15526
rect 390908 -15668 391248 -15582
rect 390908 -15724 390980 -15668
rect 391036 -15724 391122 -15668
rect 391178 -15724 391248 -15668
rect 390908 -15810 391248 -15724
rect 390908 -15866 390980 -15810
rect 391036 -15866 391122 -15810
rect 391178 -15866 391248 -15810
rect 390908 -15952 391248 -15866
rect 390908 -16008 390980 -15952
rect 391036 -16008 391122 -15952
rect 391178 -16008 391248 -15952
rect 390908 -16094 391248 -16008
rect 390908 -16150 390980 -16094
rect 391036 -16150 391122 -16094
rect 391178 -16150 391248 -16094
rect 390908 -16236 391248 -16150
rect 390908 -16292 390980 -16236
rect 391036 -16292 391122 -16236
rect 391178 -16292 391248 -16236
rect 390908 -16378 391248 -16292
rect 390908 -16434 390980 -16378
rect 391036 -16434 391122 -16378
rect 391178 -16434 391248 -16378
rect 390908 -16520 391248 -16434
rect 390908 -16576 390980 -16520
rect 391036 -16576 391122 -16520
rect 391178 -16576 391248 -16520
rect 390908 -16662 391248 -16576
rect 390908 -16718 390980 -16662
rect 391036 -16718 391122 -16662
rect 391178 -16718 391248 -16662
rect 390908 -16804 391248 -16718
rect 390908 -16860 390980 -16804
rect 391036 -16860 391122 -16804
rect 391178 -16860 391248 -16804
rect 390908 -16946 391248 -16860
rect 390908 -17002 390980 -16946
rect 391036 -17002 391122 -16946
rect 391178 -17002 391248 -16946
rect 390908 -17088 391248 -17002
rect 390908 -17144 390980 -17088
rect 391036 -17144 391122 -17088
rect 391178 -17144 391248 -17088
rect 390908 -17230 391248 -17144
rect 390908 -17286 390980 -17230
rect 391036 -17286 391122 -17230
rect 391178 -17286 391248 -17230
rect 390908 -17372 391248 -17286
rect 390908 -17428 390980 -17372
rect 391036 -17428 391122 -17372
rect 391178 -17428 391248 -17372
rect 390908 -17514 391248 -17428
rect 390908 -17570 390980 -17514
rect 391036 -17570 391122 -17514
rect 391178 -17570 391248 -17514
rect 390908 -17656 391248 -17570
rect 390908 -17712 390980 -17656
rect 391036 -17712 391122 -17656
rect 391178 -17712 391248 -17656
rect 390908 -17798 391248 -17712
rect 390908 -17854 390980 -17798
rect 391036 -17854 391122 -17798
rect 391178 -17854 391248 -17798
rect 390908 -17940 391248 -17854
rect 390908 -17996 390980 -17940
rect 391036 -17996 391122 -17940
rect 391178 -17996 391248 -17940
rect 390908 -18082 391248 -17996
rect 390908 -18138 390980 -18082
rect 391036 -18138 391122 -18082
rect 391178 -18138 391248 -18082
rect 390908 -18224 391248 -18138
rect 390908 -18280 390980 -18224
rect 391036 -18280 391122 -18224
rect 391178 -18280 391248 -18224
rect 390908 -18366 391248 -18280
rect 390908 -18422 390980 -18366
rect 391036 -18422 391122 -18366
rect 391178 -18422 391248 -18366
rect 390908 -18508 391248 -18422
rect 390908 -18564 390980 -18508
rect 391036 -18564 391122 -18508
rect 391178 -18564 391248 -18508
rect 390908 -18650 391248 -18564
rect 390908 -18706 390980 -18650
rect 391036 -18706 391122 -18650
rect 391178 -18706 391248 -18650
rect 390908 -18792 391248 -18706
rect 390908 -18848 390980 -18792
rect 391036 -18848 391122 -18792
rect 391178 -18848 391248 -18792
rect 390908 -18934 391248 -18848
rect 390908 -18990 390980 -18934
rect 391036 -18990 391122 -18934
rect 391178 -18990 391248 -18934
rect 390908 -19076 391248 -18990
rect 390908 -19132 390980 -19076
rect 391036 -19132 391122 -19076
rect 391178 -19132 391248 -19076
rect 390908 -19218 391248 -19132
rect 390908 -19274 390980 -19218
rect 391036 -19274 391122 -19218
rect 391178 -19274 391248 -19218
rect 390908 -19360 391248 -19274
rect 390908 -19416 390980 -19360
rect 391036 -19416 391122 -19360
rect 391178 -19416 391248 -19360
rect 390908 -19502 391248 -19416
rect 390908 -19558 390980 -19502
rect 391036 -19558 391122 -19502
rect 391178 -19558 391248 -19502
rect 390908 -19644 391248 -19558
rect 390908 -19700 390980 -19644
rect 391036 -19700 391122 -19644
rect 391178 -19700 391248 -19644
rect 390908 -19786 391248 -19700
rect 390908 -19842 390980 -19786
rect 391036 -19842 391122 -19786
rect 391178 -19842 391248 -19786
rect 390908 -19928 391248 -19842
rect 390908 -19984 390980 -19928
rect 391036 -19984 391122 -19928
rect 391178 -19984 391248 -19928
rect 390908 -20070 391248 -19984
rect 390908 -20126 390980 -20070
rect 391036 -20126 391122 -20070
rect 391178 -20126 391248 -20070
rect 390908 -20212 391248 -20126
rect 390908 -20268 390980 -20212
rect 391036 -20268 391122 -20212
rect 391178 -20268 391248 -20212
rect 390908 -20354 391248 -20268
rect 390908 -20410 390980 -20354
rect 391036 -20410 391122 -20354
rect 391178 -20410 391248 -20354
rect 390908 -20496 391248 -20410
rect 390908 -20552 390980 -20496
rect 391036 -20552 391122 -20496
rect 391178 -20552 391248 -20496
rect 390908 -20638 391248 -20552
rect 390908 -20694 390980 -20638
rect 391036 -20694 391122 -20638
rect 391178 -20694 391248 -20638
rect 390908 -20780 391248 -20694
rect 390908 -20836 390980 -20780
rect 391036 -20836 391122 -20780
rect 391178 -20836 391248 -20780
rect 390908 -20922 391248 -20836
rect 390908 -20978 390980 -20922
rect 391036 -20978 391122 -20922
rect 391178 -20978 391248 -20922
rect 390908 -21064 391248 -20978
rect 390908 -21120 390980 -21064
rect 391036 -21120 391122 -21064
rect 391178 -21120 391248 -21064
rect 390908 -21206 391248 -21120
rect 390908 -21262 390980 -21206
rect 391036 -21262 391122 -21206
rect 391178 -21262 391248 -21206
rect 390908 -21348 391248 -21262
rect 390908 -21404 390980 -21348
rect 391036 -21404 391122 -21348
rect 391178 -21404 391248 -21348
rect 390908 -21490 391248 -21404
rect 390908 -21546 390980 -21490
rect 391036 -21546 391122 -21490
rect 391178 -21546 391248 -21490
rect 390908 -21632 391248 -21546
rect 390908 -21688 390980 -21632
rect 391036 -21688 391122 -21632
rect 391178 -21688 391248 -21632
rect 390908 -21774 391248 -21688
rect 390908 -21830 390980 -21774
rect 391036 -21830 391122 -21774
rect 391178 -21830 391248 -21774
rect 390908 -21916 391248 -21830
rect 390908 -21972 390980 -21916
rect 391036 -21972 391122 -21916
rect 391178 -21972 391248 -21916
rect 390908 -22058 391248 -21972
rect 390908 -22114 390980 -22058
rect 391036 -22114 391122 -22058
rect 391178 -22114 391248 -22058
rect 390908 -22200 391248 -22114
rect 390908 -22256 390980 -22200
rect 391036 -22256 391122 -22200
rect 391178 -22256 391248 -22200
rect 390908 -22342 391248 -22256
rect 390908 -22398 390980 -22342
rect 391036 -22398 391122 -22342
rect 391178 -22398 391248 -22342
rect 390908 -22484 391248 -22398
rect 390908 -22540 390980 -22484
rect 391036 -22540 391122 -22484
rect 391178 -22540 391248 -22484
rect 390908 -22626 391248 -22540
rect 390908 -22682 390980 -22626
rect 391036 -22682 391122 -22626
rect 391178 -22682 391248 -22626
rect 390908 -22768 391248 -22682
rect 390908 -22824 390980 -22768
rect 391036 -22824 391122 -22768
rect 391178 -22824 391248 -22768
rect 390908 -22910 391248 -22824
rect 390908 -22966 390980 -22910
rect 391036 -22966 391122 -22910
rect 391178 -22966 391248 -22910
rect 390908 -23052 391248 -22966
rect 390908 -23108 390980 -23052
rect 391036 -23108 391122 -23052
rect 391178 -23108 391248 -23052
rect 390908 -23194 391248 -23108
rect 390908 -23250 390980 -23194
rect 391036 -23250 391122 -23194
rect 391178 -23250 391248 -23194
rect 390908 -23336 391248 -23250
rect 390908 -23392 390980 -23336
rect 391036 -23392 391122 -23336
rect 391178 -23392 391248 -23336
rect 390908 -23478 391248 -23392
rect 390908 -23534 390980 -23478
rect 391036 -23534 391122 -23478
rect 391178 -23534 391248 -23478
rect 390908 -23620 391248 -23534
rect 390908 -23676 390980 -23620
rect 391036 -23676 391122 -23620
rect 391178 -23676 391248 -23620
rect 390908 -23762 391248 -23676
rect 390908 -23818 390980 -23762
rect 391036 -23818 391122 -23762
rect 391178 -23818 391248 -23762
rect 390908 -23904 391248 -23818
rect 390908 -23960 390980 -23904
rect 391036 -23960 391122 -23904
rect 391178 -23960 391248 -23904
rect 390908 -24046 391248 -23960
rect 390908 -24102 390980 -24046
rect 391036 -24102 391122 -24046
rect 391178 -24102 391248 -24046
rect 390908 -24188 391248 -24102
rect 390908 -24244 390980 -24188
rect 391036 -24244 391122 -24188
rect 391178 -24244 391248 -24188
rect 390908 -24330 391248 -24244
rect 390908 -24386 390980 -24330
rect 391036 -24386 391122 -24330
rect 391178 -24386 391248 -24330
rect 390908 -24472 391248 -24386
rect 390908 -24528 390980 -24472
rect 391036 -24528 391122 -24472
rect 391178 -24528 391248 -24472
rect 390908 -24614 391248 -24528
rect 390908 -24670 390980 -24614
rect 391036 -24670 391122 -24614
rect 391178 -24670 391248 -24614
rect 390908 -24756 391248 -24670
rect 390908 -24812 390980 -24756
rect 391036 -24812 391122 -24756
rect 391178 -24812 391248 -24756
rect 390908 -24898 391248 -24812
rect 390908 -24954 390980 -24898
rect 391036 -24954 391122 -24898
rect 391178 -24954 391248 -24898
rect 390908 -25040 391248 -24954
rect 390908 -25096 390980 -25040
rect 391036 -25096 391122 -25040
rect 391178 -25096 391248 -25040
rect 390908 -25182 391248 -25096
rect 390908 -25238 390980 -25182
rect 391036 -25238 391122 -25182
rect 391178 -25238 391248 -25182
rect 390908 -25324 391248 -25238
rect 390908 -25380 390980 -25324
rect 391036 -25380 391122 -25324
rect 391178 -25380 391248 -25324
rect 390908 -25466 391248 -25380
rect 390908 -25522 390980 -25466
rect 391036 -25522 391122 -25466
rect 391178 -25522 391248 -25466
rect 390908 -25532 391248 -25522
rect 391308 -13680 391648 -13670
rect 391308 -13736 391376 -13680
rect 391432 -13736 391518 -13680
rect 391574 -13736 391648 -13680
rect 391308 -13822 391648 -13736
rect 391308 -13878 391376 -13822
rect 391432 -13878 391518 -13822
rect 391574 -13878 391648 -13822
rect 391308 -13964 391648 -13878
rect 391308 -14020 391376 -13964
rect 391432 -14020 391518 -13964
rect 391574 -14020 391648 -13964
rect 391308 -14106 391648 -14020
rect 391308 -14162 391376 -14106
rect 391432 -14162 391518 -14106
rect 391574 -14162 391648 -14106
rect 391308 -14248 391648 -14162
rect 391308 -14304 391376 -14248
rect 391432 -14304 391518 -14248
rect 391574 -14304 391648 -14248
rect 391308 -14390 391648 -14304
rect 391308 -14446 391376 -14390
rect 391432 -14446 391518 -14390
rect 391574 -14446 391648 -14390
rect 391308 -14532 391648 -14446
rect 391308 -14588 391376 -14532
rect 391432 -14588 391518 -14532
rect 391574 -14588 391648 -14532
rect 391308 -14674 391648 -14588
rect 391308 -14730 391376 -14674
rect 391432 -14730 391518 -14674
rect 391574 -14730 391648 -14674
rect 391308 -14816 391648 -14730
rect 391308 -14872 391376 -14816
rect 391432 -14872 391518 -14816
rect 391574 -14872 391648 -14816
rect 391308 -14958 391648 -14872
rect 391308 -15014 391376 -14958
rect 391432 -15014 391518 -14958
rect 391574 -15014 391648 -14958
rect 391308 -15100 391648 -15014
rect 391308 -15156 391376 -15100
rect 391432 -15156 391518 -15100
rect 391574 -15156 391648 -15100
rect 391308 -15242 391648 -15156
rect 391308 -15298 391376 -15242
rect 391432 -15298 391518 -15242
rect 391574 -15298 391648 -15242
rect 391308 -15384 391648 -15298
rect 391308 -15440 391376 -15384
rect 391432 -15440 391518 -15384
rect 391574 -15440 391648 -15384
rect 391308 -15526 391648 -15440
rect 391308 -15582 391376 -15526
rect 391432 -15582 391518 -15526
rect 391574 -15582 391648 -15526
rect 391308 -15668 391648 -15582
rect 391308 -15724 391376 -15668
rect 391432 -15724 391518 -15668
rect 391574 -15724 391648 -15668
rect 391308 -15810 391648 -15724
rect 391308 -15866 391376 -15810
rect 391432 -15866 391518 -15810
rect 391574 -15866 391648 -15810
rect 391308 -15952 391648 -15866
rect 391308 -16008 391376 -15952
rect 391432 -16008 391518 -15952
rect 391574 -16008 391648 -15952
rect 391308 -16094 391648 -16008
rect 391308 -16150 391376 -16094
rect 391432 -16150 391518 -16094
rect 391574 -16150 391648 -16094
rect 391308 -16236 391648 -16150
rect 391308 -16292 391376 -16236
rect 391432 -16292 391518 -16236
rect 391574 -16292 391648 -16236
rect 391308 -16378 391648 -16292
rect 391308 -16434 391376 -16378
rect 391432 -16434 391518 -16378
rect 391574 -16434 391648 -16378
rect 391308 -16520 391648 -16434
rect 391308 -16576 391376 -16520
rect 391432 -16576 391518 -16520
rect 391574 -16576 391648 -16520
rect 391308 -16662 391648 -16576
rect 391308 -16718 391376 -16662
rect 391432 -16718 391518 -16662
rect 391574 -16718 391648 -16662
rect 391308 -16804 391648 -16718
rect 391308 -16860 391376 -16804
rect 391432 -16860 391518 -16804
rect 391574 -16860 391648 -16804
rect 391308 -16946 391648 -16860
rect 391308 -17002 391376 -16946
rect 391432 -17002 391518 -16946
rect 391574 -17002 391648 -16946
rect 391308 -17088 391648 -17002
rect 391308 -17144 391376 -17088
rect 391432 -17144 391518 -17088
rect 391574 -17144 391648 -17088
rect 391308 -17230 391648 -17144
rect 391308 -17286 391376 -17230
rect 391432 -17286 391518 -17230
rect 391574 -17286 391648 -17230
rect 391308 -17372 391648 -17286
rect 391308 -17428 391376 -17372
rect 391432 -17428 391518 -17372
rect 391574 -17428 391648 -17372
rect 391308 -17514 391648 -17428
rect 391308 -17570 391376 -17514
rect 391432 -17570 391518 -17514
rect 391574 -17570 391648 -17514
rect 391308 -17656 391648 -17570
rect 391308 -17712 391376 -17656
rect 391432 -17712 391518 -17656
rect 391574 -17712 391648 -17656
rect 391308 -17798 391648 -17712
rect 391308 -17854 391376 -17798
rect 391432 -17854 391518 -17798
rect 391574 -17854 391648 -17798
rect 391308 -17940 391648 -17854
rect 391308 -17996 391376 -17940
rect 391432 -17996 391518 -17940
rect 391574 -17996 391648 -17940
rect 391308 -18082 391648 -17996
rect 391308 -18138 391376 -18082
rect 391432 -18138 391518 -18082
rect 391574 -18138 391648 -18082
rect 391308 -18224 391648 -18138
rect 391308 -18280 391376 -18224
rect 391432 -18280 391518 -18224
rect 391574 -18280 391648 -18224
rect 391308 -18366 391648 -18280
rect 391308 -18422 391376 -18366
rect 391432 -18422 391518 -18366
rect 391574 -18422 391648 -18366
rect 391308 -18508 391648 -18422
rect 391308 -18564 391376 -18508
rect 391432 -18564 391518 -18508
rect 391574 -18564 391648 -18508
rect 391308 -18650 391648 -18564
rect 391308 -18706 391376 -18650
rect 391432 -18706 391518 -18650
rect 391574 -18706 391648 -18650
rect 391308 -18792 391648 -18706
rect 391308 -18848 391376 -18792
rect 391432 -18848 391518 -18792
rect 391574 -18848 391648 -18792
rect 391308 -18934 391648 -18848
rect 391308 -18990 391376 -18934
rect 391432 -18990 391518 -18934
rect 391574 -18990 391648 -18934
rect 391308 -19076 391648 -18990
rect 391308 -19132 391376 -19076
rect 391432 -19132 391518 -19076
rect 391574 -19132 391648 -19076
rect 391308 -19218 391648 -19132
rect 391308 -19274 391376 -19218
rect 391432 -19274 391518 -19218
rect 391574 -19274 391648 -19218
rect 391308 -19360 391648 -19274
rect 391308 -19416 391376 -19360
rect 391432 -19416 391518 -19360
rect 391574 -19416 391648 -19360
rect 391308 -19502 391648 -19416
rect 391308 -19558 391376 -19502
rect 391432 -19558 391518 -19502
rect 391574 -19558 391648 -19502
rect 391308 -19644 391648 -19558
rect 391308 -19700 391376 -19644
rect 391432 -19700 391518 -19644
rect 391574 -19700 391648 -19644
rect 391308 -19786 391648 -19700
rect 391308 -19842 391376 -19786
rect 391432 -19842 391518 -19786
rect 391574 -19842 391648 -19786
rect 391308 -19928 391648 -19842
rect 391308 -19984 391376 -19928
rect 391432 -19984 391518 -19928
rect 391574 -19984 391648 -19928
rect 391308 -20070 391648 -19984
rect 391308 -20126 391376 -20070
rect 391432 -20126 391518 -20070
rect 391574 -20126 391648 -20070
rect 391308 -20212 391648 -20126
rect 391308 -20268 391376 -20212
rect 391432 -20268 391518 -20212
rect 391574 -20268 391648 -20212
rect 391308 -20354 391648 -20268
rect 391308 -20410 391376 -20354
rect 391432 -20410 391518 -20354
rect 391574 -20410 391648 -20354
rect 391308 -20496 391648 -20410
rect 391308 -20552 391376 -20496
rect 391432 -20552 391518 -20496
rect 391574 -20552 391648 -20496
rect 391308 -20638 391648 -20552
rect 391308 -20694 391376 -20638
rect 391432 -20694 391518 -20638
rect 391574 -20694 391648 -20638
rect 391308 -20780 391648 -20694
rect 391308 -20836 391376 -20780
rect 391432 -20836 391518 -20780
rect 391574 -20836 391648 -20780
rect 391308 -20922 391648 -20836
rect 391308 -20978 391376 -20922
rect 391432 -20978 391518 -20922
rect 391574 -20978 391648 -20922
rect 391308 -21064 391648 -20978
rect 391308 -21120 391376 -21064
rect 391432 -21120 391518 -21064
rect 391574 -21120 391648 -21064
rect 391308 -21206 391648 -21120
rect 391308 -21262 391376 -21206
rect 391432 -21262 391518 -21206
rect 391574 -21262 391648 -21206
rect 391308 -21348 391648 -21262
rect 391308 -21404 391376 -21348
rect 391432 -21404 391518 -21348
rect 391574 -21404 391648 -21348
rect 391308 -21490 391648 -21404
rect 391308 -21546 391376 -21490
rect 391432 -21546 391518 -21490
rect 391574 -21546 391648 -21490
rect 391308 -21632 391648 -21546
rect 391308 -21688 391376 -21632
rect 391432 -21688 391518 -21632
rect 391574 -21688 391648 -21632
rect 391308 -21774 391648 -21688
rect 391308 -21830 391376 -21774
rect 391432 -21830 391518 -21774
rect 391574 -21830 391648 -21774
rect 391308 -21916 391648 -21830
rect 391308 -21972 391376 -21916
rect 391432 -21972 391518 -21916
rect 391574 -21972 391648 -21916
rect 391308 -22058 391648 -21972
rect 391308 -22114 391376 -22058
rect 391432 -22114 391518 -22058
rect 391574 -22114 391648 -22058
rect 391308 -22200 391648 -22114
rect 391308 -22256 391376 -22200
rect 391432 -22256 391518 -22200
rect 391574 -22256 391648 -22200
rect 391308 -22342 391648 -22256
rect 391308 -22398 391376 -22342
rect 391432 -22398 391518 -22342
rect 391574 -22398 391648 -22342
rect 391308 -22484 391648 -22398
rect 391308 -22540 391376 -22484
rect 391432 -22540 391518 -22484
rect 391574 -22540 391648 -22484
rect 391308 -22626 391648 -22540
rect 391308 -22682 391376 -22626
rect 391432 -22682 391518 -22626
rect 391574 -22682 391648 -22626
rect 391308 -22768 391648 -22682
rect 391308 -22824 391376 -22768
rect 391432 -22824 391518 -22768
rect 391574 -22824 391648 -22768
rect 391308 -22910 391648 -22824
rect 391308 -22966 391376 -22910
rect 391432 -22966 391518 -22910
rect 391574 -22966 391648 -22910
rect 391308 -23052 391648 -22966
rect 391308 -23108 391376 -23052
rect 391432 -23108 391518 -23052
rect 391574 -23108 391648 -23052
rect 391308 -23194 391648 -23108
rect 391308 -23250 391376 -23194
rect 391432 -23250 391518 -23194
rect 391574 -23250 391648 -23194
rect 391308 -23336 391648 -23250
rect 391308 -23392 391376 -23336
rect 391432 -23392 391518 -23336
rect 391574 -23392 391648 -23336
rect 391308 -23478 391648 -23392
rect 391308 -23534 391376 -23478
rect 391432 -23534 391518 -23478
rect 391574 -23534 391648 -23478
rect 391308 -23620 391648 -23534
rect 391308 -23676 391376 -23620
rect 391432 -23676 391518 -23620
rect 391574 -23676 391648 -23620
rect 391308 -23762 391648 -23676
rect 391308 -23818 391376 -23762
rect 391432 -23818 391518 -23762
rect 391574 -23818 391648 -23762
rect 391308 -23904 391648 -23818
rect 391308 -23960 391376 -23904
rect 391432 -23960 391518 -23904
rect 391574 -23960 391648 -23904
rect 391308 -24046 391648 -23960
rect 391308 -24102 391376 -24046
rect 391432 -24102 391518 -24046
rect 391574 -24102 391648 -24046
rect 391308 -24188 391648 -24102
rect 391308 -24244 391376 -24188
rect 391432 -24244 391518 -24188
rect 391574 -24244 391648 -24188
rect 391308 -24330 391648 -24244
rect 391308 -24386 391376 -24330
rect 391432 -24386 391518 -24330
rect 391574 -24386 391648 -24330
rect 391308 -24472 391648 -24386
rect 391308 -24528 391376 -24472
rect 391432 -24528 391518 -24472
rect 391574 -24528 391648 -24472
rect 391308 -24614 391648 -24528
rect 391308 -24670 391376 -24614
rect 391432 -24670 391518 -24614
rect 391574 -24670 391648 -24614
rect 391308 -24756 391648 -24670
rect 391308 -24812 391376 -24756
rect 391432 -24812 391518 -24756
rect 391574 -24812 391648 -24756
rect 391308 -24898 391648 -24812
rect 391308 -24954 391376 -24898
rect 391432 -24954 391518 -24898
rect 391574 -24954 391648 -24898
rect 391308 -25040 391648 -24954
rect 391308 -25096 391376 -25040
rect 391432 -25096 391518 -25040
rect 391574 -25096 391648 -25040
rect 391308 -25182 391648 -25096
rect 391308 -25238 391376 -25182
rect 391432 -25238 391518 -25182
rect 391574 -25238 391648 -25182
rect 391308 -25324 391648 -25238
rect 391308 -25380 391376 -25324
rect 391432 -25380 391518 -25324
rect 391574 -25380 391648 -25324
rect 391308 -25466 391648 -25380
rect 391308 -25522 391376 -25466
rect 391432 -25522 391518 -25466
rect 391574 -25522 391648 -25466
rect 391308 -25532 391648 -25522
rect 391708 -13680 392048 -13670
rect 391708 -13736 391776 -13680
rect 391832 -13736 391918 -13680
rect 391974 -13736 392048 -13680
rect 391708 -13822 392048 -13736
rect 391708 -13878 391776 -13822
rect 391832 -13878 391918 -13822
rect 391974 -13878 392048 -13822
rect 391708 -13964 392048 -13878
rect 391708 -14020 391776 -13964
rect 391832 -14020 391918 -13964
rect 391974 -14020 392048 -13964
rect 391708 -14106 392048 -14020
rect 391708 -14162 391776 -14106
rect 391832 -14162 391918 -14106
rect 391974 -14162 392048 -14106
rect 391708 -14248 392048 -14162
rect 391708 -14304 391776 -14248
rect 391832 -14304 391918 -14248
rect 391974 -14304 392048 -14248
rect 391708 -14390 392048 -14304
rect 391708 -14446 391776 -14390
rect 391832 -14446 391918 -14390
rect 391974 -14446 392048 -14390
rect 391708 -14532 392048 -14446
rect 391708 -14588 391776 -14532
rect 391832 -14588 391918 -14532
rect 391974 -14588 392048 -14532
rect 391708 -14674 392048 -14588
rect 391708 -14730 391776 -14674
rect 391832 -14730 391918 -14674
rect 391974 -14730 392048 -14674
rect 391708 -14816 392048 -14730
rect 391708 -14872 391776 -14816
rect 391832 -14872 391918 -14816
rect 391974 -14872 392048 -14816
rect 391708 -14958 392048 -14872
rect 391708 -15014 391776 -14958
rect 391832 -15014 391918 -14958
rect 391974 -15014 392048 -14958
rect 391708 -15100 392048 -15014
rect 391708 -15156 391776 -15100
rect 391832 -15156 391918 -15100
rect 391974 -15156 392048 -15100
rect 391708 -15242 392048 -15156
rect 391708 -15298 391776 -15242
rect 391832 -15298 391918 -15242
rect 391974 -15298 392048 -15242
rect 391708 -15384 392048 -15298
rect 391708 -15440 391776 -15384
rect 391832 -15440 391918 -15384
rect 391974 -15440 392048 -15384
rect 391708 -15526 392048 -15440
rect 391708 -15582 391776 -15526
rect 391832 -15582 391918 -15526
rect 391974 -15582 392048 -15526
rect 391708 -15668 392048 -15582
rect 391708 -15724 391776 -15668
rect 391832 -15724 391918 -15668
rect 391974 -15724 392048 -15668
rect 391708 -15810 392048 -15724
rect 391708 -15866 391776 -15810
rect 391832 -15866 391918 -15810
rect 391974 -15866 392048 -15810
rect 391708 -15952 392048 -15866
rect 391708 -16008 391776 -15952
rect 391832 -16008 391918 -15952
rect 391974 -16008 392048 -15952
rect 391708 -16094 392048 -16008
rect 391708 -16150 391776 -16094
rect 391832 -16150 391918 -16094
rect 391974 -16150 392048 -16094
rect 391708 -16236 392048 -16150
rect 391708 -16292 391776 -16236
rect 391832 -16292 391918 -16236
rect 391974 -16292 392048 -16236
rect 391708 -16378 392048 -16292
rect 391708 -16434 391776 -16378
rect 391832 -16434 391918 -16378
rect 391974 -16434 392048 -16378
rect 391708 -16520 392048 -16434
rect 391708 -16576 391776 -16520
rect 391832 -16576 391918 -16520
rect 391974 -16576 392048 -16520
rect 391708 -16662 392048 -16576
rect 391708 -16718 391776 -16662
rect 391832 -16718 391918 -16662
rect 391974 -16718 392048 -16662
rect 391708 -16804 392048 -16718
rect 391708 -16860 391776 -16804
rect 391832 -16860 391918 -16804
rect 391974 -16860 392048 -16804
rect 391708 -16946 392048 -16860
rect 391708 -17002 391776 -16946
rect 391832 -17002 391918 -16946
rect 391974 -17002 392048 -16946
rect 391708 -17088 392048 -17002
rect 391708 -17144 391776 -17088
rect 391832 -17144 391918 -17088
rect 391974 -17144 392048 -17088
rect 391708 -17230 392048 -17144
rect 391708 -17286 391776 -17230
rect 391832 -17286 391918 -17230
rect 391974 -17286 392048 -17230
rect 391708 -17372 392048 -17286
rect 391708 -17428 391776 -17372
rect 391832 -17428 391918 -17372
rect 391974 -17428 392048 -17372
rect 391708 -17514 392048 -17428
rect 391708 -17570 391776 -17514
rect 391832 -17570 391918 -17514
rect 391974 -17570 392048 -17514
rect 391708 -17656 392048 -17570
rect 391708 -17712 391776 -17656
rect 391832 -17712 391918 -17656
rect 391974 -17712 392048 -17656
rect 391708 -17798 392048 -17712
rect 391708 -17854 391776 -17798
rect 391832 -17854 391918 -17798
rect 391974 -17854 392048 -17798
rect 391708 -17940 392048 -17854
rect 391708 -17996 391776 -17940
rect 391832 -17996 391918 -17940
rect 391974 -17996 392048 -17940
rect 391708 -18082 392048 -17996
rect 391708 -18138 391776 -18082
rect 391832 -18138 391918 -18082
rect 391974 -18138 392048 -18082
rect 391708 -18224 392048 -18138
rect 391708 -18280 391776 -18224
rect 391832 -18280 391918 -18224
rect 391974 -18280 392048 -18224
rect 391708 -18366 392048 -18280
rect 391708 -18422 391776 -18366
rect 391832 -18422 391918 -18366
rect 391974 -18422 392048 -18366
rect 391708 -18508 392048 -18422
rect 391708 -18564 391776 -18508
rect 391832 -18564 391918 -18508
rect 391974 -18564 392048 -18508
rect 391708 -18650 392048 -18564
rect 391708 -18706 391776 -18650
rect 391832 -18706 391918 -18650
rect 391974 -18706 392048 -18650
rect 391708 -18792 392048 -18706
rect 391708 -18848 391776 -18792
rect 391832 -18848 391918 -18792
rect 391974 -18848 392048 -18792
rect 391708 -18934 392048 -18848
rect 391708 -18990 391776 -18934
rect 391832 -18990 391918 -18934
rect 391974 -18990 392048 -18934
rect 391708 -19076 392048 -18990
rect 391708 -19132 391776 -19076
rect 391832 -19132 391918 -19076
rect 391974 -19132 392048 -19076
rect 391708 -19218 392048 -19132
rect 391708 -19274 391776 -19218
rect 391832 -19274 391918 -19218
rect 391974 -19274 392048 -19218
rect 391708 -19360 392048 -19274
rect 391708 -19416 391776 -19360
rect 391832 -19416 391918 -19360
rect 391974 -19416 392048 -19360
rect 391708 -19502 392048 -19416
rect 391708 -19558 391776 -19502
rect 391832 -19558 391918 -19502
rect 391974 -19558 392048 -19502
rect 391708 -19644 392048 -19558
rect 391708 -19700 391776 -19644
rect 391832 -19700 391918 -19644
rect 391974 -19700 392048 -19644
rect 391708 -19786 392048 -19700
rect 391708 -19842 391776 -19786
rect 391832 -19842 391918 -19786
rect 391974 -19842 392048 -19786
rect 391708 -19928 392048 -19842
rect 391708 -19984 391776 -19928
rect 391832 -19984 391918 -19928
rect 391974 -19984 392048 -19928
rect 391708 -20070 392048 -19984
rect 391708 -20126 391776 -20070
rect 391832 -20126 391918 -20070
rect 391974 -20126 392048 -20070
rect 391708 -20212 392048 -20126
rect 391708 -20268 391776 -20212
rect 391832 -20268 391918 -20212
rect 391974 -20268 392048 -20212
rect 391708 -20354 392048 -20268
rect 391708 -20410 391776 -20354
rect 391832 -20410 391918 -20354
rect 391974 -20410 392048 -20354
rect 391708 -20496 392048 -20410
rect 391708 -20552 391776 -20496
rect 391832 -20552 391918 -20496
rect 391974 -20552 392048 -20496
rect 391708 -20638 392048 -20552
rect 391708 -20694 391776 -20638
rect 391832 -20694 391918 -20638
rect 391974 -20694 392048 -20638
rect 391708 -20780 392048 -20694
rect 391708 -20836 391776 -20780
rect 391832 -20836 391918 -20780
rect 391974 -20836 392048 -20780
rect 391708 -20922 392048 -20836
rect 391708 -20978 391776 -20922
rect 391832 -20978 391918 -20922
rect 391974 -20978 392048 -20922
rect 391708 -21064 392048 -20978
rect 391708 -21120 391776 -21064
rect 391832 -21120 391918 -21064
rect 391974 -21120 392048 -21064
rect 391708 -21206 392048 -21120
rect 391708 -21262 391776 -21206
rect 391832 -21262 391918 -21206
rect 391974 -21262 392048 -21206
rect 391708 -21348 392048 -21262
rect 391708 -21404 391776 -21348
rect 391832 -21404 391918 -21348
rect 391974 -21404 392048 -21348
rect 391708 -21490 392048 -21404
rect 391708 -21546 391776 -21490
rect 391832 -21546 391918 -21490
rect 391974 -21546 392048 -21490
rect 391708 -21632 392048 -21546
rect 391708 -21688 391776 -21632
rect 391832 -21688 391918 -21632
rect 391974 -21688 392048 -21632
rect 391708 -21774 392048 -21688
rect 391708 -21830 391776 -21774
rect 391832 -21830 391918 -21774
rect 391974 -21830 392048 -21774
rect 391708 -21916 392048 -21830
rect 391708 -21972 391776 -21916
rect 391832 -21972 391918 -21916
rect 391974 -21972 392048 -21916
rect 391708 -22058 392048 -21972
rect 391708 -22114 391776 -22058
rect 391832 -22114 391918 -22058
rect 391974 -22114 392048 -22058
rect 391708 -22200 392048 -22114
rect 391708 -22256 391776 -22200
rect 391832 -22256 391918 -22200
rect 391974 -22256 392048 -22200
rect 391708 -22342 392048 -22256
rect 391708 -22398 391776 -22342
rect 391832 -22398 391918 -22342
rect 391974 -22398 392048 -22342
rect 391708 -22484 392048 -22398
rect 391708 -22540 391776 -22484
rect 391832 -22540 391918 -22484
rect 391974 -22540 392048 -22484
rect 391708 -22626 392048 -22540
rect 391708 -22682 391776 -22626
rect 391832 -22682 391918 -22626
rect 391974 -22682 392048 -22626
rect 391708 -22768 392048 -22682
rect 391708 -22824 391776 -22768
rect 391832 -22824 391918 -22768
rect 391974 -22824 392048 -22768
rect 391708 -22910 392048 -22824
rect 391708 -22966 391776 -22910
rect 391832 -22966 391918 -22910
rect 391974 -22966 392048 -22910
rect 391708 -23052 392048 -22966
rect 391708 -23108 391776 -23052
rect 391832 -23108 391918 -23052
rect 391974 -23108 392048 -23052
rect 391708 -23194 392048 -23108
rect 391708 -23250 391776 -23194
rect 391832 -23250 391918 -23194
rect 391974 -23250 392048 -23194
rect 391708 -23336 392048 -23250
rect 391708 -23392 391776 -23336
rect 391832 -23392 391918 -23336
rect 391974 -23392 392048 -23336
rect 391708 -23478 392048 -23392
rect 391708 -23534 391776 -23478
rect 391832 -23534 391918 -23478
rect 391974 -23534 392048 -23478
rect 391708 -23620 392048 -23534
rect 391708 -23676 391776 -23620
rect 391832 -23676 391918 -23620
rect 391974 -23676 392048 -23620
rect 391708 -23762 392048 -23676
rect 391708 -23818 391776 -23762
rect 391832 -23818 391918 -23762
rect 391974 -23818 392048 -23762
rect 391708 -23904 392048 -23818
rect 391708 -23960 391776 -23904
rect 391832 -23960 391918 -23904
rect 391974 -23960 392048 -23904
rect 391708 -24046 392048 -23960
rect 391708 -24102 391776 -24046
rect 391832 -24102 391918 -24046
rect 391974 -24102 392048 -24046
rect 391708 -24188 392048 -24102
rect 391708 -24244 391776 -24188
rect 391832 -24244 391918 -24188
rect 391974 -24244 392048 -24188
rect 391708 -24330 392048 -24244
rect 391708 -24386 391776 -24330
rect 391832 -24386 391918 -24330
rect 391974 -24386 392048 -24330
rect 391708 -24472 392048 -24386
rect 391708 -24528 391776 -24472
rect 391832 -24528 391918 -24472
rect 391974 -24528 392048 -24472
rect 391708 -24614 392048 -24528
rect 391708 -24670 391776 -24614
rect 391832 -24670 391918 -24614
rect 391974 -24670 392048 -24614
rect 391708 -24756 392048 -24670
rect 391708 -24812 391776 -24756
rect 391832 -24812 391918 -24756
rect 391974 -24812 392048 -24756
rect 391708 -24898 392048 -24812
rect 391708 -24954 391776 -24898
rect 391832 -24954 391918 -24898
rect 391974 -24954 392048 -24898
rect 391708 -25040 392048 -24954
rect 391708 -25096 391776 -25040
rect 391832 -25096 391918 -25040
rect 391974 -25096 392048 -25040
rect 391708 -25182 392048 -25096
rect 391708 -25238 391776 -25182
rect 391832 -25238 391918 -25182
rect 391974 -25238 392048 -25182
rect 391708 -25324 392048 -25238
rect 391708 -25380 391776 -25324
rect 391832 -25380 391918 -25324
rect 391974 -25380 392048 -25324
rect 391708 -25466 392048 -25380
rect 391708 -25522 391776 -25466
rect 391832 -25522 391918 -25466
rect 391974 -25522 392048 -25466
rect 391708 -25532 392048 -25522
rect 392108 -13680 392448 -13670
rect 392108 -13736 392173 -13680
rect 392229 -13736 392315 -13680
rect 392371 -13736 392448 -13680
rect 392108 -13822 392448 -13736
rect 392108 -13878 392173 -13822
rect 392229 -13878 392315 -13822
rect 392371 -13878 392448 -13822
rect 392108 -13964 392448 -13878
rect 392108 -14020 392173 -13964
rect 392229 -14020 392315 -13964
rect 392371 -14020 392448 -13964
rect 392108 -14106 392448 -14020
rect 392108 -14162 392173 -14106
rect 392229 -14162 392315 -14106
rect 392371 -14162 392448 -14106
rect 392108 -14248 392448 -14162
rect 392108 -14304 392173 -14248
rect 392229 -14304 392315 -14248
rect 392371 -14304 392448 -14248
rect 392108 -14390 392448 -14304
rect 392108 -14446 392173 -14390
rect 392229 -14446 392315 -14390
rect 392371 -14446 392448 -14390
rect 392108 -14532 392448 -14446
rect 392108 -14588 392173 -14532
rect 392229 -14588 392315 -14532
rect 392371 -14588 392448 -14532
rect 392108 -14674 392448 -14588
rect 392108 -14730 392173 -14674
rect 392229 -14730 392315 -14674
rect 392371 -14730 392448 -14674
rect 392108 -14816 392448 -14730
rect 392108 -14872 392173 -14816
rect 392229 -14872 392315 -14816
rect 392371 -14872 392448 -14816
rect 392108 -14958 392448 -14872
rect 392108 -15014 392173 -14958
rect 392229 -15014 392315 -14958
rect 392371 -15014 392448 -14958
rect 392108 -15100 392448 -15014
rect 392108 -15156 392173 -15100
rect 392229 -15156 392315 -15100
rect 392371 -15156 392448 -15100
rect 392108 -15242 392448 -15156
rect 392108 -15298 392173 -15242
rect 392229 -15298 392315 -15242
rect 392371 -15298 392448 -15242
rect 392108 -15384 392448 -15298
rect 392108 -15440 392173 -15384
rect 392229 -15440 392315 -15384
rect 392371 -15440 392448 -15384
rect 392108 -15526 392448 -15440
rect 392108 -15582 392173 -15526
rect 392229 -15582 392315 -15526
rect 392371 -15582 392448 -15526
rect 392108 -15668 392448 -15582
rect 392108 -15724 392173 -15668
rect 392229 -15724 392315 -15668
rect 392371 -15724 392448 -15668
rect 392108 -15810 392448 -15724
rect 392108 -15866 392173 -15810
rect 392229 -15866 392315 -15810
rect 392371 -15866 392448 -15810
rect 392108 -15952 392448 -15866
rect 392108 -16008 392173 -15952
rect 392229 -16008 392315 -15952
rect 392371 -16008 392448 -15952
rect 392108 -16094 392448 -16008
rect 392108 -16150 392173 -16094
rect 392229 -16150 392315 -16094
rect 392371 -16150 392448 -16094
rect 392108 -16236 392448 -16150
rect 392108 -16292 392173 -16236
rect 392229 -16292 392315 -16236
rect 392371 -16292 392448 -16236
rect 392108 -16378 392448 -16292
rect 392108 -16434 392173 -16378
rect 392229 -16434 392315 -16378
rect 392371 -16434 392448 -16378
rect 392108 -16520 392448 -16434
rect 392108 -16576 392173 -16520
rect 392229 -16576 392315 -16520
rect 392371 -16576 392448 -16520
rect 392108 -16662 392448 -16576
rect 392108 -16718 392173 -16662
rect 392229 -16718 392315 -16662
rect 392371 -16718 392448 -16662
rect 392108 -16804 392448 -16718
rect 392108 -16860 392173 -16804
rect 392229 -16860 392315 -16804
rect 392371 -16860 392448 -16804
rect 392108 -16946 392448 -16860
rect 392108 -17002 392173 -16946
rect 392229 -17002 392315 -16946
rect 392371 -17002 392448 -16946
rect 392108 -17088 392448 -17002
rect 392108 -17144 392173 -17088
rect 392229 -17144 392315 -17088
rect 392371 -17144 392448 -17088
rect 392108 -17230 392448 -17144
rect 392108 -17286 392173 -17230
rect 392229 -17286 392315 -17230
rect 392371 -17286 392448 -17230
rect 392108 -17372 392448 -17286
rect 392108 -17428 392173 -17372
rect 392229 -17428 392315 -17372
rect 392371 -17428 392448 -17372
rect 392108 -17514 392448 -17428
rect 392108 -17570 392173 -17514
rect 392229 -17570 392315 -17514
rect 392371 -17570 392448 -17514
rect 392108 -17656 392448 -17570
rect 392108 -17712 392173 -17656
rect 392229 -17712 392315 -17656
rect 392371 -17712 392448 -17656
rect 392108 -17798 392448 -17712
rect 392108 -17854 392173 -17798
rect 392229 -17854 392315 -17798
rect 392371 -17854 392448 -17798
rect 392108 -17940 392448 -17854
rect 392108 -17996 392173 -17940
rect 392229 -17996 392315 -17940
rect 392371 -17996 392448 -17940
rect 392108 -18082 392448 -17996
rect 392108 -18138 392173 -18082
rect 392229 -18138 392315 -18082
rect 392371 -18138 392448 -18082
rect 392108 -18224 392448 -18138
rect 392108 -18280 392173 -18224
rect 392229 -18280 392315 -18224
rect 392371 -18280 392448 -18224
rect 392108 -18366 392448 -18280
rect 392108 -18422 392173 -18366
rect 392229 -18422 392315 -18366
rect 392371 -18422 392448 -18366
rect 392108 -18508 392448 -18422
rect 392108 -18564 392173 -18508
rect 392229 -18564 392315 -18508
rect 392371 -18564 392448 -18508
rect 392108 -18650 392448 -18564
rect 392108 -18706 392173 -18650
rect 392229 -18706 392315 -18650
rect 392371 -18706 392448 -18650
rect 392108 -18792 392448 -18706
rect 392108 -18848 392173 -18792
rect 392229 -18848 392315 -18792
rect 392371 -18848 392448 -18792
rect 392108 -18934 392448 -18848
rect 392108 -18990 392173 -18934
rect 392229 -18990 392315 -18934
rect 392371 -18990 392448 -18934
rect 392108 -19076 392448 -18990
rect 392108 -19132 392173 -19076
rect 392229 -19132 392315 -19076
rect 392371 -19132 392448 -19076
rect 392108 -19218 392448 -19132
rect 392108 -19274 392173 -19218
rect 392229 -19274 392315 -19218
rect 392371 -19274 392448 -19218
rect 392108 -19360 392448 -19274
rect 392108 -19416 392173 -19360
rect 392229 -19416 392315 -19360
rect 392371 -19416 392448 -19360
rect 392108 -19502 392448 -19416
rect 392108 -19558 392173 -19502
rect 392229 -19558 392315 -19502
rect 392371 -19558 392448 -19502
rect 392108 -19644 392448 -19558
rect 392108 -19700 392173 -19644
rect 392229 -19700 392315 -19644
rect 392371 -19700 392448 -19644
rect 392108 -19786 392448 -19700
rect 392108 -19842 392173 -19786
rect 392229 -19842 392315 -19786
rect 392371 -19842 392448 -19786
rect 392108 -19928 392448 -19842
rect 392108 -19984 392173 -19928
rect 392229 -19984 392315 -19928
rect 392371 -19984 392448 -19928
rect 392108 -20070 392448 -19984
rect 392108 -20126 392173 -20070
rect 392229 -20126 392315 -20070
rect 392371 -20126 392448 -20070
rect 392108 -20212 392448 -20126
rect 392108 -20268 392173 -20212
rect 392229 -20268 392315 -20212
rect 392371 -20268 392448 -20212
rect 392108 -20354 392448 -20268
rect 392108 -20410 392173 -20354
rect 392229 -20410 392315 -20354
rect 392371 -20410 392448 -20354
rect 392108 -20496 392448 -20410
rect 392108 -20552 392173 -20496
rect 392229 -20552 392315 -20496
rect 392371 -20552 392448 -20496
rect 392108 -20638 392448 -20552
rect 392108 -20694 392173 -20638
rect 392229 -20694 392315 -20638
rect 392371 -20694 392448 -20638
rect 392108 -20780 392448 -20694
rect 392108 -20836 392173 -20780
rect 392229 -20836 392315 -20780
rect 392371 -20836 392448 -20780
rect 392108 -20922 392448 -20836
rect 392108 -20978 392173 -20922
rect 392229 -20978 392315 -20922
rect 392371 -20978 392448 -20922
rect 392108 -21064 392448 -20978
rect 392108 -21120 392173 -21064
rect 392229 -21120 392315 -21064
rect 392371 -21120 392448 -21064
rect 392108 -21206 392448 -21120
rect 392108 -21262 392173 -21206
rect 392229 -21262 392315 -21206
rect 392371 -21262 392448 -21206
rect 392108 -21348 392448 -21262
rect 392108 -21404 392173 -21348
rect 392229 -21404 392315 -21348
rect 392371 -21404 392448 -21348
rect 392108 -21490 392448 -21404
rect 392108 -21546 392173 -21490
rect 392229 -21546 392315 -21490
rect 392371 -21546 392448 -21490
rect 392108 -21632 392448 -21546
rect 392108 -21688 392173 -21632
rect 392229 -21688 392315 -21632
rect 392371 -21688 392448 -21632
rect 392108 -21774 392448 -21688
rect 392108 -21830 392173 -21774
rect 392229 -21830 392315 -21774
rect 392371 -21830 392448 -21774
rect 392108 -21916 392448 -21830
rect 392108 -21972 392173 -21916
rect 392229 -21972 392315 -21916
rect 392371 -21972 392448 -21916
rect 392108 -22058 392448 -21972
rect 392108 -22114 392173 -22058
rect 392229 -22114 392315 -22058
rect 392371 -22114 392448 -22058
rect 392108 -22200 392448 -22114
rect 392108 -22256 392173 -22200
rect 392229 -22256 392315 -22200
rect 392371 -22256 392448 -22200
rect 392108 -22342 392448 -22256
rect 392108 -22398 392173 -22342
rect 392229 -22398 392315 -22342
rect 392371 -22398 392448 -22342
rect 392108 -22484 392448 -22398
rect 392108 -22540 392173 -22484
rect 392229 -22540 392315 -22484
rect 392371 -22540 392448 -22484
rect 392108 -22626 392448 -22540
rect 392108 -22682 392173 -22626
rect 392229 -22682 392315 -22626
rect 392371 -22682 392448 -22626
rect 392108 -22768 392448 -22682
rect 392108 -22824 392173 -22768
rect 392229 -22824 392315 -22768
rect 392371 -22824 392448 -22768
rect 392108 -22910 392448 -22824
rect 392108 -22966 392173 -22910
rect 392229 -22966 392315 -22910
rect 392371 -22966 392448 -22910
rect 392108 -23052 392448 -22966
rect 392108 -23108 392173 -23052
rect 392229 -23108 392315 -23052
rect 392371 -23108 392448 -23052
rect 392108 -23194 392448 -23108
rect 392108 -23250 392173 -23194
rect 392229 -23250 392315 -23194
rect 392371 -23250 392448 -23194
rect 392108 -23336 392448 -23250
rect 392108 -23392 392173 -23336
rect 392229 -23392 392315 -23336
rect 392371 -23392 392448 -23336
rect 392108 -23478 392448 -23392
rect 392108 -23534 392173 -23478
rect 392229 -23534 392315 -23478
rect 392371 -23534 392448 -23478
rect 392108 -23620 392448 -23534
rect 392108 -23676 392173 -23620
rect 392229 -23676 392315 -23620
rect 392371 -23676 392448 -23620
rect 392108 -23762 392448 -23676
rect 392108 -23818 392173 -23762
rect 392229 -23818 392315 -23762
rect 392371 -23818 392448 -23762
rect 392108 -23904 392448 -23818
rect 392108 -23960 392173 -23904
rect 392229 -23960 392315 -23904
rect 392371 -23960 392448 -23904
rect 392108 -24046 392448 -23960
rect 392108 -24102 392173 -24046
rect 392229 -24102 392315 -24046
rect 392371 -24102 392448 -24046
rect 392108 -24188 392448 -24102
rect 392108 -24244 392173 -24188
rect 392229 -24244 392315 -24188
rect 392371 -24244 392448 -24188
rect 392108 -24330 392448 -24244
rect 392108 -24386 392173 -24330
rect 392229 -24386 392315 -24330
rect 392371 -24386 392448 -24330
rect 392108 -24472 392448 -24386
rect 392108 -24528 392173 -24472
rect 392229 -24528 392315 -24472
rect 392371 -24528 392448 -24472
rect 392108 -24614 392448 -24528
rect 392108 -24670 392173 -24614
rect 392229 -24670 392315 -24614
rect 392371 -24670 392448 -24614
rect 392108 -24756 392448 -24670
rect 392108 -24812 392173 -24756
rect 392229 -24812 392315 -24756
rect 392371 -24812 392448 -24756
rect 392108 -24898 392448 -24812
rect 392108 -24954 392173 -24898
rect 392229 -24954 392315 -24898
rect 392371 -24954 392448 -24898
rect 392108 -25040 392448 -24954
rect 392108 -25096 392173 -25040
rect 392229 -25096 392315 -25040
rect 392371 -25096 392448 -25040
rect 392108 -25182 392448 -25096
rect 392108 -25238 392173 -25182
rect 392229 -25238 392315 -25182
rect 392371 -25238 392448 -25182
rect 392108 -25324 392448 -25238
rect 392108 -25380 392173 -25324
rect 392229 -25380 392315 -25324
rect 392371 -25380 392448 -25324
rect 392108 -25466 392448 -25380
rect 392108 -25522 392173 -25466
rect 392229 -25522 392315 -25466
rect 392371 -25522 392448 -25466
rect 392108 -25532 392448 -25522
rect 392508 -13680 392848 -13670
rect 392508 -13736 392578 -13680
rect 392634 -13736 392720 -13680
rect 392776 -13736 392848 -13680
rect 392508 -13822 392848 -13736
rect 392508 -13878 392578 -13822
rect 392634 -13878 392720 -13822
rect 392776 -13878 392848 -13822
rect 392508 -13964 392848 -13878
rect 392508 -14020 392578 -13964
rect 392634 -14020 392720 -13964
rect 392776 -14020 392848 -13964
rect 392508 -14106 392848 -14020
rect 392508 -14162 392578 -14106
rect 392634 -14162 392720 -14106
rect 392776 -14162 392848 -14106
rect 392508 -14248 392848 -14162
rect 392508 -14304 392578 -14248
rect 392634 -14304 392720 -14248
rect 392776 -14304 392848 -14248
rect 392508 -14390 392848 -14304
rect 392508 -14446 392578 -14390
rect 392634 -14446 392720 -14390
rect 392776 -14446 392848 -14390
rect 392508 -14532 392848 -14446
rect 392508 -14588 392578 -14532
rect 392634 -14588 392720 -14532
rect 392776 -14588 392848 -14532
rect 392508 -14674 392848 -14588
rect 392508 -14730 392578 -14674
rect 392634 -14730 392720 -14674
rect 392776 -14730 392848 -14674
rect 392508 -14816 392848 -14730
rect 392508 -14872 392578 -14816
rect 392634 -14872 392720 -14816
rect 392776 -14872 392848 -14816
rect 392508 -14958 392848 -14872
rect 392508 -15014 392578 -14958
rect 392634 -15014 392720 -14958
rect 392776 -15014 392848 -14958
rect 392508 -15100 392848 -15014
rect 392508 -15156 392578 -15100
rect 392634 -15156 392720 -15100
rect 392776 -15156 392848 -15100
rect 392508 -15242 392848 -15156
rect 392508 -15298 392578 -15242
rect 392634 -15298 392720 -15242
rect 392776 -15298 392848 -15242
rect 392508 -15384 392848 -15298
rect 392508 -15440 392578 -15384
rect 392634 -15440 392720 -15384
rect 392776 -15440 392848 -15384
rect 392508 -15526 392848 -15440
rect 392508 -15582 392578 -15526
rect 392634 -15582 392720 -15526
rect 392776 -15582 392848 -15526
rect 392508 -15668 392848 -15582
rect 392508 -15724 392578 -15668
rect 392634 -15724 392720 -15668
rect 392776 -15724 392848 -15668
rect 392508 -15810 392848 -15724
rect 392508 -15866 392578 -15810
rect 392634 -15866 392720 -15810
rect 392776 -15866 392848 -15810
rect 392508 -15952 392848 -15866
rect 392508 -16008 392578 -15952
rect 392634 -16008 392720 -15952
rect 392776 -16008 392848 -15952
rect 392508 -16094 392848 -16008
rect 392508 -16150 392578 -16094
rect 392634 -16150 392720 -16094
rect 392776 -16150 392848 -16094
rect 392508 -16236 392848 -16150
rect 392508 -16292 392578 -16236
rect 392634 -16292 392720 -16236
rect 392776 -16292 392848 -16236
rect 392508 -16378 392848 -16292
rect 392508 -16434 392578 -16378
rect 392634 -16434 392720 -16378
rect 392776 -16434 392848 -16378
rect 392508 -16520 392848 -16434
rect 392508 -16576 392578 -16520
rect 392634 -16576 392720 -16520
rect 392776 -16576 392848 -16520
rect 392508 -16662 392848 -16576
rect 392508 -16718 392578 -16662
rect 392634 -16718 392720 -16662
rect 392776 -16718 392848 -16662
rect 392508 -16804 392848 -16718
rect 392508 -16860 392578 -16804
rect 392634 -16860 392720 -16804
rect 392776 -16860 392848 -16804
rect 392508 -16946 392848 -16860
rect 392508 -17002 392578 -16946
rect 392634 -17002 392720 -16946
rect 392776 -17002 392848 -16946
rect 392508 -17088 392848 -17002
rect 392508 -17144 392578 -17088
rect 392634 -17144 392720 -17088
rect 392776 -17144 392848 -17088
rect 392508 -17230 392848 -17144
rect 392508 -17286 392578 -17230
rect 392634 -17286 392720 -17230
rect 392776 -17286 392848 -17230
rect 392508 -17372 392848 -17286
rect 392508 -17428 392578 -17372
rect 392634 -17428 392720 -17372
rect 392776 -17428 392848 -17372
rect 392508 -17514 392848 -17428
rect 392508 -17570 392578 -17514
rect 392634 -17570 392720 -17514
rect 392776 -17570 392848 -17514
rect 392508 -17656 392848 -17570
rect 392508 -17712 392578 -17656
rect 392634 -17712 392720 -17656
rect 392776 -17712 392848 -17656
rect 392508 -17798 392848 -17712
rect 392508 -17854 392578 -17798
rect 392634 -17854 392720 -17798
rect 392776 -17854 392848 -17798
rect 392508 -17940 392848 -17854
rect 392508 -17996 392578 -17940
rect 392634 -17996 392720 -17940
rect 392776 -17996 392848 -17940
rect 392508 -18082 392848 -17996
rect 392508 -18138 392578 -18082
rect 392634 -18138 392720 -18082
rect 392776 -18138 392848 -18082
rect 392508 -18224 392848 -18138
rect 392508 -18280 392578 -18224
rect 392634 -18280 392720 -18224
rect 392776 -18280 392848 -18224
rect 392508 -18366 392848 -18280
rect 392508 -18422 392578 -18366
rect 392634 -18422 392720 -18366
rect 392776 -18422 392848 -18366
rect 392508 -18508 392848 -18422
rect 392508 -18564 392578 -18508
rect 392634 -18564 392720 -18508
rect 392776 -18564 392848 -18508
rect 392508 -18650 392848 -18564
rect 392508 -18706 392578 -18650
rect 392634 -18706 392720 -18650
rect 392776 -18706 392848 -18650
rect 392508 -18792 392848 -18706
rect 392508 -18848 392578 -18792
rect 392634 -18848 392720 -18792
rect 392776 -18848 392848 -18792
rect 392508 -18934 392848 -18848
rect 392508 -18990 392578 -18934
rect 392634 -18990 392720 -18934
rect 392776 -18990 392848 -18934
rect 392508 -19076 392848 -18990
rect 392508 -19132 392578 -19076
rect 392634 -19132 392720 -19076
rect 392776 -19132 392848 -19076
rect 392508 -19218 392848 -19132
rect 392508 -19274 392578 -19218
rect 392634 -19274 392720 -19218
rect 392776 -19274 392848 -19218
rect 392508 -19360 392848 -19274
rect 392508 -19416 392578 -19360
rect 392634 -19416 392720 -19360
rect 392776 -19416 392848 -19360
rect 392508 -19502 392848 -19416
rect 392508 -19558 392578 -19502
rect 392634 -19558 392720 -19502
rect 392776 -19558 392848 -19502
rect 392508 -19644 392848 -19558
rect 392508 -19700 392578 -19644
rect 392634 -19700 392720 -19644
rect 392776 -19700 392848 -19644
rect 392508 -19786 392848 -19700
rect 392508 -19842 392578 -19786
rect 392634 -19842 392720 -19786
rect 392776 -19842 392848 -19786
rect 392508 -19928 392848 -19842
rect 392508 -19984 392578 -19928
rect 392634 -19984 392720 -19928
rect 392776 -19984 392848 -19928
rect 392508 -20070 392848 -19984
rect 392508 -20126 392578 -20070
rect 392634 -20126 392720 -20070
rect 392776 -20126 392848 -20070
rect 392508 -20212 392848 -20126
rect 392508 -20268 392578 -20212
rect 392634 -20268 392720 -20212
rect 392776 -20268 392848 -20212
rect 392508 -20354 392848 -20268
rect 392508 -20410 392578 -20354
rect 392634 -20410 392720 -20354
rect 392776 -20410 392848 -20354
rect 392508 -20496 392848 -20410
rect 392508 -20552 392578 -20496
rect 392634 -20552 392720 -20496
rect 392776 -20552 392848 -20496
rect 392508 -20638 392848 -20552
rect 392508 -20694 392578 -20638
rect 392634 -20694 392720 -20638
rect 392776 -20694 392848 -20638
rect 392508 -20780 392848 -20694
rect 392508 -20836 392578 -20780
rect 392634 -20836 392720 -20780
rect 392776 -20836 392848 -20780
rect 392508 -20922 392848 -20836
rect 392508 -20978 392578 -20922
rect 392634 -20978 392720 -20922
rect 392776 -20978 392848 -20922
rect 392508 -21064 392848 -20978
rect 392508 -21120 392578 -21064
rect 392634 -21120 392720 -21064
rect 392776 -21120 392848 -21064
rect 392508 -21206 392848 -21120
rect 392508 -21262 392578 -21206
rect 392634 -21262 392720 -21206
rect 392776 -21262 392848 -21206
rect 392508 -21348 392848 -21262
rect 392508 -21404 392578 -21348
rect 392634 -21404 392720 -21348
rect 392776 -21404 392848 -21348
rect 392508 -21490 392848 -21404
rect 392508 -21546 392578 -21490
rect 392634 -21546 392720 -21490
rect 392776 -21546 392848 -21490
rect 392508 -21632 392848 -21546
rect 392508 -21688 392578 -21632
rect 392634 -21688 392720 -21632
rect 392776 -21688 392848 -21632
rect 392508 -21774 392848 -21688
rect 392508 -21830 392578 -21774
rect 392634 -21830 392720 -21774
rect 392776 -21830 392848 -21774
rect 392508 -21916 392848 -21830
rect 392508 -21972 392578 -21916
rect 392634 -21972 392720 -21916
rect 392776 -21972 392848 -21916
rect 392508 -22058 392848 -21972
rect 392508 -22114 392578 -22058
rect 392634 -22114 392720 -22058
rect 392776 -22114 392848 -22058
rect 392508 -22200 392848 -22114
rect 392508 -22256 392578 -22200
rect 392634 -22256 392720 -22200
rect 392776 -22256 392848 -22200
rect 392508 -22342 392848 -22256
rect 392508 -22398 392578 -22342
rect 392634 -22398 392720 -22342
rect 392776 -22398 392848 -22342
rect 392508 -22484 392848 -22398
rect 392508 -22540 392578 -22484
rect 392634 -22540 392720 -22484
rect 392776 -22540 392848 -22484
rect 392508 -22626 392848 -22540
rect 392508 -22682 392578 -22626
rect 392634 -22682 392720 -22626
rect 392776 -22682 392848 -22626
rect 392508 -22768 392848 -22682
rect 392508 -22824 392578 -22768
rect 392634 -22824 392720 -22768
rect 392776 -22824 392848 -22768
rect 392508 -22910 392848 -22824
rect 392508 -22966 392578 -22910
rect 392634 -22966 392720 -22910
rect 392776 -22966 392848 -22910
rect 392508 -23052 392848 -22966
rect 392508 -23108 392578 -23052
rect 392634 -23108 392720 -23052
rect 392776 -23108 392848 -23052
rect 392508 -23194 392848 -23108
rect 392508 -23250 392578 -23194
rect 392634 -23250 392720 -23194
rect 392776 -23250 392848 -23194
rect 392508 -23336 392848 -23250
rect 392508 -23392 392578 -23336
rect 392634 -23392 392720 -23336
rect 392776 -23392 392848 -23336
rect 392508 -23478 392848 -23392
rect 392508 -23534 392578 -23478
rect 392634 -23534 392720 -23478
rect 392776 -23534 392848 -23478
rect 392508 -23620 392848 -23534
rect 392508 -23676 392578 -23620
rect 392634 -23676 392720 -23620
rect 392776 -23676 392848 -23620
rect 392508 -23762 392848 -23676
rect 392508 -23818 392578 -23762
rect 392634 -23818 392720 -23762
rect 392776 -23818 392848 -23762
rect 392508 -23904 392848 -23818
rect 392508 -23960 392578 -23904
rect 392634 -23960 392720 -23904
rect 392776 -23960 392848 -23904
rect 392508 -24046 392848 -23960
rect 392508 -24102 392578 -24046
rect 392634 -24102 392720 -24046
rect 392776 -24102 392848 -24046
rect 392508 -24188 392848 -24102
rect 392508 -24244 392578 -24188
rect 392634 -24244 392720 -24188
rect 392776 -24244 392848 -24188
rect 392508 -24330 392848 -24244
rect 392508 -24386 392578 -24330
rect 392634 -24386 392720 -24330
rect 392776 -24386 392848 -24330
rect 392508 -24472 392848 -24386
rect 392508 -24528 392578 -24472
rect 392634 -24528 392720 -24472
rect 392776 -24528 392848 -24472
rect 392508 -24614 392848 -24528
rect 392508 -24670 392578 -24614
rect 392634 -24670 392720 -24614
rect 392776 -24670 392848 -24614
rect 392508 -24756 392848 -24670
rect 392508 -24812 392578 -24756
rect 392634 -24812 392720 -24756
rect 392776 -24812 392848 -24756
rect 392508 -24898 392848 -24812
rect 392508 -24954 392578 -24898
rect 392634 -24954 392720 -24898
rect 392776 -24954 392848 -24898
rect 392508 -25040 392848 -24954
rect 392508 -25096 392578 -25040
rect 392634 -25096 392720 -25040
rect 392776 -25096 392848 -25040
rect 392508 -25182 392848 -25096
rect 392508 -25238 392578 -25182
rect 392634 -25238 392720 -25182
rect 392776 -25238 392848 -25182
rect 392508 -25324 392848 -25238
rect 392508 -25380 392578 -25324
rect 392634 -25380 392720 -25324
rect 392776 -25380 392848 -25324
rect 392508 -25466 392848 -25380
rect 392508 -25522 392578 -25466
rect 392634 -25522 392720 -25466
rect 392776 -25522 392848 -25466
rect 392508 -25532 392848 -25522
rect 392908 -13680 393248 -13670
rect 392908 -13736 392978 -13680
rect 393034 -13736 393120 -13680
rect 393176 -13736 393248 -13680
rect 392908 -13822 393248 -13736
rect 392908 -13878 392978 -13822
rect 393034 -13878 393120 -13822
rect 393176 -13878 393248 -13822
rect 392908 -13964 393248 -13878
rect 392908 -14020 392978 -13964
rect 393034 -14020 393120 -13964
rect 393176 -14020 393248 -13964
rect 392908 -14106 393248 -14020
rect 392908 -14162 392978 -14106
rect 393034 -14162 393120 -14106
rect 393176 -14162 393248 -14106
rect 392908 -14248 393248 -14162
rect 392908 -14304 392978 -14248
rect 393034 -14304 393120 -14248
rect 393176 -14304 393248 -14248
rect 392908 -14390 393248 -14304
rect 392908 -14446 392978 -14390
rect 393034 -14446 393120 -14390
rect 393176 -14446 393248 -14390
rect 392908 -14532 393248 -14446
rect 392908 -14588 392978 -14532
rect 393034 -14588 393120 -14532
rect 393176 -14588 393248 -14532
rect 392908 -14674 393248 -14588
rect 392908 -14730 392978 -14674
rect 393034 -14730 393120 -14674
rect 393176 -14730 393248 -14674
rect 392908 -14816 393248 -14730
rect 392908 -14872 392978 -14816
rect 393034 -14872 393120 -14816
rect 393176 -14872 393248 -14816
rect 392908 -14958 393248 -14872
rect 392908 -15014 392978 -14958
rect 393034 -15014 393120 -14958
rect 393176 -15014 393248 -14958
rect 392908 -15100 393248 -15014
rect 392908 -15156 392978 -15100
rect 393034 -15156 393120 -15100
rect 393176 -15156 393248 -15100
rect 392908 -15242 393248 -15156
rect 392908 -15298 392978 -15242
rect 393034 -15298 393120 -15242
rect 393176 -15298 393248 -15242
rect 392908 -15384 393248 -15298
rect 392908 -15440 392978 -15384
rect 393034 -15440 393120 -15384
rect 393176 -15440 393248 -15384
rect 392908 -15526 393248 -15440
rect 392908 -15582 392978 -15526
rect 393034 -15582 393120 -15526
rect 393176 -15582 393248 -15526
rect 392908 -15668 393248 -15582
rect 392908 -15724 392978 -15668
rect 393034 -15724 393120 -15668
rect 393176 -15724 393248 -15668
rect 392908 -15810 393248 -15724
rect 392908 -15866 392978 -15810
rect 393034 -15866 393120 -15810
rect 393176 -15866 393248 -15810
rect 392908 -15952 393248 -15866
rect 392908 -16008 392978 -15952
rect 393034 -16008 393120 -15952
rect 393176 -16008 393248 -15952
rect 392908 -16094 393248 -16008
rect 392908 -16150 392978 -16094
rect 393034 -16150 393120 -16094
rect 393176 -16150 393248 -16094
rect 392908 -16236 393248 -16150
rect 392908 -16292 392978 -16236
rect 393034 -16292 393120 -16236
rect 393176 -16292 393248 -16236
rect 392908 -16378 393248 -16292
rect 392908 -16434 392978 -16378
rect 393034 -16434 393120 -16378
rect 393176 -16434 393248 -16378
rect 392908 -16520 393248 -16434
rect 392908 -16576 392978 -16520
rect 393034 -16576 393120 -16520
rect 393176 -16576 393248 -16520
rect 392908 -16662 393248 -16576
rect 392908 -16718 392978 -16662
rect 393034 -16718 393120 -16662
rect 393176 -16718 393248 -16662
rect 392908 -16804 393248 -16718
rect 392908 -16860 392978 -16804
rect 393034 -16860 393120 -16804
rect 393176 -16860 393248 -16804
rect 392908 -16946 393248 -16860
rect 392908 -17002 392978 -16946
rect 393034 -17002 393120 -16946
rect 393176 -17002 393248 -16946
rect 392908 -17088 393248 -17002
rect 392908 -17144 392978 -17088
rect 393034 -17144 393120 -17088
rect 393176 -17144 393248 -17088
rect 392908 -17230 393248 -17144
rect 392908 -17286 392978 -17230
rect 393034 -17286 393120 -17230
rect 393176 -17286 393248 -17230
rect 392908 -17372 393248 -17286
rect 392908 -17428 392978 -17372
rect 393034 -17428 393120 -17372
rect 393176 -17428 393248 -17372
rect 392908 -17514 393248 -17428
rect 392908 -17570 392978 -17514
rect 393034 -17570 393120 -17514
rect 393176 -17570 393248 -17514
rect 392908 -17656 393248 -17570
rect 392908 -17712 392978 -17656
rect 393034 -17712 393120 -17656
rect 393176 -17712 393248 -17656
rect 392908 -17798 393248 -17712
rect 392908 -17854 392978 -17798
rect 393034 -17854 393120 -17798
rect 393176 -17854 393248 -17798
rect 392908 -17940 393248 -17854
rect 392908 -17996 392978 -17940
rect 393034 -17996 393120 -17940
rect 393176 -17996 393248 -17940
rect 392908 -18082 393248 -17996
rect 392908 -18138 392978 -18082
rect 393034 -18138 393120 -18082
rect 393176 -18138 393248 -18082
rect 392908 -18224 393248 -18138
rect 392908 -18280 392978 -18224
rect 393034 -18280 393120 -18224
rect 393176 -18280 393248 -18224
rect 392908 -18366 393248 -18280
rect 392908 -18422 392978 -18366
rect 393034 -18422 393120 -18366
rect 393176 -18422 393248 -18366
rect 392908 -18508 393248 -18422
rect 392908 -18564 392978 -18508
rect 393034 -18564 393120 -18508
rect 393176 -18564 393248 -18508
rect 392908 -18650 393248 -18564
rect 392908 -18706 392978 -18650
rect 393034 -18706 393120 -18650
rect 393176 -18706 393248 -18650
rect 392908 -18792 393248 -18706
rect 392908 -18848 392978 -18792
rect 393034 -18848 393120 -18792
rect 393176 -18848 393248 -18792
rect 392908 -18934 393248 -18848
rect 392908 -18990 392978 -18934
rect 393034 -18990 393120 -18934
rect 393176 -18990 393248 -18934
rect 392908 -19076 393248 -18990
rect 392908 -19132 392978 -19076
rect 393034 -19132 393120 -19076
rect 393176 -19132 393248 -19076
rect 392908 -19218 393248 -19132
rect 392908 -19274 392978 -19218
rect 393034 -19274 393120 -19218
rect 393176 -19274 393248 -19218
rect 392908 -19360 393248 -19274
rect 392908 -19416 392978 -19360
rect 393034 -19416 393120 -19360
rect 393176 -19416 393248 -19360
rect 392908 -19502 393248 -19416
rect 392908 -19558 392978 -19502
rect 393034 -19558 393120 -19502
rect 393176 -19558 393248 -19502
rect 392908 -19644 393248 -19558
rect 392908 -19700 392978 -19644
rect 393034 -19700 393120 -19644
rect 393176 -19700 393248 -19644
rect 392908 -19786 393248 -19700
rect 392908 -19842 392978 -19786
rect 393034 -19842 393120 -19786
rect 393176 -19842 393248 -19786
rect 392908 -19928 393248 -19842
rect 392908 -19984 392978 -19928
rect 393034 -19984 393120 -19928
rect 393176 -19984 393248 -19928
rect 392908 -20070 393248 -19984
rect 392908 -20126 392978 -20070
rect 393034 -20126 393120 -20070
rect 393176 -20126 393248 -20070
rect 392908 -20212 393248 -20126
rect 392908 -20268 392978 -20212
rect 393034 -20268 393120 -20212
rect 393176 -20268 393248 -20212
rect 392908 -20354 393248 -20268
rect 392908 -20410 392978 -20354
rect 393034 -20410 393120 -20354
rect 393176 -20410 393248 -20354
rect 392908 -20496 393248 -20410
rect 392908 -20552 392978 -20496
rect 393034 -20552 393120 -20496
rect 393176 -20552 393248 -20496
rect 392908 -20638 393248 -20552
rect 392908 -20694 392978 -20638
rect 393034 -20694 393120 -20638
rect 393176 -20694 393248 -20638
rect 392908 -20780 393248 -20694
rect 392908 -20836 392978 -20780
rect 393034 -20836 393120 -20780
rect 393176 -20836 393248 -20780
rect 392908 -20922 393248 -20836
rect 392908 -20978 392978 -20922
rect 393034 -20978 393120 -20922
rect 393176 -20978 393248 -20922
rect 392908 -21064 393248 -20978
rect 392908 -21120 392978 -21064
rect 393034 -21120 393120 -21064
rect 393176 -21120 393248 -21064
rect 392908 -21206 393248 -21120
rect 392908 -21262 392978 -21206
rect 393034 -21262 393120 -21206
rect 393176 -21262 393248 -21206
rect 392908 -21348 393248 -21262
rect 392908 -21404 392978 -21348
rect 393034 -21404 393120 -21348
rect 393176 -21404 393248 -21348
rect 392908 -21490 393248 -21404
rect 392908 -21546 392978 -21490
rect 393034 -21546 393120 -21490
rect 393176 -21546 393248 -21490
rect 392908 -21632 393248 -21546
rect 392908 -21688 392978 -21632
rect 393034 -21688 393120 -21632
rect 393176 -21688 393248 -21632
rect 392908 -21774 393248 -21688
rect 392908 -21830 392978 -21774
rect 393034 -21830 393120 -21774
rect 393176 -21830 393248 -21774
rect 392908 -21916 393248 -21830
rect 392908 -21972 392978 -21916
rect 393034 -21972 393120 -21916
rect 393176 -21972 393248 -21916
rect 392908 -22058 393248 -21972
rect 392908 -22114 392978 -22058
rect 393034 -22114 393120 -22058
rect 393176 -22114 393248 -22058
rect 392908 -22200 393248 -22114
rect 392908 -22256 392978 -22200
rect 393034 -22256 393120 -22200
rect 393176 -22256 393248 -22200
rect 392908 -22342 393248 -22256
rect 392908 -22398 392978 -22342
rect 393034 -22398 393120 -22342
rect 393176 -22398 393248 -22342
rect 392908 -22484 393248 -22398
rect 392908 -22540 392978 -22484
rect 393034 -22540 393120 -22484
rect 393176 -22540 393248 -22484
rect 392908 -22626 393248 -22540
rect 392908 -22682 392978 -22626
rect 393034 -22682 393120 -22626
rect 393176 -22682 393248 -22626
rect 392908 -22768 393248 -22682
rect 392908 -22824 392978 -22768
rect 393034 -22824 393120 -22768
rect 393176 -22824 393248 -22768
rect 392908 -22910 393248 -22824
rect 392908 -22966 392978 -22910
rect 393034 -22966 393120 -22910
rect 393176 -22966 393248 -22910
rect 392908 -23052 393248 -22966
rect 392908 -23108 392978 -23052
rect 393034 -23108 393120 -23052
rect 393176 -23108 393248 -23052
rect 392908 -23194 393248 -23108
rect 392908 -23250 392978 -23194
rect 393034 -23250 393120 -23194
rect 393176 -23250 393248 -23194
rect 392908 -23336 393248 -23250
rect 392908 -23392 392978 -23336
rect 393034 -23392 393120 -23336
rect 393176 -23392 393248 -23336
rect 392908 -23478 393248 -23392
rect 392908 -23534 392978 -23478
rect 393034 -23534 393120 -23478
rect 393176 -23534 393248 -23478
rect 392908 -23620 393248 -23534
rect 392908 -23676 392978 -23620
rect 393034 -23676 393120 -23620
rect 393176 -23676 393248 -23620
rect 392908 -23762 393248 -23676
rect 392908 -23818 392978 -23762
rect 393034 -23818 393120 -23762
rect 393176 -23818 393248 -23762
rect 392908 -23904 393248 -23818
rect 392908 -23960 392978 -23904
rect 393034 -23960 393120 -23904
rect 393176 -23960 393248 -23904
rect 392908 -24046 393248 -23960
rect 392908 -24102 392978 -24046
rect 393034 -24102 393120 -24046
rect 393176 -24102 393248 -24046
rect 392908 -24188 393248 -24102
rect 392908 -24244 392978 -24188
rect 393034 -24244 393120 -24188
rect 393176 -24244 393248 -24188
rect 392908 -24330 393248 -24244
rect 392908 -24386 392978 -24330
rect 393034 -24386 393120 -24330
rect 393176 -24386 393248 -24330
rect 392908 -24472 393248 -24386
rect 392908 -24528 392978 -24472
rect 393034 -24528 393120 -24472
rect 393176 -24528 393248 -24472
rect 392908 -24614 393248 -24528
rect 392908 -24670 392978 -24614
rect 393034 -24670 393120 -24614
rect 393176 -24670 393248 -24614
rect 392908 -24756 393248 -24670
rect 392908 -24812 392978 -24756
rect 393034 -24812 393120 -24756
rect 393176 -24812 393248 -24756
rect 392908 -24898 393248 -24812
rect 392908 -24954 392978 -24898
rect 393034 -24954 393120 -24898
rect 393176 -24954 393248 -24898
rect 392908 -25040 393248 -24954
rect 392908 -25096 392978 -25040
rect 393034 -25096 393120 -25040
rect 393176 -25096 393248 -25040
rect 392908 -25182 393248 -25096
rect 392908 -25238 392978 -25182
rect 393034 -25238 393120 -25182
rect 393176 -25238 393248 -25182
rect 392908 -25324 393248 -25238
rect 392908 -25380 392978 -25324
rect 393034 -25380 393120 -25324
rect 393176 -25380 393248 -25324
rect 392908 -25466 393248 -25380
rect 392908 -25522 392978 -25466
rect 393034 -25522 393120 -25466
rect 393176 -25522 393248 -25466
rect 392908 -25532 393248 -25522
rect 393308 -13680 393648 -13670
rect 393308 -13736 393383 -13680
rect 393439 -13736 393525 -13680
rect 393581 -13736 393648 -13680
rect 393308 -13822 393648 -13736
rect 393308 -13878 393383 -13822
rect 393439 -13878 393525 -13822
rect 393581 -13878 393648 -13822
rect 393308 -13964 393648 -13878
rect 393308 -14020 393383 -13964
rect 393439 -14020 393525 -13964
rect 393581 -14020 393648 -13964
rect 393308 -14106 393648 -14020
rect 393308 -14162 393383 -14106
rect 393439 -14162 393525 -14106
rect 393581 -14162 393648 -14106
rect 393308 -14248 393648 -14162
rect 393308 -14304 393383 -14248
rect 393439 -14304 393525 -14248
rect 393581 -14304 393648 -14248
rect 393308 -14390 393648 -14304
rect 393308 -14446 393383 -14390
rect 393439 -14446 393525 -14390
rect 393581 -14446 393648 -14390
rect 393308 -14532 393648 -14446
rect 393308 -14588 393383 -14532
rect 393439 -14588 393525 -14532
rect 393581 -14588 393648 -14532
rect 393308 -14674 393648 -14588
rect 393308 -14730 393383 -14674
rect 393439 -14730 393525 -14674
rect 393581 -14730 393648 -14674
rect 393308 -14816 393648 -14730
rect 393308 -14872 393383 -14816
rect 393439 -14872 393525 -14816
rect 393581 -14872 393648 -14816
rect 393308 -14958 393648 -14872
rect 393308 -15014 393383 -14958
rect 393439 -15014 393525 -14958
rect 393581 -15014 393648 -14958
rect 393308 -15100 393648 -15014
rect 393308 -15156 393383 -15100
rect 393439 -15156 393525 -15100
rect 393581 -15156 393648 -15100
rect 393308 -15242 393648 -15156
rect 393308 -15298 393383 -15242
rect 393439 -15298 393525 -15242
rect 393581 -15298 393648 -15242
rect 393308 -15384 393648 -15298
rect 393308 -15440 393383 -15384
rect 393439 -15440 393525 -15384
rect 393581 -15440 393648 -15384
rect 393308 -15526 393648 -15440
rect 393308 -15582 393383 -15526
rect 393439 -15582 393525 -15526
rect 393581 -15582 393648 -15526
rect 393308 -15668 393648 -15582
rect 393308 -15724 393383 -15668
rect 393439 -15724 393525 -15668
rect 393581 -15724 393648 -15668
rect 393308 -15810 393648 -15724
rect 393308 -15866 393383 -15810
rect 393439 -15866 393525 -15810
rect 393581 -15866 393648 -15810
rect 393308 -15952 393648 -15866
rect 393308 -16008 393383 -15952
rect 393439 -16008 393525 -15952
rect 393581 -16008 393648 -15952
rect 393308 -16094 393648 -16008
rect 393308 -16150 393383 -16094
rect 393439 -16150 393525 -16094
rect 393581 -16150 393648 -16094
rect 393308 -16236 393648 -16150
rect 393308 -16292 393383 -16236
rect 393439 -16292 393525 -16236
rect 393581 -16292 393648 -16236
rect 393308 -16378 393648 -16292
rect 393308 -16434 393383 -16378
rect 393439 -16434 393525 -16378
rect 393581 -16434 393648 -16378
rect 393308 -16520 393648 -16434
rect 393308 -16576 393383 -16520
rect 393439 -16576 393525 -16520
rect 393581 -16576 393648 -16520
rect 393308 -16662 393648 -16576
rect 393308 -16718 393383 -16662
rect 393439 -16718 393525 -16662
rect 393581 -16718 393648 -16662
rect 393308 -16804 393648 -16718
rect 393308 -16860 393383 -16804
rect 393439 -16860 393525 -16804
rect 393581 -16860 393648 -16804
rect 393308 -16946 393648 -16860
rect 393308 -17002 393383 -16946
rect 393439 -17002 393525 -16946
rect 393581 -17002 393648 -16946
rect 393308 -17088 393648 -17002
rect 393308 -17144 393383 -17088
rect 393439 -17144 393525 -17088
rect 393581 -17144 393648 -17088
rect 393308 -17230 393648 -17144
rect 393308 -17286 393383 -17230
rect 393439 -17286 393525 -17230
rect 393581 -17286 393648 -17230
rect 393308 -17372 393648 -17286
rect 393308 -17428 393383 -17372
rect 393439 -17428 393525 -17372
rect 393581 -17428 393648 -17372
rect 393308 -17514 393648 -17428
rect 393308 -17570 393383 -17514
rect 393439 -17570 393525 -17514
rect 393581 -17570 393648 -17514
rect 393308 -17656 393648 -17570
rect 393308 -17712 393383 -17656
rect 393439 -17712 393525 -17656
rect 393581 -17712 393648 -17656
rect 393308 -17798 393648 -17712
rect 393308 -17854 393383 -17798
rect 393439 -17854 393525 -17798
rect 393581 -17854 393648 -17798
rect 393308 -17940 393648 -17854
rect 393308 -17996 393383 -17940
rect 393439 -17996 393525 -17940
rect 393581 -17996 393648 -17940
rect 393308 -18082 393648 -17996
rect 393308 -18138 393383 -18082
rect 393439 -18138 393525 -18082
rect 393581 -18138 393648 -18082
rect 393308 -18224 393648 -18138
rect 393308 -18280 393383 -18224
rect 393439 -18280 393525 -18224
rect 393581 -18280 393648 -18224
rect 393308 -18366 393648 -18280
rect 393308 -18422 393383 -18366
rect 393439 -18422 393525 -18366
rect 393581 -18422 393648 -18366
rect 393308 -18508 393648 -18422
rect 393308 -18564 393383 -18508
rect 393439 -18564 393525 -18508
rect 393581 -18564 393648 -18508
rect 393308 -18650 393648 -18564
rect 393308 -18706 393383 -18650
rect 393439 -18706 393525 -18650
rect 393581 -18706 393648 -18650
rect 393308 -18792 393648 -18706
rect 393308 -18848 393383 -18792
rect 393439 -18848 393525 -18792
rect 393581 -18848 393648 -18792
rect 393308 -18934 393648 -18848
rect 393308 -18990 393383 -18934
rect 393439 -18990 393525 -18934
rect 393581 -18990 393648 -18934
rect 393308 -19076 393648 -18990
rect 393308 -19132 393383 -19076
rect 393439 -19132 393525 -19076
rect 393581 -19132 393648 -19076
rect 393308 -19218 393648 -19132
rect 393308 -19274 393383 -19218
rect 393439 -19274 393525 -19218
rect 393581 -19274 393648 -19218
rect 393308 -19360 393648 -19274
rect 393308 -19416 393383 -19360
rect 393439 -19416 393525 -19360
rect 393581 -19416 393648 -19360
rect 393308 -19502 393648 -19416
rect 393308 -19558 393383 -19502
rect 393439 -19558 393525 -19502
rect 393581 -19558 393648 -19502
rect 393308 -19644 393648 -19558
rect 393308 -19700 393383 -19644
rect 393439 -19700 393525 -19644
rect 393581 -19700 393648 -19644
rect 393308 -19786 393648 -19700
rect 393308 -19842 393383 -19786
rect 393439 -19842 393525 -19786
rect 393581 -19842 393648 -19786
rect 393308 -19928 393648 -19842
rect 393308 -19984 393383 -19928
rect 393439 -19984 393525 -19928
rect 393581 -19984 393648 -19928
rect 393308 -20070 393648 -19984
rect 393308 -20126 393383 -20070
rect 393439 -20126 393525 -20070
rect 393581 -20126 393648 -20070
rect 393308 -20212 393648 -20126
rect 393308 -20268 393383 -20212
rect 393439 -20268 393525 -20212
rect 393581 -20268 393648 -20212
rect 393308 -20354 393648 -20268
rect 393308 -20410 393383 -20354
rect 393439 -20410 393525 -20354
rect 393581 -20410 393648 -20354
rect 393308 -20496 393648 -20410
rect 393308 -20552 393383 -20496
rect 393439 -20552 393525 -20496
rect 393581 -20552 393648 -20496
rect 393308 -20638 393648 -20552
rect 393308 -20694 393383 -20638
rect 393439 -20694 393525 -20638
rect 393581 -20694 393648 -20638
rect 393308 -20780 393648 -20694
rect 393308 -20836 393383 -20780
rect 393439 -20836 393525 -20780
rect 393581 -20836 393648 -20780
rect 393308 -20922 393648 -20836
rect 393308 -20978 393383 -20922
rect 393439 -20978 393525 -20922
rect 393581 -20978 393648 -20922
rect 393308 -21064 393648 -20978
rect 393308 -21120 393383 -21064
rect 393439 -21120 393525 -21064
rect 393581 -21120 393648 -21064
rect 393308 -21206 393648 -21120
rect 393308 -21262 393383 -21206
rect 393439 -21262 393525 -21206
rect 393581 -21262 393648 -21206
rect 393308 -21348 393648 -21262
rect 393308 -21404 393383 -21348
rect 393439 -21404 393525 -21348
rect 393581 -21404 393648 -21348
rect 393308 -21490 393648 -21404
rect 393308 -21546 393383 -21490
rect 393439 -21546 393525 -21490
rect 393581 -21546 393648 -21490
rect 393308 -21632 393648 -21546
rect 393308 -21688 393383 -21632
rect 393439 -21688 393525 -21632
rect 393581 -21688 393648 -21632
rect 393308 -21774 393648 -21688
rect 393308 -21830 393383 -21774
rect 393439 -21830 393525 -21774
rect 393581 -21830 393648 -21774
rect 393308 -21916 393648 -21830
rect 393308 -21972 393383 -21916
rect 393439 -21972 393525 -21916
rect 393581 -21972 393648 -21916
rect 393308 -22058 393648 -21972
rect 393308 -22114 393383 -22058
rect 393439 -22114 393525 -22058
rect 393581 -22114 393648 -22058
rect 393308 -22200 393648 -22114
rect 393308 -22256 393383 -22200
rect 393439 -22256 393525 -22200
rect 393581 -22256 393648 -22200
rect 393308 -22342 393648 -22256
rect 393308 -22398 393383 -22342
rect 393439 -22398 393525 -22342
rect 393581 -22398 393648 -22342
rect 393308 -22484 393648 -22398
rect 393308 -22540 393383 -22484
rect 393439 -22540 393525 -22484
rect 393581 -22540 393648 -22484
rect 393308 -22626 393648 -22540
rect 393308 -22682 393383 -22626
rect 393439 -22682 393525 -22626
rect 393581 -22682 393648 -22626
rect 393308 -22768 393648 -22682
rect 393308 -22824 393383 -22768
rect 393439 -22824 393525 -22768
rect 393581 -22824 393648 -22768
rect 393308 -22910 393648 -22824
rect 393308 -22966 393383 -22910
rect 393439 -22966 393525 -22910
rect 393581 -22966 393648 -22910
rect 393308 -23052 393648 -22966
rect 393308 -23108 393383 -23052
rect 393439 -23108 393525 -23052
rect 393581 -23108 393648 -23052
rect 393308 -23194 393648 -23108
rect 393308 -23250 393383 -23194
rect 393439 -23250 393525 -23194
rect 393581 -23250 393648 -23194
rect 393308 -23336 393648 -23250
rect 393308 -23392 393383 -23336
rect 393439 -23392 393525 -23336
rect 393581 -23392 393648 -23336
rect 393308 -23478 393648 -23392
rect 393308 -23534 393383 -23478
rect 393439 -23534 393525 -23478
rect 393581 -23534 393648 -23478
rect 393308 -23620 393648 -23534
rect 393308 -23676 393383 -23620
rect 393439 -23676 393525 -23620
rect 393581 -23676 393648 -23620
rect 393308 -23762 393648 -23676
rect 393308 -23818 393383 -23762
rect 393439 -23818 393525 -23762
rect 393581 -23818 393648 -23762
rect 393308 -23904 393648 -23818
rect 393308 -23960 393383 -23904
rect 393439 -23960 393525 -23904
rect 393581 -23960 393648 -23904
rect 393308 -24046 393648 -23960
rect 393308 -24102 393383 -24046
rect 393439 -24102 393525 -24046
rect 393581 -24102 393648 -24046
rect 393308 -24188 393648 -24102
rect 393308 -24244 393383 -24188
rect 393439 -24244 393525 -24188
rect 393581 -24244 393648 -24188
rect 393308 -24330 393648 -24244
rect 393308 -24386 393383 -24330
rect 393439 -24386 393525 -24330
rect 393581 -24386 393648 -24330
rect 393308 -24472 393648 -24386
rect 393308 -24528 393383 -24472
rect 393439 -24528 393525 -24472
rect 393581 -24528 393648 -24472
rect 393308 -24614 393648 -24528
rect 393308 -24670 393383 -24614
rect 393439 -24670 393525 -24614
rect 393581 -24670 393648 -24614
rect 393308 -24756 393648 -24670
rect 393308 -24812 393383 -24756
rect 393439 -24812 393525 -24756
rect 393581 -24812 393648 -24756
rect 393308 -24898 393648 -24812
rect 393308 -24954 393383 -24898
rect 393439 -24954 393525 -24898
rect 393581 -24954 393648 -24898
rect 393308 -25040 393648 -24954
rect 393308 -25096 393383 -25040
rect 393439 -25096 393525 -25040
rect 393581 -25096 393648 -25040
rect 393308 -25182 393648 -25096
rect 393308 -25238 393383 -25182
rect 393439 -25238 393525 -25182
rect 393581 -25238 393648 -25182
rect 393308 -25324 393648 -25238
rect 393308 -25380 393383 -25324
rect 393439 -25380 393525 -25324
rect 393581 -25380 393648 -25324
rect 393308 -25466 393648 -25380
rect 393308 -25522 393383 -25466
rect 393439 -25522 393525 -25466
rect 393581 -25522 393648 -25466
rect 393308 -25532 393648 -25522
rect 393708 -13680 394048 -13670
rect 393708 -13736 393780 -13680
rect 393836 -13736 393922 -13680
rect 393978 -13736 394048 -13680
rect 393708 -13822 394048 -13736
rect 393708 -13878 393780 -13822
rect 393836 -13878 393922 -13822
rect 393978 -13878 394048 -13822
rect 393708 -13964 394048 -13878
rect 393708 -14020 393780 -13964
rect 393836 -14020 393922 -13964
rect 393978 -14020 394048 -13964
rect 393708 -14106 394048 -14020
rect 393708 -14162 393780 -14106
rect 393836 -14162 393922 -14106
rect 393978 -14162 394048 -14106
rect 393708 -14248 394048 -14162
rect 393708 -14304 393780 -14248
rect 393836 -14304 393922 -14248
rect 393978 -14304 394048 -14248
rect 393708 -14390 394048 -14304
rect 393708 -14446 393780 -14390
rect 393836 -14446 393922 -14390
rect 393978 -14446 394048 -14390
rect 393708 -14532 394048 -14446
rect 393708 -14588 393780 -14532
rect 393836 -14588 393922 -14532
rect 393978 -14588 394048 -14532
rect 393708 -14674 394048 -14588
rect 393708 -14730 393780 -14674
rect 393836 -14730 393922 -14674
rect 393978 -14730 394048 -14674
rect 393708 -14816 394048 -14730
rect 393708 -14872 393780 -14816
rect 393836 -14872 393922 -14816
rect 393978 -14872 394048 -14816
rect 393708 -14958 394048 -14872
rect 393708 -15014 393780 -14958
rect 393836 -15014 393922 -14958
rect 393978 -15014 394048 -14958
rect 393708 -15100 394048 -15014
rect 393708 -15156 393780 -15100
rect 393836 -15156 393922 -15100
rect 393978 -15156 394048 -15100
rect 393708 -15242 394048 -15156
rect 393708 -15298 393780 -15242
rect 393836 -15298 393922 -15242
rect 393978 -15298 394048 -15242
rect 393708 -15384 394048 -15298
rect 393708 -15440 393780 -15384
rect 393836 -15440 393922 -15384
rect 393978 -15440 394048 -15384
rect 393708 -15526 394048 -15440
rect 393708 -15582 393780 -15526
rect 393836 -15582 393922 -15526
rect 393978 -15582 394048 -15526
rect 393708 -15668 394048 -15582
rect 393708 -15724 393780 -15668
rect 393836 -15724 393922 -15668
rect 393978 -15724 394048 -15668
rect 393708 -15810 394048 -15724
rect 393708 -15866 393780 -15810
rect 393836 -15866 393922 -15810
rect 393978 -15866 394048 -15810
rect 393708 -15952 394048 -15866
rect 393708 -16008 393780 -15952
rect 393836 -16008 393922 -15952
rect 393978 -16008 394048 -15952
rect 393708 -16094 394048 -16008
rect 393708 -16150 393780 -16094
rect 393836 -16150 393922 -16094
rect 393978 -16150 394048 -16094
rect 393708 -16236 394048 -16150
rect 393708 -16292 393780 -16236
rect 393836 -16292 393922 -16236
rect 393978 -16292 394048 -16236
rect 393708 -16378 394048 -16292
rect 393708 -16434 393780 -16378
rect 393836 -16434 393922 -16378
rect 393978 -16434 394048 -16378
rect 393708 -16520 394048 -16434
rect 393708 -16576 393780 -16520
rect 393836 -16576 393922 -16520
rect 393978 -16576 394048 -16520
rect 393708 -16662 394048 -16576
rect 393708 -16718 393780 -16662
rect 393836 -16718 393922 -16662
rect 393978 -16718 394048 -16662
rect 393708 -16804 394048 -16718
rect 393708 -16860 393780 -16804
rect 393836 -16860 393922 -16804
rect 393978 -16860 394048 -16804
rect 393708 -16946 394048 -16860
rect 393708 -17002 393780 -16946
rect 393836 -17002 393922 -16946
rect 393978 -17002 394048 -16946
rect 393708 -17088 394048 -17002
rect 393708 -17144 393780 -17088
rect 393836 -17144 393922 -17088
rect 393978 -17144 394048 -17088
rect 393708 -17230 394048 -17144
rect 393708 -17286 393780 -17230
rect 393836 -17286 393922 -17230
rect 393978 -17286 394048 -17230
rect 393708 -17372 394048 -17286
rect 393708 -17428 393780 -17372
rect 393836 -17428 393922 -17372
rect 393978 -17428 394048 -17372
rect 393708 -17514 394048 -17428
rect 393708 -17570 393780 -17514
rect 393836 -17570 393922 -17514
rect 393978 -17570 394048 -17514
rect 393708 -17656 394048 -17570
rect 393708 -17712 393780 -17656
rect 393836 -17712 393922 -17656
rect 393978 -17712 394048 -17656
rect 393708 -17798 394048 -17712
rect 393708 -17854 393780 -17798
rect 393836 -17854 393922 -17798
rect 393978 -17854 394048 -17798
rect 393708 -17940 394048 -17854
rect 393708 -17996 393780 -17940
rect 393836 -17996 393922 -17940
rect 393978 -17996 394048 -17940
rect 393708 -18082 394048 -17996
rect 393708 -18138 393780 -18082
rect 393836 -18138 393922 -18082
rect 393978 -18138 394048 -18082
rect 393708 -18224 394048 -18138
rect 393708 -18280 393780 -18224
rect 393836 -18280 393922 -18224
rect 393978 -18280 394048 -18224
rect 393708 -18366 394048 -18280
rect 393708 -18422 393780 -18366
rect 393836 -18422 393922 -18366
rect 393978 -18422 394048 -18366
rect 393708 -18508 394048 -18422
rect 393708 -18564 393780 -18508
rect 393836 -18564 393922 -18508
rect 393978 -18564 394048 -18508
rect 393708 -18650 394048 -18564
rect 393708 -18706 393780 -18650
rect 393836 -18706 393922 -18650
rect 393978 -18706 394048 -18650
rect 393708 -18792 394048 -18706
rect 393708 -18848 393780 -18792
rect 393836 -18848 393922 -18792
rect 393978 -18848 394048 -18792
rect 393708 -18934 394048 -18848
rect 393708 -18990 393780 -18934
rect 393836 -18990 393922 -18934
rect 393978 -18990 394048 -18934
rect 393708 -19076 394048 -18990
rect 393708 -19132 393780 -19076
rect 393836 -19132 393922 -19076
rect 393978 -19132 394048 -19076
rect 393708 -19218 394048 -19132
rect 393708 -19274 393780 -19218
rect 393836 -19274 393922 -19218
rect 393978 -19274 394048 -19218
rect 393708 -19360 394048 -19274
rect 393708 -19416 393780 -19360
rect 393836 -19416 393922 -19360
rect 393978 -19416 394048 -19360
rect 393708 -19502 394048 -19416
rect 393708 -19558 393780 -19502
rect 393836 -19558 393922 -19502
rect 393978 -19558 394048 -19502
rect 393708 -19644 394048 -19558
rect 393708 -19700 393780 -19644
rect 393836 -19700 393922 -19644
rect 393978 -19700 394048 -19644
rect 393708 -19786 394048 -19700
rect 393708 -19842 393780 -19786
rect 393836 -19842 393922 -19786
rect 393978 -19842 394048 -19786
rect 393708 -19928 394048 -19842
rect 393708 -19984 393780 -19928
rect 393836 -19984 393922 -19928
rect 393978 -19984 394048 -19928
rect 393708 -20070 394048 -19984
rect 393708 -20126 393780 -20070
rect 393836 -20126 393922 -20070
rect 393978 -20126 394048 -20070
rect 393708 -20212 394048 -20126
rect 393708 -20268 393780 -20212
rect 393836 -20268 393922 -20212
rect 393978 -20268 394048 -20212
rect 393708 -20354 394048 -20268
rect 393708 -20410 393780 -20354
rect 393836 -20410 393922 -20354
rect 393978 -20410 394048 -20354
rect 393708 -20496 394048 -20410
rect 393708 -20552 393780 -20496
rect 393836 -20552 393922 -20496
rect 393978 -20552 394048 -20496
rect 393708 -20638 394048 -20552
rect 393708 -20694 393780 -20638
rect 393836 -20694 393922 -20638
rect 393978 -20694 394048 -20638
rect 393708 -20780 394048 -20694
rect 393708 -20836 393780 -20780
rect 393836 -20836 393922 -20780
rect 393978 -20836 394048 -20780
rect 393708 -20922 394048 -20836
rect 393708 -20978 393780 -20922
rect 393836 -20978 393922 -20922
rect 393978 -20978 394048 -20922
rect 393708 -21064 394048 -20978
rect 393708 -21120 393780 -21064
rect 393836 -21120 393922 -21064
rect 393978 -21120 394048 -21064
rect 393708 -21206 394048 -21120
rect 393708 -21262 393780 -21206
rect 393836 -21262 393922 -21206
rect 393978 -21262 394048 -21206
rect 393708 -21348 394048 -21262
rect 393708 -21404 393780 -21348
rect 393836 -21404 393922 -21348
rect 393978 -21404 394048 -21348
rect 393708 -21490 394048 -21404
rect 393708 -21546 393780 -21490
rect 393836 -21546 393922 -21490
rect 393978 -21546 394048 -21490
rect 393708 -21632 394048 -21546
rect 393708 -21688 393780 -21632
rect 393836 -21688 393922 -21632
rect 393978 -21688 394048 -21632
rect 393708 -21774 394048 -21688
rect 393708 -21830 393780 -21774
rect 393836 -21830 393922 -21774
rect 393978 -21830 394048 -21774
rect 393708 -21916 394048 -21830
rect 393708 -21972 393780 -21916
rect 393836 -21972 393922 -21916
rect 393978 -21972 394048 -21916
rect 393708 -22058 394048 -21972
rect 393708 -22114 393780 -22058
rect 393836 -22114 393922 -22058
rect 393978 -22114 394048 -22058
rect 393708 -22200 394048 -22114
rect 393708 -22256 393780 -22200
rect 393836 -22256 393922 -22200
rect 393978 -22256 394048 -22200
rect 393708 -22342 394048 -22256
rect 393708 -22398 393780 -22342
rect 393836 -22398 393922 -22342
rect 393978 -22398 394048 -22342
rect 393708 -22484 394048 -22398
rect 393708 -22540 393780 -22484
rect 393836 -22540 393922 -22484
rect 393978 -22540 394048 -22484
rect 393708 -22626 394048 -22540
rect 393708 -22682 393780 -22626
rect 393836 -22682 393922 -22626
rect 393978 -22682 394048 -22626
rect 393708 -22768 394048 -22682
rect 393708 -22824 393780 -22768
rect 393836 -22824 393922 -22768
rect 393978 -22824 394048 -22768
rect 393708 -22910 394048 -22824
rect 393708 -22966 393780 -22910
rect 393836 -22966 393922 -22910
rect 393978 -22966 394048 -22910
rect 393708 -23052 394048 -22966
rect 393708 -23108 393780 -23052
rect 393836 -23108 393922 -23052
rect 393978 -23108 394048 -23052
rect 393708 -23194 394048 -23108
rect 393708 -23250 393780 -23194
rect 393836 -23250 393922 -23194
rect 393978 -23250 394048 -23194
rect 393708 -23336 394048 -23250
rect 393708 -23392 393780 -23336
rect 393836 -23392 393922 -23336
rect 393978 -23392 394048 -23336
rect 393708 -23478 394048 -23392
rect 393708 -23534 393780 -23478
rect 393836 -23534 393922 -23478
rect 393978 -23534 394048 -23478
rect 393708 -23620 394048 -23534
rect 393708 -23676 393780 -23620
rect 393836 -23676 393922 -23620
rect 393978 -23676 394048 -23620
rect 393708 -23762 394048 -23676
rect 393708 -23818 393780 -23762
rect 393836 -23818 393922 -23762
rect 393978 -23818 394048 -23762
rect 393708 -23904 394048 -23818
rect 393708 -23960 393780 -23904
rect 393836 -23960 393922 -23904
rect 393978 -23960 394048 -23904
rect 393708 -24046 394048 -23960
rect 393708 -24102 393780 -24046
rect 393836 -24102 393922 -24046
rect 393978 -24102 394048 -24046
rect 393708 -24188 394048 -24102
rect 393708 -24244 393780 -24188
rect 393836 -24244 393922 -24188
rect 393978 -24244 394048 -24188
rect 393708 -24330 394048 -24244
rect 393708 -24386 393780 -24330
rect 393836 -24386 393922 -24330
rect 393978 -24386 394048 -24330
rect 393708 -24472 394048 -24386
rect 393708 -24528 393780 -24472
rect 393836 -24528 393922 -24472
rect 393978 -24528 394048 -24472
rect 393708 -24614 394048 -24528
rect 393708 -24670 393780 -24614
rect 393836 -24670 393922 -24614
rect 393978 -24670 394048 -24614
rect 393708 -24756 394048 -24670
rect 393708 -24812 393780 -24756
rect 393836 -24812 393922 -24756
rect 393978 -24812 394048 -24756
rect 393708 -24898 394048 -24812
rect 393708 -24954 393780 -24898
rect 393836 -24954 393922 -24898
rect 393978 -24954 394048 -24898
rect 393708 -25040 394048 -24954
rect 393708 -25096 393780 -25040
rect 393836 -25096 393922 -25040
rect 393978 -25096 394048 -25040
rect 393708 -25182 394048 -25096
rect 393708 -25238 393780 -25182
rect 393836 -25238 393922 -25182
rect 393978 -25238 394048 -25182
rect 393708 -25324 394048 -25238
rect 393708 -25380 393780 -25324
rect 393836 -25380 393922 -25324
rect 393978 -25380 394048 -25324
rect 393708 -25466 394048 -25380
rect 393708 -25522 393780 -25466
rect 393836 -25522 393922 -25466
rect 393978 -25522 394048 -25466
rect 393708 -25532 394048 -25522
rect 394108 -13680 394448 -13670
rect 394108 -13736 394177 -13680
rect 394233 -13736 394319 -13680
rect 394375 -13736 394448 -13680
rect 394108 -13822 394448 -13736
rect 394108 -13878 394177 -13822
rect 394233 -13878 394319 -13822
rect 394375 -13878 394448 -13822
rect 394108 -13964 394448 -13878
rect 394108 -14020 394177 -13964
rect 394233 -14020 394319 -13964
rect 394375 -14020 394448 -13964
rect 394108 -14106 394448 -14020
rect 394108 -14162 394177 -14106
rect 394233 -14162 394319 -14106
rect 394375 -14162 394448 -14106
rect 394108 -14248 394448 -14162
rect 394108 -14304 394177 -14248
rect 394233 -14304 394319 -14248
rect 394375 -14304 394448 -14248
rect 394108 -14390 394448 -14304
rect 394108 -14446 394177 -14390
rect 394233 -14446 394319 -14390
rect 394375 -14446 394448 -14390
rect 394108 -14532 394448 -14446
rect 394108 -14588 394177 -14532
rect 394233 -14588 394319 -14532
rect 394375 -14588 394448 -14532
rect 394108 -14674 394448 -14588
rect 394108 -14730 394177 -14674
rect 394233 -14730 394319 -14674
rect 394375 -14730 394448 -14674
rect 394108 -14816 394448 -14730
rect 394108 -14872 394177 -14816
rect 394233 -14872 394319 -14816
rect 394375 -14872 394448 -14816
rect 394108 -14958 394448 -14872
rect 394108 -15014 394177 -14958
rect 394233 -15014 394319 -14958
rect 394375 -15014 394448 -14958
rect 394108 -15100 394448 -15014
rect 394108 -15156 394177 -15100
rect 394233 -15156 394319 -15100
rect 394375 -15156 394448 -15100
rect 394108 -15242 394448 -15156
rect 394108 -15298 394177 -15242
rect 394233 -15298 394319 -15242
rect 394375 -15298 394448 -15242
rect 394108 -15384 394448 -15298
rect 394108 -15440 394177 -15384
rect 394233 -15440 394319 -15384
rect 394375 -15440 394448 -15384
rect 394108 -15526 394448 -15440
rect 394108 -15582 394177 -15526
rect 394233 -15582 394319 -15526
rect 394375 -15582 394448 -15526
rect 394108 -15668 394448 -15582
rect 394108 -15724 394177 -15668
rect 394233 -15724 394319 -15668
rect 394375 -15724 394448 -15668
rect 394108 -15810 394448 -15724
rect 394108 -15866 394177 -15810
rect 394233 -15866 394319 -15810
rect 394375 -15866 394448 -15810
rect 394108 -15952 394448 -15866
rect 394108 -16008 394177 -15952
rect 394233 -16008 394319 -15952
rect 394375 -16008 394448 -15952
rect 394108 -16094 394448 -16008
rect 394108 -16150 394177 -16094
rect 394233 -16150 394319 -16094
rect 394375 -16150 394448 -16094
rect 394108 -16236 394448 -16150
rect 394108 -16292 394177 -16236
rect 394233 -16292 394319 -16236
rect 394375 -16292 394448 -16236
rect 394108 -16378 394448 -16292
rect 394108 -16434 394177 -16378
rect 394233 -16434 394319 -16378
rect 394375 -16434 394448 -16378
rect 394108 -16520 394448 -16434
rect 394108 -16576 394177 -16520
rect 394233 -16576 394319 -16520
rect 394375 -16576 394448 -16520
rect 394108 -16662 394448 -16576
rect 394108 -16718 394177 -16662
rect 394233 -16718 394319 -16662
rect 394375 -16718 394448 -16662
rect 394108 -16804 394448 -16718
rect 394108 -16860 394177 -16804
rect 394233 -16860 394319 -16804
rect 394375 -16860 394448 -16804
rect 394108 -16946 394448 -16860
rect 394108 -17002 394177 -16946
rect 394233 -17002 394319 -16946
rect 394375 -17002 394448 -16946
rect 394108 -17088 394448 -17002
rect 394108 -17144 394177 -17088
rect 394233 -17144 394319 -17088
rect 394375 -17144 394448 -17088
rect 394108 -17230 394448 -17144
rect 394108 -17286 394177 -17230
rect 394233 -17286 394319 -17230
rect 394375 -17286 394448 -17230
rect 394108 -17372 394448 -17286
rect 394108 -17428 394177 -17372
rect 394233 -17428 394319 -17372
rect 394375 -17428 394448 -17372
rect 394108 -17514 394448 -17428
rect 394108 -17570 394177 -17514
rect 394233 -17570 394319 -17514
rect 394375 -17570 394448 -17514
rect 394108 -17656 394448 -17570
rect 394108 -17712 394177 -17656
rect 394233 -17712 394319 -17656
rect 394375 -17712 394448 -17656
rect 394108 -17798 394448 -17712
rect 394108 -17854 394177 -17798
rect 394233 -17854 394319 -17798
rect 394375 -17854 394448 -17798
rect 394108 -17940 394448 -17854
rect 394108 -17996 394177 -17940
rect 394233 -17996 394319 -17940
rect 394375 -17996 394448 -17940
rect 394108 -18082 394448 -17996
rect 394108 -18138 394177 -18082
rect 394233 -18138 394319 -18082
rect 394375 -18138 394448 -18082
rect 394108 -18224 394448 -18138
rect 394108 -18280 394177 -18224
rect 394233 -18280 394319 -18224
rect 394375 -18280 394448 -18224
rect 394108 -18366 394448 -18280
rect 394108 -18422 394177 -18366
rect 394233 -18422 394319 -18366
rect 394375 -18422 394448 -18366
rect 394108 -18508 394448 -18422
rect 394108 -18564 394177 -18508
rect 394233 -18564 394319 -18508
rect 394375 -18564 394448 -18508
rect 394108 -18650 394448 -18564
rect 394108 -18706 394177 -18650
rect 394233 -18706 394319 -18650
rect 394375 -18706 394448 -18650
rect 394108 -18792 394448 -18706
rect 394108 -18848 394177 -18792
rect 394233 -18848 394319 -18792
rect 394375 -18848 394448 -18792
rect 394108 -18934 394448 -18848
rect 394108 -18990 394177 -18934
rect 394233 -18990 394319 -18934
rect 394375 -18990 394448 -18934
rect 394108 -19076 394448 -18990
rect 394108 -19132 394177 -19076
rect 394233 -19132 394319 -19076
rect 394375 -19132 394448 -19076
rect 394108 -19218 394448 -19132
rect 394108 -19274 394177 -19218
rect 394233 -19274 394319 -19218
rect 394375 -19274 394448 -19218
rect 394108 -19360 394448 -19274
rect 394108 -19416 394177 -19360
rect 394233 -19416 394319 -19360
rect 394375 -19416 394448 -19360
rect 394108 -19502 394448 -19416
rect 394108 -19558 394177 -19502
rect 394233 -19558 394319 -19502
rect 394375 -19558 394448 -19502
rect 394108 -19644 394448 -19558
rect 394108 -19700 394177 -19644
rect 394233 -19700 394319 -19644
rect 394375 -19700 394448 -19644
rect 394108 -19786 394448 -19700
rect 394108 -19842 394177 -19786
rect 394233 -19842 394319 -19786
rect 394375 -19842 394448 -19786
rect 394108 -19928 394448 -19842
rect 394108 -19984 394177 -19928
rect 394233 -19984 394319 -19928
rect 394375 -19984 394448 -19928
rect 394108 -20070 394448 -19984
rect 394108 -20126 394177 -20070
rect 394233 -20126 394319 -20070
rect 394375 -20126 394448 -20070
rect 394108 -20212 394448 -20126
rect 394108 -20268 394177 -20212
rect 394233 -20268 394319 -20212
rect 394375 -20268 394448 -20212
rect 394108 -20354 394448 -20268
rect 394108 -20410 394177 -20354
rect 394233 -20410 394319 -20354
rect 394375 -20410 394448 -20354
rect 394108 -20496 394448 -20410
rect 394108 -20552 394177 -20496
rect 394233 -20552 394319 -20496
rect 394375 -20552 394448 -20496
rect 394108 -20638 394448 -20552
rect 394108 -20694 394177 -20638
rect 394233 -20694 394319 -20638
rect 394375 -20694 394448 -20638
rect 394108 -20780 394448 -20694
rect 394108 -20836 394177 -20780
rect 394233 -20836 394319 -20780
rect 394375 -20836 394448 -20780
rect 394108 -20922 394448 -20836
rect 394108 -20978 394177 -20922
rect 394233 -20978 394319 -20922
rect 394375 -20978 394448 -20922
rect 394108 -21064 394448 -20978
rect 394108 -21120 394177 -21064
rect 394233 -21120 394319 -21064
rect 394375 -21120 394448 -21064
rect 394108 -21206 394448 -21120
rect 394108 -21262 394177 -21206
rect 394233 -21262 394319 -21206
rect 394375 -21262 394448 -21206
rect 394108 -21348 394448 -21262
rect 394108 -21404 394177 -21348
rect 394233 -21404 394319 -21348
rect 394375 -21404 394448 -21348
rect 394108 -21490 394448 -21404
rect 394108 -21546 394177 -21490
rect 394233 -21546 394319 -21490
rect 394375 -21546 394448 -21490
rect 394108 -21632 394448 -21546
rect 394108 -21688 394177 -21632
rect 394233 -21688 394319 -21632
rect 394375 -21688 394448 -21632
rect 394108 -21774 394448 -21688
rect 394108 -21830 394177 -21774
rect 394233 -21830 394319 -21774
rect 394375 -21830 394448 -21774
rect 394108 -21916 394448 -21830
rect 394108 -21972 394177 -21916
rect 394233 -21972 394319 -21916
rect 394375 -21972 394448 -21916
rect 394108 -22058 394448 -21972
rect 394108 -22114 394177 -22058
rect 394233 -22114 394319 -22058
rect 394375 -22114 394448 -22058
rect 394108 -22200 394448 -22114
rect 394108 -22256 394177 -22200
rect 394233 -22256 394319 -22200
rect 394375 -22256 394448 -22200
rect 394108 -22342 394448 -22256
rect 394108 -22398 394177 -22342
rect 394233 -22398 394319 -22342
rect 394375 -22398 394448 -22342
rect 394108 -22484 394448 -22398
rect 394108 -22540 394177 -22484
rect 394233 -22540 394319 -22484
rect 394375 -22540 394448 -22484
rect 394108 -22626 394448 -22540
rect 394108 -22682 394177 -22626
rect 394233 -22682 394319 -22626
rect 394375 -22682 394448 -22626
rect 394108 -22768 394448 -22682
rect 394108 -22824 394177 -22768
rect 394233 -22824 394319 -22768
rect 394375 -22824 394448 -22768
rect 394108 -22910 394448 -22824
rect 394108 -22966 394177 -22910
rect 394233 -22966 394319 -22910
rect 394375 -22966 394448 -22910
rect 394108 -23052 394448 -22966
rect 394108 -23108 394177 -23052
rect 394233 -23108 394319 -23052
rect 394375 -23108 394448 -23052
rect 394108 -23194 394448 -23108
rect 394108 -23250 394177 -23194
rect 394233 -23250 394319 -23194
rect 394375 -23250 394448 -23194
rect 394108 -23336 394448 -23250
rect 394108 -23392 394177 -23336
rect 394233 -23392 394319 -23336
rect 394375 -23392 394448 -23336
rect 394108 -23478 394448 -23392
rect 394108 -23534 394177 -23478
rect 394233 -23534 394319 -23478
rect 394375 -23534 394448 -23478
rect 394108 -23620 394448 -23534
rect 394108 -23676 394177 -23620
rect 394233 -23676 394319 -23620
rect 394375 -23676 394448 -23620
rect 394108 -23762 394448 -23676
rect 394108 -23818 394177 -23762
rect 394233 -23818 394319 -23762
rect 394375 -23818 394448 -23762
rect 394108 -23904 394448 -23818
rect 394108 -23960 394177 -23904
rect 394233 -23960 394319 -23904
rect 394375 -23960 394448 -23904
rect 394108 -24046 394448 -23960
rect 394108 -24102 394177 -24046
rect 394233 -24102 394319 -24046
rect 394375 -24102 394448 -24046
rect 394108 -24188 394448 -24102
rect 394108 -24244 394177 -24188
rect 394233 -24244 394319 -24188
rect 394375 -24244 394448 -24188
rect 394108 -24330 394448 -24244
rect 394108 -24386 394177 -24330
rect 394233 -24386 394319 -24330
rect 394375 -24386 394448 -24330
rect 394108 -24472 394448 -24386
rect 394108 -24528 394177 -24472
rect 394233 -24528 394319 -24472
rect 394375 -24528 394448 -24472
rect 394108 -24614 394448 -24528
rect 394108 -24670 394177 -24614
rect 394233 -24670 394319 -24614
rect 394375 -24670 394448 -24614
rect 394108 -24756 394448 -24670
rect 394108 -24812 394177 -24756
rect 394233 -24812 394319 -24756
rect 394375 -24812 394448 -24756
rect 394108 -24898 394448 -24812
rect 394108 -24954 394177 -24898
rect 394233 -24954 394319 -24898
rect 394375 -24954 394448 -24898
rect 394108 -25040 394448 -24954
rect 394108 -25096 394177 -25040
rect 394233 -25096 394319 -25040
rect 394375 -25096 394448 -25040
rect 394108 -25182 394448 -25096
rect 394108 -25238 394177 -25182
rect 394233 -25238 394319 -25182
rect 394375 -25238 394448 -25182
rect 394108 -25324 394448 -25238
rect 394108 -25380 394177 -25324
rect 394233 -25380 394319 -25324
rect 394375 -25380 394448 -25324
rect 394108 -25466 394448 -25380
rect 394108 -25522 394177 -25466
rect 394233 -25522 394319 -25466
rect 394375 -25522 394448 -25466
rect 394108 -25532 394448 -25522
rect 394508 -13680 394848 -13670
rect 394508 -13736 394580 -13680
rect 394636 -13736 394722 -13680
rect 394778 -13736 394848 -13680
rect 394508 -13822 394848 -13736
rect 394508 -13878 394580 -13822
rect 394636 -13878 394722 -13822
rect 394778 -13878 394848 -13822
rect 394508 -13964 394848 -13878
rect 394508 -14020 394580 -13964
rect 394636 -14020 394722 -13964
rect 394778 -14020 394848 -13964
rect 394508 -14106 394848 -14020
rect 394508 -14162 394580 -14106
rect 394636 -14162 394722 -14106
rect 394778 -14162 394848 -14106
rect 394508 -14248 394848 -14162
rect 394508 -14304 394580 -14248
rect 394636 -14304 394722 -14248
rect 394778 -14304 394848 -14248
rect 394508 -14390 394848 -14304
rect 394508 -14446 394580 -14390
rect 394636 -14446 394722 -14390
rect 394778 -14446 394848 -14390
rect 394508 -14532 394848 -14446
rect 394508 -14588 394580 -14532
rect 394636 -14588 394722 -14532
rect 394778 -14588 394848 -14532
rect 394508 -14674 394848 -14588
rect 394508 -14730 394580 -14674
rect 394636 -14730 394722 -14674
rect 394778 -14730 394848 -14674
rect 394508 -14816 394848 -14730
rect 394508 -14872 394580 -14816
rect 394636 -14872 394722 -14816
rect 394778 -14872 394848 -14816
rect 394508 -14958 394848 -14872
rect 394508 -15014 394580 -14958
rect 394636 -15014 394722 -14958
rect 394778 -15014 394848 -14958
rect 394508 -15100 394848 -15014
rect 394508 -15156 394580 -15100
rect 394636 -15156 394722 -15100
rect 394778 -15156 394848 -15100
rect 394508 -15242 394848 -15156
rect 394508 -15298 394580 -15242
rect 394636 -15298 394722 -15242
rect 394778 -15298 394848 -15242
rect 394508 -15384 394848 -15298
rect 394508 -15440 394580 -15384
rect 394636 -15440 394722 -15384
rect 394778 -15440 394848 -15384
rect 394508 -15526 394848 -15440
rect 394508 -15582 394580 -15526
rect 394636 -15582 394722 -15526
rect 394778 -15582 394848 -15526
rect 394508 -15668 394848 -15582
rect 394508 -15724 394580 -15668
rect 394636 -15724 394722 -15668
rect 394778 -15724 394848 -15668
rect 394508 -15810 394848 -15724
rect 394508 -15866 394580 -15810
rect 394636 -15866 394722 -15810
rect 394778 -15866 394848 -15810
rect 394508 -15952 394848 -15866
rect 394508 -16008 394580 -15952
rect 394636 -16008 394722 -15952
rect 394778 -16008 394848 -15952
rect 394508 -16094 394848 -16008
rect 394508 -16150 394580 -16094
rect 394636 -16150 394722 -16094
rect 394778 -16150 394848 -16094
rect 394508 -16236 394848 -16150
rect 394508 -16292 394580 -16236
rect 394636 -16292 394722 -16236
rect 394778 -16292 394848 -16236
rect 394508 -16378 394848 -16292
rect 394508 -16434 394580 -16378
rect 394636 -16434 394722 -16378
rect 394778 -16434 394848 -16378
rect 394508 -16520 394848 -16434
rect 394508 -16576 394580 -16520
rect 394636 -16576 394722 -16520
rect 394778 -16576 394848 -16520
rect 394508 -16662 394848 -16576
rect 394508 -16718 394580 -16662
rect 394636 -16718 394722 -16662
rect 394778 -16718 394848 -16662
rect 394508 -16804 394848 -16718
rect 394508 -16860 394580 -16804
rect 394636 -16860 394722 -16804
rect 394778 -16860 394848 -16804
rect 394508 -16946 394848 -16860
rect 394508 -17002 394580 -16946
rect 394636 -17002 394722 -16946
rect 394778 -17002 394848 -16946
rect 394508 -17088 394848 -17002
rect 394508 -17144 394580 -17088
rect 394636 -17144 394722 -17088
rect 394778 -17144 394848 -17088
rect 394508 -17230 394848 -17144
rect 394508 -17286 394580 -17230
rect 394636 -17286 394722 -17230
rect 394778 -17286 394848 -17230
rect 394508 -17372 394848 -17286
rect 394508 -17428 394580 -17372
rect 394636 -17428 394722 -17372
rect 394778 -17428 394848 -17372
rect 394508 -17514 394848 -17428
rect 394508 -17570 394580 -17514
rect 394636 -17570 394722 -17514
rect 394778 -17570 394848 -17514
rect 394508 -17656 394848 -17570
rect 394508 -17712 394580 -17656
rect 394636 -17712 394722 -17656
rect 394778 -17712 394848 -17656
rect 394508 -17798 394848 -17712
rect 394508 -17854 394580 -17798
rect 394636 -17854 394722 -17798
rect 394778 -17854 394848 -17798
rect 394508 -17940 394848 -17854
rect 394508 -17996 394580 -17940
rect 394636 -17996 394722 -17940
rect 394778 -17996 394848 -17940
rect 394508 -18082 394848 -17996
rect 394508 -18138 394580 -18082
rect 394636 -18138 394722 -18082
rect 394778 -18138 394848 -18082
rect 394508 -18224 394848 -18138
rect 394508 -18280 394580 -18224
rect 394636 -18280 394722 -18224
rect 394778 -18280 394848 -18224
rect 394508 -18366 394848 -18280
rect 394508 -18422 394580 -18366
rect 394636 -18422 394722 -18366
rect 394778 -18422 394848 -18366
rect 394508 -18508 394848 -18422
rect 394508 -18564 394580 -18508
rect 394636 -18564 394722 -18508
rect 394778 -18564 394848 -18508
rect 394508 -18650 394848 -18564
rect 394508 -18706 394580 -18650
rect 394636 -18706 394722 -18650
rect 394778 -18706 394848 -18650
rect 394508 -18792 394848 -18706
rect 394508 -18848 394580 -18792
rect 394636 -18848 394722 -18792
rect 394778 -18848 394848 -18792
rect 394508 -18934 394848 -18848
rect 394508 -18990 394580 -18934
rect 394636 -18990 394722 -18934
rect 394778 -18990 394848 -18934
rect 394508 -19076 394848 -18990
rect 394508 -19132 394580 -19076
rect 394636 -19132 394722 -19076
rect 394778 -19132 394848 -19076
rect 394508 -19218 394848 -19132
rect 394508 -19274 394580 -19218
rect 394636 -19274 394722 -19218
rect 394778 -19274 394848 -19218
rect 394508 -19360 394848 -19274
rect 394508 -19416 394580 -19360
rect 394636 -19416 394722 -19360
rect 394778 -19416 394848 -19360
rect 394508 -19502 394848 -19416
rect 394508 -19558 394580 -19502
rect 394636 -19558 394722 -19502
rect 394778 -19558 394848 -19502
rect 394508 -19644 394848 -19558
rect 394508 -19700 394580 -19644
rect 394636 -19700 394722 -19644
rect 394778 -19700 394848 -19644
rect 394508 -19786 394848 -19700
rect 394508 -19842 394580 -19786
rect 394636 -19842 394722 -19786
rect 394778 -19842 394848 -19786
rect 394508 -19928 394848 -19842
rect 394508 -19984 394580 -19928
rect 394636 -19984 394722 -19928
rect 394778 -19984 394848 -19928
rect 394508 -20070 394848 -19984
rect 394508 -20126 394580 -20070
rect 394636 -20126 394722 -20070
rect 394778 -20126 394848 -20070
rect 394508 -20212 394848 -20126
rect 394508 -20268 394580 -20212
rect 394636 -20268 394722 -20212
rect 394778 -20268 394848 -20212
rect 394508 -20354 394848 -20268
rect 394508 -20410 394580 -20354
rect 394636 -20410 394722 -20354
rect 394778 -20410 394848 -20354
rect 394508 -20496 394848 -20410
rect 394508 -20552 394580 -20496
rect 394636 -20552 394722 -20496
rect 394778 -20552 394848 -20496
rect 394508 -20638 394848 -20552
rect 394508 -20694 394580 -20638
rect 394636 -20694 394722 -20638
rect 394778 -20694 394848 -20638
rect 394508 -20780 394848 -20694
rect 394508 -20836 394580 -20780
rect 394636 -20836 394722 -20780
rect 394778 -20836 394848 -20780
rect 394508 -20922 394848 -20836
rect 394508 -20978 394580 -20922
rect 394636 -20978 394722 -20922
rect 394778 -20978 394848 -20922
rect 394508 -21064 394848 -20978
rect 394508 -21120 394580 -21064
rect 394636 -21120 394722 -21064
rect 394778 -21120 394848 -21064
rect 394508 -21206 394848 -21120
rect 394508 -21262 394580 -21206
rect 394636 -21262 394722 -21206
rect 394778 -21262 394848 -21206
rect 394508 -21348 394848 -21262
rect 394508 -21404 394580 -21348
rect 394636 -21404 394722 -21348
rect 394778 -21404 394848 -21348
rect 394508 -21490 394848 -21404
rect 394508 -21546 394580 -21490
rect 394636 -21546 394722 -21490
rect 394778 -21546 394848 -21490
rect 394508 -21632 394848 -21546
rect 394508 -21688 394580 -21632
rect 394636 -21688 394722 -21632
rect 394778 -21688 394848 -21632
rect 394508 -21774 394848 -21688
rect 394508 -21830 394580 -21774
rect 394636 -21830 394722 -21774
rect 394778 -21830 394848 -21774
rect 394508 -21916 394848 -21830
rect 394508 -21972 394580 -21916
rect 394636 -21972 394722 -21916
rect 394778 -21972 394848 -21916
rect 394508 -22058 394848 -21972
rect 394508 -22114 394580 -22058
rect 394636 -22114 394722 -22058
rect 394778 -22114 394848 -22058
rect 394508 -22200 394848 -22114
rect 394508 -22256 394580 -22200
rect 394636 -22256 394722 -22200
rect 394778 -22256 394848 -22200
rect 394508 -22342 394848 -22256
rect 394508 -22398 394580 -22342
rect 394636 -22398 394722 -22342
rect 394778 -22398 394848 -22342
rect 394508 -22484 394848 -22398
rect 394508 -22540 394580 -22484
rect 394636 -22540 394722 -22484
rect 394778 -22540 394848 -22484
rect 394508 -22626 394848 -22540
rect 394508 -22682 394580 -22626
rect 394636 -22682 394722 -22626
rect 394778 -22682 394848 -22626
rect 394508 -22768 394848 -22682
rect 394508 -22824 394580 -22768
rect 394636 -22824 394722 -22768
rect 394778 -22824 394848 -22768
rect 394508 -22910 394848 -22824
rect 394508 -22966 394580 -22910
rect 394636 -22966 394722 -22910
rect 394778 -22966 394848 -22910
rect 394508 -23052 394848 -22966
rect 394508 -23108 394580 -23052
rect 394636 -23108 394722 -23052
rect 394778 -23108 394848 -23052
rect 394508 -23194 394848 -23108
rect 394508 -23250 394580 -23194
rect 394636 -23250 394722 -23194
rect 394778 -23250 394848 -23194
rect 394508 -23336 394848 -23250
rect 394508 -23392 394580 -23336
rect 394636 -23392 394722 -23336
rect 394778 -23392 394848 -23336
rect 394508 -23478 394848 -23392
rect 394508 -23534 394580 -23478
rect 394636 -23534 394722 -23478
rect 394778 -23534 394848 -23478
rect 394508 -23620 394848 -23534
rect 394508 -23676 394580 -23620
rect 394636 -23676 394722 -23620
rect 394778 -23676 394848 -23620
rect 394508 -23762 394848 -23676
rect 394508 -23818 394580 -23762
rect 394636 -23818 394722 -23762
rect 394778 -23818 394848 -23762
rect 394508 -23904 394848 -23818
rect 394508 -23960 394580 -23904
rect 394636 -23960 394722 -23904
rect 394778 -23960 394848 -23904
rect 394508 -24046 394848 -23960
rect 394508 -24102 394580 -24046
rect 394636 -24102 394722 -24046
rect 394778 -24102 394848 -24046
rect 394508 -24188 394848 -24102
rect 394508 -24244 394580 -24188
rect 394636 -24244 394722 -24188
rect 394778 -24244 394848 -24188
rect 394508 -24330 394848 -24244
rect 394508 -24386 394580 -24330
rect 394636 -24386 394722 -24330
rect 394778 -24386 394848 -24330
rect 394508 -24472 394848 -24386
rect 394508 -24528 394580 -24472
rect 394636 -24528 394722 -24472
rect 394778 -24528 394848 -24472
rect 394508 -24614 394848 -24528
rect 394508 -24670 394580 -24614
rect 394636 -24670 394722 -24614
rect 394778 -24670 394848 -24614
rect 394508 -24756 394848 -24670
rect 394508 -24812 394580 -24756
rect 394636 -24812 394722 -24756
rect 394778 -24812 394848 -24756
rect 394508 -24898 394848 -24812
rect 394508 -24954 394580 -24898
rect 394636 -24954 394722 -24898
rect 394778 -24954 394848 -24898
rect 394508 -25040 394848 -24954
rect 394508 -25096 394580 -25040
rect 394636 -25096 394722 -25040
rect 394778 -25096 394848 -25040
rect 394508 -25182 394848 -25096
rect 394508 -25238 394580 -25182
rect 394636 -25238 394722 -25182
rect 394778 -25238 394848 -25182
rect 394508 -25324 394848 -25238
rect 394508 -25380 394580 -25324
rect 394636 -25380 394722 -25324
rect 394778 -25380 394848 -25324
rect 394508 -25466 394848 -25380
rect 394508 -25522 394580 -25466
rect 394636 -25522 394722 -25466
rect 394778 -25522 394848 -25466
rect 394508 -25532 394848 -25522
rect 394908 -13680 395248 -13670
rect 394908 -13736 394982 -13680
rect 395038 -13736 395124 -13680
rect 395180 -13736 395248 -13680
rect 394908 -13822 395248 -13736
rect 394908 -13878 394982 -13822
rect 395038 -13878 395124 -13822
rect 395180 -13878 395248 -13822
rect 394908 -13964 395248 -13878
rect 394908 -14020 394982 -13964
rect 395038 -14020 395124 -13964
rect 395180 -14020 395248 -13964
rect 394908 -14106 395248 -14020
rect 394908 -14162 394982 -14106
rect 395038 -14162 395124 -14106
rect 395180 -14162 395248 -14106
rect 394908 -14248 395248 -14162
rect 394908 -14304 394982 -14248
rect 395038 -14304 395124 -14248
rect 395180 -14304 395248 -14248
rect 394908 -14390 395248 -14304
rect 394908 -14446 394982 -14390
rect 395038 -14446 395124 -14390
rect 395180 -14446 395248 -14390
rect 394908 -14532 395248 -14446
rect 394908 -14588 394982 -14532
rect 395038 -14588 395124 -14532
rect 395180 -14588 395248 -14532
rect 394908 -14674 395248 -14588
rect 394908 -14730 394982 -14674
rect 395038 -14730 395124 -14674
rect 395180 -14730 395248 -14674
rect 394908 -14816 395248 -14730
rect 394908 -14872 394982 -14816
rect 395038 -14872 395124 -14816
rect 395180 -14872 395248 -14816
rect 394908 -14958 395248 -14872
rect 394908 -15014 394982 -14958
rect 395038 -15014 395124 -14958
rect 395180 -15014 395248 -14958
rect 394908 -15100 395248 -15014
rect 394908 -15156 394982 -15100
rect 395038 -15156 395124 -15100
rect 395180 -15156 395248 -15100
rect 394908 -15242 395248 -15156
rect 394908 -15298 394982 -15242
rect 395038 -15298 395124 -15242
rect 395180 -15298 395248 -15242
rect 394908 -15384 395248 -15298
rect 394908 -15440 394982 -15384
rect 395038 -15440 395124 -15384
rect 395180 -15440 395248 -15384
rect 394908 -15526 395248 -15440
rect 394908 -15582 394982 -15526
rect 395038 -15582 395124 -15526
rect 395180 -15582 395248 -15526
rect 394908 -15668 395248 -15582
rect 394908 -15724 394982 -15668
rect 395038 -15724 395124 -15668
rect 395180 -15724 395248 -15668
rect 394908 -15810 395248 -15724
rect 394908 -15866 394982 -15810
rect 395038 -15866 395124 -15810
rect 395180 -15866 395248 -15810
rect 394908 -15952 395248 -15866
rect 394908 -16008 394982 -15952
rect 395038 -16008 395124 -15952
rect 395180 -16008 395248 -15952
rect 394908 -16094 395248 -16008
rect 394908 -16150 394982 -16094
rect 395038 -16150 395124 -16094
rect 395180 -16150 395248 -16094
rect 394908 -16236 395248 -16150
rect 394908 -16292 394982 -16236
rect 395038 -16292 395124 -16236
rect 395180 -16292 395248 -16236
rect 394908 -16378 395248 -16292
rect 394908 -16434 394982 -16378
rect 395038 -16434 395124 -16378
rect 395180 -16434 395248 -16378
rect 394908 -16520 395248 -16434
rect 394908 -16576 394982 -16520
rect 395038 -16576 395124 -16520
rect 395180 -16576 395248 -16520
rect 394908 -16662 395248 -16576
rect 394908 -16718 394982 -16662
rect 395038 -16718 395124 -16662
rect 395180 -16718 395248 -16662
rect 394908 -16804 395248 -16718
rect 394908 -16860 394982 -16804
rect 395038 -16860 395124 -16804
rect 395180 -16860 395248 -16804
rect 394908 -16946 395248 -16860
rect 394908 -17002 394982 -16946
rect 395038 -17002 395124 -16946
rect 395180 -17002 395248 -16946
rect 394908 -17088 395248 -17002
rect 394908 -17144 394982 -17088
rect 395038 -17144 395124 -17088
rect 395180 -17144 395248 -17088
rect 394908 -17230 395248 -17144
rect 394908 -17286 394982 -17230
rect 395038 -17286 395124 -17230
rect 395180 -17286 395248 -17230
rect 394908 -17372 395248 -17286
rect 394908 -17428 394982 -17372
rect 395038 -17428 395124 -17372
rect 395180 -17428 395248 -17372
rect 394908 -17514 395248 -17428
rect 394908 -17570 394982 -17514
rect 395038 -17570 395124 -17514
rect 395180 -17570 395248 -17514
rect 394908 -17656 395248 -17570
rect 394908 -17712 394982 -17656
rect 395038 -17712 395124 -17656
rect 395180 -17712 395248 -17656
rect 394908 -17798 395248 -17712
rect 394908 -17854 394982 -17798
rect 395038 -17854 395124 -17798
rect 395180 -17854 395248 -17798
rect 394908 -17940 395248 -17854
rect 394908 -17996 394982 -17940
rect 395038 -17996 395124 -17940
rect 395180 -17996 395248 -17940
rect 394908 -18082 395248 -17996
rect 394908 -18138 394982 -18082
rect 395038 -18138 395124 -18082
rect 395180 -18138 395248 -18082
rect 394908 -18224 395248 -18138
rect 394908 -18280 394982 -18224
rect 395038 -18280 395124 -18224
rect 395180 -18280 395248 -18224
rect 394908 -18366 395248 -18280
rect 394908 -18422 394982 -18366
rect 395038 -18422 395124 -18366
rect 395180 -18422 395248 -18366
rect 394908 -18508 395248 -18422
rect 394908 -18564 394982 -18508
rect 395038 -18564 395124 -18508
rect 395180 -18564 395248 -18508
rect 394908 -18650 395248 -18564
rect 394908 -18706 394982 -18650
rect 395038 -18706 395124 -18650
rect 395180 -18706 395248 -18650
rect 394908 -18792 395248 -18706
rect 394908 -18848 394982 -18792
rect 395038 -18848 395124 -18792
rect 395180 -18848 395248 -18792
rect 394908 -18934 395248 -18848
rect 394908 -18990 394982 -18934
rect 395038 -18990 395124 -18934
rect 395180 -18990 395248 -18934
rect 394908 -19076 395248 -18990
rect 394908 -19132 394982 -19076
rect 395038 -19132 395124 -19076
rect 395180 -19132 395248 -19076
rect 394908 -19218 395248 -19132
rect 394908 -19274 394982 -19218
rect 395038 -19274 395124 -19218
rect 395180 -19274 395248 -19218
rect 394908 -19360 395248 -19274
rect 394908 -19416 394982 -19360
rect 395038 -19416 395124 -19360
rect 395180 -19416 395248 -19360
rect 394908 -19502 395248 -19416
rect 394908 -19558 394982 -19502
rect 395038 -19558 395124 -19502
rect 395180 -19558 395248 -19502
rect 394908 -19644 395248 -19558
rect 394908 -19700 394982 -19644
rect 395038 -19700 395124 -19644
rect 395180 -19700 395248 -19644
rect 394908 -19786 395248 -19700
rect 394908 -19842 394982 -19786
rect 395038 -19842 395124 -19786
rect 395180 -19842 395248 -19786
rect 394908 -19928 395248 -19842
rect 394908 -19984 394982 -19928
rect 395038 -19984 395124 -19928
rect 395180 -19984 395248 -19928
rect 394908 -20070 395248 -19984
rect 394908 -20126 394982 -20070
rect 395038 -20126 395124 -20070
rect 395180 -20126 395248 -20070
rect 394908 -20212 395248 -20126
rect 394908 -20268 394982 -20212
rect 395038 -20268 395124 -20212
rect 395180 -20268 395248 -20212
rect 394908 -20354 395248 -20268
rect 394908 -20410 394982 -20354
rect 395038 -20410 395124 -20354
rect 395180 -20410 395248 -20354
rect 394908 -20496 395248 -20410
rect 394908 -20552 394982 -20496
rect 395038 -20552 395124 -20496
rect 395180 -20552 395248 -20496
rect 394908 -20638 395248 -20552
rect 394908 -20694 394982 -20638
rect 395038 -20694 395124 -20638
rect 395180 -20694 395248 -20638
rect 394908 -20780 395248 -20694
rect 394908 -20836 394982 -20780
rect 395038 -20836 395124 -20780
rect 395180 -20836 395248 -20780
rect 394908 -20922 395248 -20836
rect 394908 -20978 394982 -20922
rect 395038 -20978 395124 -20922
rect 395180 -20978 395248 -20922
rect 394908 -21064 395248 -20978
rect 394908 -21120 394982 -21064
rect 395038 -21120 395124 -21064
rect 395180 -21120 395248 -21064
rect 394908 -21206 395248 -21120
rect 394908 -21262 394982 -21206
rect 395038 -21262 395124 -21206
rect 395180 -21262 395248 -21206
rect 394908 -21348 395248 -21262
rect 394908 -21404 394982 -21348
rect 395038 -21404 395124 -21348
rect 395180 -21404 395248 -21348
rect 394908 -21490 395248 -21404
rect 394908 -21546 394982 -21490
rect 395038 -21546 395124 -21490
rect 395180 -21546 395248 -21490
rect 394908 -21632 395248 -21546
rect 394908 -21688 394982 -21632
rect 395038 -21688 395124 -21632
rect 395180 -21688 395248 -21632
rect 394908 -21774 395248 -21688
rect 394908 -21830 394982 -21774
rect 395038 -21830 395124 -21774
rect 395180 -21830 395248 -21774
rect 394908 -21916 395248 -21830
rect 394908 -21972 394982 -21916
rect 395038 -21972 395124 -21916
rect 395180 -21972 395248 -21916
rect 394908 -22058 395248 -21972
rect 394908 -22114 394982 -22058
rect 395038 -22114 395124 -22058
rect 395180 -22114 395248 -22058
rect 394908 -22200 395248 -22114
rect 394908 -22256 394982 -22200
rect 395038 -22256 395124 -22200
rect 395180 -22256 395248 -22200
rect 394908 -22342 395248 -22256
rect 394908 -22398 394982 -22342
rect 395038 -22398 395124 -22342
rect 395180 -22398 395248 -22342
rect 394908 -22484 395248 -22398
rect 394908 -22540 394982 -22484
rect 395038 -22540 395124 -22484
rect 395180 -22540 395248 -22484
rect 394908 -22626 395248 -22540
rect 394908 -22682 394982 -22626
rect 395038 -22682 395124 -22626
rect 395180 -22682 395248 -22626
rect 394908 -22768 395248 -22682
rect 394908 -22824 394982 -22768
rect 395038 -22824 395124 -22768
rect 395180 -22824 395248 -22768
rect 394908 -22910 395248 -22824
rect 394908 -22966 394982 -22910
rect 395038 -22966 395124 -22910
rect 395180 -22966 395248 -22910
rect 394908 -23052 395248 -22966
rect 394908 -23108 394982 -23052
rect 395038 -23108 395124 -23052
rect 395180 -23108 395248 -23052
rect 394908 -23194 395248 -23108
rect 394908 -23250 394982 -23194
rect 395038 -23250 395124 -23194
rect 395180 -23250 395248 -23194
rect 394908 -23336 395248 -23250
rect 394908 -23392 394982 -23336
rect 395038 -23392 395124 -23336
rect 395180 -23392 395248 -23336
rect 394908 -23478 395248 -23392
rect 394908 -23534 394982 -23478
rect 395038 -23534 395124 -23478
rect 395180 -23534 395248 -23478
rect 394908 -23620 395248 -23534
rect 394908 -23676 394982 -23620
rect 395038 -23676 395124 -23620
rect 395180 -23676 395248 -23620
rect 394908 -23762 395248 -23676
rect 394908 -23818 394982 -23762
rect 395038 -23818 395124 -23762
rect 395180 -23818 395248 -23762
rect 394908 -23904 395248 -23818
rect 394908 -23960 394982 -23904
rect 395038 -23960 395124 -23904
rect 395180 -23960 395248 -23904
rect 394908 -24046 395248 -23960
rect 394908 -24102 394982 -24046
rect 395038 -24102 395124 -24046
rect 395180 -24102 395248 -24046
rect 394908 -24188 395248 -24102
rect 394908 -24244 394982 -24188
rect 395038 -24244 395124 -24188
rect 395180 -24244 395248 -24188
rect 394908 -24330 395248 -24244
rect 394908 -24386 394982 -24330
rect 395038 -24386 395124 -24330
rect 395180 -24386 395248 -24330
rect 394908 -24472 395248 -24386
rect 394908 -24528 394982 -24472
rect 395038 -24528 395124 -24472
rect 395180 -24528 395248 -24472
rect 394908 -24614 395248 -24528
rect 394908 -24670 394982 -24614
rect 395038 -24670 395124 -24614
rect 395180 -24670 395248 -24614
rect 394908 -24756 395248 -24670
rect 394908 -24812 394982 -24756
rect 395038 -24812 395124 -24756
rect 395180 -24812 395248 -24756
rect 394908 -24898 395248 -24812
rect 394908 -24954 394982 -24898
rect 395038 -24954 395124 -24898
rect 395180 -24954 395248 -24898
rect 394908 -25040 395248 -24954
rect 394908 -25096 394982 -25040
rect 395038 -25096 395124 -25040
rect 395180 -25096 395248 -25040
rect 394908 -25182 395248 -25096
rect 394908 -25238 394982 -25182
rect 395038 -25238 395124 -25182
rect 395180 -25238 395248 -25182
rect 394908 -25324 395248 -25238
rect 394908 -25380 394982 -25324
rect 395038 -25380 395124 -25324
rect 395180 -25380 395248 -25324
rect 394908 -25466 395248 -25380
rect 394908 -25522 394982 -25466
rect 395038 -25522 395124 -25466
rect 395180 -25522 395248 -25466
rect 394908 -25532 395248 -25522
rect 395308 -13680 395648 -13670
rect 395308 -13736 395385 -13680
rect 395441 -13736 395527 -13680
rect 395583 -13736 395648 -13680
rect 395308 -13822 395648 -13736
rect 395308 -13878 395385 -13822
rect 395441 -13878 395527 -13822
rect 395583 -13878 395648 -13822
rect 395308 -13964 395648 -13878
rect 395308 -14020 395385 -13964
rect 395441 -14020 395527 -13964
rect 395583 -14020 395648 -13964
rect 395308 -14106 395648 -14020
rect 395308 -14162 395385 -14106
rect 395441 -14162 395527 -14106
rect 395583 -14162 395648 -14106
rect 395308 -14248 395648 -14162
rect 395308 -14304 395385 -14248
rect 395441 -14304 395527 -14248
rect 395583 -14304 395648 -14248
rect 395308 -14390 395648 -14304
rect 395308 -14446 395385 -14390
rect 395441 -14446 395527 -14390
rect 395583 -14446 395648 -14390
rect 395308 -14532 395648 -14446
rect 395308 -14588 395385 -14532
rect 395441 -14588 395527 -14532
rect 395583 -14588 395648 -14532
rect 395308 -14674 395648 -14588
rect 395308 -14730 395385 -14674
rect 395441 -14730 395527 -14674
rect 395583 -14730 395648 -14674
rect 395308 -14816 395648 -14730
rect 395308 -14872 395385 -14816
rect 395441 -14872 395527 -14816
rect 395583 -14872 395648 -14816
rect 395308 -14958 395648 -14872
rect 395308 -15014 395385 -14958
rect 395441 -15014 395527 -14958
rect 395583 -15014 395648 -14958
rect 395308 -15100 395648 -15014
rect 395308 -15156 395385 -15100
rect 395441 -15156 395527 -15100
rect 395583 -15156 395648 -15100
rect 395308 -15242 395648 -15156
rect 395308 -15298 395385 -15242
rect 395441 -15298 395527 -15242
rect 395583 -15298 395648 -15242
rect 395308 -15384 395648 -15298
rect 395308 -15440 395385 -15384
rect 395441 -15440 395527 -15384
rect 395583 -15440 395648 -15384
rect 395308 -15526 395648 -15440
rect 395308 -15582 395385 -15526
rect 395441 -15582 395527 -15526
rect 395583 -15582 395648 -15526
rect 395308 -15668 395648 -15582
rect 395308 -15724 395385 -15668
rect 395441 -15724 395527 -15668
rect 395583 -15724 395648 -15668
rect 395308 -15810 395648 -15724
rect 395308 -15866 395385 -15810
rect 395441 -15866 395527 -15810
rect 395583 -15866 395648 -15810
rect 395308 -15952 395648 -15866
rect 395308 -16008 395385 -15952
rect 395441 -16008 395527 -15952
rect 395583 -16008 395648 -15952
rect 395308 -16094 395648 -16008
rect 395308 -16150 395385 -16094
rect 395441 -16150 395527 -16094
rect 395583 -16150 395648 -16094
rect 395308 -16236 395648 -16150
rect 395308 -16292 395385 -16236
rect 395441 -16292 395527 -16236
rect 395583 -16292 395648 -16236
rect 395308 -16378 395648 -16292
rect 395308 -16434 395385 -16378
rect 395441 -16434 395527 -16378
rect 395583 -16434 395648 -16378
rect 395308 -16520 395648 -16434
rect 395308 -16576 395385 -16520
rect 395441 -16576 395527 -16520
rect 395583 -16576 395648 -16520
rect 395308 -16662 395648 -16576
rect 395308 -16718 395385 -16662
rect 395441 -16718 395527 -16662
rect 395583 -16718 395648 -16662
rect 395308 -16804 395648 -16718
rect 395308 -16860 395385 -16804
rect 395441 -16860 395527 -16804
rect 395583 -16860 395648 -16804
rect 395308 -16946 395648 -16860
rect 395308 -17002 395385 -16946
rect 395441 -17002 395527 -16946
rect 395583 -17002 395648 -16946
rect 395308 -17088 395648 -17002
rect 395308 -17144 395385 -17088
rect 395441 -17144 395527 -17088
rect 395583 -17144 395648 -17088
rect 395308 -17230 395648 -17144
rect 395308 -17286 395385 -17230
rect 395441 -17286 395527 -17230
rect 395583 -17286 395648 -17230
rect 395308 -17372 395648 -17286
rect 395308 -17428 395385 -17372
rect 395441 -17428 395527 -17372
rect 395583 -17428 395648 -17372
rect 395308 -17514 395648 -17428
rect 395308 -17570 395385 -17514
rect 395441 -17570 395527 -17514
rect 395583 -17570 395648 -17514
rect 395308 -17656 395648 -17570
rect 395308 -17712 395385 -17656
rect 395441 -17712 395527 -17656
rect 395583 -17712 395648 -17656
rect 395308 -17798 395648 -17712
rect 395308 -17854 395385 -17798
rect 395441 -17854 395527 -17798
rect 395583 -17854 395648 -17798
rect 395308 -17940 395648 -17854
rect 395308 -17996 395385 -17940
rect 395441 -17996 395527 -17940
rect 395583 -17996 395648 -17940
rect 395308 -18082 395648 -17996
rect 395308 -18138 395385 -18082
rect 395441 -18138 395527 -18082
rect 395583 -18138 395648 -18082
rect 395308 -18224 395648 -18138
rect 395308 -18280 395385 -18224
rect 395441 -18280 395527 -18224
rect 395583 -18280 395648 -18224
rect 395308 -18366 395648 -18280
rect 395308 -18422 395385 -18366
rect 395441 -18422 395527 -18366
rect 395583 -18422 395648 -18366
rect 395308 -18508 395648 -18422
rect 395308 -18564 395385 -18508
rect 395441 -18564 395527 -18508
rect 395583 -18564 395648 -18508
rect 395308 -18650 395648 -18564
rect 395308 -18706 395385 -18650
rect 395441 -18706 395527 -18650
rect 395583 -18706 395648 -18650
rect 395308 -18792 395648 -18706
rect 395308 -18848 395385 -18792
rect 395441 -18848 395527 -18792
rect 395583 -18848 395648 -18792
rect 395308 -18934 395648 -18848
rect 395308 -18990 395385 -18934
rect 395441 -18990 395527 -18934
rect 395583 -18990 395648 -18934
rect 395308 -19076 395648 -18990
rect 395308 -19132 395385 -19076
rect 395441 -19132 395527 -19076
rect 395583 -19132 395648 -19076
rect 395308 -19218 395648 -19132
rect 395308 -19274 395385 -19218
rect 395441 -19274 395527 -19218
rect 395583 -19274 395648 -19218
rect 395308 -19360 395648 -19274
rect 395308 -19416 395385 -19360
rect 395441 -19416 395527 -19360
rect 395583 -19416 395648 -19360
rect 395308 -19502 395648 -19416
rect 395308 -19558 395385 -19502
rect 395441 -19558 395527 -19502
rect 395583 -19558 395648 -19502
rect 395308 -19644 395648 -19558
rect 395308 -19700 395385 -19644
rect 395441 -19700 395527 -19644
rect 395583 -19700 395648 -19644
rect 395308 -19786 395648 -19700
rect 395308 -19842 395385 -19786
rect 395441 -19842 395527 -19786
rect 395583 -19842 395648 -19786
rect 395308 -19928 395648 -19842
rect 395308 -19984 395385 -19928
rect 395441 -19984 395527 -19928
rect 395583 -19984 395648 -19928
rect 395308 -20070 395648 -19984
rect 395308 -20126 395385 -20070
rect 395441 -20126 395527 -20070
rect 395583 -20126 395648 -20070
rect 395308 -20212 395648 -20126
rect 395308 -20268 395385 -20212
rect 395441 -20268 395527 -20212
rect 395583 -20268 395648 -20212
rect 395308 -20354 395648 -20268
rect 395308 -20410 395385 -20354
rect 395441 -20410 395527 -20354
rect 395583 -20410 395648 -20354
rect 395308 -20496 395648 -20410
rect 395308 -20552 395385 -20496
rect 395441 -20552 395527 -20496
rect 395583 -20552 395648 -20496
rect 395308 -20638 395648 -20552
rect 395308 -20694 395385 -20638
rect 395441 -20694 395527 -20638
rect 395583 -20694 395648 -20638
rect 395308 -20780 395648 -20694
rect 395308 -20836 395385 -20780
rect 395441 -20836 395527 -20780
rect 395583 -20836 395648 -20780
rect 395308 -20922 395648 -20836
rect 395308 -20978 395385 -20922
rect 395441 -20978 395527 -20922
rect 395583 -20978 395648 -20922
rect 395308 -21064 395648 -20978
rect 395308 -21120 395385 -21064
rect 395441 -21120 395527 -21064
rect 395583 -21120 395648 -21064
rect 395308 -21206 395648 -21120
rect 395308 -21262 395385 -21206
rect 395441 -21262 395527 -21206
rect 395583 -21262 395648 -21206
rect 395308 -21348 395648 -21262
rect 395308 -21404 395385 -21348
rect 395441 -21404 395527 -21348
rect 395583 -21404 395648 -21348
rect 395308 -21490 395648 -21404
rect 395308 -21546 395385 -21490
rect 395441 -21546 395527 -21490
rect 395583 -21546 395648 -21490
rect 395308 -21632 395648 -21546
rect 395308 -21688 395385 -21632
rect 395441 -21688 395527 -21632
rect 395583 -21688 395648 -21632
rect 395308 -21774 395648 -21688
rect 395308 -21830 395385 -21774
rect 395441 -21830 395527 -21774
rect 395583 -21830 395648 -21774
rect 395308 -21916 395648 -21830
rect 395308 -21972 395385 -21916
rect 395441 -21972 395527 -21916
rect 395583 -21972 395648 -21916
rect 395308 -22058 395648 -21972
rect 395308 -22114 395385 -22058
rect 395441 -22114 395527 -22058
rect 395583 -22114 395648 -22058
rect 395308 -22200 395648 -22114
rect 395308 -22256 395385 -22200
rect 395441 -22256 395527 -22200
rect 395583 -22256 395648 -22200
rect 395308 -22342 395648 -22256
rect 395308 -22398 395385 -22342
rect 395441 -22398 395527 -22342
rect 395583 -22398 395648 -22342
rect 395308 -22484 395648 -22398
rect 395308 -22540 395385 -22484
rect 395441 -22540 395527 -22484
rect 395583 -22540 395648 -22484
rect 395308 -22626 395648 -22540
rect 395308 -22682 395385 -22626
rect 395441 -22682 395527 -22626
rect 395583 -22682 395648 -22626
rect 395308 -22768 395648 -22682
rect 395308 -22824 395385 -22768
rect 395441 -22824 395527 -22768
rect 395583 -22824 395648 -22768
rect 395308 -22910 395648 -22824
rect 395308 -22966 395385 -22910
rect 395441 -22966 395527 -22910
rect 395583 -22966 395648 -22910
rect 395308 -23052 395648 -22966
rect 395308 -23108 395385 -23052
rect 395441 -23108 395527 -23052
rect 395583 -23108 395648 -23052
rect 395308 -23194 395648 -23108
rect 395308 -23250 395385 -23194
rect 395441 -23250 395527 -23194
rect 395583 -23250 395648 -23194
rect 395308 -23336 395648 -23250
rect 395308 -23392 395385 -23336
rect 395441 -23392 395527 -23336
rect 395583 -23392 395648 -23336
rect 395308 -23478 395648 -23392
rect 395308 -23534 395385 -23478
rect 395441 -23534 395527 -23478
rect 395583 -23534 395648 -23478
rect 395308 -23620 395648 -23534
rect 395308 -23676 395385 -23620
rect 395441 -23676 395527 -23620
rect 395583 -23676 395648 -23620
rect 395308 -23762 395648 -23676
rect 395308 -23818 395385 -23762
rect 395441 -23818 395527 -23762
rect 395583 -23818 395648 -23762
rect 395308 -23904 395648 -23818
rect 395308 -23960 395385 -23904
rect 395441 -23960 395527 -23904
rect 395583 -23960 395648 -23904
rect 395308 -24046 395648 -23960
rect 395308 -24102 395385 -24046
rect 395441 -24102 395527 -24046
rect 395583 -24102 395648 -24046
rect 395308 -24188 395648 -24102
rect 395308 -24244 395385 -24188
rect 395441 -24244 395527 -24188
rect 395583 -24244 395648 -24188
rect 395308 -24330 395648 -24244
rect 395308 -24386 395385 -24330
rect 395441 -24386 395527 -24330
rect 395583 -24386 395648 -24330
rect 395308 -24472 395648 -24386
rect 395308 -24528 395385 -24472
rect 395441 -24528 395527 -24472
rect 395583 -24528 395648 -24472
rect 395308 -24614 395648 -24528
rect 395308 -24670 395385 -24614
rect 395441 -24670 395527 -24614
rect 395583 -24670 395648 -24614
rect 395308 -24756 395648 -24670
rect 395308 -24812 395385 -24756
rect 395441 -24812 395527 -24756
rect 395583 -24812 395648 -24756
rect 395308 -24898 395648 -24812
rect 395308 -24954 395385 -24898
rect 395441 -24954 395527 -24898
rect 395583 -24954 395648 -24898
rect 395308 -25040 395648 -24954
rect 395308 -25096 395385 -25040
rect 395441 -25096 395527 -25040
rect 395583 -25096 395648 -25040
rect 395308 -25182 395648 -25096
rect 395308 -25238 395385 -25182
rect 395441 -25238 395527 -25182
rect 395583 -25238 395648 -25182
rect 395308 -25324 395648 -25238
rect 395308 -25380 395385 -25324
rect 395441 -25380 395527 -25324
rect 395583 -25380 395648 -25324
rect 395308 -25466 395648 -25380
rect 395308 -25522 395385 -25466
rect 395441 -25522 395527 -25466
rect 395583 -25522 395648 -25466
rect 395308 -25532 395648 -25522
rect 395708 -13680 396048 -13670
rect 395708 -13736 395779 -13680
rect 395835 -13736 395921 -13680
rect 395977 -13736 396048 -13680
rect 395708 -13822 396048 -13736
rect 395708 -13878 395779 -13822
rect 395835 -13878 395921 -13822
rect 395977 -13878 396048 -13822
rect 395708 -13964 396048 -13878
rect 395708 -14020 395779 -13964
rect 395835 -14020 395921 -13964
rect 395977 -14020 396048 -13964
rect 395708 -14106 396048 -14020
rect 395708 -14162 395779 -14106
rect 395835 -14162 395921 -14106
rect 395977 -14162 396048 -14106
rect 395708 -14248 396048 -14162
rect 395708 -14304 395779 -14248
rect 395835 -14304 395921 -14248
rect 395977 -14304 396048 -14248
rect 395708 -14390 396048 -14304
rect 395708 -14446 395779 -14390
rect 395835 -14446 395921 -14390
rect 395977 -14446 396048 -14390
rect 395708 -14532 396048 -14446
rect 395708 -14588 395779 -14532
rect 395835 -14588 395921 -14532
rect 395977 -14588 396048 -14532
rect 395708 -14674 396048 -14588
rect 395708 -14730 395779 -14674
rect 395835 -14730 395921 -14674
rect 395977 -14730 396048 -14674
rect 395708 -14816 396048 -14730
rect 395708 -14872 395779 -14816
rect 395835 -14872 395921 -14816
rect 395977 -14872 396048 -14816
rect 395708 -14958 396048 -14872
rect 395708 -15014 395779 -14958
rect 395835 -15014 395921 -14958
rect 395977 -15014 396048 -14958
rect 395708 -15100 396048 -15014
rect 395708 -15156 395779 -15100
rect 395835 -15156 395921 -15100
rect 395977 -15156 396048 -15100
rect 395708 -15242 396048 -15156
rect 395708 -15298 395779 -15242
rect 395835 -15298 395921 -15242
rect 395977 -15298 396048 -15242
rect 395708 -15384 396048 -15298
rect 395708 -15440 395779 -15384
rect 395835 -15440 395921 -15384
rect 395977 -15440 396048 -15384
rect 395708 -15526 396048 -15440
rect 395708 -15582 395779 -15526
rect 395835 -15582 395921 -15526
rect 395977 -15582 396048 -15526
rect 395708 -15668 396048 -15582
rect 395708 -15724 395779 -15668
rect 395835 -15724 395921 -15668
rect 395977 -15724 396048 -15668
rect 395708 -15810 396048 -15724
rect 395708 -15866 395779 -15810
rect 395835 -15866 395921 -15810
rect 395977 -15866 396048 -15810
rect 395708 -15952 396048 -15866
rect 395708 -16008 395779 -15952
rect 395835 -16008 395921 -15952
rect 395977 -16008 396048 -15952
rect 395708 -16094 396048 -16008
rect 395708 -16150 395779 -16094
rect 395835 -16150 395921 -16094
rect 395977 -16150 396048 -16094
rect 395708 -16236 396048 -16150
rect 395708 -16292 395779 -16236
rect 395835 -16292 395921 -16236
rect 395977 -16292 396048 -16236
rect 395708 -16378 396048 -16292
rect 395708 -16434 395779 -16378
rect 395835 -16434 395921 -16378
rect 395977 -16434 396048 -16378
rect 395708 -16520 396048 -16434
rect 395708 -16576 395779 -16520
rect 395835 -16576 395921 -16520
rect 395977 -16576 396048 -16520
rect 395708 -16662 396048 -16576
rect 395708 -16718 395779 -16662
rect 395835 -16718 395921 -16662
rect 395977 -16718 396048 -16662
rect 395708 -16804 396048 -16718
rect 395708 -16860 395779 -16804
rect 395835 -16860 395921 -16804
rect 395977 -16860 396048 -16804
rect 395708 -16946 396048 -16860
rect 395708 -17002 395779 -16946
rect 395835 -17002 395921 -16946
rect 395977 -17002 396048 -16946
rect 395708 -17088 396048 -17002
rect 395708 -17144 395779 -17088
rect 395835 -17144 395921 -17088
rect 395977 -17144 396048 -17088
rect 395708 -17230 396048 -17144
rect 395708 -17286 395779 -17230
rect 395835 -17286 395921 -17230
rect 395977 -17286 396048 -17230
rect 395708 -17372 396048 -17286
rect 395708 -17428 395779 -17372
rect 395835 -17428 395921 -17372
rect 395977 -17428 396048 -17372
rect 395708 -17514 396048 -17428
rect 395708 -17570 395779 -17514
rect 395835 -17570 395921 -17514
rect 395977 -17570 396048 -17514
rect 395708 -17656 396048 -17570
rect 395708 -17712 395779 -17656
rect 395835 -17712 395921 -17656
rect 395977 -17712 396048 -17656
rect 395708 -17798 396048 -17712
rect 395708 -17854 395779 -17798
rect 395835 -17854 395921 -17798
rect 395977 -17854 396048 -17798
rect 395708 -17940 396048 -17854
rect 395708 -17996 395779 -17940
rect 395835 -17996 395921 -17940
rect 395977 -17996 396048 -17940
rect 395708 -18082 396048 -17996
rect 395708 -18138 395779 -18082
rect 395835 -18138 395921 -18082
rect 395977 -18138 396048 -18082
rect 395708 -18224 396048 -18138
rect 395708 -18280 395779 -18224
rect 395835 -18280 395921 -18224
rect 395977 -18280 396048 -18224
rect 395708 -18366 396048 -18280
rect 395708 -18422 395779 -18366
rect 395835 -18422 395921 -18366
rect 395977 -18422 396048 -18366
rect 395708 -18508 396048 -18422
rect 395708 -18564 395779 -18508
rect 395835 -18564 395921 -18508
rect 395977 -18564 396048 -18508
rect 395708 -18650 396048 -18564
rect 395708 -18706 395779 -18650
rect 395835 -18706 395921 -18650
rect 395977 -18706 396048 -18650
rect 395708 -18792 396048 -18706
rect 395708 -18848 395779 -18792
rect 395835 -18848 395921 -18792
rect 395977 -18848 396048 -18792
rect 395708 -18934 396048 -18848
rect 395708 -18990 395779 -18934
rect 395835 -18990 395921 -18934
rect 395977 -18990 396048 -18934
rect 395708 -19076 396048 -18990
rect 395708 -19132 395779 -19076
rect 395835 -19132 395921 -19076
rect 395977 -19132 396048 -19076
rect 395708 -19218 396048 -19132
rect 395708 -19274 395779 -19218
rect 395835 -19274 395921 -19218
rect 395977 -19274 396048 -19218
rect 395708 -19360 396048 -19274
rect 395708 -19416 395779 -19360
rect 395835 -19416 395921 -19360
rect 395977 -19416 396048 -19360
rect 395708 -19502 396048 -19416
rect 395708 -19558 395779 -19502
rect 395835 -19558 395921 -19502
rect 395977 -19558 396048 -19502
rect 395708 -19644 396048 -19558
rect 395708 -19700 395779 -19644
rect 395835 -19700 395921 -19644
rect 395977 -19700 396048 -19644
rect 395708 -19786 396048 -19700
rect 395708 -19842 395779 -19786
rect 395835 -19842 395921 -19786
rect 395977 -19842 396048 -19786
rect 395708 -19928 396048 -19842
rect 395708 -19984 395779 -19928
rect 395835 -19984 395921 -19928
rect 395977 -19984 396048 -19928
rect 395708 -20070 396048 -19984
rect 395708 -20126 395779 -20070
rect 395835 -20126 395921 -20070
rect 395977 -20126 396048 -20070
rect 395708 -20212 396048 -20126
rect 395708 -20268 395779 -20212
rect 395835 -20268 395921 -20212
rect 395977 -20268 396048 -20212
rect 395708 -20354 396048 -20268
rect 395708 -20410 395779 -20354
rect 395835 -20410 395921 -20354
rect 395977 -20410 396048 -20354
rect 395708 -20496 396048 -20410
rect 395708 -20552 395779 -20496
rect 395835 -20552 395921 -20496
rect 395977 -20552 396048 -20496
rect 395708 -20638 396048 -20552
rect 395708 -20694 395779 -20638
rect 395835 -20694 395921 -20638
rect 395977 -20694 396048 -20638
rect 395708 -20780 396048 -20694
rect 395708 -20836 395779 -20780
rect 395835 -20836 395921 -20780
rect 395977 -20836 396048 -20780
rect 395708 -20922 396048 -20836
rect 395708 -20978 395779 -20922
rect 395835 -20978 395921 -20922
rect 395977 -20978 396048 -20922
rect 395708 -21064 396048 -20978
rect 395708 -21120 395779 -21064
rect 395835 -21120 395921 -21064
rect 395977 -21120 396048 -21064
rect 395708 -21206 396048 -21120
rect 395708 -21262 395779 -21206
rect 395835 -21262 395921 -21206
rect 395977 -21262 396048 -21206
rect 395708 -21348 396048 -21262
rect 395708 -21404 395779 -21348
rect 395835 -21404 395921 -21348
rect 395977 -21404 396048 -21348
rect 395708 -21490 396048 -21404
rect 395708 -21546 395779 -21490
rect 395835 -21546 395921 -21490
rect 395977 -21546 396048 -21490
rect 395708 -21632 396048 -21546
rect 395708 -21688 395779 -21632
rect 395835 -21688 395921 -21632
rect 395977 -21688 396048 -21632
rect 395708 -21774 396048 -21688
rect 395708 -21830 395779 -21774
rect 395835 -21830 395921 -21774
rect 395977 -21830 396048 -21774
rect 395708 -21916 396048 -21830
rect 395708 -21972 395779 -21916
rect 395835 -21972 395921 -21916
rect 395977 -21972 396048 -21916
rect 395708 -22058 396048 -21972
rect 395708 -22114 395779 -22058
rect 395835 -22114 395921 -22058
rect 395977 -22114 396048 -22058
rect 395708 -22200 396048 -22114
rect 395708 -22256 395779 -22200
rect 395835 -22256 395921 -22200
rect 395977 -22256 396048 -22200
rect 395708 -22342 396048 -22256
rect 395708 -22398 395779 -22342
rect 395835 -22398 395921 -22342
rect 395977 -22398 396048 -22342
rect 395708 -22484 396048 -22398
rect 395708 -22540 395779 -22484
rect 395835 -22540 395921 -22484
rect 395977 -22540 396048 -22484
rect 395708 -22626 396048 -22540
rect 395708 -22682 395779 -22626
rect 395835 -22682 395921 -22626
rect 395977 -22682 396048 -22626
rect 395708 -22768 396048 -22682
rect 395708 -22824 395779 -22768
rect 395835 -22824 395921 -22768
rect 395977 -22824 396048 -22768
rect 395708 -22910 396048 -22824
rect 395708 -22966 395779 -22910
rect 395835 -22966 395921 -22910
rect 395977 -22966 396048 -22910
rect 395708 -23052 396048 -22966
rect 395708 -23108 395779 -23052
rect 395835 -23108 395921 -23052
rect 395977 -23108 396048 -23052
rect 395708 -23194 396048 -23108
rect 395708 -23250 395779 -23194
rect 395835 -23250 395921 -23194
rect 395977 -23250 396048 -23194
rect 395708 -23336 396048 -23250
rect 395708 -23392 395779 -23336
rect 395835 -23392 395921 -23336
rect 395977 -23392 396048 -23336
rect 395708 -23478 396048 -23392
rect 395708 -23534 395779 -23478
rect 395835 -23534 395921 -23478
rect 395977 -23534 396048 -23478
rect 395708 -23620 396048 -23534
rect 395708 -23676 395779 -23620
rect 395835 -23676 395921 -23620
rect 395977 -23676 396048 -23620
rect 395708 -23762 396048 -23676
rect 395708 -23818 395779 -23762
rect 395835 -23818 395921 -23762
rect 395977 -23818 396048 -23762
rect 395708 -23904 396048 -23818
rect 395708 -23960 395779 -23904
rect 395835 -23960 395921 -23904
rect 395977 -23960 396048 -23904
rect 395708 -24046 396048 -23960
rect 395708 -24102 395779 -24046
rect 395835 -24102 395921 -24046
rect 395977 -24102 396048 -24046
rect 395708 -24188 396048 -24102
rect 395708 -24244 395779 -24188
rect 395835 -24244 395921 -24188
rect 395977 -24244 396048 -24188
rect 395708 -24330 396048 -24244
rect 395708 -24386 395779 -24330
rect 395835 -24386 395921 -24330
rect 395977 -24386 396048 -24330
rect 395708 -24472 396048 -24386
rect 395708 -24528 395779 -24472
rect 395835 -24528 395921 -24472
rect 395977 -24528 396048 -24472
rect 395708 -24614 396048 -24528
rect 395708 -24670 395779 -24614
rect 395835 -24670 395921 -24614
rect 395977 -24670 396048 -24614
rect 395708 -24756 396048 -24670
rect 395708 -24812 395779 -24756
rect 395835 -24812 395921 -24756
rect 395977 -24812 396048 -24756
rect 395708 -24898 396048 -24812
rect 395708 -24954 395779 -24898
rect 395835 -24954 395921 -24898
rect 395977 -24954 396048 -24898
rect 395708 -25040 396048 -24954
rect 395708 -25096 395779 -25040
rect 395835 -25096 395921 -25040
rect 395977 -25096 396048 -25040
rect 395708 -25182 396048 -25096
rect 395708 -25238 395779 -25182
rect 395835 -25238 395921 -25182
rect 395977 -25238 396048 -25182
rect 395708 -25324 396048 -25238
rect 395708 -25380 395779 -25324
rect 395835 -25380 395921 -25324
rect 395977 -25380 396048 -25324
rect 395708 -25466 396048 -25380
rect 395708 -25522 395779 -25466
rect 395835 -25522 395921 -25466
rect 395977 -25522 396048 -25466
rect 395708 -25532 396048 -25522
rect 396108 -13680 396448 -13670
rect 396108 -13736 396180 -13680
rect 396236 -13736 396322 -13680
rect 396378 -13736 396448 -13680
rect 396108 -13822 396448 -13736
rect 396108 -13878 396180 -13822
rect 396236 -13878 396322 -13822
rect 396378 -13878 396448 -13822
rect 396108 -13964 396448 -13878
rect 396108 -14020 396180 -13964
rect 396236 -14020 396322 -13964
rect 396378 -14020 396448 -13964
rect 396108 -14106 396448 -14020
rect 396108 -14162 396180 -14106
rect 396236 -14162 396322 -14106
rect 396378 -14162 396448 -14106
rect 396108 -14248 396448 -14162
rect 396108 -14304 396180 -14248
rect 396236 -14304 396322 -14248
rect 396378 -14304 396448 -14248
rect 396108 -14390 396448 -14304
rect 396108 -14446 396180 -14390
rect 396236 -14446 396322 -14390
rect 396378 -14446 396448 -14390
rect 396108 -14532 396448 -14446
rect 396108 -14588 396180 -14532
rect 396236 -14588 396322 -14532
rect 396378 -14588 396448 -14532
rect 396108 -14674 396448 -14588
rect 396108 -14730 396180 -14674
rect 396236 -14730 396322 -14674
rect 396378 -14730 396448 -14674
rect 396108 -14816 396448 -14730
rect 396108 -14872 396180 -14816
rect 396236 -14872 396322 -14816
rect 396378 -14872 396448 -14816
rect 396108 -14958 396448 -14872
rect 396108 -15014 396180 -14958
rect 396236 -15014 396322 -14958
rect 396378 -15014 396448 -14958
rect 396108 -15100 396448 -15014
rect 396108 -15156 396180 -15100
rect 396236 -15156 396322 -15100
rect 396378 -15156 396448 -15100
rect 396108 -15242 396448 -15156
rect 396108 -15298 396180 -15242
rect 396236 -15298 396322 -15242
rect 396378 -15298 396448 -15242
rect 396108 -15384 396448 -15298
rect 396108 -15440 396180 -15384
rect 396236 -15440 396322 -15384
rect 396378 -15440 396448 -15384
rect 396108 -15526 396448 -15440
rect 396108 -15582 396180 -15526
rect 396236 -15582 396322 -15526
rect 396378 -15582 396448 -15526
rect 396108 -15668 396448 -15582
rect 396108 -15724 396180 -15668
rect 396236 -15724 396322 -15668
rect 396378 -15724 396448 -15668
rect 396108 -15810 396448 -15724
rect 396108 -15866 396180 -15810
rect 396236 -15866 396322 -15810
rect 396378 -15866 396448 -15810
rect 396108 -15952 396448 -15866
rect 396108 -16008 396180 -15952
rect 396236 -16008 396322 -15952
rect 396378 -16008 396448 -15952
rect 396108 -16094 396448 -16008
rect 396108 -16150 396180 -16094
rect 396236 -16150 396322 -16094
rect 396378 -16150 396448 -16094
rect 396108 -16236 396448 -16150
rect 396108 -16292 396180 -16236
rect 396236 -16292 396322 -16236
rect 396378 -16292 396448 -16236
rect 396108 -16378 396448 -16292
rect 396108 -16434 396180 -16378
rect 396236 -16434 396322 -16378
rect 396378 -16434 396448 -16378
rect 396108 -16520 396448 -16434
rect 396108 -16576 396180 -16520
rect 396236 -16576 396322 -16520
rect 396378 -16576 396448 -16520
rect 396108 -16662 396448 -16576
rect 396108 -16718 396180 -16662
rect 396236 -16718 396322 -16662
rect 396378 -16718 396448 -16662
rect 396108 -16804 396448 -16718
rect 396108 -16860 396180 -16804
rect 396236 -16860 396322 -16804
rect 396378 -16860 396448 -16804
rect 396108 -16946 396448 -16860
rect 396108 -17002 396180 -16946
rect 396236 -17002 396322 -16946
rect 396378 -17002 396448 -16946
rect 396108 -17088 396448 -17002
rect 396108 -17144 396180 -17088
rect 396236 -17144 396322 -17088
rect 396378 -17144 396448 -17088
rect 396108 -17230 396448 -17144
rect 396108 -17286 396180 -17230
rect 396236 -17286 396322 -17230
rect 396378 -17286 396448 -17230
rect 396108 -17372 396448 -17286
rect 396108 -17428 396180 -17372
rect 396236 -17428 396322 -17372
rect 396378 -17428 396448 -17372
rect 396108 -17514 396448 -17428
rect 396108 -17570 396180 -17514
rect 396236 -17570 396322 -17514
rect 396378 -17570 396448 -17514
rect 396108 -17656 396448 -17570
rect 396108 -17712 396180 -17656
rect 396236 -17712 396322 -17656
rect 396378 -17712 396448 -17656
rect 396108 -17798 396448 -17712
rect 396108 -17854 396180 -17798
rect 396236 -17854 396322 -17798
rect 396378 -17854 396448 -17798
rect 396108 -17940 396448 -17854
rect 396108 -17996 396180 -17940
rect 396236 -17996 396322 -17940
rect 396378 -17996 396448 -17940
rect 396108 -18082 396448 -17996
rect 396108 -18138 396180 -18082
rect 396236 -18138 396322 -18082
rect 396378 -18138 396448 -18082
rect 396108 -18224 396448 -18138
rect 396108 -18280 396180 -18224
rect 396236 -18280 396322 -18224
rect 396378 -18280 396448 -18224
rect 396108 -18366 396448 -18280
rect 396108 -18422 396180 -18366
rect 396236 -18422 396322 -18366
rect 396378 -18422 396448 -18366
rect 396108 -18508 396448 -18422
rect 396108 -18564 396180 -18508
rect 396236 -18564 396322 -18508
rect 396378 -18564 396448 -18508
rect 396108 -18650 396448 -18564
rect 396108 -18706 396180 -18650
rect 396236 -18706 396322 -18650
rect 396378 -18706 396448 -18650
rect 396108 -18792 396448 -18706
rect 396108 -18848 396180 -18792
rect 396236 -18848 396322 -18792
rect 396378 -18848 396448 -18792
rect 396108 -18934 396448 -18848
rect 396108 -18990 396180 -18934
rect 396236 -18990 396322 -18934
rect 396378 -18990 396448 -18934
rect 396108 -19076 396448 -18990
rect 396108 -19132 396180 -19076
rect 396236 -19132 396322 -19076
rect 396378 -19132 396448 -19076
rect 396108 -19218 396448 -19132
rect 396108 -19274 396180 -19218
rect 396236 -19274 396322 -19218
rect 396378 -19274 396448 -19218
rect 396108 -19360 396448 -19274
rect 396108 -19416 396180 -19360
rect 396236 -19416 396322 -19360
rect 396378 -19416 396448 -19360
rect 396108 -19502 396448 -19416
rect 396108 -19558 396180 -19502
rect 396236 -19558 396322 -19502
rect 396378 -19558 396448 -19502
rect 396108 -19644 396448 -19558
rect 396108 -19700 396180 -19644
rect 396236 -19700 396322 -19644
rect 396378 -19700 396448 -19644
rect 396108 -19786 396448 -19700
rect 396108 -19842 396180 -19786
rect 396236 -19842 396322 -19786
rect 396378 -19842 396448 -19786
rect 396108 -19928 396448 -19842
rect 396108 -19984 396180 -19928
rect 396236 -19984 396322 -19928
rect 396378 -19984 396448 -19928
rect 396108 -20070 396448 -19984
rect 396108 -20126 396180 -20070
rect 396236 -20126 396322 -20070
rect 396378 -20126 396448 -20070
rect 396108 -20212 396448 -20126
rect 396108 -20268 396180 -20212
rect 396236 -20268 396322 -20212
rect 396378 -20268 396448 -20212
rect 396108 -20354 396448 -20268
rect 396108 -20410 396180 -20354
rect 396236 -20410 396322 -20354
rect 396378 -20410 396448 -20354
rect 396108 -20496 396448 -20410
rect 396108 -20552 396180 -20496
rect 396236 -20552 396322 -20496
rect 396378 -20552 396448 -20496
rect 396108 -20638 396448 -20552
rect 396108 -20694 396180 -20638
rect 396236 -20694 396322 -20638
rect 396378 -20694 396448 -20638
rect 396108 -20780 396448 -20694
rect 396108 -20836 396180 -20780
rect 396236 -20836 396322 -20780
rect 396378 -20836 396448 -20780
rect 396108 -20922 396448 -20836
rect 396108 -20978 396180 -20922
rect 396236 -20978 396322 -20922
rect 396378 -20978 396448 -20922
rect 396108 -21064 396448 -20978
rect 396108 -21120 396180 -21064
rect 396236 -21120 396322 -21064
rect 396378 -21120 396448 -21064
rect 396108 -21206 396448 -21120
rect 396108 -21262 396180 -21206
rect 396236 -21262 396322 -21206
rect 396378 -21262 396448 -21206
rect 396108 -21348 396448 -21262
rect 396108 -21404 396180 -21348
rect 396236 -21404 396322 -21348
rect 396378 -21404 396448 -21348
rect 396108 -21490 396448 -21404
rect 396108 -21546 396180 -21490
rect 396236 -21546 396322 -21490
rect 396378 -21546 396448 -21490
rect 396108 -21632 396448 -21546
rect 396108 -21688 396180 -21632
rect 396236 -21688 396322 -21632
rect 396378 -21688 396448 -21632
rect 396108 -21774 396448 -21688
rect 396108 -21830 396180 -21774
rect 396236 -21830 396322 -21774
rect 396378 -21830 396448 -21774
rect 396108 -21916 396448 -21830
rect 396108 -21972 396180 -21916
rect 396236 -21972 396322 -21916
rect 396378 -21972 396448 -21916
rect 396108 -22058 396448 -21972
rect 396108 -22114 396180 -22058
rect 396236 -22114 396322 -22058
rect 396378 -22114 396448 -22058
rect 396108 -22200 396448 -22114
rect 396108 -22256 396180 -22200
rect 396236 -22256 396322 -22200
rect 396378 -22256 396448 -22200
rect 396108 -22342 396448 -22256
rect 396108 -22398 396180 -22342
rect 396236 -22398 396322 -22342
rect 396378 -22398 396448 -22342
rect 396108 -22484 396448 -22398
rect 396108 -22540 396180 -22484
rect 396236 -22540 396322 -22484
rect 396378 -22540 396448 -22484
rect 396108 -22626 396448 -22540
rect 396108 -22682 396180 -22626
rect 396236 -22682 396322 -22626
rect 396378 -22682 396448 -22626
rect 396108 -22768 396448 -22682
rect 396108 -22824 396180 -22768
rect 396236 -22824 396322 -22768
rect 396378 -22824 396448 -22768
rect 396108 -22910 396448 -22824
rect 396108 -22966 396180 -22910
rect 396236 -22966 396322 -22910
rect 396378 -22966 396448 -22910
rect 396108 -23052 396448 -22966
rect 396108 -23108 396180 -23052
rect 396236 -23108 396322 -23052
rect 396378 -23108 396448 -23052
rect 396108 -23194 396448 -23108
rect 396108 -23250 396180 -23194
rect 396236 -23250 396322 -23194
rect 396378 -23250 396448 -23194
rect 396108 -23336 396448 -23250
rect 396108 -23392 396180 -23336
rect 396236 -23392 396322 -23336
rect 396378 -23392 396448 -23336
rect 396108 -23478 396448 -23392
rect 396108 -23534 396180 -23478
rect 396236 -23534 396322 -23478
rect 396378 -23534 396448 -23478
rect 396108 -23620 396448 -23534
rect 396108 -23676 396180 -23620
rect 396236 -23676 396322 -23620
rect 396378 -23676 396448 -23620
rect 396108 -23762 396448 -23676
rect 396108 -23818 396180 -23762
rect 396236 -23818 396322 -23762
rect 396378 -23818 396448 -23762
rect 396108 -23904 396448 -23818
rect 396108 -23960 396180 -23904
rect 396236 -23960 396322 -23904
rect 396378 -23960 396448 -23904
rect 396108 -24046 396448 -23960
rect 396108 -24102 396180 -24046
rect 396236 -24102 396322 -24046
rect 396378 -24102 396448 -24046
rect 396108 -24188 396448 -24102
rect 396108 -24244 396180 -24188
rect 396236 -24244 396322 -24188
rect 396378 -24244 396448 -24188
rect 396108 -24330 396448 -24244
rect 396108 -24386 396180 -24330
rect 396236 -24386 396322 -24330
rect 396378 -24386 396448 -24330
rect 396108 -24472 396448 -24386
rect 396108 -24528 396180 -24472
rect 396236 -24528 396322 -24472
rect 396378 -24528 396448 -24472
rect 396108 -24614 396448 -24528
rect 396108 -24670 396180 -24614
rect 396236 -24670 396322 -24614
rect 396378 -24670 396448 -24614
rect 396108 -24756 396448 -24670
rect 396108 -24812 396180 -24756
rect 396236 -24812 396322 -24756
rect 396378 -24812 396448 -24756
rect 396108 -24898 396448 -24812
rect 396108 -24954 396180 -24898
rect 396236 -24954 396322 -24898
rect 396378 -24954 396448 -24898
rect 396108 -25040 396448 -24954
rect 396108 -25096 396180 -25040
rect 396236 -25096 396322 -25040
rect 396378 -25096 396448 -25040
rect 396108 -25182 396448 -25096
rect 396108 -25238 396180 -25182
rect 396236 -25238 396322 -25182
rect 396378 -25238 396448 -25182
rect 396108 -25324 396448 -25238
rect 396108 -25380 396180 -25324
rect 396236 -25380 396322 -25324
rect 396378 -25380 396448 -25324
rect 396108 -25466 396448 -25380
rect 396108 -25522 396180 -25466
rect 396236 -25522 396322 -25466
rect 396378 -25522 396448 -25466
rect 396108 -25532 396448 -25522
rect 396508 -13680 396848 -13670
rect 396508 -13736 396580 -13680
rect 396636 -13736 396722 -13680
rect 396778 -13736 396848 -13680
rect 396508 -13822 396848 -13736
rect 396508 -13878 396580 -13822
rect 396636 -13878 396722 -13822
rect 396778 -13878 396848 -13822
rect 396508 -13964 396848 -13878
rect 396508 -14020 396580 -13964
rect 396636 -14020 396722 -13964
rect 396778 -14020 396848 -13964
rect 396508 -14106 396848 -14020
rect 396508 -14162 396580 -14106
rect 396636 -14162 396722 -14106
rect 396778 -14162 396848 -14106
rect 396508 -14248 396848 -14162
rect 396508 -14304 396580 -14248
rect 396636 -14304 396722 -14248
rect 396778 -14304 396848 -14248
rect 396508 -14390 396848 -14304
rect 396508 -14446 396580 -14390
rect 396636 -14446 396722 -14390
rect 396778 -14446 396848 -14390
rect 396508 -14532 396848 -14446
rect 396508 -14588 396580 -14532
rect 396636 -14588 396722 -14532
rect 396778 -14588 396848 -14532
rect 396508 -14674 396848 -14588
rect 396508 -14730 396580 -14674
rect 396636 -14730 396722 -14674
rect 396778 -14730 396848 -14674
rect 396508 -14816 396848 -14730
rect 396508 -14872 396580 -14816
rect 396636 -14872 396722 -14816
rect 396778 -14872 396848 -14816
rect 396508 -14958 396848 -14872
rect 396508 -15014 396580 -14958
rect 396636 -15014 396722 -14958
rect 396778 -15014 396848 -14958
rect 396508 -15100 396848 -15014
rect 396508 -15156 396580 -15100
rect 396636 -15156 396722 -15100
rect 396778 -15156 396848 -15100
rect 396508 -15242 396848 -15156
rect 396508 -15298 396580 -15242
rect 396636 -15298 396722 -15242
rect 396778 -15298 396848 -15242
rect 396508 -15384 396848 -15298
rect 396508 -15440 396580 -15384
rect 396636 -15440 396722 -15384
rect 396778 -15440 396848 -15384
rect 396508 -15526 396848 -15440
rect 396508 -15582 396580 -15526
rect 396636 -15582 396722 -15526
rect 396778 -15582 396848 -15526
rect 396508 -15668 396848 -15582
rect 396508 -15724 396580 -15668
rect 396636 -15724 396722 -15668
rect 396778 -15724 396848 -15668
rect 396508 -15810 396848 -15724
rect 396508 -15866 396580 -15810
rect 396636 -15866 396722 -15810
rect 396778 -15866 396848 -15810
rect 396508 -15952 396848 -15866
rect 396508 -16008 396580 -15952
rect 396636 -16008 396722 -15952
rect 396778 -16008 396848 -15952
rect 396508 -16094 396848 -16008
rect 396508 -16150 396580 -16094
rect 396636 -16150 396722 -16094
rect 396778 -16150 396848 -16094
rect 396508 -16236 396848 -16150
rect 396508 -16292 396580 -16236
rect 396636 -16292 396722 -16236
rect 396778 -16292 396848 -16236
rect 396508 -16378 396848 -16292
rect 396508 -16434 396580 -16378
rect 396636 -16434 396722 -16378
rect 396778 -16434 396848 -16378
rect 396508 -16520 396848 -16434
rect 396508 -16576 396580 -16520
rect 396636 -16576 396722 -16520
rect 396778 -16576 396848 -16520
rect 396508 -16662 396848 -16576
rect 396508 -16718 396580 -16662
rect 396636 -16718 396722 -16662
rect 396778 -16718 396848 -16662
rect 396508 -16804 396848 -16718
rect 396508 -16860 396580 -16804
rect 396636 -16860 396722 -16804
rect 396778 -16860 396848 -16804
rect 396508 -16946 396848 -16860
rect 396508 -17002 396580 -16946
rect 396636 -17002 396722 -16946
rect 396778 -17002 396848 -16946
rect 396508 -17088 396848 -17002
rect 396508 -17144 396580 -17088
rect 396636 -17144 396722 -17088
rect 396778 -17144 396848 -17088
rect 396508 -17230 396848 -17144
rect 396508 -17286 396580 -17230
rect 396636 -17286 396722 -17230
rect 396778 -17286 396848 -17230
rect 396508 -17372 396848 -17286
rect 396508 -17428 396580 -17372
rect 396636 -17428 396722 -17372
rect 396778 -17428 396848 -17372
rect 396508 -17514 396848 -17428
rect 396508 -17570 396580 -17514
rect 396636 -17570 396722 -17514
rect 396778 -17570 396848 -17514
rect 396508 -17656 396848 -17570
rect 396508 -17712 396580 -17656
rect 396636 -17712 396722 -17656
rect 396778 -17712 396848 -17656
rect 396508 -17798 396848 -17712
rect 396508 -17854 396580 -17798
rect 396636 -17854 396722 -17798
rect 396778 -17854 396848 -17798
rect 396508 -17940 396848 -17854
rect 396508 -17996 396580 -17940
rect 396636 -17996 396722 -17940
rect 396778 -17996 396848 -17940
rect 396508 -18082 396848 -17996
rect 396508 -18138 396580 -18082
rect 396636 -18138 396722 -18082
rect 396778 -18138 396848 -18082
rect 396508 -18224 396848 -18138
rect 396508 -18280 396580 -18224
rect 396636 -18280 396722 -18224
rect 396778 -18280 396848 -18224
rect 396508 -18366 396848 -18280
rect 396508 -18422 396580 -18366
rect 396636 -18422 396722 -18366
rect 396778 -18422 396848 -18366
rect 396508 -18508 396848 -18422
rect 396508 -18564 396580 -18508
rect 396636 -18564 396722 -18508
rect 396778 -18564 396848 -18508
rect 396508 -18650 396848 -18564
rect 396508 -18706 396580 -18650
rect 396636 -18706 396722 -18650
rect 396778 -18706 396848 -18650
rect 396508 -18792 396848 -18706
rect 396508 -18848 396580 -18792
rect 396636 -18848 396722 -18792
rect 396778 -18848 396848 -18792
rect 396508 -18934 396848 -18848
rect 396508 -18990 396580 -18934
rect 396636 -18990 396722 -18934
rect 396778 -18990 396848 -18934
rect 396508 -19076 396848 -18990
rect 396508 -19132 396580 -19076
rect 396636 -19132 396722 -19076
rect 396778 -19132 396848 -19076
rect 396508 -19218 396848 -19132
rect 396508 -19274 396580 -19218
rect 396636 -19274 396722 -19218
rect 396778 -19274 396848 -19218
rect 396508 -19360 396848 -19274
rect 396508 -19416 396580 -19360
rect 396636 -19416 396722 -19360
rect 396778 -19416 396848 -19360
rect 396508 -19502 396848 -19416
rect 396508 -19558 396580 -19502
rect 396636 -19558 396722 -19502
rect 396778 -19558 396848 -19502
rect 396508 -19644 396848 -19558
rect 396508 -19700 396580 -19644
rect 396636 -19700 396722 -19644
rect 396778 -19700 396848 -19644
rect 396508 -19786 396848 -19700
rect 396508 -19842 396580 -19786
rect 396636 -19842 396722 -19786
rect 396778 -19842 396848 -19786
rect 396508 -19928 396848 -19842
rect 396508 -19984 396580 -19928
rect 396636 -19984 396722 -19928
rect 396778 -19984 396848 -19928
rect 396508 -20070 396848 -19984
rect 396508 -20126 396580 -20070
rect 396636 -20126 396722 -20070
rect 396778 -20126 396848 -20070
rect 396508 -20212 396848 -20126
rect 396508 -20268 396580 -20212
rect 396636 -20268 396722 -20212
rect 396778 -20268 396848 -20212
rect 396508 -20354 396848 -20268
rect 396508 -20410 396580 -20354
rect 396636 -20410 396722 -20354
rect 396778 -20410 396848 -20354
rect 396508 -20496 396848 -20410
rect 396508 -20552 396580 -20496
rect 396636 -20552 396722 -20496
rect 396778 -20552 396848 -20496
rect 396508 -20638 396848 -20552
rect 396508 -20694 396580 -20638
rect 396636 -20694 396722 -20638
rect 396778 -20694 396848 -20638
rect 396508 -20780 396848 -20694
rect 396508 -20836 396580 -20780
rect 396636 -20836 396722 -20780
rect 396778 -20836 396848 -20780
rect 396508 -20922 396848 -20836
rect 396508 -20978 396580 -20922
rect 396636 -20978 396722 -20922
rect 396778 -20978 396848 -20922
rect 396508 -21064 396848 -20978
rect 396508 -21120 396580 -21064
rect 396636 -21120 396722 -21064
rect 396778 -21120 396848 -21064
rect 396508 -21206 396848 -21120
rect 396508 -21262 396580 -21206
rect 396636 -21262 396722 -21206
rect 396778 -21262 396848 -21206
rect 396508 -21348 396848 -21262
rect 396508 -21404 396580 -21348
rect 396636 -21404 396722 -21348
rect 396778 -21404 396848 -21348
rect 396508 -21490 396848 -21404
rect 396508 -21546 396580 -21490
rect 396636 -21546 396722 -21490
rect 396778 -21546 396848 -21490
rect 396508 -21632 396848 -21546
rect 396508 -21688 396580 -21632
rect 396636 -21688 396722 -21632
rect 396778 -21688 396848 -21632
rect 396508 -21774 396848 -21688
rect 396508 -21830 396580 -21774
rect 396636 -21830 396722 -21774
rect 396778 -21830 396848 -21774
rect 396508 -21916 396848 -21830
rect 396508 -21972 396580 -21916
rect 396636 -21972 396722 -21916
rect 396778 -21972 396848 -21916
rect 396508 -22058 396848 -21972
rect 396508 -22114 396580 -22058
rect 396636 -22114 396722 -22058
rect 396778 -22114 396848 -22058
rect 396508 -22200 396848 -22114
rect 396508 -22256 396580 -22200
rect 396636 -22256 396722 -22200
rect 396778 -22256 396848 -22200
rect 396508 -22342 396848 -22256
rect 396508 -22398 396580 -22342
rect 396636 -22398 396722 -22342
rect 396778 -22398 396848 -22342
rect 396508 -22484 396848 -22398
rect 396508 -22540 396580 -22484
rect 396636 -22540 396722 -22484
rect 396778 -22540 396848 -22484
rect 396508 -22626 396848 -22540
rect 396508 -22682 396580 -22626
rect 396636 -22682 396722 -22626
rect 396778 -22682 396848 -22626
rect 396508 -22768 396848 -22682
rect 396508 -22824 396580 -22768
rect 396636 -22824 396722 -22768
rect 396778 -22824 396848 -22768
rect 396508 -22910 396848 -22824
rect 396508 -22966 396580 -22910
rect 396636 -22966 396722 -22910
rect 396778 -22966 396848 -22910
rect 396508 -23052 396848 -22966
rect 396508 -23108 396580 -23052
rect 396636 -23108 396722 -23052
rect 396778 -23108 396848 -23052
rect 396508 -23194 396848 -23108
rect 396508 -23250 396580 -23194
rect 396636 -23250 396722 -23194
rect 396778 -23250 396848 -23194
rect 396508 -23336 396848 -23250
rect 396508 -23392 396580 -23336
rect 396636 -23392 396722 -23336
rect 396778 -23392 396848 -23336
rect 396508 -23478 396848 -23392
rect 396508 -23534 396580 -23478
rect 396636 -23534 396722 -23478
rect 396778 -23534 396848 -23478
rect 396508 -23620 396848 -23534
rect 396508 -23676 396580 -23620
rect 396636 -23676 396722 -23620
rect 396778 -23676 396848 -23620
rect 396508 -23762 396848 -23676
rect 396508 -23818 396580 -23762
rect 396636 -23818 396722 -23762
rect 396778 -23818 396848 -23762
rect 396508 -23904 396848 -23818
rect 396508 -23960 396580 -23904
rect 396636 -23960 396722 -23904
rect 396778 -23960 396848 -23904
rect 396508 -24046 396848 -23960
rect 396508 -24102 396580 -24046
rect 396636 -24102 396722 -24046
rect 396778 -24102 396848 -24046
rect 396508 -24188 396848 -24102
rect 396508 -24244 396580 -24188
rect 396636 -24244 396722 -24188
rect 396778 -24244 396848 -24188
rect 396508 -24330 396848 -24244
rect 396508 -24386 396580 -24330
rect 396636 -24386 396722 -24330
rect 396778 -24386 396848 -24330
rect 396508 -24472 396848 -24386
rect 396508 -24528 396580 -24472
rect 396636 -24528 396722 -24472
rect 396778 -24528 396848 -24472
rect 396508 -24614 396848 -24528
rect 396508 -24670 396580 -24614
rect 396636 -24670 396722 -24614
rect 396778 -24670 396848 -24614
rect 396508 -24756 396848 -24670
rect 396508 -24812 396580 -24756
rect 396636 -24812 396722 -24756
rect 396778 -24812 396848 -24756
rect 396508 -24898 396848 -24812
rect 396508 -24954 396580 -24898
rect 396636 -24954 396722 -24898
rect 396778 -24954 396848 -24898
rect 396508 -25040 396848 -24954
rect 396508 -25096 396580 -25040
rect 396636 -25096 396722 -25040
rect 396778 -25096 396848 -25040
rect 396508 -25182 396848 -25096
rect 396508 -25238 396580 -25182
rect 396636 -25238 396722 -25182
rect 396778 -25238 396848 -25182
rect 396508 -25324 396848 -25238
rect 396508 -25380 396580 -25324
rect 396636 -25380 396722 -25324
rect 396778 -25380 396848 -25324
rect 396508 -25466 396848 -25380
rect 396508 -25522 396580 -25466
rect 396636 -25522 396722 -25466
rect 396778 -25522 396848 -25466
rect 396508 -25532 396848 -25522
rect 396908 -13680 397248 -13670
rect 396908 -13736 396977 -13680
rect 397033 -13736 397119 -13680
rect 397175 -13736 397248 -13680
rect 396908 -13822 397248 -13736
rect 396908 -13878 396977 -13822
rect 397033 -13878 397119 -13822
rect 397175 -13878 397248 -13822
rect 396908 -13964 397248 -13878
rect 396908 -14020 396977 -13964
rect 397033 -14020 397119 -13964
rect 397175 -14020 397248 -13964
rect 396908 -14106 397248 -14020
rect 396908 -14162 396977 -14106
rect 397033 -14162 397119 -14106
rect 397175 -14162 397248 -14106
rect 396908 -14248 397248 -14162
rect 396908 -14304 396977 -14248
rect 397033 -14304 397119 -14248
rect 397175 -14304 397248 -14248
rect 396908 -14390 397248 -14304
rect 396908 -14446 396977 -14390
rect 397033 -14446 397119 -14390
rect 397175 -14446 397248 -14390
rect 396908 -14532 397248 -14446
rect 396908 -14588 396977 -14532
rect 397033 -14588 397119 -14532
rect 397175 -14588 397248 -14532
rect 396908 -14674 397248 -14588
rect 396908 -14730 396977 -14674
rect 397033 -14730 397119 -14674
rect 397175 -14730 397248 -14674
rect 396908 -14816 397248 -14730
rect 396908 -14872 396977 -14816
rect 397033 -14872 397119 -14816
rect 397175 -14872 397248 -14816
rect 396908 -14958 397248 -14872
rect 396908 -15014 396977 -14958
rect 397033 -15014 397119 -14958
rect 397175 -15014 397248 -14958
rect 396908 -15100 397248 -15014
rect 396908 -15156 396977 -15100
rect 397033 -15156 397119 -15100
rect 397175 -15156 397248 -15100
rect 396908 -15242 397248 -15156
rect 396908 -15298 396977 -15242
rect 397033 -15298 397119 -15242
rect 397175 -15298 397248 -15242
rect 396908 -15384 397248 -15298
rect 396908 -15440 396977 -15384
rect 397033 -15440 397119 -15384
rect 397175 -15440 397248 -15384
rect 396908 -15526 397248 -15440
rect 396908 -15582 396977 -15526
rect 397033 -15582 397119 -15526
rect 397175 -15582 397248 -15526
rect 396908 -15668 397248 -15582
rect 396908 -15724 396977 -15668
rect 397033 -15724 397119 -15668
rect 397175 -15724 397248 -15668
rect 396908 -15810 397248 -15724
rect 396908 -15866 396977 -15810
rect 397033 -15866 397119 -15810
rect 397175 -15866 397248 -15810
rect 396908 -15952 397248 -15866
rect 396908 -16008 396977 -15952
rect 397033 -16008 397119 -15952
rect 397175 -16008 397248 -15952
rect 396908 -16094 397248 -16008
rect 396908 -16150 396977 -16094
rect 397033 -16150 397119 -16094
rect 397175 -16150 397248 -16094
rect 396908 -16236 397248 -16150
rect 396908 -16292 396977 -16236
rect 397033 -16292 397119 -16236
rect 397175 -16292 397248 -16236
rect 396908 -16378 397248 -16292
rect 396908 -16434 396977 -16378
rect 397033 -16434 397119 -16378
rect 397175 -16434 397248 -16378
rect 396908 -16520 397248 -16434
rect 396908 -16576 396977 -16520
rect 397033 -16576 397119 -16520
rect 397175 -16576 397248 -16520
rect 396908 -16662 397248 -16576
rect 396908 -16718 396977 -16662
rect 397033 -16718 397119 -16662
rect 397175 -16718 397248 -16662
rect 396908 -16804 397248 -16718
rect 396908 -16860 396977 -16804
rect 397033 -16860 397119 -16804
rect 397175 -16860 397248 -16804
rect 396908 -16946 397248 -16860
rect 396908 -17002 396977 -16946
rect 397033 -17002 397119 -16946
rect 397175 -17002 397248 -16946
rect 396908 -17088 397248 -17002
rect 396908 -17144 396977 -17088
rect 397033 -17144 397119 -17088
rect 397175 -17144 397248 -17088
rect 396908 -17230 397248 -17144
rect 396908 -17286 396977 -17230
rect 397033 -17286 397119 -17230
rect 397175 -17286 397248 -17230
rect 396908 -17372 397248 -17286
rect 396908 -17428 396977 -17372
rect 397033 -17428 397119 -17372
rect 397175 -17428 397248 -17372
rect 396908 -17514 397248 -17428
rect 396908 -17570 396977 -17514
rect 397033 -17570 397119 -17514
rect 397175 -17570 397248 -17514
rect 396908 -17656 397248 -17570
rect 396908 -17712 396977 -17656
rect 397033 -17712 397119 -17656
rect 397175 -17712 397248 -17656
rect 396908 -17798 397248 -17712
rect 396908 -17854 396977 -17798
rect 397033 -17854 397119 -17798
rect 397175 -17854 397248 -17798
rect 396908 -17940 397248 -17854
rect 396908 -17996 396977 -17940
rect 397033 -17996 397119 -17940
rect 397175 -17996 397248 -17940
rect 396908 -18082 397248 -17996
rect 396908 -18138 396977 -18082
rect 397033 -18138 397119 -18082
rect 397175 -18138 397248 -18082
rect 396908 -18224 397248 -18138
rect 396908 -18280 396977 -18224
rect 397033 -18280 397119 -18224
rect 397175 -18280 397248 -18224
rect 396908 -18366 397248 -18280
rect 396908 -18422 396977 -18366
rect 397033 -18422 397119 -18366
rect 397175 -18422 397248 -18366
rect 396908 -18508 397248 -18422
rect 396908 -18564 396977 -18508
rect 397033 -18564 397119 -18508
rect 397175 -18564 397248 -18508
rect 396908 -18650 397248 -18564
rect 396908 -18706 396977 -18650
rect 397033 -18706 397119 -18650
rect 397175 -18706 397248 -18650
rect 396908 -18792 397248 -18706
rect 396908 -18848 396977 -18792
rect 397033 -18848 397119 -18792
rect 397175 -18848 397248 -18792
rect 396908 -18934 397248 -18848
rect 396908 -18990 396977 -18934
rect 397033 -18990 397119 -18934
rect 397175 -18990 397248 -18934
rect 396908 -19076 397248 -18990
rect 396908 -19132 396977 -19076
rect 397033 -19132 397119 -19076
rect 397175 -19132 397248 -19076
rect 396908 -19218 397248 -19132
rect 396908 -19274 396977 -19218
rect 397033 -19274 397119 -19218
rect 397175 -19274 397248 -19218
rect 396908 -19360 397248 -19274
rect 396908 -19416 396977 -19360
rect 397033 -19416 397119 -19360
rect 397175 -19416 397248 -19360
rect 396908 -19502 397248 -19416
rect 396908 -19558 396977 -19502
rect 397033 -19558 397119 -19502
rect 397175 -19558 397248 -19502
rect 396908 -19644 397248 -19558
rect 396908 -19700 396977 -19644
rect 397033 -19700 397119 -19644
rect 397175 -19700 397248 -19644
rect 396908 -19786 397248 -19700
rect 396908 -19842 396977 -19786
rect 397033 -19842 397119 -19786
rect 397175 -19842 397248 -19786
rect 396908 -19928 397248 -19842
rect 396908 -19984 396977 -19928
rect 397033 -19984 397119 -19928
rect 397175 -19984 397248 -19928
rect 396908 -20070 397248 -19984
rect 396908 -20126 396977 -20070
rect 397033 -20126 397119 -20070
rect 397175 -20126 397248 -20070
rect 396908 -20212 397248 -20126
rect 396908 -20268 396977 -20212
rect 397033 -20268 397119 -20212
rect 397175 -20268 397248 -20212
rect 396908 -20354 397248 -20268
rect 396908 -20410 396977 -20354
rect 397033 -20410 397119 -20354
rect 397175 -20410 397248 -20354
rect 396908 -20496 397248 -20410
rect 396908 -20552 396977 -20496
rect 397033 -20552 397119 -20496
rect 397175 -20552 397248 -20496
rect 396908 -20638 397248 -20552
rect 396908 -20694 396977 -20638
rect 397033 -20694 397119 -20638
rect 397175 -20694 397248 -20638
rect 396908 -20780 397248 -20694
rect 396908 -20836 396977 -20780
rect 397033 -20836 397119 -20780
rect 397175 -20836 397248 -20780
rect 396908 -20922 397248 -20836
rect 396908 -20978 396977 -20922
rect 397033 -20978 397119 -20922
rect 397175 -20978 397248 -20922
rect 396908 -21064 397248 -20978
rect 396908 -21120 396977 -21064
rect 397033 -21120 397119 -21064
rect 397175 -21120 397248 -21064
rect 396908 -21206 397248 -21120
rect 396908 -21262 396977 -21206
rect 397033 -21262 397119 -21206
rect 397175 -21262 397248 -21206
rect 396908 -21348 397248 -21262
rect 396908 -21404 396977 -21348
rect 397033 -21404 397119 -21348
rect 397175 -21404 397248 -21348
rect 396908 -21490 397248 -21404
rect 396908 -21546 396977 -21490
rect 397033 -21546 397119 -21490
rect 397175 -21546 397248 -21490
rect 396908 -21632 397248 -21546
rect 396908 -21688 396977 -21632
rect 397033 -21688 397119 -21632
rect 397175 -21688 397248 -21632
rect 396908 -21774 397248 -21688
rect 396908 -21830 396977 -21774
rect 397033 -21830 397119 -21774
rect 397175 -21830 397248 -21774
rect 396908 -21916 397248 -21830
rect 396908 -21972 396977 -21916
rect 397033 -21972 397119 -21916
rect 397175 -21972 397248 -21916
rect 396908 -22058 397248 -21972
rect 396908 -22114 396977 -22058
rect 397033 -22114 397119 -22058
rect 397175 -22114 397248 -22058
rect 396908 -22200 397248 -22114
rect 396908 -22256 396977 -22200
rect 397033 -22256 397119 -22200
rect 397175 -22256 397248 -22200
rect 396908 -22342 397248 -22256
rect 396908 -22398 396977 -22342
rect 397033 -22398 397119 -22342
rect 397175 -22398 397248 -22342
rect 396908 -22484 397248 -22398
rect 396908 -22540 396977 -22484
rect 397033 -22540 397119 -22484
rect 397175 -22540 397248 -22484
rect 396908 -22626 397248 -22540
rect 396908 -22682 396977 -22626
rect 397033 -22682 397119 -22626
rect 397175 -22682 397248 -22626
rect 396908 -22768 397248 -22682
rect 396908 -22824 396977 -22768
rect 397033 -22824 397119 -22768
rect 397175 -22824 397248 -22768
rect 396908 -22910 397248 -22824
rect 396908 -22966 396977 -22910
rect 397033 -22966 397119 -22910
rect 397175 -22966 397248 -22910
rect 396908 -23052 397248 -22966
rect 396908 -23108 396977 -23052
rect 397033 -23108 397119 -23052
rect 397175 -23108 397248 -23052
rect 396908 -23194 397248 -23108
rect 396908 -23250 396977 -23194
rect 397033 -23250 397119 -23194
rect 397175 -23250 397248 -23194
rect 396908 -23336 397248 -23250
rect 396908 -23392 396977 -23336
rect 397033 -23392 397119 -23336
rect 397175 -23392 397248 -23336
rect 396908 -23478 397248 -23392
rect 396908 -23534 396977 -23478
rect 397033 -23534 397119 -23478
rect 397175 -23534 397248 -23478
rect 396908 -23620 397248 -23534
rect 396908 -23676 396977 -23620
rect 397033 -23676 397119 -23620
rect 397175 -23676 397248 -23620
rect 396908 -23762 397248 -23676
rect 396908 -23818 396977 -23762
rect 397033 -23818 397119 -23762
rect 397175 -23818 397248 -23762
rect 396908 -23904 397248 -23818
rect 396908 -23960 396977 -23904
rect 397033 -23960 397119 -23904
rect 397175 -23960 397248 -23904
rect 396908 -24046 397248 -23960
rect 396908 -24102 396977 -24046
rect 397033 -24102 397119 -24046
rect 397175 -24102 397248 -24046
rect 396908 -24188 397248 -24102
rect 396908 -24244 396977 -24188
rect 397033 -24244 397119 -24188
rect 397175 -24244 397248 -24188
rect 396908 -24330 397248 -24244
rect 396908 -24386 396977 -24330
rect 397033 -24386 397119 -24330
rect 397175 -24386 397248 -24330
rect 396908 -24472 397248 -24386
rect 396908 -24528 396977 -24472
rect 397033 -24528 397119 -24472
rect 397175 -24528 397248 -24472
rect 396908 -24614 397248 -24528
rect 396908 -24670 396977 -24614
rect 397033 -24670 397119 -24614
rect 397175 -24670 397248 -24614
rect 396908 -24756 397248 -24670
rect 396908 -24812 396977 -24756
rect 397033 -24812 397119 -24756
rect 397175 -24812 397248 -24756
rect 396908 -24898 397248 -24812
rect 396908 -24954 396977 -24898
rect 397033 -24954 397119 -24898
rect 397175 -24954 397248 -24898
rect 396908 -25040 397248 -24954
rect 396908 -25096 396977 -25040
rect 397033 -25096 397119 -25040
rect 397175 -25096 397248 -25040
rect 396908 -25182 397248 -25096
rect 396908 -25238 396977 -25182
rect 397033 -25238 397119 -25182
rect 397175 -25238 397248 -25182
rect 396908 -25324 397248 -25238
rect 396908 -25380 396977 -25324
rect 397033 -25380 397119 -25324
rect 397175 -25380 397248 -25324
rect 396908 -25466 397248 -25380
rect 396908 -25522 396977 -25466
rect 397033 -25522 397119 -25466
rect 397175 -25522 397248 -25466
rect 396908 -25532 397248 -25522
rect 397308 -13680 397648 -13670
rect 397308 -13736 397374 -13680
rect 397430 -13736 397516 -13680
rect 397572 -13736 397648 -13680
rect 397308 -13822 397648 -13736
rect 397308 -13878 397374 -13822
rect 397430 -13878 397516 -13822
rect 397572 -13878 397648 -13822
rect 397308 -13964 397648 -13878
rect 397308 -14020 397374 -13964
rect 397430 -14020 397516 -13964
rect 397572 -14020 397648 -13964
rect 397308 -14106 397648 -14020
rect 397308 -14162 397374 -14106
rect 397430 -14162 397516 -14106
rect 397572 -14162 397648 -14106
rect 397308 -14248 397648 -14162
rect 397308 -14304 397374 -14248
rect 397430 -14304 397516 -14248
rect 397572 -14304 397648 -14248
rect 397308 -14390 397648 -14304
rect 397308 -14446 397374 -14390
rect 397430 -14446 397516 -14390
rect 397572 -14446 397648 -14390
rect 397308 -14532 397648 -14446
rect 397308 -14588 397374 -14532
rect 397430 -14588 397516 -14532
rect 397572 -14588 397648 -14532
rect 397308 -14674 397648 -14588
rect 397308 -14730 397374 -14674
rect 397430 -14730 397516 -14674
rect 397572 -14730 397648 -14674
rect 397308 -14816 397648 -14730
rect 397308 -14872 397374 -14816
rect 397430 -14872 397516 -14816
rect 397572 -14872 397648 -14816
rect 397308 -14958 397648 -14872
rect 397308 -15014 397374 -14958
rect 397430 -15014 397516 -14958
rect 397572 -15014 397648 -14958
rect 397308 -15100 397648 -15014
rect 397308 -15156 397374 -15100
rect 397430 -15156 397516 -15100
rect 397572 -15156 397648 -15100
rect 397308 -15242 397648 -15156
rect 397308 -15298 397374 -15242
rect 397430 -15298 397516 -15242
rect 397572 -15298 397648 -15242
rect 397308 -15384 397648 -15298
rect 397308 -15440 397374 -15384
rect 397430 -15440 397516 -15384
rect 397572 -15440 397648 -15384
rect 397308 -15526 397648 -15440
rect 397308 -15582 397374 -15526
rect 397430 -15582 397516 -15526
rect 397572 -15582 397648 -15526
rect 397308 -15668 397648 -15582
rect 397308 -15724 397374 -15668
rect 397430 -15724 397516 -15668
rect 397572 -15724 397648 -15668
rect 397308 -15810 397648 -15724
rect 397308 -15866 397374 -15810
rect 397430 -15866 397516 -15810
rect 397572 -15866 397648 -15810
rect 397308 -15952 397648 -15866
rect 397308 -16008 397374 -15952
rect 397430 -16008 397516 -15952
rect 397572 -16008 397648 -15952
rect 397308 -16094 397648 -16008
rect 397308 -16150 397374 -16094
rect 397430 -16150 397516 -16094
rect 397572 -16150 397648 -16094
rect 397308 -16236 397648 -16150
rect 397308 -16292 397374 -16236
rect 397430 -16292 397516 -16236
rect 397572 -16292 397648 -16236
rect 397308 -16378 397648 -16292
rect 397308 -16434 397374 -16378
rect 397430 -16434 397516 -16378
rect 397572 -16434 397648 -16378
rect 397308 -16520 397648 -16434
rect 397308 -16576 397374 -16520
rect 397430 -16576 397516 -16520
rect 397572 -16576 397648 -16520
rect 397308 -16662 397648 -16576
rect 397308 -16718 397374 -16662
rect 397430 -16718 397516 -16662
rect 397572 -16718 397648 -16662
rect 397308 -16804 397648 -16718
rect 397308 -16860 397374 -16804
rect 397430 -16860 397516 -16804
rect 397572 -16860 397648 -16804
rect 397308 -16946 397648 -16860
rect 397308 -17002 397374 -16946
rect 397430 -17002 397516 -16946
rect 397572 -17002 397648 -16946
rect 397308 -17088 397648 -17002
rect 397308 -17144 397374 -17088
rect 397430 -17144 397516 -17088
rect 397572 -17144 397648 -17088
rect 397308 -17230 397648 -17144
rect 397308 -17286 397374 -17230
rect 397430 -17286 397516 -17230
rect 397572 -17286 397648 -17230
rect 397308 -17372 397648 -17286
rect 397308 -17428 397374 -17372
rect 397430 -17428 397516 -17372
rect 397572 -17428 397648 -17372
rect 397308 -17514 397648 -17428
rect 397308 -17570 397374 -17514
rect 397430 -17570 397516 -17514
rect 397572 -17570 397648 -17514
rect 397308 -17656 397648 -17570
rect 397308 -17712 397374 -17656
rect 397430 -17712 397516 -17656
rect 397572 -17712 397648 -17656
rect 397308 -17798 397648 -17712
rect 397308 -17854 397374 -17798
rect 397430 -17854 397516 -17798
rect 397572 -17854 397648 -17798
rect 397308 -17940 397648 -17854
rect 397308 -17996 397374 -17940
rect 397430 -17996 397516 -17940
rect 397572 -17996 397648 -17940
rect 397308 -18082 397648 -17996
rect 397308 -18138 397374 -18082
rect 397430 -18138 397516 -18082
rect 397572 -18138 397648 -18082
rect 397308 -18224 397648 -18138
rect 397308 -18280 397374 -18224
rect 397430 -18280 397516 -18224
rect 397572 -18280 397648 -18224
rect 397308 -18366 397648 -18280
rect 397308 -18422 397374 -18366
rect 397430 -18422 397516 -18366
rect 397572 -18422 397648 -18366
rect 397308 -18508 397648 -18422
rect 397308 -18564 397374 -18508
rect 397430 -18564 397516 -18508
rect 397572 -18564 397648 -18508
rect 397308 -18650 397648 -18564
rect 397308 -18706 397374 -18650
rect 397430 -18706 397516 -18650
rect 397572 -18706 397648 -18650
rect 397308 -18792 397648 -18706
rect 397308 -18848 397374 -18792
rect 397430 -18848 397516 -18792
rect 397572 -18848 397648 -18792
rect 397308 -18934 397648 -18848
rect 397308 -18990 397374 -18934
rect 397430 -18990 397516 -18934
rect 397572 -18990 397648 -18934
rect 397308 -19076 397648 -18990
rect 397308 -19132 397374 -19076
rect 397430 -19132 397516 -19076
rect 397572 -19132 397648 -19076
rect 397308 -19218 397648 -19132
rect 397308 -19274 397374 -19218
rect 397430 -19274 397516 -19218
rect 397572 -19274 397648 -19218
rect 397308 -19360 397648 -19274
rect 397308 -19416 397374 -19360
rect 397430 -19416 397516 -19360
rect 397572 -19416 397648 -19360
rect 397308 -19502 397648 -19416
rect 397308 -19558 397374 -19502
rect 397430 -19558 397516 -19502
rect 397572 -19558 397648 -19502
rect 397308 -19644 397648 -19558
rect 397308 -19700 397374 -19644
rect 397430 -19700 397516 -19644
rect 397572 -19700 397648 -19644
rect 397308 -19786 397648 -19700
rect 397308 -19842 397374 -19786
rect 397430 -19842 397516 -19786
rect 397572 -19842 397648 -19786
rect 397308 -19928 397648 -19842
rect 397308 -19984 397374 -19928
rect 397430 -19984 397516 -19928
rect 397572 -19984 397648 -19928
rect 397308 -20070 397648 -19984
rect 397308 -20126 397374 -20070
rect 397430 -20126 397516 -20070
rect 397572 -20126 397648 -20070
rect 397308 -20212 397648 -20126
rect 397308 -20268 397374 -20212
rect 397430 -20268 397516 -20212
rect 397572 -20268 397648 -20212
rect 397308 -20354 397648 -20268
rect 397308 -20410 397374 -20354
rect 397430 -20410 397516 -20354
rect 397572 -20410 397648 -20354
rect 397308 -20496 397648 -20410
rect 397308 -20552 397374 -20496
rect 397430 -20552 397516 -20496
rect 397572 -20552 397648 -20496
rect 397308 -20638 397648 -20552
rect 397308 -20694 397374 -20638
rect 397430 -20694 397516 -20638
rect 397572 -20694 397648 -20638
rect 397308 -20780 397648 -20694
rect 397308 -20836 397374 -20780
rect 397430 -20836 397516 -20780
rect 397572 -20836 397648 -20780
rect 397308 -20922 397648 -20836
rect 397308 -20978 397374 -20922
rect 397430 -20978 397516 -20922
rect 397572 -20978 397648 -20922
rect 397308 -21064 397648 -20978
rect 397308 -21120 397374 -21064
rect 397430 -21120 397516 -21064
rect 397572 -21120 397648 -21064
rect 397308 -21206 397648 -21120
rect 397308 -21262 397374 -21206
rect 397430 -21262 397516 -21206
rect 397572 -21262 397648 -21206
rect 397308 -21348 397648 -21262
rect 397308 -21404 397374 -21348
rect 397430 -21404 397516 -21348
rect 397572 -21404 397648 -21348
rect 397308 -21490 397648 -21404
rect 397308 -21546 397374 -21490
rect 397430 -21546 397516 -21490
rect 397572 -21546 397648 -21490
rect 397308 -21632 397648 -21546
rect 397308 -21688 397374 -21632
rect 397430 -21688 397516 -21632
rect 397572 -21688 397648 -21632
rect 397308 -21774 397648 -21688
rect 397308 -21830 397374 -21774
rect 397430 -21830 397516 -21774
rect 397572 -21830 397648 -21774
rect 397308 -21916 397648 -21830
rect 397308 -21972 397374 -21916
rect 397430 -21972 397516 -21916
rect 397572 -21972 397648 -21916
rect 397308 -22058 397648 -21972
rect 397308 -22114 397374 -22058
rect 397430 -22114 397516 -22058
rect 397572 -22114 397648 -22058
rect 397308 -22200 397648 -22114
rect 397308 -22256 397374 -22200
rect 397430 -22256 397516 -22200
rect 397572 -22256 397648 -22200
rect 397308 -22342 397648 -22256
rect 397308 -22398 397374 -22342
rect 397430 -22398 397516 -22342
rect 397572 -22398 397648 -22342
rect 397308 -22484 397648 -22398
rect 397308 -22540 397374 -22484
rect 397430 -22540 397516 -22484
rect 397572 -22540 397648 -22484
rect 397308 -22626 397648 -22540
rect 397308 -22682 397374 -22626
rect 397430 -22682 397516 -22626
rect 397572 -22682 397648 -22626
rect 397308 -22768 397648 -22682
rect 397308 -22824 397374 -22768
rect 397430 -22824 397516 -22768
rect 397572 -22824 397648 -22768
rect 397308 -22910 397648 -22824
rect 397308 -22966 397374 -22910
rect 397430 -22966 397516 -22910
rect 397572 -22966 397648 -22910
rect 397308 -23052 397648 -22966
rect 397308 -23108 397374 -23052
rect 397430 -23108 397516 -23052
rect 397572 -23108 397648 -23052
rect 397308 -23194 397648 -23108
rect 397308 -23250 397374 -23194
rect 397430 -23250 397516 -23194
rect 397572 -23250 397648 -23194
rect 397308 -23336 397648 -23250
rect 397308 -23392 397374 -23336
rect 397430 -23392 397516 -23336
rect 397572 -23392 397648 -23336
rect 397308 -23478 397648 -23392
rect 397308 -23534 397374 -23478
rect 397430 -23534 397516 -23478
rect 397572 -23534 397648 -23478
rect 397308 -23620 397648 -23534
rect 397308 -23676 397374 -23620
rect 397430 -23676 397516 -23620
rect 397572 -23676 397648 -23620
rect 397308 -23762 397648 -23676
rect 397308 -23818 397374 -23762
rect 397430 -23818 397516 -23762
rect 397572 -23818 397648 -23762
rect 397308 -23904 397648 -23818
rect 397308 -23960 397374 -23904
rect 397430 -23960 397516 -23904
rect 397572 -23960 397648 -23904
rect 397308 -24046 397648 -23960
rect 397308 -24102 397374 -24046
rect 397430 -24102 397516 -24046
rect 397572 -24102 397648 -24046
rect 397308 -24188 397648 -24102
rect 397308 -24244 397374 -24188
rect 397430 -24244 397516 -24188
rect 397572 -24244 397648 -24188
rect 397308 -24330 397648 -24244
rect 397308 -24386 397374 -24330
rect 397430 -24386 397516 -24330
rect 397572 -24386 397648 -24330
rect 397308 -24472 397648 -24386
rect 397308 -24528 397374 -24472
rect 397430 -24528 397516 -24472
rect 397572 -24528 397648 -24472
rect 397308 -24614 397648 -24528
rect 397308 -24670 397374 -24614
rect 397430 -24670 397516 -24614
rect 397572 -24670 397648 -24614
rect 397308 -24756 397648 -24670
rect 397308 -24812 397374 -24756
rect 397430 -24812 397516 -24756
rect 397572 -24812 397648 -24756
rect 397308 -24898 397648 -24812
rect 397308 -24954 397374 -24898
rect 397430 -24954 397516 -24898
rect 397572 -24954 397648 -24898
rect 397308 -25040 397648 -24954
rect 397308 -25096 397374 -25040
rect 397430 -25096 397516 -25040
rect 397572 -25096 397648 -25040
rect 397308 -25182 397648 -25096
rect 397308 -25238 397374 -25182
rect 397430 -25238 397516 -25182
rect 397572 -25238 397648 -25182
rect 397308 -25324 397648 -25238
rect 397308 -25380 397374 -25324
rect 397430 -25380 397516 -25324
rect 397572 -25380 397648 -25324
rect 397308 -25466 397648 -25380
rect 397308 -25522 397374 -25466
rect 397430 -25522 397516 -25466
rect 397572 -25522 397648 -25466
rect 397308 -25532 397648 -25522
rect 397708 -13680 398048 -13670
rect 397708 -13736 397778 -13680
rect 397834 -13736 397920 -13680
rect 397976 -13736 398048 -13680
rect 397708 -13822 398048 -13736
rect 397708 -13878 397778 -13822
rect 397834 -13878 397920 -13822
rect 397976 -13878 398048 -13822
rect 397708 -13964 398048 -13878
rect 397708 -14020 397778 -13964
rect 397834 -14020 397920 -13964
rect 397976 -14020 398048 -13964
rect 397708 -14106 398048 -14020
rect 397708 -14162 397778 -14106
rect 397834 -14162 397920 -14106
rect 397976 -14162 398048 -14106
rect 397708 -14248 398048 -14162
rect 397708 -14304 397778 -14248
rect 397834 -14304 397920 -14248
rect 397976 -14304 398048 -14248
rect 397708 -14390 398048 -14304
rect 397708 -14446 397778 -14390
rect 397834 -14446 397920 -14390
rect 397976 -14446 398048 -14390
rect 397708 -14532 398048 -14446
rect 397708 -14588 397778 -14532
rect 397834 -14588 397920 -14532
rect 397976 -14588 398048 -14532
rect 397708 -14674 398048 -14588
rect 397708 -14730 397778 -14674
rect 397834 -14730 397920 -14674
rect 397976 -14730 398048 -14674
rect 397708 -14816 398048 -14730
rect 397708 -14872 397778 -14816
rect 397834 -14872 397920 -14816
rect 397976 -14872 398048 -14816
rect 397708 -14958 398048 -14872
rect 397708 -15014 397778 -14958
rect 397834 -15014 397920 -14958
rect 397976 -15014 398048 -14958
rect 397708 -15100 398048 -15014
rect 397708 -15156 397778 -15100
rect 397834 -15156 397920 -15100
rect 397976 -15156 398048 -15100
rect 397708 -15242 398048 -15156
rect 397708 -15298 397778 -15242
rect 397834 -15298 397920 -15242
rect 397976 -15298 398048 -15242
rect 397708 -15384 398048 -15298
rect 397708 -15440 397778 -15384
rect 397834 -15440 397920 -15384
rect 397976 -15440 398048 -15384
rect 397708 -15526 398048 -15440
rect 397708 -15582 397778 -15526
rect 397834 -15582 397920 -15526
rect 397976 -15582 398048 -15526
rect 397708 -15668 398048 -15582
rect 397708 -15724 397778 -15668
rect 397834 -15724 397920 -15668
rect 397976 -15724 398048 -15668
rect 397708 -15810 398048 -15724
rect 397708 -15866 397778 -15810
rect 397834 -15866 397920 -15810
rect 397976 -15866 398048 -15810
rect 397708 -15952 398048 -15866
rect 397708 -16008 397778 -15952
rect 397834 -16008 397920 -15952
rect 397976 -16008 398048 -15952
rect 397708 -16094 398048 -16008
rect 397708 -16150 397778 -16094
rect 397834 -16150 397920 -16094
rect 397976 -16150 398048 -16094
rect 397708 -16236 398048 -16150
rect 397708 -16292 397778 -16236
rect 397834 -16292 397920 -16236
rect 397976 -16292 398048 -16236
rect 397708 -16378 398048 -16292
rect 397708 -16434 397778 -16378
rect 397834 -16434 397920 -16378
rect 397976 -16434 398048 -16378
rect 397708 -16520 398048 -16434
rect 397708 -16576 397778 -16520
rect 397834 -16576 397920 -16520
rect 397976 -16576 398048 -16520
rect 397708 -16662 398048 -16576
rect 397708 -16718 397778 -16662
rect 397834 -16718 397920 -16662
rect 397976 -16718 398048 -16662
rect 397708 -16804 398048 -16718
rect 397708 -16860 397778 -16804
rect 397834 -16860 397920 -16804
rect 397976 -16860 398048 -16804
rect 397708 -16946 398048 -16860
rect 397708 -17002 397778 -16946
rect 397834 -17002 397920 -16946
rect 397976 -17002 398048 -16946
rect 397708 -17088 398048 -17002
rect 397708 -17144 397778 -17088
rect 397834 -17144 397920 -17088
rect 397976 -17144 398048 -17088
rect 397708 -17230 398048 -17144
rect 397708 -17286 397778 -17230
rect 397834 -17286 397920 -17230
rect 397976 -17286 398048 -17230
rect 397708 -17372 398048 -17286
rect 397708 -17428 397778 -17372
rect 397834 -17428 397920 -17372
rect 397976 -17428 398048 -17372
rect 397708 -17514 398048 -17428
rect 397708 -17570 397778 -17514
rect 397834 -17570 397920 -17514
rect 397976 -17570 398048 -17514
rect 397708 -17656 398048 -17570
rect 397708 -17712 397778 -17656
rect 397834 -17712 397920 -17656
rect 397976 -17712 398048 -17656
rect 397708 -17798 398048 -17712
rect 397708 -17854 397778 -17798
rect 397834 -17854 397920 -17798
rect 397976 -17854 398048 -17798
rect 397708 -17940 398048 -17854
rect 397708 -17996 397778 -17940
rect 397834 -17996 397920 -17940
rect 397976 -17996 398048 -17940
rect 397708 -18082 398048 -17996
rect 397708 -18138 397778 -18082
rect 397834 -18138 397920 -18082
rect 397976 -18138 398048 -18082
rect 397708 -18224 398048 -18138
rect 397708 -18280 397778 -18224
rect 397834 -18280 397920 -18224
rect 397976 -18280 398048 -18224
rect 397708 -18366 398048 -18280
rect 397708 -18422 397778 -18366
rect 397834 -18422 397920 -18366
rect 397976 -18422 398048 -18366
rect 397708 -18508 398048 -18422
rect 397708 -18564 397778 -18508
rect 397834 -18564 397920 -18508
rect 397976 -18564 398048 -18508
rect 397708 -18650 398048 -18564
rect 397708 -18706 397778 -18650
rect 397834 -18706 397920 -18650
rect 397976 -18706 398048 -18650
rect 397708 -18792 398048 -18706
rect 397708 -18848 397778 -18792
rect 397834 -18848 397920 -18792
rect 397976 -18848 398048 -18792
rect 397708 -18934 398048 -18848
rect 397708 -18990 397778 -18934
rect 397834 -18990 397920 -18934
rect 397976 -18990 398048 -18934
rect 397708 -19076 398048 -18990
rect 397708 -19132 397778 -19076
rect 397834 -19132 397920 -19076
rect 397976 -19132 398048 -19076
rect 397708 -19218 398048 -19132
rect 397708 -19274 397778 -19218
rect 397834 -19274 397920 -19218
rect 397976 -19274 398048 -19218
rect 397708 -19360 398048 -19274
rect 397708 -19416 397778 -19360
rect 397834 -19416 397920 -19360
rect 397976 -19416 398048 -19360
rect 397708 -19502 398048 -19416
rect 397708 -19558 397778 -19502
rect 397834 -19558 397920 -19502
rect 397976 -19558 398048 -19502
rect 397708 -19644 398048 -19558
rect 397708 -19700 397778 -19644
rect 397834 -19700 397920 -19644
rect 397976 -19700 398048 -19644
rect 397708 -19786 398048 -19700
rect 397708 -19842 397778 -19786
rect 397834 -19842 397920 -19786
rect 397976 -19842 398048 -19786
rect 397708 -19928 398048 -19842
rect 397708 -19984 397778 -19928
rect 397834 -19984 397920 -19928
rect 397976 -19984 398048 -19928
rect 397708 -20070 398048 -19984
rect 397708 -20126 397778 -20070
rect 397834 -20126 397920 -20070
rect 397976 -20126 398048 -20070
rect 397708 -20212 398048 -20126
rect 397708 -20268 397778 -20212
rect 397834 -20268 397920 -20212
rect 397976 -20268 398048 -20212
rect 397708 -20354 398048 -20268
rect 397708 -20410 397778 -20354
rect 397834 -20410 397920 -20354
rect 397976 -20410 398048 -20354
rect 397708 -20496 398048 -20410
rect 397708 -20552 397778 -20496
rect 397834 -20552 397920 -20496
rect 397976 -20552 398048 -20496
rect 397708 -20638 398048 -20552
rect 397708 -20694 397778 -20638
rect 397834 -20694 397920 -20638
rect 397976 -20694 398048 -20638
rect 397708 -20780 398048 -20694
rect 397708 -20836 397778 -20780
rect 397834 -20836 397920 -20780
rect 397976 -20836 398048 -20780
rect 397708 -20922 398048 -20836
rect 397708 -20978 397778 -20922
rect 397834 -20978 397920 -20922
rect 397976 -20978 398048 -20922
rect 397708 -21064 398048 -20978
rect 397708 -21120 397778 -21064
rect 397834 -21120 397920 -21064
rect 397976 -21120 398048 -21064
rect 397708 -21206 398048 -21120
rect 397708 -21262 397778 -21206
rect 397834 -21262 397920 -21206
rect 397976 -21262 398048 -21206
rect 397708 -21348 398048 -21262
rect 397708 -21404 397778 -21348
rect 397834 -21404 397920 -21348
rect 397976 -21404 398048 -21348
rect 397708 -21490 398048 -21404
rect 397708 -21546 397778 -21490
rect 397834 -21546 397920 -21490
rect 397976 -21546 398048 -21490
rect 397708 -21632 398048 -21546
rect 397708 -21688 397778 -21632
rect 397834 -21688 397920 -21632
rect 397976 -21688 398048 -21632
rect 397708 -21774 398048 -21688
rect 397708 -21830 397778 -21774
rect 397834 -21830 397920 -21774
rect 397976 -21830 398048 -21774
rect 397708 -21916 398048 -21830
rect 397708 -21972 397778 -21916
rect 397834 -21972 397920 -21916
rect 397976 -21972 398048 -21916
rect 397708 -22058 398048 -21972
rect 397708 -22114 397778 -22058
rect 397834 -22114 397920 -22058
rect 397976 -22114 398048 -22058
rect 397708 -22200 398048 -22114
rect 397708 -22256 397778 -22200
rect 397834 -22256 397920 -22200
rect 397976 -22256 398048 -22200
rect 397708 -22342 398048 -22256
rect 397708 -22398 397778 -22342
rect 397834 -22398 397920 -22342
rect 397976 -22398 398048 -22342
rect 397708 -22484 398048 -22398
rect 397708 -22540 397778 -22484
rect 397834 -22540 397920 -22484
rect 397976 -22540 398048 -22484
rect 397708 -22626 398048 -22540
rect 397708 -22682 397778 -22626
rect 397834 -22682 397920 -22626
rect 397976 -22682 398048 -22626
rect 397708 -22768 398048 -22682
rect 397708 -22824 397778 -22768
rect 397834 -22824 397920 -22768
rect 397976 -22824 398048 -22768
rect 397708 -22910 398048 -22824
rect 397708 -22966 397778 -22910
rect 397834 -22966 397920 -22910
rect 397976 -22966 398048 -22910
rect 397708 -23052 398048 -22966
rect 397708 -23108 397778 -23052
rect 397834 -23108 397920 -23052
rect 397976 -23108 398048 -23052
rect 397708 -23194 398048 -23108
rect 397708 -23250 397778 -23194
rect 397834 -23250 397920 -23194
rect 397976 -23250 398048 -23194
rect 397708 -23336 398048 -23250
rect 397708 -23392 397778 -23336
rect 397834 -23392 397920 -23336
rect 397976 -23392 398048 -23336
rect 397708 -23478 398048 -23392
rect 397708 -23534 397778 -23478
rect 397834 -23534 397920 -23478
rect 397976 -23534 398048 -23478
rect 397708 -23620 398048 -23534
rect 397708 -23676 397778 -23620
rect 397834 -23676 397920 -23620
rect 397976 -23676 398048 -23620
rect 397708 -23762 398048 -23676
rect 397708 -23818 397778 -23762
rect 397834 -23818 397920 -23762
rect 397976 -23818 398048 -23762
rect 397708 -23904 398048 -23818
rect 397708 -23960 397778 -23904
rect 397834 -23960 397920 -23904
rect 397976 -23960 398048 -23904
rect 397708 -24046 398048 -23960
rect 397708 -24102 397778 -24046
rect 397834 -24102 397920 -24046
rect 397976 -24102 398048 -24046
rect 397708 -24188 398048 -24102
rect 397708 -24244 397778 -24188
rect 397834 -24244 397920 -24188
rect 397976 -24244 398048 -24188
rect 397708 -24330 398048 -24244
rect 397708 -24386 397778 -24330
rect 397834 -24386 397920 -24330
rect 397976 -24386 398048 -24330
rect 397708 -24472 398048 -24386
rect 397708 -24528 397778 -24472
rect 397834 -24528 397920 -24472
rect 397976 -24528 398048 -24472
rect 397708 -24614 398048 -24528
rect 397708 -24670 397778 -24614
rect 397834 -24670 397920 -24614
rect 397976 -24670 398048 -24614
rect 397708 -24756 398048 -24670
rect 397708 -24812 397778 -24756
rect 397834 -24812 397920 -24756
rect 397976 -24812 398048 -24756
rect 397708 -24898 398048 -24812
rect 397708 -24954 397778 -24898
rect 397834 -24954 397920 -24898
rect 397976 -24954 398048 -24898
rect 397708 -25040 398048 -24954
rect 397708 -25096 397778 -25040
rect 397834 -25096 397920 -25040
rect 397976 -25096 398048 -25040
rect 397708 -25182 398048 -25096
rect 397708 -25238 397778 -25182
rect 397834 -25238 397920 -25182
rect 397976 -25238 398048 -25182
rect 397708 -25324 398048 -25238
rect 397708 -25380 397778 -25324
rect 397834 -25380 397920 -25324
rect 397976 -25380 398048 -25324
rect 397708 -25466 398048 -25380
rect 397708 -25522 397778 -25466
rect 397834 -25522 397920 -25466
rect 397976 -25522 398048 -25466
rect 397708 -25532 398048 -25522
rect 398108 -13680 398448 -13670
rect 398108 -13736 398174 -13680
rect 398230 -13736 398316 -13680
rect 398372 -13736 398448 -13680
rect 398108 -13822 398448 -13736
rect 398108 -13878 398174 -13822
rect 398230 -13878 398316 -13822
rect 398372 -13878 398448 -13822
rect 398108 -13964 398448 -13878
rect 398108 -14020 398174 -13964
rect 398230 -14020 398316 -13964
rect 398372 -14020 398448 -13964
rect 398108 -14106 398448 -14020
rect 398108 -14162 398174 -14106
rect 398230 -14162 398316 -14106
rect 398372 -14162 398448 -14106
rect 398108 -14248 398448 -14162
rect 398108 -14304 398174 -14248
rect 398230 -14304 398316 -14248
rect 398372 -14304 398448 -14248
rect 398108 -14390 398448 -14304
rect 398108 -14446 398174 -14390
rect 398230 -14446 398316 -14390
rect 398372 -14446 398448 -14390
rect 398108 -14532 398448 -14446
rect 398108 -14588 398174 -14532
rect 398230 -14588 398316 -14532
rect 398372 -14588 398448 -14532
rect 398108 -14674 398448 -14588
rect 398108 -14730 398174 -14674
rect 398230 -14730 398316 -14674
rect 398372 -14730 398448 -14674
rect 398108 -14816 398448 -14730
rect 398108 -14872 398174 -14816
rect 398230 -14872 398316 -14816
rect 398372 -14872 398448 -14816
rect 398108 -14958 398448 -14872
rect 398108 -15014 398174 -14958
rect 398230 -15014 398316 -14958
rect 398372 -15014 398448 -14958
rect 398108 -15100 398448 -15014
rect 398108 -15156 398174 -15100
rect 398230 -15156 398316 -15100
rect 398372 -15156 398448 -15100
rect 398108 -15242 398448 -15156
rect 398108 -15298 398174 -15242
rect 398230 -15298 398316 -15242
rect 398372 -15298 398448 -15242
rect 398108 -15384 398448 -15298
rect 398108 -15440 398174 -15384
rect 398230 -15440 398316 -15384
rect 398372 -15440 398448 -15384
rect 398108 -15526 398448 -15440
rect 398108 -15582 398174 -15526
rect 398230 -15582 398316 -15526
rect 398372 -15582 398448 -15526
rect 398108 -15668 398448 -15582
rect 398108 -15724 398174 -15668
rect 398230 -15724 398316 -15668
rect 398372 -15724 398448 -15668
rect 398108 -15810 398448 -15724
rect 398108 -15866 398174 -15810
rect 398230 -15866 398316 -15810
rect 398372 -15866 398448 -15810
rect 398108 -15952 398448 -15866
rect 398108 -16008 398174 -15952
rect 398230 -16008 398316 -15952
rect 398372 -16008 398448 -15952
rect 398108 -16094 398448 -16008
rect 398108 -16150 398174 -16094
rect 398230 -16150 398316 -16094
rect 398372 -16150 398448 -16094
rect 398108 -16236 398448 -16150
rect 398108 -16292 398174 -16236
rect 398230 -16292 398316 -16236
rect 398372 -16292 398448 -16236
rect 398108 -16378 398448 -16292
rect 398108 -16434 398174 -16378
rect 398230 -16434 398316 -16378
rect 398372 -16434 398448 -16378
rect 398108 -16520 398448 -16434
rect 398108 -16576 398174 -16520
rect 398230 -16576 398316 -16520
rect 398372 -16576 398448 -16520
rect 398108 -16662 398448 -16576
rect 398108 -16718 398174 -16662
rect 398230 -16718 398316 -16662
rect 398372 -16718 398448 -16662
rect 398108 -16804 398448 -16718
rect 398108 -16860 398174 -16804
rect 398230 -16860 398316 -16804
rect 398372 -16860 398448 -16804
rect 398108 -16946 398448 -16860
rect 398108 -17002 398174 -16946
rect 398230 -17002 398316 -16946
rect 398372 -17002 398448 -16946
rect 398108 -17088 398448 -17002
rect 398108 -17144 398174 -17088
rect 398230 -17144 398316 -17088
rect 398372 -17144 398448 -17088
rect 398108 -17230 398448 -17144
rect 398108 -17286 398174 -17230
rect 398230 -17286 398316 -17230
rect 398372 -17286 398448 -17230
rect 398108 -17372 398448 -17286
rect 398108 -17428 398174 -17372
rect 398230 -17428 398316 -17372
rect 398372 -17428 398448 -17372
rect 398108 -17514 398448 -17428
rect 398108 -17570 398174 -17514
rect 398230 -17570 398316 -17514
rect 398372 -17570 398448 -17514
rect 398108 -17656 398448 -17570
rect 398108 -17712 398174 -17656
rect 398230 -17712 398316 -17656
rect 398372 -17712 398448 -17656
rect 398108 -17798 398448 -17712
rect 398108 -17854 398174 -17798
rect 398230 -17854 398316 -17798
rect 398372 -17854 398448 -17798
rect 398108 -17940 398448 -17854
rect 398108 -17996 398174 -17940
rect 398230 -17996 398316 -17940
rect 398372 -17996 398448 -17940
rect 398108 -18082 398448 -17996
rect 398108 -18138 398174 -18082
rect 398230 -18138 398316 -18082
rect 398372 -18138 398448 -18082
rect 398108 -18224 398448 -18138
rect 398108 -18280 398174 -18224
rect 398230 -18280 398316 -18224
rect 398372 -18280 398448 -18224
rect 398108 -18366 398448 -18280
rect 398108 -18422 398174 -18366
rect 398230 -18422 398316 -18366
rect 398372 -18422 398448 -18366
rect 398108 -18508 398448 -18422
rect 398108 -18564 398174 -18508
rect 398230 -18564 398316 -18508
rect 398372 -18564 398448 -18508
rect 398108 -18650 398448 -18564
rect 398108 -18706 398174 -18650
rect 398230 -18706 398316 -18650
rect 398372 -18706 398448 -18650
rect 398108 -18792 398448 -18706
rect 398108 -18848 398174 -18792
rect 398230 -18848 398316 -18792
rect 398372 -18848 398448 -18792
rect 398108 -18934 398448 -18848
rect 398108 -18990 398174 -18934
rect 398230 -18990 398316 -18934
rect 398372 -18990 398448 -18934
rect 398108 -19076 398448 -18990
rect 398108 -19132 398174 -19076
rect 398230 -19132 398316 -19076
rect 398372 -19132 398448 -19076
rect 398108 -19218 398448 -19132
rect 398108 -19274 398174 -19218
rect 398230 -19274 398316 -19218
rect 398372 -19274 398448 -19218
rect 398108 -19360 398448 -19274
rect 398108 -19416 398174 -19360
rect 398230 -19416 398316 -19360
rect 398372 -19416 398448 -19360
rect 398108 -19502 398448 -19416
rect 398108 -19558 398174 -19502
rect 398230 -19558 398316 -19502
rect 398372 -19558 398448 -19502
rect 398108 -19644 398448 -19558
rect 398108 -19700 398174 -19644
rect 398230 -19700 398316 -19644
rect 398372 -19700 398448 -19644
rect 398108 -19786 398448 -19700
rect 398108 -19842 398174 -19786
rect 398230 -19842 398316 -19786
rect 398372 -19842 398448 -19786
rect 398108 -19928 398448 -19842
rect 398108 -19984 398174 -19928
rect 398230 -19984 398316 -19928
rect 398372 -19984 398448 -19928
rect 398108 -20070 398448 -19984
rect 398108 -20126 398174 -20070
rect 398230 -20126 398316 -20070
rect 398372 -20126 398448 -20070
rect 398108 -20212 398448 -20126
rect 398108 -20268 398174 -20212
rect 398230 -20268 398316 -20212
rect 398372 -20268 398448 -20212
rect 398108 -20354 398448 -20268
rect 398108 -20410 398174 -20354
rect 398230 -20410 398316 -20354
rect 398372 -20410 398448 -20354
rect 398108 -20496 398448 -20410
rect 398108 -20552 398174 -20496
rect 398230 -20552 398316 -20496
rect 398372 -20552 398448 -20496
rect 398108 -20638 398448 -20552
rect 398108 -20694 398174 -20638
rect 398230 -20694 398316 -20638
rect 398372 -20694 398448 -20638
rect 398108 -20780 398448 -20694
rect 398108 -20836 398174 -20780
rect 398230 -20836 398316 -20780
rect 398372 -20836 398448 -20780
rect 398108 -20922 398448 -20836
rect 398108 -20978 398174 -20922
rect 398230 -20978 398316 -20922
rect 398372 -20978 398448 -20922
rect 398108 -21064 398448 -20978
rect 398108 -21120 398174 -21064
rect 398230 -21120 398316 -21064
rect 398372 -21120 398448 -21064
rect 398108 -21206 398448 -21120
rect 398108 -21262 398174 -21206
rect 398230 -21262 398316 -21206
rect 398372 -21262 398448 -21206
rect 398108 -21348 398448 -21262
rect 398108 -21404 398174 -21348
rect 398230 -21404 398316 -21348
rect 398372 -21404 398448 -21348
rect 398108 -21490 398448 -21404
rect 398108 -21546 398174 -21490
rect 398230 -21546 398316 -21490
rect 398372 -21546 398448 -21490
rect 398108 -21632 398448 -21546
rect 398108 -21688 398174 -21632
rect 398230 -21688 398316 -21632
rect 398372 -21688 398448 -21632
rect 398108 -21774 398448 -21688
rect 398108 -21830 398174 -21774
rect 398230 -21830 398316 -21774
rect 398372 -21830 398448 -21774
rect 398108 -21916 398448 -21830
rect 398108 -21972 398174 -21916
rect 398230 -21972 398316 -21916
rect 398372 -21972 398448 -21916
rect 398108 -22058 398448 -21972
rect 398108 -22114 398174 -22058
rect 398230 -22114 398316 -22058
rect 398372 -22114 398448 -22058
rect 398108 -22200 398448 -22114
rect 398108 -22256 398174 -22200
rect 398230 -22256 398316 -22200
rect 398372 -22256 398448 -22200
rect 398108 -22342 398448 -22256
rect 398108 -22398 398174 -22342
rect 398230 -22398 398316 -22342
rect 398372 -22398 398448 -22342
rect 398108 -22484 398448 -22398
rect 398108 -22540 398174 -22484
rect 398230 -22540 398316 -22484
rect 398372 -22540 398448 -22484
rect 398108 -22626 398448 -22540
rect 398108 -22682 398174 -22626
rect 398230 -22682 398316 -22626
rect 398372 -22682 398448 -22626
rect 398108 -22768 398448 -22682
rect 398108 -22824 398174 -22768
rect 398230 -22824 398316 -22768
rect 398372 -22824 398448 -22768
rect 398108 -22910 398448 -22824
rect 398108 -22966 398174 -22910
rect 398230 -22966 398316 -22910
rect 398372 -22966 398448 -22910
rect 398108 -23052 398448 -22966
rect 398108 -23108 398174 -23052
rect 398230 -23108 398316 -23052
rect 398372 -23108 398448 -23052
rect 398108 -23194 398448 -23108
rect 398108 -23250 398174 -23194
rect 398230 -23250 398316 -23194
rect 398372 -23250 398448 -23194
rect 398108 -23336 398448 -23250
rect 398108 -23392 398174 -23336
rect 398230 -23392 398316 -23336
rect 398372 -23392 398448 -23336
rect 398108 -23478 398448 -23392
rect 398108 -23534 398174 -23478
rect 398230 -23534 398316 -23478
rect 398372 -23534 398448 -23478
rect 398108 -23620 398448 -23534
rect 398108 -23676 398174 -23620
rect 398230 -23676 398316 -23620
rect 398372 -23676 398448 -23620
rect 398108 -23762 398448 -23676
rect 398108 -23818 398174 -23762
rect 398230 -23818 398316 -23762
rect 398372 -23818 398448 -23762
rect 398108 -23904 398448 -23818
rect 398108 -23960 398174 -23904
rect 398230 -23960 398316 -23904
rect 398372 -23960 398448 -23904
rect 398108 -24046 398448 -23960
rect 398108 -24102 398174 -24046
rect 398230 -24102 398316 -24046
rect 398372 -24102 398448 -24046
rect 398108 -24188 398448 -24102
rect 398108 -24244 398174 -24188
rect 398230 -24244 398316 -24188
rect 398372 -24244 398448 -24188
rect 398108 -24330 398448 -24244
rect 398108 -24386 398174 -24330
rect 398230 -24386 398316 -24330
rect 398372 -24386 398448 -24330
rect 398108 -24472 398448 -24386
rect 398108 -24528 398174 -24472
rect 398230 -24528 398316 -24472
rect 398372 -24528 398448 -24472
rect 398108 -24614 398448 -24528
rect 398108 -24670 398174 -24614
rect 398230 -24670 398316 -24614
rect 398372 -24670 398448 -24614
rect 398108 -24756 398448 -24670
rect 398108 -24812 398174 -24756
rect 398230 -24812 398316 -24756
rect 398372 -24812 398448 -24756
rect 398108 -24898 398448 -24812
rect 398108 -24954 398174 -24898
rect 398230 -24954 398316 -24898
rect 398372 -24954 398448 -24898
rect 398108 -25040 398448 -24954
rect 398108 -25096 398174 -25040
rect 398230 -25096 398316 -25040
rect 398372 -25096 398448 -25040
rect 398108 -25182 398448 -25096
rect 398108 -25238 398174 -25182
rect 398230 -25238 398316 -25182
rect 398372 -25238 398448 -25182
rect 398108 -25324 398448 -25238
rect 398108 -25380 398174 -25324
rect 398230 -25380 398316 -25324
rect 398372 -25380 398448 -25324
rect 398108 -25466 398448 -25380
rect 398108 -25522 398174 -25466
rect 398230 -25522 398316 -25466
rect 398372 -25522 398448 -25466
rect 398108 -25532 398448 -25522
rect 398508 -13680 398848 -13670
rect 398508 -13736 398574 -13680
rect 398630 -13736 398716 -13680
rect 398772 -13736 398848 -13680
rect 398508 -13822 398848 -13736
rect 398508 -13878 398574 -13822
rect 398630 -13878 398716 -13822
rect 398772 -13878 398848 -13822
rect 398508 -13964 398848 -13878
rect 398508 -14020 398574 -13964
rect 398630 -14020 398716 -13964
rect 398772 -14020 398848 -13964
rect 398508 -14106 398848 -14020
rect 398508 -14162 398574 -14106
rect 398630 -14162 398716 -14106
rect 398772 -14162 398848 -14106
rect 398508 -14248 398848 -14162
rect 398508 -14304 398574 -14248
rect 398630 -14304 398716 -14248
rect 398772 -14304 398848 -14248
rect 398508 -14390 398848 -14304
rect 398508 -14446 398574 -14390
rect 398630 -14446 398716 -14390
rect 398772 -14446 398848 -14390
rect 398508 -14532 398848 -14446
rect 398508 -14588 398574 -14532
rect 398630 -14588 398716 -14532
rect 398772 -14588 398848 -14532
rect 398508 -14674 398848 -14588
rect 398508 -14730 398574 -14674
rect 398630 -14730 398716 -14674
rect 398772 -14730 398848 -14674
rect 398508 -14816 398848 -14730
rect 398508 -14872 398574 -14816
rect 398630 -14872 398716 -14816
rect 398772 -14872 398848 -14816
rect 398508 -14958 398848 -14872
rect 398508 -15014 398574 -14958
rect 398630 -15014 398716 -14958
rect 398772 -15014 398848 -14958
rect 398508 -15100 398848 -15014
rect 398508 -15156 398574 -15100
rect 398630 -15156 398716 -15100
rect 398772 -15156 398848 -15100
rect 398508 -15242 398848 -15156
rect 398508 -15298 398574 -15242
rect 398630 -15298 398716 -15242
rect 398772 -15298 398848 -15242
rect 398508 -15384 398848 -15298
rect 398508 -15440 398574 -15384
rect 398630 -15440 398716 -15384
rect 398772 -15440 398848 -15384
rect 398508 -15526 398848 -15440
rect 398508 -15582 398574 -15526
rect 398630 -15582 398716 -15526
rect 398772 -15582 398848 -15526
rect 398508 -15668 398848 -15582
rect 398508 -15724 398574 -15668
rect 398630 -15724 398716 -15668
rect 398772 -15724 398848 -15668
rect 398508 -15810 398848 -15724
rect 398508 -15866 398574 -15810
rect 398630 -15866 398716 -15810
rect 398772 -15866 398848 -15810
rect 398508 -15952 398848 -15866
rect 398508 -16008 398574 -15952
rect 398630 -16008 398716 -15952
rect 398772 -16008 398848 -15952
rect 398508 -16094 398848 -16008
rect 398508 -16150 398574 -16094
rect 398630 -16150 398716 -16094
rect 398772 -16150 398848 -16094
rect 398508 -16236 398848 -16150
rect 398508 -16292 398574 -16236
rect 398630 -16292 398716 -16236
rect 398772 -16292 398848 -16236
rect 398508 -16378 398848 -16292
rect 398508 -16434 398574 -16378
rect 398630 -16434 398716 -16378
rect 398772 -16434 398848 -16378
rect 398508 -16520 398848 -16434
rect 398508 -16576 398574 -16520
rect 398630 -16576 398716 -16520
rect 398772 -16576 398848 -16520
rect 398508 -16662 398848 -16576
rect 398508 -16718 398574 -16662
rect 398630 -16718 398716 -16662
rect 398772 -16718 398848 -16662
rect 398508 -16804 398848 -16718
rect 398508 -16860 398574 -16804
rect 398630 -16860 398716 -16804
rect 398772 -16860 398848 -16804
rect 398508 -16946 398848 -16860
rect 398508 -17002 398574 -16946
rect 398630 -17002 398716 -16946
rect 398772 -17002 398848 -16946
rect 398508 -17088 398848 -17002
rect 398508 -17144 398574 -17088
rect 398630 -17144 398716 -17088
rect 398772 -17144 398848 -17088
rect 398508 -17230 398848 -17144
rect 398508 -17286 398574 -17230
rect 398630 -17286 398716 -17230
rect 398772 -17286 398848 -17230
rect 398508 -17372 398848 -17286
rect 398508 -17428 398574 -17372
rect 398630 -17428 398716 -17372
rect 398772 -17428 398848 -17372
rect 398508 -17514 398848 -17428
rect 398508 -17570 398574 -17514
rect 398630 -17570 398716 -17514
rect 398772 -17570 398848 -17514
rect 398508 -17656 398848 -17570
rect 398508 -17712 398574 -17656
rect 398630 -17712 398716 -17656
rect 398772 -17712 398848 -17656
rect 398508 -17798 398848 -17712
rect 398508 -17854 398574 -17798
rect 398630 -17854 398716 -17798
rect 398772 -17854 398848 -17798
rect 398508 -17940 398848 -17854
rect 398508 -17996 398574 -17940
rect 398630 -17996 398716 -17940
rect 398772 -17996 398848 -17940
rect 398508 -18082 398848 -17996
rect 398508 -18138 398574 -18082
rect 398630 -18138 398716 -18082
rect 398772 -18138 398848 -18082
rect 398508 -18224 398848 -18138
rect 398508 -18280 398574 -18224
rect 398630 -18280 398716 -18224
rect 398772 -18280 398848 -18224
rect 398508 -18366 398848 -18280
rect 398508 -18422 398574 -18366
rect 398630 -18422 398716 -18366
rect 398772 -18422 398848 -18366
rect 398508 -18508 398848 -18422
rect 398508 -18564 398574 -18508
rect 398630 -18564 398716 -18508
rect 398772 -18564 398848 -18508
rect 398508 -18650 398848 -18564
rect 398508 -18706 398574 -18650
rect 398630 -18706 398716 -18650
rect 398772 -18706 398848 -18650
rect 398508 -18792 398848 -18706
rect 398508 -18848 398574 -18792
rect 398630 -18848 398716 -18792
rect 398772 -18848 398848 -18792
rect 398508 -18934 398848 -18848
rect 398508 -18990 398574 -18934
rect 398630 -18990 398716 -18934
rect 398772 -18990 398848 -18934
rect 398508 -19076 398848 -18990
rect 398508 -19132 398574 -19076
rect 398630 -19132 398716 -19076
rect 398772 -19132 398848 -19076
rect 398508 -19218 398848 -19132
rect 398508 -19274 398574 -19218
rect 398630 -19274 398716 -19218
rect 398772 -19274 398848 -19218
rect 398508 -19360 398848 -19274
rect 398508 -19416 398574 -19360
rect 398630 -19416 398716 -19360
rect 398772 -19416 398848 -19360
rect 398508 -19502 398848 -19416
rect 398508 -19558 398574 -19502
rect 398630 -19558 398716 -19502
rect 398772 -19558 398848 -19502
rect 398508 -19644 398848 -19558
rect 398508 -19700 398574 -19644
rect 398630 -19700 398716 -19644
rect 398772 -19700 398848 -19644
rect 398508 -19786 398848 -19700
rect 398508 -19842 398574 -19786
rect 398630 -19842 398716 -19786
rect 398772 -19842 398848 -19786
rect 398508 -19928 398848 -19842
rect 398508 -19984 398574 -19928
rect 398630 -19984 398716 -19928
rect 398772 -19984 398848 -19928
rect 398508 -20070 398848 -19984
rect 398508 -20126 398574 -20070
rect 398630 -20126 398716 -20070
rect 398772 -20126 398848 -20070
rect 398508 -20212 398848 -20126
rect 398508 -20268 398574 -20212
rect 398630 -20268 398716 -20212
rect 398772 -20268 398848 -20212
rect 398508 -20354 398848 -20268
rect 398508 -20410 398574 -20354
rect 398630 -20410 398716 -20354
rect 398772 -20410 398848 -20354
rect 398508 -20496 398848 -20410
rect 398508 -20552 398574 -20496
rect 398630 -20552 398716 -20496
rect 398772 -20552 398848 -20496
rect 398508 -20638 398848 -20552
rect 398508 -20694 398574 -20638
rect 398630 -20694 398716 -20638
rect 398772 -20694 398848 -20638
rect 398508 -20780 398848 -20694
rect 398508 -20836 398574 -20780
rect 398630 -20836 398716 -20780
rect 398772 -20836 398848 -20780
rect 398508 -20922 398848 -20836
rect 398508 -20978 398574 -20922
rect 398630 -20978 398716 -20922
rect 398772 -20978 398848 -20922
rect 398508 -21064 398848 -20978
rect 398508 -21120 398574 -21064
rect 398630 -21120 398716 -21064
rect 398772 -21120 398848 -21064
rect 398508 -21206 398848 -21120
rect 398508 -21262 398574 -21206
rect 398630 -21262 398716 -21206
rect 398772 -21262 398848 -21206
rect 398508 -21348 398848 -21262
rect 398508 -21404 398574 -21348
rect 398630 -21404 398716 -21348
rect 398772 -21404 398848 -21348
rect 398508 -21490 398848 -21404
rect 398508 -21546 398574 -21490
rect 398630 -21546 398716 -21490
rect 398772 -21546 398848 -21490
rect 398508 -21632 398848 -21546
rect 398508 -21688 398574 -21632
rect 398630 -21688 398716 -21632
rect 398772 -21688 398848 -21632
rect 398508 -21774 398848 -21688
rect 398508 -21830 398574 -21774
rect 398630 -21830 398716 -21774
rect 398772 -21830 398848 -21774
rect 398508 -21916 398848 -21830
rect 398508 -21972 398574 -21916
rect 398630 -21972 398716 -21916
rect 398772 -21972 398848 -21916
rect 398508 -22058 398848 -21972
rect 398508 -22114 398574 -22058
rect 398630 -22114 398716 -22058
rect 398772 -22114 398848 -22058
rect 398508 -22200 398848 -22114
rect 398508 -22256 398574 -22200
rect 398630 -22256 398716 -22200
rect 398772 -22256 398848 -22200
rect 398508 -22342 398848 -22256
rect 398508 -22398 398574 -22342
rect 398630 -22398 398716 -22342
rect 398772 -22398 398848 -22342
rect 398508 -22484 398848 -22398
rect 398508 -22540 398574 -22484
rect 398630 -22540 398716 -22484
rect 398772 -22540 398848 -22484
rect 398508 -22626 398848 -22540
rect 398508 -22682 398574 -22626
rect 398630 -22682 398716 -22626
rect 398772 -22682 398848 -22626
rect 398508 -22768 398848 -22682
rect 398508 -22824 398574 -22768
rect 398630 -22824 398716 -22768
rect 398772 -22824 398848 -22768
rect 398508 -22910 398848 -22824
rect 398508 -22966 398574 -22910
rect 398630 -22966 398716 -22910
rect 398772 -22966 398848 -22910
rect 398508 -23052 398848 -22966
rect 398508 -23108 398574 -23052
rect 398630 -23108 398716 -23052
rect 398772 -23108 398848 -23052
rect 398508 -23194 398848 -23108
rect 398508 -23250 398574 -23194
rect 398630 -23250 398716 -23194
rect 398772 -23250 398848 -23194
rect 398508 -23336 398848 -23250
rect 398508 -23392 398574 -23336
rect 398630 -23392 398716 -23336
rect 398772 -23392 398848 -23336
rect 398508 -23478 398848 -23392
rect 398508 -23534 398574 -23478
rect 398630 -23534 398716 -23478
rect 398772 -23534 398848 -23478
rect 398508 -23620 398848 -23534
rect 398508 -23676 398574 -23620
rect 398630 -23676 398716 -23620
rect 398772 -23676 398848 -23620
rect 398508 -23762 398848 -23676
rect 398508 -23818 398574 -23762
rect 398630 -23818 398716 -23762
rect 398772 -23818 398848 -23762
rect 398508 -23904 398848 -23818
rect 398508 -23960 398574 -23904
rect 398630 -23960 398716 -23904
rect 398772 -23960 398848 -23904
rect 398508 -24046 398848 -23960
rect 398508 -24102 398574 -24046
rect 398630 -24102 398716 -24046
rect 398772 -24102 398848 -24046
rect 398508 -24188 398848 -24102
rect 398508 -24244 398574 -24188
rect 398630 -24244 398716 -24188
rect 398772 -24244 398848 -24188
rect 398508 -24330 398848 -24244
rect 398508 -24386 398574 -24330
rect 398630 -24386 398716 -24330
rect 398772 -24386 398848 -24330
rect 398508 -24472 398848 -24386
rect 398508 -24528 398574 -24472
rect 398630 -24528 398716 -24472
rect 398772 -24528 398848 -24472
rect 398508 -24614 398848 -24528
rect 398508 -24670 398574 -24614
rect 398630 -24670 398716 -24614
rect 398772 -24670 398848 -24614
rect 398508 -24756 398848 -24670
rect 398508 -24812 398574 -24756
rect 398630 -24812 398716 -24756
rect 398772 -24812 398848 -24756
rect 398508 -24898 398848 -24812
rect 398508 -24954 398574 -24898
rect 398630 -24954 398716 -24898
rect 398772 -24954 398848 -24898
rect 398508 -25040 398848 -24954
rect 398508 -25096 398574 -25040
rect 398630 -25096 398716 -25040
rect 398772 -25096 398848 -25040
rect 398508 -25182 398848 -25096
rect 398508 -25238 398574 -25182
rect 398630 -25238 398716 -25182
rect 398772 -25238 398848 -25182
rect 398508 -25324 398848 -25238
rect 398508 -25380 398574 -25324
rect 398630 -25380 398716 -25324
rect 398772 -25380 398848 -25324
rect 398508 -25466 398848 -25380
rect 398508 -25522 398574 -25466
rect 398630 -25522 398716 -25466
rect 398772 -25522 398848 -25466
rect 398508 -25532 398848 -25522
rect 398908 -13680 399248 -13670
rect 398908 -13736 398971 -13680
rect 399027 -13736 399113 -13680
rect 399169 -13736 399248 -13680
rect 398908 -13822 399248 -13736
rect 398908 -13878 398971 -13822
rect 399027 -13878 399113 -13822
rect 399169 -13878 399248 -13822
rect 398908 -13964 399248 -13878
rect 398908 -14020 398971 -13964
rect 399027 -14020 399113 -13964
rect 399169 -14020 399248 -13964
rect 398908 -14106 399248 -14020
rect 398908 -14162 398971 -14106
rect 399027 -14162 399113 -14106
rect 399169 -14162 399248 -14106
rect 398908 -14248 399248 -14162
rect 398908 -14304 398971 -14248
rect 399027 -14304 399113 -14248
rect 399169 -14304 399248 -14248
rect 398908 -14390 399248 -14304
rect 398908 -14446 398971 -14390
rect 399027 -14446 399113 -14390
rect 399169 -14446 399248 -14390
rect 398908 -14532 399248 -14446
rect 398908 -14588 398971 -14532
rect 399027 -14588 399113 -14532
rect 399169 -14588 399248 -14532
rect 398908 -14674 399248 -14588
rect 398908 -14730 398971 -14674
rect 399027 -14730 399113 -14674
rect 399169 -14730 399248 -14674
rect 398908 -14816 399248 -14730
rect 398908 -14872 398971 -14816
rect 399027 -14872 399113 -14816
rect 399169 -14872 399248 -14816
rect 398908 -14958 399248 -14872
rect 398908 -15014 398971 -14958
rect 399027 -15014 399113 -14958
rect 399169 -15014 399248 -14958
rect 398908 -15100 399248 -15014
rect 398908 -15156 398971 -15100
rect 399027 -15156 399113 -15100
rect 399169 -15156 399248 -15100
rect 398908 -15242 399248 -15156
rect 398908 -15298 398971 -15242
rect 399027 -15298 399113 -15242
rect 399169 -15298 399248 -15242
rect 398908 -15384 399248 -15298
rect 398908 -15440 398971 -15384
rect 399027 -15440 399113 -15384
rect 399169 -15440 399248 -15384
rect 398908 -15526 399248 -15440
rect 398908 -15582 398971 -15526
rect 399027 -15582 399113 -15526
rect 399169 -15582 399248 -15526
rect 398908 -15668 399248 -15582
rect 398908 -15724 398971 -15668
rect 399027 -15724 399113 -15668
rect 399169 -15724 399248 -15668
rect 398908 -15810 399248 -15724
rect 398908 -15866 398971 -15810
rect 399027 -15866 399113 -15810
rect 399169 -15866 399248 -15810
rect 398908 -15952 399248 -15866
rect 398908 -16008 398971 -15952
rect 399027 -16008 399113 -15952
rect 399169 -16008 399248 -15952
rect 398908 -16094 399248 -16008
rect 398908 -16150 398971 -16094
rect 399027 -16150 399113 -16094
rect 399169 -16150 399248 -16094
rect 398908 -16236 399248 -16150
rect 398908 -16292 398971 -16236
rect 399027 -16292 399113 -16236
rect 399169 -16292 399248 -16236
rect 398908 -16378 399248 -16292
rect 398908 -16434 398971 -16378
rect 399027 -16434 399113 -16378
rect 399169 -16434 399248 -16378
rect 398908 -16520 399248 -16434
rect 398908 -16576 398971 -16520
rect 399027 -16576 399113 -16520
rect 399169 -16576 399248 -16520
rect 398908 -16662 399248 -16576
rect 398908 -16718 398971 -16662
rect 399027 -16718 399113 -16662
rect 399169 -16718 399248 -16662
rect 398908 -16804 399248 -16718
rect 398908 -16860 398971 -16804
rect 399027 -16860 399113 -16804
rect 399169 -16860 399248 -16804
rect 398908 -16946 399248 -16860
rect 398908 -17002 398971 -16946
rect 399027 -17002 399113 -16946
rect 399169 -17002 399248 -16946
rect 398908 -17088 399248 -17002
rect 398908 -17144 398971 -17088
rect 399027 -17144 399113 -17088
rect 399169 -17144 399248 -17088
rect 398908 -17230 399248 -17144
rect 398908 -17286 398971 -17230
rect 399027 -17286 399113 -17230
rect 399169 -17286 399248 -17230
rect 398908 -17372 399248 -17286
rect 398908 -17428 398971 -17372
rect 399027 -17428 399113 -17372
rect 399169 -17428 399248 -17372
rect 398908 -17514 399248 -17428
rect 398908 -17570 398971 -17514
rect 399027 -17570 399113 -17514
rect 399169 -17570 399248 -17514
rect 398908 -17656 399248 -17570
rect 398908 -17712 398971 -17656
rect 399027 -17712 399113 -17656
rect 399169 -17712 399248 -17656
rect 398908 -17798 399248 -17712
rect 398908 -17854 398971 -17798
rect 399027 -17854 399113 -17798
rect 399169 -17854 399248 -17798
rect 398908 -17940 399248 -17854
rect 398908 -17996 398971 -17940
rect 399027 -17996 399113 -17940
rect 399169 -17996 399248 -17940
rect 398908 -18082 399248 -17996
rect 398908 -18138 398971 -18082
rect 399027 -18138 399113 -18082
rect 399169 -18138 399248 -18082
rect 398908 -18224 399248 -18138
rect 398908 -18280 398971 -18224
rect 399027 -18280 399113 -18224
rect 399169 -18280 399248 -18224
rect 398908 -18366 399248 -18280
rect 398908 -18422 398971 -18366
rect 399027 -18422 399113 -18366
rect 399169 -18422 399248 -18366
rect 398908 -18508 399248 -18422
rect 398908 -18564 398971 -18508
rect 399027 -18564 399113 -18508
rect 399169 -18564 399248 -18508
rect 398908 -18650 399248 -18564
rect 398908 -18706 398971 -18650
rect 399027 -18706 399113 -18650
rect 399169 -18706 399248 -18650
rect 398908 -18792 399248 -18706
rect 398908 -18848 398971 -18792
rect 399027 -18848 399113 -18792
rect 399169 -18848 399248 -18792
rect 398908 -18934 399248 -18848
rect 398908 -18990 398971 -18934
rect 399027 -18990 399113 -18934
rect 399169 -18990 399248 -18934
rect 398908 -19076 399248 -18990
rect 398908 -19132 398971 -19076
rect 399027 -19132 399113 -19076
rect 399169 -19132 399248 -19076
rect 398908 -19218 399248 -19132
rect 398908 -19274 398971 -19218
rect 399027 -19274 399113 -19218
rect 399169 -19274 399248 -19218
rect 398908 -19360 399248 -19274
rect 398908 -19416 398971 -19360
rect 399027 -19416 399113 -19360
rect 399169 -19416 399248 -19360
rect 398908 -19502 399248 -19416
rect 398908 -19558 398971 -19502
rect 399027 -19558 399113 -19502
rect 399169 -19558 399248 -19502
rect 398908 -19644 399248 -19558
rect 398908 -19700 398971 -19644
rect 399027 -19700 399113 -19644
rect 399169 -19700 399248 -19644
rect 398908 -19786 399248 -19700
rect 398908 -19842 398971 -19786
rect 399027 -19842 399113 -19786
rect 399169 -19842 399248 -19786
rect 398908 -19928 399248 -19842
rect 398908 -19984 398971 -19928
rect 399027 -19984 399113 -19928
rect 399169 -19984 399248 -19928
rect 398908 -20070 399248 -19984
rect 398908 -20126 398971 -20070
rect 399027 -20126 399113 -20070
rect 399169 -20126 399248 -20070
rect 398908 -20212 399248 -20126
rect 398908 -20268 398971 -20212
rect 399027 -20268 399113 -20212
rect 399169 -20268 399248 -20212
rect 398908 -20354 399248 -20268
rect 398908 -20410 398971 -20354
rect 399027 -20410 399113 -20354
rect 399169 -20410 399248 -20354
rect 398908 -20496 399248 -20410
rect 398908 -20552 398971 -20496
rect 399027 -20552 399113 -20496
rect 399169 -20552 399248 -20496
rect 398908 -20638 399248 -20552
rect 398908 -20694 398971 -20638
rect 399027 -20694 399113 -20638
rect 399169 -20694 399248 -20638
rect 398908 -20780 399248 -20694
rect 398908 -20836 398971 -20780
rect 399027 -20836 399113 -20780
rect 399169 -20836 399248 -20780
rect 398908 -20922 399248 -20836
rect 398908 -20978 398971 -20922
rect 399027 -20978 399113 -20922
rect 399169 -20978 399248 -20922
rect 398908 -21064 399248 -20978
rect 398908 -21120 398971 -21064
rect 399027 -21120 399113 -21064
rect 399169 -21120 399248 -21064
rect 398908 -21206 399248 -21120
rect 398908 -21262 398971 -21206
rect 399027 -21262 399113 -21206
rect 399169 -21262 399248 -21206
rect 398908 -21348 399248 -21262
rect 398908 -21404 398971 -21348
rect 399027 -21404 399113 -21348
rect 399169 -21404 399248 -21348
rect 398908 -21490 399248 -21404
rect 398908 -21546 398971 -21490
rect 399027 -21546 399113 -21490
rect 399169 -21546 399248 -21490
rect 398908 -21632 399248 -21546
rect 398908 -21688 398971 -21632
rect 399027 -21688 399113 -21632
rect 399169 -21688 399248 -21632
rect 398908 -21774 399248 -21688
rect 398908 -21830 398971 -21774
rect 399027 -21830 399113 -21774
rect 399169 -21830 399248 -21774
rect 398908 -21916 399248 -21830
rect 398908 -21972 398971 -21916
rect 399027 -21972 399113 -21916
rect 399169 -21972 399248 -21916
rect 398908 -22058 399248 -21972
rect 398908 -22114 398971 -22058
rect 399027 -22114 399113 -22058
rect 399169 -22114 399248 -22058
rect 398908 -22200 399248 -22114
rect 398908 -22256 398971 -22200
rect 399027 -22256 399113 -22200
rect 399169 -22256 399248 -22200
rect 398908 -22342 399248 -22256
rect 398908 -22398 398971 -22342
rect 399027 -22398 399113 -22342
rect 399169 -22398 399248 -22342
rect 398908 -22484 399248 -22398
rect 398908 -22540 398971 -22484
rect 399027 -22540 399113 -22484
rect 399169 -22540 399248 -22484
rect 398908 -22626 399248 -22540
rect 398908 -22682 398971 -22626
rect 399027 -22682 399113 -22626
rect 399169 -22682 399248 -22626
rect 398908 -22768 399248 -22682
rect 398908 -22824 398971 -22768
rect 399027 -22824 399113 -22768
rect 399169 -22824 399248 -22768
rect 398908 -22910 399248 -22824
rect 398908 -22966 398971 -22910
rect 399027 -22966 399113 -22910
rect 399169 -22966 399248 -22910
rect 398908 -23052 399248 -22966
rect 398908 -23108 398971 -23052
rect 399027 -23108 399113 -23052
rect 399169 -23108 399248 -23052
rect 398908 -23194 399248 -23108
rect 398908 -23250 398971 -23194
rect 399027 -23250 399113 -23194
rect 399169 -23250 399248 -23194
rect 398908 -23336 399248 -23250
rect 398908 -23392 398971 -23336
rect 399027 -23392 399113 -23336
rect 399169 -23392 399248 -23336
rect 398908 -23478 399248 -23392
rect 398908 -23534 398971 -23478
rect 399027 -23534 399113 -23478
rect 399169 -23534 399248 -23478
rect 398908 -23620 399248 -23534
rect 398908 -23676 398971 -23620
rect 399027 -23676 399113 -23620
rect 399169 -23676 399248 -23620
rect 398908 -23762 399248 -23676
rect 398908 -23818 398971 -23762
rect 399027 -23818 399113 -23762
rect 399169 -23818 399248 -23762
rect 398908 -23904 399248 -23818
rect 398908 -23960 398971 -23904
rect 399027 -23960 399113 -23904
rect 399169 -23960 399248 -23904
rect 398908 -24046 399248 -23960
rect 398908 -24102 398971 -24046
rect 399027 -24102 399113 -24046
rect 399169 -24102 399248 -24046
rect 398908 -24188 399248 -24102
rect 398908 -24244 398971 -24188
rect 399027 -24244 399113 -24188
rect 399169 -24244 399248 -24188
rect 398908 -24330 399248 -24244
rect 398908 -24386 398971 -24330
rect 399027 -24386 399113 -24330
rect 399169 -24386 399248 -24330
rect 398908 -24472 399248 -24386
rect 398908 -24528 398971 -24472
rect 399027 -24528 399113 -24472
rect 399169 -24528 399248 -24472
rect 398908 -24614 399248 -24528
rect 398908 -24670 398971 -24614
rect 399027 -24670 399113 -24614
rect 399169 -24670 399248 -24614
rect 398908 -24756 399248 -24670
rect 398908 -24812 398971 -24756
rect 399027 -24812 399113 -24756
rect 399169 -24812 399248 -24756
rect 398908 -24898 399248 -24812
rect 398908 -24954 398971 -24898
rect 399027 -24954 399113 -24898
rect 399169 -24954 399248 -24898
rect 398908 -25040 399248 -24954
rect 398908 -25096 398971 -25040
rect 399027 -25096 399113 -25040
rect 399169 -25096 399248 -25040
rect 398908 -25182 399248 -25096
rect 398908 -25238 398971 -25182
rect 399027 -25238 399113 -25182
rect 399169 -25238 399248 -25182
rect 398908 -25324 399248 -25238
rect 398908 -25380 398971 -25324
rect 399027 -25380 399113 -25324
rect 399169 -25380 399248 -25324
rect 398908 -25466 399248 -25380
rect 398908 -25522 398971 -25466
rect 399027 -25522 399113 -25466
rect 399169 -25522 399248 -25466
rect 398908 -25532 399248 -25522
rect 399308 -13680 399648 -13670
rect 399308 -13736 399376 -13680
rect 399432 -13736 399518 -13680
rect 399574 -13736 399648 -13680
rect 399308 -13822 399648 -13736
rect 399308 -13878 399376 -13822
rect 399432 -13878 399518 -13822
rect 399574 -13878 399648 -13822
rect 399308 -13964 399648 -13878
rect 399308 -14020 399376 -13964
rect 399432 -14020 399518 -13964
rect 399574 -14020 399648 -13964
rect 399308 -14106 399648 -14020
rect 399308 -14162 399376 -14106
rect 399432 -14162 399518 -14106
rect 399574 -14162 399648 -14106
rect 399308 -14248 399648 -14162
rect 399308 -14304 399376 -14248
rect 399432 -14304 399518 -14248
rect 399574 -14304 399648 -14248
rect 399308 -14390 399648 -14304
rect 399308 -14446 399376 -14390
rect 399432 -14446 399518 -14390
rect 399574 -14446 399648 -14390
rect 399308 -14532 399648 -14446
rect 399308 -14588 399376 -14532
rect 399432 -14588 399518 -14532
rect 399574 -14588 399648 -14532
rect 399308 -14674 399648 -14588
rect 399308 -14730 399376 -14674
rect 399432 -14730 399518 -14674
rect 399574 -14730 399648 -14674
rect 399308 -14816 399648 -14730
rect 399308 -14872 399376 -14816
rect 399432 -14872 399518 -14816
rect 399574 -14872 399648 -14816
rect 399308 -14958 399648 -14872
rect 399308 -15014 399376 -14958
rect 399432 -15014 399518 -14958
rect 399574 -15014 399648 -14958
rect 399308 -15100 399648 -15014
rect 399308 -15156 399376 -15100
rect 399432 -15156 399518 -15100
rect 399574 -15156 399648 -15100
rect 399308 -15242 399648 -15156
rect 399308 -15298 399376 -15242
rect 399432 -15298 399518 -15242
rect 399574 -15298 399648 -15242
rect 399308 -15384 399648 -15298
rect 399308 -15440 399376 -15384
rect 399432 -15440 399518 -15384
rect 399574 -15440 399648 -15384
rect 399308 -15526 399648 -15440
rect 399308 -15582 399376 -15526
rect 399432 -15582 399518 -15526
rect 399574 -15582 399648 -15526
rect 399308 -15668 399648 -15582
rect 399308 -15724 399376 -15668
rect 399432 -15724 399518 -15668
rect 399574 -15724 399648 -15668
rect 399308 -15810 399648 -15724
rect 399308 -15866 399376 -15810
rect 399432 -15866 399518 -15810
rect 399574 -15866 399648 -15810
rect 399308 -15952 399648 -15866
rect 399308 -16008 399376 -15952
rect 399432 -16008 399518 -15952
rect 399574 -16008 399648 -15952
rect 399308 -16094 399648 -16008
rect 399308 -16150 399376 -16094
rect 399432 -16150 399518 -16094
rect 399574 -16150 399648 -16094
rect 399308 -16236 399648 -16150
rect 399308 -16292 399376 -16236
rect 399432 -16292 399518 -16236
rect 399574 -16292 399648 -16236
rect 399308 -16378 399648 -16292
rect 399308 -16434 399376 -16378
rect 399432 -16434 399518 -16378
rect 399574 -16434 399648 -16378
rect 399308 -16520 399648 -16434
rect 399308 -16576 399376 -16520
rect 399432 -16576 399518 -16520
rect 399574 -16576 399648 -16520
rect 399308 -16662 399648 -16576
rect 399308 -16718 399376 -16662
rect 399432 -16718 399518 -16662
rect 399574 -16718 399648 -16662
rect 399308 -16804 399648 -16718
rect 399308 -16860 399376 -16804
rect 399432 -16860 399518 -16804
rect 399574 -16860 399648 -16804
rect 399308 -16946 399648 -16860
rect 399308 -17002 399376 -16946
rect 399432 -17002 399518 -16946
rect 399574 -17002 399648 -16946
rect 399308 -17088 399648 -17002
rect 399308 -17144 399376 -17088
rect 399432 -17144 399518 -17088
rect 399574 -17144 399648 -17088
rect 399308 -17230 399648 -17144
rect 399308 -17286 399376 -17230
rect 399432 -17286 399518 -17230
rect 399574 -17286 399648 -17230
rect 399308 -17372 399648 -17286
rect 399308 -17428 399376 -17372
rect 399432 -17428 399518 -17372
rect 399574 -17428 399648 -17372
rect 399308 -17514 399648 -17428
rect 399308 -17570 399376 -17514
rect 399432 -17570 399518 -17514
rect 399574 -17570 399648 -17514
rect 399308 -17656 399648 -17570
rect 399308 -17712 399376 -17656
rect 399432 -17712 399518 -17656
rect 399574 -17712 399648 -17656
rect 399308 -17798 399648 -17712
rect 399308 -17854 399376 -17798
rect 399432 -17854 399518 -17798
rect 399574 -17854 399648 -17798
rect 399308 -17940 399648 -17854
rect 399308 -17996 399376 -17940
rect 399432 -17996 399518 -17940
rect 399574 -17996 399648 -17940
rect 399308 -18082 399648 -17996
rect 399308 -18138 399376 -18082
rect 399432 -18138 399518 -18082
rect 399574 -18138 399648 -18082
rect 399308 -18224 399648 -18138
rect 399308 -18280 399376 -18224
rect 399432 -18280 399518 -18224
rect 399574 -18280 399648 -18224
rect 399308 -18366 399648 -18280
rect 399308 -18422 399376 -18366
rect 399432 -18422 399518 -18366
rect 399574 -18422 399648 -18366
rect 399308 -18508 399648 -18422
rect 399308 -18564 399376 -18508
rect 399432 -18564 399518 -18508
rect 399574 -18564 399648 -18508
rect 399308 -18650 399648 -18564
rect 399308 -18706 399376 -18650
rect 399432 -18706 399518 -18650
rect 399574 -18706 399648 -18650
rect 399308 -18792 399648 -18706
rect 399308 -18848 399376 -18792
rect 399432 -18848 399518 -18792
rect 399574 -18848 399648 -18792
rect 399308 -18934 399648 -18848
rect 399308 -18990 399376 -18934
rect 399432 -18990 399518 -18934
rect 399574 -18990 399648 -18934
rect 399308 -19076 399648 -18990
rect 399308 -19132 399376 -19076
rect 399432 -19132 399518 -19076
rect 399574 -19132 399648 -19076
rect 399308 -19218 399648 -19132
rect 399308 -19274 399376 -19218
rect 399432 -19274 399518 -19218
rect 399574 -19274 399648 -19218
rect 399308 -19360 399648 -19274
rect 399308 -19416 399376 -19360
rect 399432 -19416 399518 -19360
rect 399574 -19416 399648 -19360
rect 399308 -19502 399648 -19416
rect 399308 -19558 399376 -19502
rect 399432 -19558 399518 -19502
rect 399574 -19558 399648 -19502
rect 399308 -19644 399648 -19558
rect 399308 -19700 399376 -19644
rect 399432 -19700 399518 -19644
rect 399574 -19700 399648 -19644
rect 399308 -19786 399648 -19700
rect 399308 -19842 399376 -19786
rect 399432 -19842 399518 -19786
rect 399574 -19842 399648 -19786
rect 399308 -19928 399648 -19842
rect 399308 -19984 399376 -19928
rect 399432 -19984 399518 -19928
rect 399574 -19984 399648 -19928
rect 399308 -20070 399648 -19984
rect 399308 -20126 399376 -20070
rect 399432 -20126 399518 -20070
rect 399574 -20126 399648 -20070
rect 399308 -20212 399648 -20126
rect 399308 -20268 399376 -20212
rect 399432 -20268 399518 -20212
rect 399574 -20268 399648 -20212
rect 399308 -20354 399648 -20268
rect 399308 -20410 399376 -20354
rect 399432 -20410 399518 -20354
rect 399574 -20410 399648 -20354
rect 399308 -20496 399648 -20410
rect 399308 -20552 399376 -20496
rect 399432 -20552 399518 -20496
rect 399574 -20552 399648 -20496
rect 399308 -20638 399648 -20552
rect 399308 -20694 399376 -20638
rect 399432 -20694 399518 -20638
rect 399574 -20694 399648 -20638
rect 399308 -20780 399648 -20694
rect 399308 -20836 399376 -20780
rect 399432 -20836 399518 -20780
rect 399574 -20836 399648 -20780
rect 399308 -20922 399648 -20836
rect 399308 -20978 399376 -20922
rect 399432 -20978 399518 -20922
rect 399574 -20978 399648 -20922
rect 399308 -21064 399648 -20978
rect 399308 -21120 399376 -21064
rect 399432 -21120 399518 -21064
rect 399574 -21120 399648 -21064
rect 399308 -21206 399648 -21120
rect 399308 -21262 399376 -21206
rect 399432 -21262 399518 -21206
rect 399574 -21262 399648 -21206
rect 399308 -21348 399648 -21262
rect 399308 -21404 399376 -21348
rect 399432 -21404 399518 -21348
rect 399574 -21404 399648 -21348
rect 399308 -21490 399648 -21404
rect 399308 -21546 399376 -21490
rect 399432 -21546 399518 -21490
rect 399574 -21546 399648 -21490
rect 399308 -21632 399648 -21546
rect 399308 -21688 399376 -21632
rect 399432 -21688 399518 -21632
rect 399574 -21688 399648 -21632
rect 399308 -21774 399648 -21688
rect 399308 -21830 399376 -21774
rect 399432 -21830 399518 -21774
rect 399574 -21830 399648 -21774
rect 399308 -21916 399648 -21830
rect 399308 -21972 399376 -21916
rect 399432 -21972 399518 -21916
rect 399574 -21972 399648 -21916
rect 399308 -22058 399648 -21972
rect 399308 -22114 399376 -22058
rect 399432 -22114 399518 -22058
rect 399574 -22114 399648 -22058
rect 399308 -22200 399648 -22114
rect 399308 -22256 399376 -22200
rect 399432 -22256 399518 -22200
rect 399574 -22256 399648 -22200
rect 399308 -22342 399648 -22256
rect 399308 -22398 399376 -22342
rect 399432 -22398 399518 -22342
rect 399574 -22398 399648 -22342
rect 399308 -22484 399648 -22398
rect 399308 -22540 399376 -22484
rect 399432 -22540 399518 -22484
rect 399574 -22540 399648 -22484
rect 399308 -22626 399648 -22540
rect 399308 -22682 399376 -22626
rect 399432 -22682 399518 -22626
rect 399574 -22682 399648 -22626
rect 399308 -22768 399648 -22682
rect 399308 -22824 399376 -22768
rect 399432 -22824 399518 -22768
rect 399574 -22824 399648 -22768
rect 399308 -22910 399648 -22824
rect 399308 -22966 399376 -22910
rect 399432 -22966 399518 -22910
rect 399574 -22966 399648 -22910
rect 399308 -23052 399648 -22966
rect 399308 -23108 399376 -23052
rect 399432 -23108 399518 -23052
rect 399574 -23108 399648 -23052
rect 399308 -23194 399648 -23108
rect 399308 -23250 399376 -23194
rect 399432 -23250 399518 -23194
rect 399574 -23250 399648 -23194
rect 399308 -23336 399648 -23250
rect 399308 -23392 399376 -23336
rect 399432 -23392 399518 -23336
rect 399574 -23392 399648 -23336
rect 399308 -23478 399648 -23392
rect 399308 -23534 399376 -23478
rect 399432 -23534 399518 -23478
rect 399574 -23534 399648 -23478
rect 399308 -23620 399648 -23534
rect 399308 -23676 399376 -23620
rect 399432 -23676 399518 -23620
rect 399574 -23676 399648 -23620
rect 399308 -23762 399648 -23676
rect 399308 -23818 399376 -23762
rect 399432 -23818 399518 -23762
rect 399574 -23818 399648 -23762
rect 399308 -23904 399648 -23818
rect 399308 -23960 399376 -23904
rect 399432 -23960 399518 -23904
rect 399574 -23960 399648 -23904
rect 399308 -24046 399648 -23960
rect 399308 -24102 399376 -24046
rect 399432 -24102 399518 -24046
rect 399574 -24102 399648 -24046
rect 399308 -24188 399648 -24102
rect 399308 -24244 399376 -24188
rect 399432 -24244 399518 -24188
rect 399574 -24244 399648 -24188
rect 399308 -24330 399648 -24244
rect 399308 -24386 399376 -24330
rect 399432 -24386 399518 -24330
rect 399574 -24386 399648 -24330
rect 399308 -24472 399648 -24386
rect 399308 -24528 399376 -24472
rect 399432 -24528 399518 -24472
rect 399574 -24528 399648 -24472
rect 399308 -24614 399648 -24528
rect 399308 -24670 399376 -24614
rect 399432 -24670 399518 -24614
rect 399574 -24670 399648 -24614
rect 399308 -24756 399648 -24670
rect 399308 -24812 399376 -24756
rect 399432 -24812 399518 -24756
rect 399574 -24812 399648 -24756
rect 399308 -24898 399648 -24812
rect 399308 -24954 399376 -24898
rect 399432 -24954 399518 -24898
rect 399574 -24954 399648 -24898
rect 399308 -25040 399648 -24954
rect 399308 -25096 399376 -25040
rect 399432 -25096 399518 -25040
rect 399574 -25096 399648 -25040
rect 399308 -25182 399648 -25096
rect 399308 -25238 399376 -25182
rect 399432 -25238 399518 -25182
rect 399574 -25238 399648 -25182
rect 399308 -25324 399648 -25238
rect 399308 -25380 399376 -25324
rect 399432 -25380 399518 -25324
rect 399574 -25380 399648 -25324
rect 399308 -25466 399648 -25380
rect 399308 -25522 399376 -25466
rect 399432 -25522 399518 -25466
rect 399574 -25522 399648 -25466
rect 399308 -25532 399648 -25522
rect 399708 -13680 400048 -13670
rect 399708 -13736 399776 -13680
rect 399832 -13736 399918 -13680
rect 399974 -13736 400048 -13680
rect 399708 -13822 400048 -13736
rect 399708 -13878 399776 -13822
rect 399832 -13878 399918 -13822
rect 399974 -13878 400048 -13822
rect 399708 -13964 400048 -13878
rect 399708 -14020 399776 -13964
rect 399832 -14020 399918 -13964
rect 399974 -14020 400048 -13964
rect 399708 -14106 400048 -14020
rect 399708 -14162 399776 -14106
rect 399832 -14162 399918 -14106
rect 399974 -14162 400048 -14106
rect 399708 -14248 400048 -14162
rect 399708 -14304 399776 -14248
rect 399832 -14304 399918 -14248
rect 399974 -14304 400048 -14248
rect 399708 -14390 400048 -14304
rect 399708 -14446 399776 -14390
rect 399832 -14446 399918 -14390
rect 399974 -14446 400048 -14390
rect 399708 -14532 400048 -14446
rect 399708 -14588 399776 -14532
rect 399832 -14588 399918 -14532
rect 399974 -14588 400048 -14532
rect 399708 -14674 400048 -14588
rect 399708 -14730 399776 -14674
rect 399832 -14730 399918 -14674
rect 399974 -14730 400048 -14674
rect 399708 -14816 400048 -14730
rect 399708 -14872 399776 -14816
rect 399832 -14872 399918 -14816
rect 399974 -14872 400048 -14816
rect 399708 -14958 400048 -14872
rect 399708 -15014 399776 -14958
rect 399832 -15014 399918 -14958
rect 399974 -15014 400048 -14958
rect 399708 -15100 400048 -15014
rect 399708 -15156 399776 -15100
rect 399832 -15156 399918 -15100
rect 399974 -15156 400048 -15100
rect 399708 -15242 400048 -15156
rect 399708 -15298 399776 -15242
rect 399832 -15298 399918 -15242
rect 399974 -15298 400048 -15242
rect 399708 -15384 400048 -15298
rect 399708 -15440 399776 -15384
rect 399832 -15440 399918 -15384
rect 399974 -15440 400048 -15384
rect 399708 -15526 400048 -15440
rect 399708 -15582 399776 -15526
rect 399832 -15582 399918 -15526
rect 399974 -15582 400048 -15526
rect 399708 -15668 400048 -15582
rect 399708 -15724 399776 -15668
rect 399832 -15724 399918 -15668
rect 399974 -15724 400048 -15668
rect 399708 -15810 400048 -15724
rect 399708 -15866 399776 -15810
rect 399832 -15866 399918 -15810
rect 399974 -15866 400048 -15810
rect 399708 -15952 400048 -15866
rect 399708 -16008 399776 -15952
rect 399832 -16008 399918 -15952
rect 399974 -16008 400048 -15952
rect 399708 -16094 400048 -16008
rect 399708 -16150 399776 -16094
rect 399832 -16150 399918 -16094
rect 399974 -16150 400048 -16094
rect 399708 -16236 400048 -16150
rect 399708 -16292 399776 -16236
rect 399832 -16292 399918 -16236
rect 399974 -16292 400048 -16236
rect 399708 -16378 400048 -16292
rect 399708 -16434 399776 -16378
rect 399832 -16434 399918 -16378
rect 399974 -16434 400048 -16378
rect 399708 -16520 400048 -16434
rect 399708 -16576 399776 -16520
rect 399832 -16576 399918 -16520
rect 399974 -16576 400048 -16520
rect 399708 -16662 400048 -16576
rect 399708 -16718 399776 -16662
rect 399832 -16718 399918 -16662
rect 399974 -16718 400048 -16662
rect 399708 -16804 400048 -16718
rect 399708 -16860 399776 -16804
rect 399832 -16860 399918 -16804
rect 399974 -16860 400048 -16804
rect 399708 -16946 400048 -16860
rect 399708 -17002 399776 -16946
rect 399832 -17002 399918 -16946
rect 399974 -17002 400048 -16946
rect 399708 -17088 400048 -17002
rect 399708 -17144 399776 -17088
rect 399832 -17144 399918 -17088
rect 399974 -17144 400048 -17088
rect 399708 -17230 400048 -17144
rect 399708 -17286 399776 -17230
rect 399832 -17286 399918 -17230
rect 399974 -17286 400048 -17230
rect 399708 -17372 400048 -17286
rect 399708 -17428 399776 -17372
rect 399832 -17428 399918 -17372
rect 399974 -17428 400048 -17372
rect 399708 -17514 400048 -17428
rect 399708 -17570 399776 -17514
rect 399832 -17570 399918 -17514
rect 399974 -17570 400048 -17514
rect 399708 -17656 400048 -17570
rect 399708 -17712 399776 -17656
rect 399832 -17712 399918 -17656
rect 399974 -17712 400048 -17656
rect 399708 -17798 400048 -17712
rect 399708 -17854 399776 -17798
rect 399832 -17854 399918 -17798
rect 399974 -17854 400048 -17798
rect 399708 -17940 400048 -17854
rect 399708 -17996 399776 -17940
rect 399832 -17996 399918 -17940
rect 399974 -17996 400048 -17940
rect 399708 -18082 400048 -17996
rect 399708 -18138 399776 -18082
rect 399832 -18138 399918 -18082
rect 399974 -18138 400048 -18082
rect 399708 -18224 400048 -18138
rect 399708 -18280 399776 -18224
rect 399832 -18280 399918 -18224
rect 399974 -18280 400048 -18224
rect 399708 -18366 400048 -18280
rect 399708 -18422 399776 -18366
rect 399832 -18422 399918 -18366
rect 399974 -18422 400048 -18366
rect 399708 -18508 400048 -18422
rect 399708 -18564 399776 -18508
rect 399832 -18564 399918 -18508
rect 399974 -18564 400048 -18508
rect 399708 -18650 400048 -18564
rect 399708 -18706 399776 -18650
rect 399832 -18706 399918 -18650
rect 399974 -18706 400048 -18650
rect 399708 -18792 400048 -18706
rect 399708 -18848 399776 -18792
rect 399832 -18848 399918 -18792
rect 399974 -18848 400048 -18792
rect 399708 -18934 400048 -18848
rect 399708 -18990 399776 -18934
rect 399832 -18990 399918 -18934
rect 399974 -18990 400048 -18934
rect 399708 -19076 400048 -18990
rect 399708 -19132 399776 -19076
rect 399832 -19132 399918 -19076
rect 399974 -19132 400048 -19076
rect 399708 -19218 400048 -19132
rect 399708 -19274 399776 -19218
rect 399832 -19274 399918 -19218
rect 399974 -19274 400048 -19218
rect 399708 -19360 400048 -19274
rect 399708 -19416 399776 -19360
rect 399832 -19416 399918 -19360
rect 399974 -19416 400048 -19360
rect 399708 -19502 400048 -19416
rect 399708 -19558 399776 -19502
rect 399832 -19558 399918 -19502
rect 399974 -19558 400048 -19502
rect 399708 -19644 400048 -19558
rect 399708 -19700 399776 -19644
rect 399832 -19700 399918 -19644
rect 399974 -19700 400048 -19644
rect 399708 -19786 400048 -19700
rect 399708 -19842 399776 -19786
rect 399832 -19842 399918 -19786
rect 399974 -19842 400048 -19786
rect 399708 -19928 400048 -19842
rect 399708 -19984 399776 -19928
rect 399832 -19984 399918 -19928
rect 399974 -19984 400048 -19928
rect 399708 -20070 400048 -19984
rect 399708 -20126 399776 -20070
rect 399832 -20126 399918 -20070
rect 399974 -20126 400048 -20070
rect 399708 -20212 400048 -20126
rect 399708 -20268 399776 -20212
rect 399832 -20268 399918 -20212
rect 399974 -20268 400048 -20212
rect 399708 -20354 400048 -20268
rect 399708 -20410 399776 -20354
rect 399832 -20410 399918 -20354
rect 399974 -20410 400048 -20354
rect 399708 -20496 400048 -20410
rect 399708 -20552 399776 -20496
rect 399832 -20552 399918 -20496
rect 399974 -20552 400048 -20496
rect 399708 -20638 400048 -20552
rect 399708 -20694 399776 -20638
rect 399832 -20694 399918 -20638
rect 399974 -20694 400048 -20638
rect 399708 -20780 400048 -20694
rect 399708 -20836 399776 -20780
rect 399832 -20836 399918 -20780
rect 399974 -20836 400048 -20780
rect 399708 -20922 400048 -20836
rect 399708 -20978 399776 -20922
rect 399832 -20978 399918 -20922
rect 399974 -20978 400048 -20922
rect 399708 -21064 400048 -20978
rect 399708 -21120 399776 -21064
rect 399832 -21120 399918 -21064
rect 399974 -21120 400048 -21064
rect 399708 -21206 400048 -21120
rect 399708 -21262 399776 -21206
rect 399832 -21262 399918 -21206
rect 399974 -21262 400048 -21206
rect 399708 -21348 400048 -21262
rect 399708 -21404 399776 -21348
rect 399832 -21404 399918 -21348
rect 399974 -21404 400048 -21348
rect 399708 -21490 400048 -21404
rect 399708 -21546 399776 -21490
rect 399832 -21546 399918 -21490
rect 399974 -21546 400048 -21490
rect 399708 -21632 400048 -21546
rect 399708 -21688 399776 -21632
rect 399832 -21688 399918 -21632
rect 399974 -21688 400048 -21632
rect 399708 -21774 400048 -21688
rect 399708 -21830 399776 -21774
rect 399832 -21830 399918 -21774
rect 399974 -21830 400048 -21774
rect 399708 -21916 400048 -21830
rect 399708 -21972 399776 -21916
rect 399832 -21972 399918 -21916
rect 399974 -21972 400048 -21916
rect 399708 -22058 400048 -21972
rect 399708 -22114 399776 -22058
rect 399832 -22114 399918 -22058
rect 399974 -22114 400048 -22058
rect 399708 -22200 400048 -22114
rect 399708 -22256 399776 -22200
rect 399832 -22256 399918 -22200
rect 399974 -22256 400048 -22200
rect 399708 -22342 400048 -22256
rect 399708 -22398 399776 -22342
rect 399832 -22398 399918 -22342
rect 399974 -22398 400048 -22342
rect 399708 -22484 400048 -22398
rect 399708 -22540 399776 -22484
rect 399832 -22540 399918 -22484
rect 399974 -22540 400048 -22484
rect 399708 -22626 400048 -22540
rect 399708 -22682 399776 -22626
rect 399832 -22682 399918 -22626
rect 399974 -22682 400048 -22626
rect 399708 -22768 400048 -22682
rect 399708 -22824 399776 -22768
rect 399832 -22824 399918 -22768
rect 399974 -22824 400048 -22768
rect 399708 -22910 400048 -22824
rect 399708 -22966 399776 -22910
rect 399832 -22966 399918 -22910
rect 399974 -22966 400048 -22910
rect 399708 -23052 400048 -22966
rect 399708 -23108 399776 -23052
rect 399832 -23108 399918 -23052
rect 399974 -23108 400048 -23052
rect 399708 -23194 400048 -23108
rect 399708 -23250 399776 -23194
rect 399832 -23250 399918 -23194
rect 399974 -23250 400048 -23194
rect 399708 -23336 400048 -23250
rect 399708 -23392 399776 -23336
rect 399832 -23392 399918 -23336
rect 399974 -23392 400048 -23336
rect 399708 -23478 400048 -23392
rect 399708 -23534 399776 -23478
rect 399832 -23534 399918 -23478
rect 399974 -23534 400048 -23478
rect 399708 -23620 400048 -23534
rect 399708 -23676 399776 -23620
rect 399832 -23676 399918 -23620
rect 399974 -23676 400048 -23620
rect 399708 -23762 400048 -23676
rect 399708 -23818 399776 -23762
rect 399832 -23818 399918 -23762
rect 399974 -23818 400048 -23762
rect 399708 -23904 400048 -23818
rect 399708 -23960 399776 -23904
rect 399832 -23960 399918 -23904
rect 399974 -23960 400048 -23904
rect 399708 -24046 400048 -23960
rect 399708 -24102 399776 -24046
rect 399832 -24102 399918 -24046
rect 399974 -24102 400048 -24046
rect 399708 -24188 400048 -24102
rect 399708 -24244 399776 -24188
rect 399832 -24244 399918 -24188
rect 399974 -24244 400048 -24188
rect 399708 -24330 400048 -24244
rect 399708 -24386 399776 -24330
rect 399832 -24386 399918 -24330
rect 399974 -24386 400048 -24330
rect 399708 -24472 400048 -24386
rect 399708 -24528 399776 -24472
rect 399832 -24528 399918 -24472
rect 399974 -24528 400048 -24472
rect 399708 -24614 400048 -24528
rect 399708 -24670 399776 -24614
rect 399832 -24670 399918 -24614
rect 399974 -24670 400048 -24614
rect 399708 -24756 400048 -24670
rect 399708 -24812 399776 -24756
rect 399832 -24812 399918 -24756
rect 399974 -24812 400048 -24756
rect 399708 -24898 400048 -24812
rect 399708 -24954 399776 -24898
rect 399832 -24954 399918 -24898
rect 399974 -24954 400048 -24898
rect 399708 -25040 400048 -24954
rect 399708 -25096 399776 -25040
rect 399832 -25096 399918 -25040
rect 399974 -25096 400048 -25040
rect 399708 -25182 400048 -25096
rect 399708 -25238 399776 -25182
rect 399832 -25238 399918 -25182
rect 399974 -25238 400048 -25182
rect 399708 -25324 400048 -25238
rect 399708 -25380 399776 -25324
rect 399832 -25380 399918 -25324
rect 399974 -25380 400048 -25324
rect 399708 -25466 400048 -25380
rect 399708 -25522 399776 -25466
rect 399832 -25522 399918 -25466
rect 399974 -25522 400048 -25466
rect 399708 -25532 400048 -25522
rect 400108 -13680 400448 -13670
rect 400108 -13736 400181 -13680
rect 400237 -13736 400323 -13680
rect 400379 -13736 400448 -13680
rect 400108 -13822 400448 -13736
rect 400108 -13878 400181 -13822
rect 400237 -13878 400323 -13822
rect 400379 -13878 400448 -13822
rect 400108 -13964 400448 -13878
rect 400108 -14020 400181 -13964
rect 400237 -14020 400323 -13964
rect 400379 -14020 400448 -13964
rect 400108 -14106 400448 -14020
rect 400108 -14162 400181 -14106
rect 400237 -14162 400323 -14106
rect 400379 -14162 400448 -14106
rect 400108 -14248 400448 -14162
rect 400108 -14304 400181 -14248
rect 400237 -14304 400323 -14248
rect 400379 -14304 400448 -14248
rect 400108 -14390 400448 -14304
rect 400108 -14446 400181 -14390
rect 400237 -14446 400323 -14390
rect 400379 -14446 400448 -14390
rect 400108 -14532 400448 -14446
rect 400108 -14588 400181 -14532
rect 400237 -14588 400323 -14532
rect 400379 -14588 400448 -14532
rect 400108 -14674 400448 -14588
rect 400108 -14730 400181 -14674
rect 400237 -14730 400323 -14674
rect 400379 -14730 400448 -14674
rect 400108 -14816 400448 -14730
rect 400108 -14872 400181 -14816
rect 400237 -14872 400323 -14816
rect 400379 -14872 400448 -14816
rect 400108 -14958 400448 -14872
rect 400108 -15014 400181 -14958
rect 400237 -15014 400323 -14958
rect 400379 -15014 400448 -14958
rect 400108 -15100 400448 -15014
rect 400108 -15156 400181 -15100
rect 400237 -15156 400323 -15100
rect 400379 -15156 400448 -15100
rect 400108 -15242 400448 -15156
rect 400108 -15298 400181 -15242
rect 400237 -15298 400323 -15242
rect 400379 -15298 400448 -15242
rect 400108 -15384 400448 -15298
rect 400108 -15440 400181 -15384
rect 400237 -15440 400323 -15384
rect 400379 -15440 400448 -15384
rect 400108 -15526 400448 -15440
rect 400108 -15582 400181 -15526
rect 400237 -15582 400323 -15526
rect 400379 -15582 400448 -15526
rect 400108 -15668 400448 -15582
rect 400108 -15724 400181 -15668
rect 400237 -15724 400323 -15668
rect 400379 -15724 400448 -15668
rect 400108 -15810 400448 -15724
rect 400108 -15866 400181 -15810
rect 400237 -15866 400323 -15810
rect 400379 -15866 400448 -15810
rect 400108 -15952 400448 -15866
rect 400108 -16008 400181 -15952
rect 400237 -16008 400323 -15952
rect 400379 -16008 400448 -15952
rect 400108 -16094 400448 -16008
rect 400108 -16150 400181 -16094
rect 400237 -16150 400323 -16094
rect 400379 -16150 400448 -16094
rect 400108 -16236 400448 -16150
rect 400108 -16292 400181 -16236
rect 400237 -16292 400323 -16236
rect 400379 -16292 400448 -16236
rect 400108 -16378 400448 -16292
rect 400108 -16434 400181 -16378
rect 400237 -16434 400323 -16378
rect 400379 -16434 400448 -16378
rect 400108 -16520 400448 -16434
rect 400108 -16576 400181 -16520
rect 400237 -16576 400323 -16520
rect 400379 -16576 400448 -16520
rect 400108 -16662 400448 -16576
rect 400108 -16718 400181 -16662
rect 400237 -16718 400323 -16662
rect 400379 -16718 400448 -16662
rect 400108 -16804 400448 -16718
rect 400108 -16860 400181 -16804
rect 400237 -16860 400323 -16804
rect 400379 -16860 400448 -16804
rect 400108 -16946 400448 -16860
rect 400108 -17002 400181 -16946
rect 400237 -17002 400323 -16946
rect 400379 -17002 400448 -16946
rect 400108 -17088 400448 -17002
rect 400108 -17144 400181 -17088
rect 400237 -17144 400323 -17088
rect 400379 -17144 400448 -17088
rect 400108 -17230 400448 -17144
rect 400108 -17286 400181 -17230
rect 400237 -17286 400323 -17230
rect 400379 -17286 400448 -17230
rect 400108 -17372 400448 -17286
rect 400108 -17428 400181 -17372
rect 400237 -17428 400323 -17372
rect 400379 -17428 400448 -17372
rect 400108 -17514 400448 -17428
rect 400108 -17570 400181 -17514
rect 400237 -17570 400323 -17514
rect 400379 -17570 400448 -17514
rect 400108 -17656 400448 -17570
rect 400108 -17712 400181 -17656
rect 400237 -17712 400323 -17656
rect 400379 -17712 400448 -17656
rect 400108 -17798 400448 -17712
rect 400108 -17854 400181 -17798
rect 400237 -17854 400323 -17798
rect 400379 -17854 400448 -17798
rect 400108 -17940 400448 -17854
rect 400108 -17996 400181 -17940
rect 400237 -17996 400323 -17940
rect 400379 -17996 400448 -17940
rect 400108 -18082 400448 -17996
rect 400108 -18138 400181 -18082
rect 400237 -18138 400323 -18082
rect 400379 -18138 400448 -18082
rect 400108 -18224 400448 -18138
rect 400108 -18280 400181 -18224
rect 400237 -18280 400323 -18224
rect 400379 -18280 400448 -18224
rect 400108 -18366 400448 -18280
rect 400108 -18422 400181 -18366
rect 400237 -18422 400323 -18366
rect 400379 -18422 400448 -18366
rect 400108 -18508 400448 -18422
rect 400108 -18564 400181 -18508
rect 400237 -18564 400323 -18508
rect 400379 -18564 400448 -18508
rect 400108 -18650 400448 -18564
rect 400108 -18706 400181 -18650
rect 400237 -18706 400323 -18650
rect 400379 -18706 400448 -18650
rect 400108 -18792 400448 -18706
rect 400108 -18848 400181 -18792
rect 400237 -18848 400323 -18792
rect 400379 -18848 400448 -18792
rect 400108 -18934 400448 -18848
rect 400108 -18990 400181 -18934
rect 400237 -18990 400323 -18934
rect 400379 -18990 400448 -18934
rect 400108 -19076 400448 -18990
rect 400108 -19132 400181 -19076
rect 400237 -19132 400323 -19076
rect 400379 -19132 400448 -19076
rect 400108 -19218 400448 -19132
rect 400108 -19274 400181 -19218
rect 400237 -19274 400323 -19218
rect 400379 -19274 400448 -19218
rect 400108 -19360 400448 -19274
rect 400108 -19416 400181 -19360
rect 400237 -19416 400323 -19360
rect 400379 -19416 400448 -19360
rect 400108 -19502 400448 -19416
rect 400108 -19558 400181 -19502
rect 400237 -19558 400323 -19502
rect 400379 -19558 400448 -19502
rect 400108 -19644 400448 -19558
rect 400108 -19700 400181 -19644
rect 400237 -19700 400323 -19644
rect 400379 -19700 400448 -19644
rect 400108 -19786 400448 -19700
rect 400108 -19842 400181 -19786
rect 400237 -19842 400323 -19786
rect 400379 -19842 400448 -19786
rect 400108 -19928 400448 -19842
rect 400108 -19984 400181 -19928
rect 400237 -19984 400323 -19928
rect 400379 -19984 400448 -19928
rect 400108 -20070 400448 -19984
rect 400108 -20126 400181 -20070
rect 400237 -20126 400323 -20070
rect 400379 -20126 400448 -20070
rect 400108 -20212 400448 -20126
rect 400108 -20268 400181 -20212
rect 400237 -20268 400323 -20212
rect 400379 -20268 400448 -20212
rect 400108 -20354 400448 -20268
rect 400108 -20410 400181 -20354
rect 400237 -20410 400323 -20354
rect 400379 -20410 400448 -20354
rect 400108 -20496 400448 -20410
rect 400108 -20552 400181 -20496
rect 400237 -20552 400323 -20496
rect 400379 -20552 400448 -20496
rect 400108 -20638 400448 -20552
rect 400108 -20694 400181 -20638
rect 400237 -20694 400323 -20638
rect 400379 -20694 400448 -20638
rect 400108 -20780 400448 -20694
rect 400108 -20836 400181 -20780
rect 400237 -20836 400323 -20780
rect 400379 -20836 400448 -20780
rect 400108 -20922 400448 -20836
rect 400108 -20978 400181 -20922
rect 400237 -20978 400323 -20922
rect 400379 -20978 400448 -20922
rect 400108 -21064 400448 -20978
rect 400108 -21120 400181 -21064
rect 400237 -21120 400323 -21064
rect 400379 -21120 400448 -21064
rect 400108 -21206 400448 -21120
rect 400108 -21262 400181 -21206
rect 400237 -21262 400323 -21206
rect 400379 -21262 400448 -21206
rect 400108 -21348 400448 -21262
rect 400108 -21404 400181 -21348
rect 400237 -21404 400323 -21348
rect 400379 -21404 400448 -21348
rect 400108 -21490 400448 -21404
rect 400108 -21546 400181 -21490
rect 400237 -21546 400323 -21490
rect 400379 -21546 400448 -21490
rect 400108 -21632 400448 -21546
rect 400108 -21688 400181 -21632
rect 400237 -21688 400323 -21632
rect 400379 -21688 400448 -21632
rect 400108 -21774 400448 -21688
rect 400108 -21830 400181 -21774
rect 400237 -21830 400323 -21774
rect 400379 -21830 400448 -21774
rect 400108 -21916 400448 -21830
rect 400108 -21972 400181 -21916
rect 400237 -21972 400323 -21916
rect 400379 -21972 400448 -21916
rect 400108 -22058 400448 -21972
rect 400108 -22114 400181 -22058
rect 400237 -22114 400323 -22058
rect 400379 -22114 400448 -22058
rect 400108 -22200 400448 -22114
rect 400108 -22256 400181 -22200
rect 400237 -22256 400323 -22200
rect 400379 -22256 400448 -22200
rect 400108 -22342 400448 -22256
rect 400108 -22398 400181 -22342
rect 400237 -22398 400323 -22342
rect 400379 -22398 400448 -22342
rect 400108 -22484 400448 -22398
rect 400108 -22540 400181 -22484
rect 400237 -22540 400323 -22484
rect 400379 -22540 400448 -22484
rect 400108 -22626 400448 -22540
rect 400108 -22682 400181 -22626
rect 400237 -22682 400323 -22626
rect 400379 -22682 400448 -22626
rect 400108 -22768 400448 -22682
rect 400108 -22824 400181 -22768
rect 400237 -22824 400323 -22768
rect 400379 -22824 400448 -22768
rect 400108 -22910 400448 -22824
rect 400108 -22966 400181 -22910
rect 400237 -22966 400323 -22910
rect 400379 -22966 400448 -22910
rect 400108 -23052 400448 -22966
rect 400108 -23108 400181 -23052
rect 400237 -23108 400323 -23052
rect 400379 -23108 400448 -23052
rect 400108 -23194 400448 -23108
rect 400108 -23250 400181 -23194
rect 400237 -23250 400323 -23194
rect 400379 -23250 400448 -23194
rect 400108 -23336 400448 -23250
rect 400108 -23392 400181 -23336
rect 400237 -23392 400323 -23336
rect 400379 -23392 400448 -23336
rect 400108 -23478 400448 -23392
rect 400108 -23534 400181 -23478
rect 400237 -23534 400323 -23478
rect 400379 -23534 400448 -23478
rect 400108 -23620 400448 -23534
rect 400108 -23676 400181 -23620
rect 400237 -23676 400323 -23620
rect 400379 -23676 400448 -23620
rect 400108 -23762 400448 -23676
rect 400108 -23818 400181 -23762
rect 400237 -23818 400323 -23762
rect 400379 -23818 400448 -23762
rect 400108 -23904 400448 -23818
rect 400108 -23960 400181 -23904
rect 400237 -23960 400323 -23904
rect 400379 -23960 400448 -23904
rect 400108 -24046 400448 -23960
rect 400108 -24102 400181 -24046
rect 400237 -24102 400323 -24046
rect 400379 -24102 400448 -24046
rect 400108 -24188 400448 -24102
rect 400108 -24244 400181 -24188
rect 400237 -24244 400323 -24188
rect 400379 -24244 400448 -24188
rect 400108 -24330 400448 -24244
rect 400108 -24386 400181 -24330
rect 400237 -24386 400323 -24330
rect 400379 -24386 400448 -24330
rect 400108 -24472 400448 -24386
rect 400108 -24528 400181 -24472
rect 400237 -24528 400323 -24472
rect 400379 -24528 400448 -24472
rect 400108 -24614 400448 -24528
rect 400108 -24670 400181 -24614
rect 400237 -24670 400323 -24614
rect 400379 -24670 400448 -24614
rect 400108 -24756 400448 -24670
rect 400108 -24812 400181 -24756
rect 400237 -24812 400323 -24756
rect 400379 -24812 400448 -24756
rect 400108 -24898 400448 -24812
rect 400108 -24954 400181 -24898
rect 400237 -24954 400323 -24898
rect 400379 -24954 400448 -24898
rect 400108 -25040 400448 -24954
rect 400108 -25096 400181 -25040
rect 400237 -25096 400323 -25040
rect 400379 -25096 400448 -25040
rect 400108 -25182 400448 -25096
rect 400108 -25238 400181 -25182
rect 400237 -25238 400323 -25182
rect 400379 -25238 400448 -25182
rect 400108 -25324 400448 -25238
rect 400108 -25380 400181 -25324
rect 400237 -25380 400323 -25324
rect 400379 -25380 400448 -25324
rect 400108 -25466 400448 -25380
rect 400108 -25522 400181 -25466
rect 400237 -25522 400323 -25466
rect 400379 -25522 400448 -25466
rect 400108 -25532 400448 -25522
rect 400640 -13688 400766 -13670
rect 400822 -13688 400890 -13632
rect 400946 -13688 401014 -13632
rect 401070 -13688 401138 -13632
rect 401194 -13688 401262 -13632
rect 401318 -13688 401440 -13632
rect 400640 -13756 401440 -13688
rect 400640 -13812 400766 -13756
rect 400822 -13812 400890 -13756
rect 400946 -13812 401014 -13756
rect 401070 -13812 401138 -13756
rect 401194 -13812 401262 -13756
rect 401318 -13812 401440 -13756
rect 400640 -13880 401440 -13812
rect 400640 -13936 400766 -13880
rect 400822 -13936 400890 -13880
rect 400946 -13936 401014 -13880
rect 401070 -13936 401138 -13880
rect 401194 -13936 401262 -13880
rect 401318 -13936 401440 -13880
rect 400640 -14004 401440 -13936
rect 400640 -14060 400766 -14004
rect 400822 -14060 400890 -14004
rect 400946 -14060 401014 -14004
rect 401070 -14060 401138 -14004
rect 401194 -14060 401262 -14004
rect 401318 -14060 401440 -14004
rect 400640 -14128 401440 -14060
rect 400640 -14184 400766 -14128
rect 400822 -14184 400890 -14128
rect 400946 -14184 401014 -14128
rect 401070 -14184 401138 -14128
rect 401194 -14184 401262 -14128
rect 401318 -14184 401440 -14128
rect 400640 -14252 401440 -14184
rect 400640 -14308 400766 -14252
rect 400822 -14308 400890 -14252
rect 400946 -14308 401014 -14252
rect 401070 -14308 401138 -14252
rect 401194 -14308 401262 -14252
rect 401318 -14308 401440 -14252
rect 400640 -14376 401440 -14308
rect 400640 -14432 400766 -14376
rect 400822 -14432 400890 -14376
rect 400946 -14432 401014 -14376
rect 401070 -14432 401138 -14376
rect 401194 -14432 401262 -14376
rect 401318 -14432 401440 -14376
rect 400640 -14500 401440 -14432
rect 400640 -14556 400766 -14500
rect 400822 -14556 400890 -14500
rect 400946 -14556 401014 -14500
rect 401070 -14556 401138 -14500
rect 401194 -14556 401262 -14500
rect 401318 -14556 401440 -14500
rect 400640 -14624 401440 -14556
rect 400640 -14680 400766 -14624
rect 400822 -14680 400890 -14624
rect 400946 -14680 401014 -14624
rect 401070 -14680 401138 -14624
rect 401194 -14680 401262 -14624
rect 401318 -14680 401440 -14624
rect 400640 -14748 401440 -14680
rect 400640 -14804 400766 -14748
rect 400822 -14804 400890 -14748
rect 400946 -14804 401014 -14748
rect 401070 -14804 401138 -14748
rect 401194 -14804 401262 -14748
rect 401318 -14804 401440 -14748
rect 400640 -14872 401440 -14804
rect 400640 -14928 400766 -14872
rect 400822 -14928 400890 -14872
rect 400946 -14928 401014 -14872
rect 401070 -14928 401138 -14872
rect 401194 -14928 401262 -14872
rect 401318 -14928 401440 -14872
rect 400640 -14996 401440 -14928
rect 400640 -15052 400766 -14996
rect 400822 -15052 400890 -14996
rect 400946 -15052 401014 -14996
rect 401070 -15052 401138 -14996
rect 401194 -15052 401262 -14996
rect 401318 -15052 401440 -14996
rect 400640 -15120 401440 -15052
rect 400640 -15176 400766 -15120
rect 400822 -15176 400890 -15120
rect 400946 -15176 401014 -15120
rect 401070 -15176 401138 -15120
rect 401194 -15176 401262 -15120
rect 401318 -15176 401440 -15120
rect 400640 -15244 401440 -15176
rect 400640 -15300 400766 -15244
rect 400822 -15300 400890 -15244
rect 400946 -15300 401014 -15244
rect 401070 -15300 401138 -15244
rect 401194 -15300 401262 -15244
rect 401318 -15300 401440 -15244
rect 400640 -15368 401440 -15300
rect 400640 -15424 400766 -15368
rect 400822 -15424 400890 -15368
rect 400946 -15424 401014 -15368
rect 401070 -15424 401138 -15368
rect 401194 -15424 401262 -15368
rect 401318 -15424 401440 -15368
rect 400640 -15492 401440 -15424
rect 400640 -15548 400766 -15492
rect 400822 -15548 400890 -15492
rect 400946 -15548 401014 -15492
rect 401070 -15548 401138 -15492
rect 401194 -15548 401262 -15492
rect 401318 -15548 401440 -15492
rect 400640 -15616 401440 -15548
rect 400640 -15672 400766 -15616
rect 400822 -15672 400890 -15616
rect 400946 -15672 401014 -15616
rect 401070 -15672 401138 -15616
rect 401194 -15672 401262 -15616
rect 401318 -15672 401440 -15616
rect 400640 -15740 401440 -15672
rect 400640 -15796 400766 -15740
rect 400822 -15796 400890 -15740
rect 400946 -15796 401014 -15740
rect 401070 -15796 401138 -15740
rect 401194 -15796 401262 -15740
rect 401318 -15796 401440 -15740
rect 400640 -15864 401440 -15796
rect 400640 -15920 400766 -15864
rect 400822 -15920 400890 -15864
rect 400946 -15920 401014 -15864
rect 401070 -15920 401138 -15864
rect 401194 -15920 401262 -15864
rect 401318 -15920 401440 -15864
rect 400640 -15988 401440 -15920
rect 400640 -16044 400766 -15988
rect 400822 -16044 400890 -15988
rect 400946 -16044 401014 -15988
rect 401070 -16044 401138 -15988
rect 401194 -16044 401262 -15988
rect 401318 -16044 401440 -15988
rect 400640 -16112 401440 -16044
rect 400640 -16168 400766 -16112
rect 400822 -16168 400890 -16112
rect 400946 -16168 401014 -16112
rect 401070 -16168 401138 -16112
rect 401194 -16168 401262 -16112
rect 401318 -16168 401440 -16112
rect 400640 -16236 401440 -16168
rect 400640 -16292 400766 -16236
rect 400822 -16292 400890 -16236
rect 400946 -16292 401014 -16236
rect 401070 -16292 401138 -16236
rect 401194 -16292 401262 -16236
rect 401318 -16292 401440 -16236
rect 400640 -16360 401440 -16292
rect 400640 -16416 400766 -16360
rect 400822 -16416 400890 -16360
rect 400946 -16416 401014 -16360
rect 401070 -16416 401138 -16360
rect 401194 -16416 401262 -16360
rect 401318 -16416 401440 -16360
rect 400640 -16484 401440 -16416
rect 400640 -16540 400766 -16484
rect 400822 -16540 400890 -16484
rect 400946 -16540 401014 -16484
rect 401070 -16540 401138 -16484
rect 401194 -16540 401262 -16484
rect 401318 -16540 401440 -16484
rect 400640 -16608 401440 -16540
rect 400640 -16664 400766 -16608
rect 400822 -16664 400890 -16608
rect 400946 -16664 401014 -16608
rect 401070 -16664 401138 -16608
rect 401194 -16664 401262 -16608
rect 401318 -16664 401440 -16608
rect 400640 -16732 401440 -16664
rect 400640 -16788 400766 -16732
rect 400822 -16788 400890 -16732
rect 400946 -16788 401014 -16732
rect 401070 -16788 401138 -16732
rect 401194 -16788 401262 -16732
rect 401318 -16788 401440 -16732
rect 400640 -16856 401440 -16788
rect 400640 -16912 400766 -16856
rect 400822 -16912 400890 -16856
rect 400946 -16912 401014 -16856
rect 401070 -16912 401138 -16856
rect 401194 -16912 401262 -16856
rect 401318 -16912 401440 -16856
rect 400640 -16980 401440 -16912
rect 400640 -17036 400766 -16980
rect 400822 -17036 400890 -16980
rect 400946 -17036 401014 -16980
rect 401070 -17036 401138 -16980
rect 401194 -17036 401262 -16980
rect 401318 -17036 401440 -16980
rect 400640 -17104 401440 -17036
rect 400640 -17160 400766 -17104
rect 400822 -17160 400890 -17104
rect 400946 -17160 401014 -17104
rect 401070 -17160 401138 -17104
rect 401194 -17160 401262 -17104
rect 401318 -17160 401440 -17104
rect 400640 -17228 401440 -17160
rect 400640 -17284 400766 -17228
rect 400822 -17284 400890 -17228
rect 400946 -17284 401014 -17228
rect 401070 -17284 401138 -17228
rect 401194 -17284 401262 -17228
rect 401318 -17284 401440 -17228
rect 400640 -17352 401440 -17284
rect 400640 -17408 400766 -17352
rect 400822 -17408 400890 -17352
rect 400946 -17408 401014 -17352
rect 401070 -17408 401138 -17352
rect 401194 -17408 401262 -17352
rect 401318 -17408 401440 -17352
rect 400640 -17476 401440 -17408
rect 400640 -17532 400766 -17476
rect 400822 -17532 400890 -17476
rect 400946 -17532 401014 -17476
rect 401070 -17532 401138 -17476
rect 401194 -17532 401262 -17476
rect 401318 -17532 401440 -17476
rect 400640 -17600 401440 -17532
rect 400640 -17656 400766 -17600
rect 400822 -17656 400890 -17600
rect 400946 -17656 401014 -17600
rect 401070 -17656 401138 -17600
rect 401194 -17656 401262 -17600
rect 401318 -17656 401440 -17600
rect 400640 -17724 401440 -17656
rect 400640 -17780 400766 -17724
rect 400822 -17780 400890 -17724
rect 400946 -17780 401014 -17724
rect 401070 -17780 401138 -17724
rect 401194 -17780 401262 -17724
rect 401318 -17780 401440 -17724
rect 400640 -17848 401440 -17780
rect 400640 -17904 400766 -17848
rect 400822 -17904 400890 -17848
rect 400946 -17904 401014 -17848
rect 401070 -17904 401138 -17848
rect 401194 -17904 401262 -17848
rect 401318 -17904 401440 -17848
rect 400640 -17972 401440 -17904
rect 400640 -18028 400766 -17972
rect 400822 -18028 400890 -17972
rect 400946 -18028 401014 -17972
rect 401070 -18028 401138 -17972
rect 401194 -18028 401262 -17972
rect 401318 -18028 401440 -17972
rect 400640 -18096 401440 -18028
rect 400640 -18152 400766 -18096
rect 400822 -18152 400890 -18096
rect 400946 -18152 401014 -18096
rect 401070 -18152 401138 -18096
rect 401194 -18152 401262 -18096
rect 401318 -18152 401440 -18096
rect 400640 -18220 401440 -18152
rect 400640 -18276 400766 -18220
rect 400822 -18276 400890 -18220
rect 400946 -18276 401014 -18220
rect 401070 -18276 401138 -18220
rect 401194 -18276 401262 -18220
rect 401318 -18276 401440 -18220
rect 400640 -18344 401440 -18276
rect 400640 -18400 400766 -18344
rect 400822 -18400 400890 -18344
rect 400946 -18400 401014 -18344
rect 401070 -18400 401138 -18344
rect 401194 -18400 401262 -18344
rect 401318 -18400 401440 -18344
rect 400640 -18468 401440 -18400
rect 400640 -18524 400766 -18468
rect 400822 -18524 400890 -18468
rect 400946 -18524 401014 -18468
rect 401070 -18524 401138 -18468
rect 401194 -18524 401262 -18468
rect 401318 -18524 401440 -18468
rect 400640 -18592 401440 -18524
rect 400640 -18648 400766 -18592
rect 400822 -18648 400890 -18592
rect 400946 -18648 401014 -18592
rect 401070 -18648 401138 -18592
rect 401194 -18648 401262 -18592
rect 401318 -18648 401440 -18592
rect 400640 -18716 401440 -18648
rect 400640 -18772 400766 -18716
rect 400822 -18772 400890 -18716
rect 400946 -18772 401014 -18716
rect 401070 -18772 401138 -18716
rect 401194 -18772 401262 -18716
rect 401318 -18772 401440 -18716
rect 400640 -18840 401440 -18772
rect 400640 -18896 400766 -18840
rect 400822 -18896 400890 -18840
rect 400946 -18896 401014 -18840
rect 401070 -18896 401138 -18840
rect 401194 -18896 401262 -18840
rect 401318 -18896 401440 -18840
rect 400640 -18964 401440 -18896
rect 400640 -19020 400766 -18964
rect 400822 -19020 400890 -18964
rect 400946 -19020 401014 -18964
rect 401070 -19020 401138 -18964
rect 401194 -19020 401262 -18964
rect 401318 -19020 401440 -18964
rect 400640 -19088 401440 -19020
rect 400640 -19144 400766 -19088
rect 400822 -19144 400890 -19088
rect 400946 -19144 401014 -19088
rect 401070 -19144 401138 -19088
rect 401194 -19144 401262 -19088
rect 401318 -19144 401440 -19088
rect 400640 -19212 401440 -19144
rect 400640 -19268 400766 -19212
rect 400822 -19268 400890 -19212
rect 400946 -19268 401014 -19212
rect 401070 -19268 401138 -19212
rect 401194 -19268 401262 -19212
rect 401318 -19268 401440 -19212
rect 400640 -19336 401440 -19268
rect 400640 -19392 400766 -19336
rect 400822 -19392 400890 -19336
rect 400946 -19392 401014 -19336
rect 401070 -19392 401138 -19336
rect 401194 -19392 401262 -19336
rect 401318 -19392 401440 -19336
rect 400640 -19460 401440 -19392
rect 400640 -19516 400766 -19460
rect 400822 -19516 400890 -19460
rect 400946 -19516 401014 -19460
rect 401070 -19516 401138 -19460
rect 401194 -19516 401262 -19460
rect 401318 -19516 401440 -19460
rect 400640 -19584 401440 -19516
rect 400640 -19640 400766 -19584
rect 400822 -19640 400890 -19584
rect 400946 -19640 401014 -19584
rect 401070 -19640 401138 -19584
rect 401194 -19640 401262 -19584
rect 401318 -19640 401440 -19584
rect 400640 -19708 401440 -19640
rect 400640 -19764 400766 -19708
rect 400822 -19764 400890 -19708
rect 400946 -19764 401014 -19708
rect 401070 -19764 401138 -19708
rect 401194 -19764 401262 -19708
rect 401318 -19764 401440 -19708
rect 400640 -19832 401440 -19764
rect 400640 -19888 400766 -19832
rect 400822 -19888 400890 -19832
rect 400946 -19888 401014 -19832
rect 401070 -19888 401138 -19832
rect 401194 -19888 401262 -19832
rect 401318 -19888 401440 -19832
rect 400640 -19956 401440 -19888
rect 400640 -20012 400766 -19956
rect 400822 -20012 400890 -19956
rect 400946 -20012 401014 -19956
rect 401070 -20012 401138 -19956
rect 401194 -20012 401262 -19956
rect 401318 -20012 401440 -19956
rect 400640 -20080 401440 -20012
rect 400640 -20136 400766 -20080
rect 400822 -20136 400890 -20080
rect 400946 -20136 401014 -20080
rect 401070 -20136 401138 -20080
rect 401194 -20136 401262 -20080
rect 401318 -20136 401440 -20080
rect 400640 -20204 401440 -20136
rect 400640 -20260 400766 -20204
rect 400822 -20260 400890 -20204
rect 400946 -20260 401014 -20204
rect 401070 -20260 401138 -20204
rect 401194 -20260 401262 -20204
rect 401318 -20260 401440 -20204
rect 400640 -20328 401440 -20260
rect 400640 -20384 400766 -20328
rect 400822 -20384 400890 -20328
rect 400946 -20384 401014 -20328
rect 401070 -20384 401138 -20328
rect 401194 -20384 401262 -20328
rect 401318 -20384 401440 -20328
rect 400640 -20452 401440 -20384
rect 400640 -20508 400766 -20452
rect 400822 -20508 400890 -20452
rect 400946 -20508 401014 -20452
rect 401070 -20508 401138 -20452
rect 401194 -20508 401262 -20452
rect 401318 -20508 401440 -20452
rect 400640 -20576 401440 -20508
rect 400640 -20632 400766 -20576
rect 400822 -20632 400890 -20576
rect 400946 -20632 401014 -20576
rect 401070 -20632 401138 -20576
rect 401194 -20632 401262 -20576
rect 401318 -20632 401440 -20576
rect 400640 -20700 401440 -20632
rect 400640 -20756 400766 -20700
rect 400822 -20756 400890 -20700
rect 400946 -20756 401014 -20700
rect 401070 -20756 401138 -20700
rect 401194 -20756 401262 -20700
rect 401318 -20756 401440 -20700
rect 400640 -20824 401440 -20756
rect 400640 -20880 400766 -20824
rect 400822 -20880 400890 -20824
rect 400946 -20880 401014 -20824
rect 401070 -20880 401138 -20824
rect 401194 -20880 401262 -20824
rect 401318 -20880 401440 -20824
rect 400640 -20948 401440 -20880
rect 400640 -21004 400766 -20948
rect 400822 -21004 400890 -20948
rect 400946 -21004 401014 -20948
rect 401070 -21004 401138 -20948
rect 401194 -21004 401262 -20948
rect 401318 -21004 401440 -20948
rect 400640 -21072 401440 -21004
rect 400640 -21128 400766 -21072
rect 400822 -21128 400890 -21072
rect 400946 -21128 401014 -21072
rect 401070 -21128 401138 -21072
rect 401194 -21128 401262 -21072
rect 401318 -21128 401440 -21072
rect 400640 -21196 401440 -21128
rect 400640 -21252 400766 -21196
rect 400822 -21252 400890 -21196
rect 400946 -21252 401014 -21196
rect 401070 -21252 401138 -21196
rect 401194 -21252 401262 -21196
rect 401318 -21252 401440 -21196
rect 400640 -21320 401440 -21252
rect 400640 -21376 400766 -21320
rect 400822 -21376 400890 -21320
rect 400946 -21376 401014 -21320
rect 401070 -21376 401138 -21320
rect 401194 -21376 401262 -21320
rect 401318 -21376 401440 -21320
rect 400640 -21444 401440 -21376
rect 400640 -21500 400766 -21444
rect 400822 -21500 400890 -21444
rect 400946 -21500 401014 -21444
rect 401070 -21500 401138 -21444
rect 401194 -21500 401262 -21444
rect 401318 -21500 401440 -21444
rect 400640 -21568 401440 -21500
rect 400640 -21624 400766 -21568
rect 400822 -21624 400890 -21568
rect 400946 -21624 401014 -21568
rect 401070 -21624 401138 -21568
rect 401194 -21624 401262 -21568
rect 401318 -21624 401440 -21568
rect 400640 -21692 401440 -21624
rect 400640 -21748 400766 -21692
rect 400822 -21748 400890 -21692
rect 400946 -21748 401014 -21692
rect 401070 -21748 401138 -21692
rect 401194 -21748 401262 -21692
rect 401318 -21748 401440 -21692
rect 400640 -21816 401440 -21748
rect 400640 -21872 400766 -21816
rect 400822 -21872 400890 -21816
rect 400946 -21872 401014 -21816
rect 401070 -21872 401138 -21816
rect 401194 -21872 401262 -21816
rect 401318 -21872 401440 -21816
rect 400640 -21940 401440 -21872
rect 400640 -21996 400766 -21940
rect 400822 -21996 400890 -21940
rect 400946 -21996 401014 -21940
rect 401070 -21996 401138 -21940
rect 401194 -21996 401262 -21940
rect 401318 -21996 401440 -21940
rect 400640 -22064 401440 -21996
rect 400640 -22120 400766 -22064
rect 400822 -22120 400890 -22064
rect 400946 -22120 401014 -22064
rect 401070 -22120 401138 -22064
rect 401194 -22120 401262 -22064
rect 401318 -22120 401440 -22064
rect 400640 -22188 401440 -22120
rect 400640 -22244 400766 -22188
rect 400822 -22244 400890 -22188
rect 400946 -22244 401014 -22188
rect 401070 -22244 401138 -22188
rect 401194 -22244 401262 -22188
rect 401318 -22244 401440 -22188
rect 400640 -22312 401440 -22244
rect 400640 -22368 400766 -22312
rect 400822 -22368 400890 -22312
rect 400946 -22368 401014 -22312
rect 401070 -22368 401138 -22312
rect 401194 -22368 401262 -22312
rect 401318 -22368 401440 -22312
rect 400640 -22436 401440 -22368
rect 400640 -22492 400766 -22436
rect 400822 -22492 400890 -22436
rect 400946 -22492 401014 -22436
rect 401070 -22492 401138 -22436
rect 401194 -22492 401262 -22436
rect 401318 -22492 401440 -22436
rect 400640 -22560 401440 -22492
rect 400640 -22616 400766 -22560
rect 400822 -22616 400890 -22560
rect 400946 -22616 401014 -22560
rect 401070 -22616 401138 -22560
rect 401194 -22616 401262 -22560
rect 401318 -22616 401440 -22560
rect 400640 -22684 401440 -22616
rect 400640 -22740 400766 -22684
rect 400822 -22740 400890 -22684
rect 400946 -22740 401014 -22684
rect 401070 -22740 401138 -22684
rect 401194 -22740 401262 -22684
rect 401318 -22740 401440 -22684
rect 400640 -22808 401440 -22740
rect 400640 -22864 400766 -22808
rect 400822 -22864 400890 -22808
rect 400946 -22864 401014 -22808
rect 401070 -22864 401138 -22808
rect 401194 -22864 401262 -22808
rect 401318 -22864 401440 -22808
rect 400640 -22932 401440 -22864
rect 400640 -22988 400766 -22932
rect 400822 -22988 400890 -22932
rect 400946 -22988 401014 -22932
rect 401070 -22988 401138 -22932
rect 401194 -22988 401262 -22932
rect 401318 -22988 401440 -22932
rect 400640 -23056 401440 -22988
rect 400640 -23112 400766 -23056
rect 400822 -23112 400890 -23056
rect 400946 -23112 401014 -23056
rect 401070 -23112 401138 -23056
rect 401194 -23112 401262 -23056
rect 401318 -23112 401440 -23056
rect 400640 -23180 401440 -23112
rect 400640 -23236 400766 -23180
rect 400822 -23236 400890 -23180
rect 400946 -23236 401014 -23180
rect 401070 -23236 401138 -23180
rect 401194 -23236 401262 -23180
rect 401318 -23236 401440 -23180
rect 400640 -23304 401440 -23236
rect 400640 -23360 400766 -23304
rect 400822 -23360 400890 -23304
rect 400946 -23360 401014 -23304
rect 401070 -23360 401138 -23304
rect 401194 -23360 401262 -23304
rect 401318 -23360 401440 -23304
rect 400640 -23428 401440 -23360
rect 400640 -23484 400766 -23428
rect 400822 -23484 400890 -23428
rect 400946 -23484 401014 -23428
rect 401070 -23484 401138 -23428
rect 401194 -23484 401262 -23428
rect 401318 -23484 401440 -23428
rect 400640 -23552 401440 -23484
rect 400640 -23608 400766 -23552
rect 400822 -23608 400890 -23552
rect 400946 -23608 401014 -23552
rect 401070 -23608 401138 -23552
rect 401194 -23608 401262 -23552
rect 401318 -23608 401440 -23552
rect 400640 -23676 401440 -23608
rect 400640 -23732 400766 -23676
rect 400822 -23732 400890 -23676
rect 400946 -23732 401014 -23676
rect 401070 -23732 401138 -23676
rect 401194 -23732 401262 -23676
rect 401318 -23732 401440 -23676
rect 400640 -23800 401440 -23732
rect 400640 -23856 400766 -23800
rect 400822 -23856 400890 -23800
rect 400946 -23856 401014 -23800
rect 401070 -23856 401138 -23800
rect 401194 -23856 401262 -23800
rect 401318 -23856 401440 -23800
rect 400640 -23924 401440 -23856
rect 400640 -23980 400766 -23924
rect 400822 -23980 400890 -23924
rect 400946 -23980 401014 -23924
rect 401070 -23980 401138 -23924
rect 401194 -23980 401262 -23924
rect 401318 -23980 401440 -23924
rect 400640 -24048 401440 -23980
rect 400640 -24104 400766 -24048
rect 400822 -24104 400890 -24048
rect 400946 -24104 401014 -24048
rect 401070 -24104 401138 -24048
rect 401194 -24104 401262 -24048
rect 401318 -24104 401440 -24048
rect 400640 -24172 401440 -24104
rect 400640 -24228 400766 -24172
rect 400822 -24228 400890 -24172
rect 400946 -24228 401014 -24172
rect 401070 -24228 401138 -24172
rect 401194 -24228 401262 -24172
rect 401318 -24228 401440 -24172
rect 400640 -24296 401440 -24228
rect 400640 -24352 400766 -24296
rect 400822 -24352 400890 -24296
rect 400946 -24352 401014 -24296
rect 401070 -24352 401138 -24296
rect 401194 -24352 401262 -24296
rect 401318 -24352 401440 -24296
rect 400640 -24420 401440 -24352
rect 400640 -24476 400766 -24420
rect 400822 -24476 400890 -24420
rect 400946 -24476 401014 -24420
rect 401070 -24476 401138 -24420
rect 401194 -24476 401262 -24420
rect 401318 -24476 401440 -24420
rect 400640 -24544 401440 -24476
rect 400640 -24600 400766 -24544
rect 400822 -24600 400890 -24544
rect 400946 -24600 401014 -24544
rect 401070 -24600 401138 -24544
rect 401194 -24600 401262 -24544
rect 401318 -24600 401440 -24544
rect 400640 -24668 401440 -24600
rect 400640 -24724 400766 -24668
rect 400822 -24724 400890 -24668
rect 400946 -24724 401014 -24668
rect 401070 -24724 401138 -24668
rect 401194 -24724 401262 -24668
rect 401318 -24724 401440 -24668
rect 400640 -24792 401440 -24724
rect 400640 -24848 400766 -24792
rect 400822 -24848 400890 -24792
rect 400946 -24848 401014 -24792
rect 401070 -24848 401138 -24792
rect 401194 -24848 401262 -24792
rect 401318 -24848 401440 -24792
rect 400640 -24916 401440 -24848
rect 400640 -24972 400766 -24916
rect 400822 -24972 400890 -24916
rect 400946 -24972 401014 -24916
rect 401070 -24972 401138 -24916
rect 401194 -24972 401262 -24916
rect 401318 -24972 401440 -24916
rect 400640 -25040 401440 -24972
rect 400640 -25096 400766 -25040
rect 400822 -25096 400890 -25040
rect 400946 -25096 401014 -25040
rect 401070 -25096 401138 -25040
rect 401194 -25096 401262 -25040
rect 401318 -25096 401440 -25040
rect 400640 -25164 401440 -25096
rect 400640 -25220 400766 -25164
rect 400822 -25220 400890 -25164
rect 400946 -25220 401014 -25164
rect 401070 -25220 401138 -25164
rect 401194 -25220 401262 -25164
rect 401318 -25220 401440 -25164
rect 400640 -25288 401440 -25220
rect 400640 -25344 400766 -25288
rect 400822 -25344 400890 -25288
rect 400946 -25344 401014 -25288
rect 401070 -25344 401138 -25288
rect 401194 -25344 401262 -25288
rect 401318 -25344 401440 -25288
rect 400640 -25412 401440 -25344
rect 400640 -25468 400766 -25412
rect 400822 -25468 400890 -25412
rect 400946 -25468 401014 -25412
rect 401070 -25468 401138 -25412
rect 401194 -25468 401262 -25412
rect 401318 -25468 401440 -25412
rect 400640 -25532 401440 -25468
rect 387840 -25536 401440 -25532
rect 387840 -25592 387954 -25536
rect 388010 -25592 388078 -25536
rect 388134 -25592 388202 -25536
rect 388258 -25592 388326 -25536
rect 388382 -25592 388450 -25536
rect 388506 -25592 400766 -25536
rect 400822 -25592 400890 -25536
rect 400946 -25592 401014 -25536
rect 401070 -25592 401138 -25536
rect 401194 -25592 401262 -25536
rect 401318 -25592 401440 -25536
rect 387840 -25660 401440 -25592
rect 387840 -25716 387954 -25660
rect 388010 -25716 388078 -25660
rect 388134 -25716 388202 -25660
rect 388258 -25716 388326 -25660
rect 388382 -25716 388450 -25660
rect 388506 -25688 400766 -25660
rect 388506 -25716 388655 -25688
rect 387840 -25744 388655 -25716
rect 388711 -25744 388797 -25688
rect 388853 -25744 388939 -25688
rect 388995 -25744 389081 -25688
rect 389137 -25744 389223 -25688
rect 389279 -25744 389365 -25688
rect 389421 -25744 389507 -25688
rect 389563 -25744 389649 -25688
rect 389705 -25744 389791 -25688
rect 389847 -25744 389933 -25688
rect 389989 -25744 390075 -25688
rect 390131 -25744 390217 -25688
rect 390273 -25744 390359 -25688
rect 390415 -25744 390501 -25688
rect 390557 -25744 390643 -25688
rect 390699 -25744 390785 -25688
rect 390841 -25744 390927 -25688
rect 390983 -25744 391069 -25688
rect 391125 -25744 391211 -25688
rect 391267 -25744 391353 -25688
rect 391409 -25744 391495 -25688
rect 391551 -25744 391637 -25688
rect 391693 -25744 391779 -25688
rect 391835 -25744 391921 -25688
rect 391977 -25744 392063 -25688
rect 392119 -25744 392205 -25688
rect 392261 -25744 392347 -25688
rect 392403 -25744 392489 -25688
rect 392545 -25744 392631 -25688
rect 392687 -25744 392773 -25688
rect 392829 -25744 392915 -25688
rect 392971 -25744 393057 -25688
rect 393113 -25744 393199 -25688
rect 393255 -25744 393341 -25688
rect 393397 -25744 393483 -25688
rect 393539 -25744 393625 -25688
rect 393681 -25744 393767 -25688
rect 393823 -25744 393909 -25688
rect 393965 -25744 394051 -25688
rect 394107 -25744 394193 -25688
rect 394249 -25744 394335 -25688
rect 394391 -25744 394477 -25688
rect 394533 -25744 394619 -25688
rect 394675 -25744 394761 -25688
rect 394817 -25744 394903 -25688
rect 394959 -25744 395045 -25688
rect 395101 -25744 395187 -25688
rect 395243 -25744 395329 -25688
rect 395385 -25744 395471 -25688
rect 395527 -25744 395613 -25688
rect 395669 -25744 395755 -25688
rect 395811 -25744 395897 -25688
rect 395953 -25744 396039 -25688
rect 396095 -25744 396181 -25688
rect 396237 -25744 396323 -25688
rect 396379 -25744 396465 -25688
rect 396521 -25744 396607 -25688
rect 396663 -25744 396749 -25688
rect 396805 -25744 396891 -25688
rect 396947 -25744 397033 -25688
rect 397089 -25744 397175 -25688
rect 397231 -25744 397317 -25688
rect 397373 -25744 397459 -25688
rect 397515 -25744 397601 -25688
rect 397657 -25744 397743 -25688
rect 397799 -25744 397885 -25688
rect 397941 -25744 398027 -25688
rect 398083 -25744 398169 -25688
rect 398225 -25744 398311 -25688
rect 398367 -25744 398453 -25688
rect 398509 -25744 398595 -25688
rect 398651 -25744 398737 -25688
rect 398793 -25744 398879 -25688
rect 398935 -25744 399021 -25688
rect 399077 -25744 399163 -25688
rect 399219 -25744 399305 -25688
rect 399361 -25744 399447 -25688
rect 399503 -25744 399589 -25688
rect 399645 -25744 399731 -25688
rect 399787 -25744 399873 -25688
rect 399929 -25744 400015 -25688
rect 400071 -25744 400157 -25688
rect 400213 -25744 400299 -25688
rect 400355 -25744 400441 -25688
rect 400497 -25744 400583 -25688
rect 400639 -25716 400766 -25688
rect 400822 -25716 400890 -25660
rect 400946 -25716 401014 -25660
rect 401070 -25716 401138 -25660
rect 401194 -25716 401262 -25660
rect 401318 -25716 401440 -25660
rect 400639 -25744 401440 -25716
rect 387840 -25784 401440 -25744
rect 387840 -25840 387954 -25784
rect 388010 -25840 388078 -25784
rect 388134 -25840 388202 -25784
rect 388258 -25840 388326 -25784
rect 388382 -25840 388450 -25784
rect 388506 -25830 400766 -25784
rect 388506 -25840 388655 -25830
rect 387840 -25886 388655 -25840
rect 388711 -25886 388797 -25830
rect 388853 -25886 388939 -25830
rect 388995 -25886 389081 -25830
rect 389137 -25886 389223 -25830
rect 389279 -25886 389365 -25830
rect 389421 -25886 389507 -25830
rect 389563 -25886 389649 -25830
rect 389705 -25886 389791 -25830
rect 389847 -25886 389933 -25830
rect 389989 -25886 390075 -25830
rect 390131 -25886 390217 -25830
rect 390273 -25886 390359 -25830
rect 390415 -25886 390501 -25830
rect 390557 -25886 390643 -25830
rect 390699 -25886 390785 -25830
rect 390841 -25886 390927 -25830
rect 390983 -25886 391069 -25830
rect 391125 -25886 391211 -25830
rect 391267 -25886 391353 -25830
rect 391409 -25886 391495 -25830
rect 391551 -25886 391637 -25830
rect 391693 -25886 391779 -25830
rect 391835 -25886 391921 -25830
rect 391977 -25886 392063 -25830
rect 392119 -25886 392205 -25830
rect 392261 -25886 392347 -25830
rect 392403 -25886 392489 -25830
rect 392545 -25886 392631 -25830
rect 392687 -25886 392773 -25830
rect 392829 -25886 392915 -25830
rect 392971 -25886 393057 -25830
rect 393113 -25886 393199 -25830
rect 393255 -25886 393341 -25830
rect 393397 -25886 393483 -25830
rect 393539 -25886 393625 -25830
rect 393681 -25886 393767 -25830
rect 393823 -25886 393909 -25830
rect 393965 -25886 394051 -25830
rect 394107 -25886 394193 -25830
rect 394249 -25886 394335 -25830
rect 394391 -25886 394477 -25830
rect 394533 -25886 394619 -25830
rect 394675 -25886 394761 -25830
rect 394817 -25886 394903 -25830
rect 394959 -25886 395045 -25830
rect 395101 -25886 395187 -25830
rect 395243 -25886 395329 -25830
rect 395385 -25886 395471 -25830
rect 395527 -25886 395613 -25830
rect 395669 -25886 395755 -25830
rect 395811 -25886 395897 -25830
rect 395953 -25886 396039 -25830
rect 396095 -25886 396181 -25830
rect 396237 -25886 396323 -25830
rect 396379 -25886 396465 -25830
rect 396521 -25886 396607 -25830
rect 396663 -25886 396749 -25830
rect 396805 -25886 396891 -25830
rect 396947 -25886 397033 -25830
rect 397089 -25886 397175 -25830
rect 397231 -25886 397317 -25830
rect 397373 -25886 397459 -25830
rect 397515 -25886 397601 -25830
rect 397657 -25886 397743 -25830
rect 397799 -25886 397885 -25830
rect 397941 -25886 398027 -25830
rect 398083 -25886 398169 -25830
rect 398225 -25886 398311 -25830
rect 398367 -25886 398453 -25830
rect 398509 -25886 398595 -25830
rect 398651 -25886 398737 -25830
rect 398793 -25886 398879 -25830
rect 398935 -25886 399021 -25830
rect 399077 -25886 399163 -25830
rect 399219 -25886 399305 -25830
rect 399361 -25886 399447 -25830
rect 399503 -25886 399589 -25830
rect 399645 -25886 399731 -25830
rect 399787 -25886 399873 -25830
rect 399929 -25886 400015 -25830
rect 400071 -25886 400157 -25830
rect 400213 -25886 400299 -25830
rect 400355 -25886 400441 -25830
rect 400497 -25886 400583 -25830
rect 400639 -25840 400766 -25830
rect 400822 -25840 400890 -25784
rect 400946 -25840 401014 -25784
rect 401070 -25840 401138 -25784
rect 401194 -25840 401262 -25784
rect 401318 -25840 401440 -25784
rect 400639 -25886 401440 -25840
rect 387840 -25990 401440 -25886
<< via4 >>
rect 387986 -13097 388042 -13041
rect 388110 -13097 388166 -13041
rect 388234 -13097 388290 -13041
rect 388358 -13097 388414 -13041
rect 388482 -13097 388538 -13041
rect 388606 -13097 388662 -13041
rect 388730 -13097 388786 -13041
rect 388854 -13097 388910 -13041
rect 388978 -13097 389034 -13041
rect 389102 -13097 389158 -13041
rect 389226 -13097 389282 -13041
rect 389350 -13097 389406 -13041
rect 389474 -13097 389530 -13041
rect 389598 -13097 389654 -13041
rect 389722 -13097 389778 -13041
rect 389846 -13097 389902 -13041
rect 389970 -13097 390026 -13041
rect 390094 -13097 390150 -13041
rect 390218 -13097 390274 -13041
rect 390342 -13097 390398 -13041
rect 390466 -13097 390522 -13041
rect 390590 -13097 390646 -13041
rect 390714 -13097 390770 -13041
rect 390838 -13097 390894 -13041
rect 390962 -13097 391018 -13041
rect 391086 -13097 391142 -13041
rect 391210 -13097 391266 -13041
rect 391334 -13097 391390 -13041
rect 391458 -13097 391514 -13041
rect 391582 -13097 391638 -13041
rect 391706 -13097 391762 -13041
rect 391830 -13097 391886 -13041
rect 391954 -13097 392010 -13041
rect 392078 -13097 392134 -13041
rect 392202 -13097 392258 -13041
rect 392326 -13097 392382 -13041
rect 392450 -13097 392506 -13041
rect 392574 -13097 392630 -13041
rect 392698 -13097 392754 -13041
rect 392822 -13097 392878 -13041
rect 392946 -13097 393002 -13041
rect 393070 -13097 393126 -13041
rect 393194 -13097 393250 -13041
rect 393318 -13097 393374 -13041
rect 393442 -13097 393498 -13041
rect 393566 -13097 393622 -13041
rect 393690 -13097 393746 -13041
rect 393814 -13097 393870 -13041
rect 393938 -13097 393994 -13041
rect 394062 -13097 394118 -13041
rect 394186 -13097 394242 -13041
rect 394310 -13097 394366 -13041
rect 394434 -13097 394490 -13041
rect 394558 -13097 394614 -13041
rect 394682 -13097 394738 -13041
rect 394806 -13097 394862 -13041
rect 394930 -13097 394986 -13041
rect 395054 -13097 395110 -13041
rect 395178 -13097 395234 -13041
rect 395302 -13097 395358 -13041
rect 395426 -13097 395482 -13041
rect 395550 -13097 395606 -13041
rect 395674 -13097 395730 -13041
rect 395798 -13097 395854 -13041
rect 395922 -13097 395978 -13041
rect 396046 -13097 396102 -13041
rect 396170 -13097 396226 -13041
rect 396294 -13097 396350 -13041
rect 396418 -13097 396474 -13041
rect 396542 -13097 396598 -13041
rect 396666 -13097 396722 -13041
rect 396790 -13097 396846 -13041
rect 396914 -13097 396970 -13041
rect 397038 -13097 397094 -13041
rect 397162 -13097 397218 -13041
rect 397286 -13097 397342 -13041
rect 397410 -13097 397466 -13041
rect 397534 -13097 397590 -13041
rect 397658 -13097 397714 -13041
rect 397782 -13097 397838 -13041
rect 397906 -13097 397962 -13041
rect 398030 -13097 398086 -13041
rect 398154 -13097 398210 -13041
rect 398278 -13097 398334 -13041
rect 398402 -13097 398458 -13041
rect 398526 -13097 398582 -13041
rect 398650 -13097 398706 -13041
rect 398774 -13097 398830 -13041
rect 398898 -13097 398954 -13041
rect 399022 -13097 399078 -13041
rect 399146 -13097 399202 -13041
rect 399270 -13097 399326 -13041
rect 399394 -13097 399450 -13041
rect 399518 -13097 399574 -13041
rect 399642 -13097 399698 -13041
rect 399766 -13097 399822 -13041
rect 399890 -13097 399946 -13041
rect 400014 -13097 400070 -13041
rect 400138 -13097 400194 -13041
rect 400262 -13097 400318 -13041
rect 400386 -13097 400442 -13041
rect 400510 -13097 400566 -13041
rect 400634 -13097 400690 -13041
rect 400758 -13097 400814 -13041
rect 400882 -13097 400938 -13041
rect 401006 -13097 401062 -13041
rect 401130 -13097 401186 -13041
rect 401254 -13097 401310 -13041
rect 387986 -13221 388042 -13165
rect 388110 -13221 388166 -13165
rect 388234 -13221 388290 -13165
rect 388358 -13221 388414 -13165
rect 388482 -13221 388538 -13165
rect 388606 -13221 388662 -13165
rect 388730 -13221 388786 -13165
rect 388854 -13221 388910 -13165
rect 388978 -13221 389034 -13165
rect 389102 -13221 389158 -13165
rect 389226 -13221 389282 -13165
rect 389350 -13221 389406 -13165
rect 389474 -13221 389530 -13165
rect 389598 -13221 389654 -13165
rect 389722 -13221 389778 -13165
rect 389846 -13221 389902 -13165
rect 389970 -13221 390026 -13165
rect 390094 -13221 390150 -13165
rect 390218 -13221 390274 -13165
rect 390342 -13221 390398 -13165
rect 390466 -13221 390522 -13165
rect 390590 -13221 390646 -13165
rect 390714 -13221 390770 -13165
rect 390838 -13221 390894 -13165
rect 390962 -13221 391018 -13165
rect 391086 -13221 391142 -13165
rect 391210 -13221 391266 -13165
rect 391334 -13221 391390 -13165
rect 391458 -13221 391514 -13165
rect 391582 -13221 391638 -13165
rect 391706 -13221 391762 -13165
rect 391830 -13221 391886 -13165
rect 391954 -13221 392010 -13165
rect 392078 -13221 392134 -13165
rect 392202 -13221 392258 -13165
rect 392326 -13221 392382 -13165
rect 392450 -13221 392506 -13165
rect 392574 -13221 392630 -13165
rect 392698 -13221 392754 -13165
rect 392822 -13221 392878 -13165
rect 392946 -13221 393002 -13165
rect 393070 -13221 393126 -13165
rect 393194 -13221 393250 -13165
rect 393318 -13221 393374 -13165
rect 393442 -13221 393498 -13165
rect 393566 -13221 393622 -13165
rect 393690 -13221 393746 -13165
rect 393814 -13221 393870 -13165
rect 393938 -13221 393994 -13165
rect 394062 -13221 394118 -13165
rect 394186 -13221 394242 -13165
rect 394310 -13221 394366 -13165
rect 394434 -13221 394490 -13165
rect 394558 -13221 394614 -13165
rect 394682 -13221 394738 -13165
rect 394806 -13221 394862 -13165
rect 394930 -13221 394986 -13165
rect 395054 -13221 395110 -13165
rect 395178 -13221 395234 -13165
rect 395302 -13221 395358 -13165
rect 395426 -13221 395482 -13165
rect 395550 -13221 395606 -13165
rect 395674 -13221 395730 -13165
rect 395798 -13221 395854 -13165
rect 395922 -13221 395978 -13165
rect 396046 -13221 396102 -13165
rect 396170 -13221 396226 -13165
rect 396294 -13221 396350 -13165
rect 396418 -13221 396474 -13165
rect 396542 -13221 396598 -13165
rect 396666 -13221 396722 -13165
rect 396790 -13221 396846 -13165
rect 396914 -13221 396970 -13165
rect 397038 -13221 397094 -13165
rect 397162 -13221 397218 -13165
rect 397286 -13221 397342 -13165
rect 397410 -13221 397466 -13165
rect 397534 -13221 397590 -13165
rect 397658 -13221 397714 -13165
rect 397782 -13221 397838 -13165
rect 397906 -13221 397962 -13165
rect 398030 -13221 398086 -13165
rect 398154 -13221 398210 -13165
rect 398278 -13221 398334 -13165
rect 398402 -13221 398458 -13165
rect 398526 -13221 398582 -13165
rect 398650 -13221 398706 -13165
rect 398774 -13221 398830 -13165
rect 398898 -13221 398954 -13165
rect 399022 -13221 399078 -13165
rect 399146 -13221 399202 -13165
rect 399270 -13221 399326 -13165
rect 399394 -13221 399450 -13165
rect 399518 -13221 399574 -13165
rect 399642 -13221 399698 -13165
rect 399766 -13221 399822 -13165
rect 399890 -13221 399946 -13165
rect 400014 -13221 400070 -13165
rect 400138 -13221 400194 -13165
rect 400262 -13221 400318 -13165
rect 400386 -13221 400442 -13165
rect 400510 -13221 400566 -13165
rect 400634 -13221 400690 -13165
rect 400758 -13221 400814 -13165
rect 400882 -13221 400938 -13165
rect 401006 -13221 401062 -13165
rect 401130 -13221 401186 -13165
rect 401254 -13221 401310 -13165
rect 387986 -13345 388042 -13289
rect 388110 -13345 388166 -13289
rect 388234 -13345 388290 -13289
rect 388358 -13345 388414 -13289
rect 388482 -13345 388538 -13289
rect 388606 -13345 388662 -13289
rect 388730 -13345 388786 -13289
rect 388854 -13345 388910 -13289
rect 388978 -13345 389034 -13289
rect 389102 -13345 389158 -13289
rect 389226 -13345 389282 -13289
rect 389350 -13345 389406 -13289
rect 389474 -13345 389530 -13289
rect 389598 -13345 389654 -13289
rect 389722 -13345 389778 -13289
rect 389846 -13345 389902 -13289
rect 389970 -13345 390026 -13289
rect 390094 -13345 390150 -13289
rect 390218 -13345 390274 -13289
rect 390342 -13345 390398 -13289
rect 390466 -13345 390522 -13289
rect 390590 -13345 390646 -13289
rect 390714 -13345 390770 -13289
rect 390838 -13345 390894 -13289
rect 390962 -13345 391018 -13289
rect 391086 -13345 391142 -13289
rect 391210 -13345 391266 -13289
rect 391334 -13345 391390 -13289
rect 391458 -13345 391514 -13289
rect 391582 -13345 391638 -13289
rect 391706 -13345 391762 -13289
rect 391830 -13345 391886 -13289
rect 391954 -13345 392010 -13289
rect 392078 -13345 392134 -13289
rect 392202 -13345 392258 -13289
rect 392326 -13345 392382 -13289
rect 392450 -13345 392506 -13289
rect 392574 -13345 392630 -13289
rect 392698 -13345 392754 -13289
rect 392822 -13345 392878 -13289
rect 392946 -13345 393002 -13289
rect 393070 -13345 393126 -13289
rect 393194 -13345 393250 -13289
rect 393318 -13345 393374 -13289
rect 393442 -13345 393498 -13289
rect 393566 -13345 393622 -13289
rect 393690 -13345 393746 -13289
rect 393814 -13345 393870 -13289
rect 393938 -13345 393994 -13289
rect 394062 -13345 394118 -13289
rect 394186 -13345 394242 -13289
rect 394310 -13345 394366 -13289
rect 394434 -13345 394490 -13289
rect 394558 -13345 394614 -13289
rect 394682 -13345 394738 -13289
rect 394806 -13345 394862 -13289
rect 394930 -13345 394986 -13289
rect 395054 -13345 395110 -13289
rect 395178 -13345 395234 -13289
rect 395302 -13345 395358 -13289
rect 395426 -13345 395482 -13289
rect 395550 -13345 395606 -13289
rect 395674 -13345 395730 -13289
rect 395798 -13345 395854 -13289
rect 395922 -13345 395978 -13289
rect 396046 -13345 396102 -13289
rect 396170 -13345 396226 -13289
rect 396294 -13345 396350 -13289
rect 396418 -13345 396474 -13289
rect 396542 -13345 396598 -13289
rect 396666 -13345 396722 -13289
rect 396790 -13345 396846 -13289
rect 396914 -13345 396970 -13289
rect 397038 -13345 397094 -13289
rect 397162 -13345 397218 -13289
rect 397286 -13345 397342 -13289
rect 397410 -13345 397466 -13289
rect 397534 -13345 397590 -13289
rect 397658 -13345 397714 -13289
rect 397782 -13345 397838 -13289
rect 397906 -13345 397962 -13289
rect 398030 -13345 398086 -13289
rect 398154 -13345 398210 -13289
rect 398278 -13345 398334 -13289
rect 398402 -13345 398458 -13289
rect 398526 -13345 398582 -13289
rect 398650 -13345 398706 -13289
rect 398774 -13345 398830 -13289
rect 398898 -13345 398954 -13289
rect 399022 -13345 399078 -13289
rect 399146 -13345 399202 -13289
rect 399270 -13345 399326 -13289
rect 399394 -13345 399450 -13289
rect 399518 -13345 399574 -13289
rect 399642 -13345 399698 -13289
rect 399766 -13345 399822 -13289
rect 399890 -13345 399946 -13289
rect 400014 -13345 400070 -13289
rect 400138 -13345 400194 -13289
rect 400262 -13345 400318 -13289
rect 400386 -13345 400442 -13289
rect 400510 -13345 400566 -13289
rect 400634 -13345 400690 -13289
rect 400758 -13345 400814 -13289
rect 400882 -13345 400938 -13289
rect 401006 -13345 401062 -13289
rect 401130 -13345 401186 -13289
rect 401254 -13345 401310 -13289
rect 387986 -13469 388042 -13413
rect 388110 -13469 388166 -13413
rect 388234 -13469 388290 -13413
rect 388358 -13469 388414 -13413
rect 388482 -13469 388538 -13413
rect 388606 -13469 388662 -13413
rect 388730 -13469 388786 -13413
rect 388854 -13469 388910 -13413
rect 388978 -13469 389034 -13413
rect 389102 -13469 389158 -13413
rect 389226 -13469 389282 -13413
rect 389350 -13469 389406 -13413
rect 389474 -13469 389530 -13413
rect 389598 -13469 389654 -13413
rect 389722 -13469 389778 -13413
rect 389846 -13469 389902 -13413
rect 389970 -13469 390026 -13413
rect 390094 -13469 390150 -13413
rect 390218 -13469 390274 -13413
rect 390342 -13469 390398 -13413
rect 390466 -13469 390522 -13413
rect 390590 -13469 390646 -13413
rect 390714 -13469 390770 -13413
rect 390838 -13469 390894 -13413
rect 390962 -13469 391018 -13413
rect 391086 -13469 391142 -13413
rect 391210 -13469 391266 -13413
rect 391334 -13469 391390 -13413
rect 391458 -13469 391514 -13413
rect 391582 -13469 391638 -13413
rect 391706 -13469 391762 -13413
rect 391830 -13469 391886 -13413
rect 391954 -13469 392010 -13413
rect 392078 -13469 392134 -13413
rect 392202 -13469 392258 -13413
rect 392326 -13469 392382 -13413
rect 392450 -13469 392506 -13413
rect 392574 -13469 392630 -13413
rect 392698 -13469 392754 -13413
rect 392822 -13469 392878 -13413
rect 392946 -13469 393002 -13413
rect 393070 -13469 393126 -13413
rect 393194 -13469 393250 -13413
rect 393318 -13469 393374 -13413
rect 393442 -13469 393498 -13413
rect 393566 -13469 393622 -13413
rect 393690 -13469 393746 -13413
rect 393814 -13469 393870 -13413
rect 393938 -13469 393994 -13413
rect 394062 -13469 394118 -13413
rect 394186 -13469 394242 -13413
rect 394310 -13469 394366 -13413
rect 394434 -13469 394490 -13413
rect 394558 -13469 394614 -13413
rect 394682 -13469 394738 -13413
rect 394806 -13469 394862 -13413
rect 394930 -13469 394986 -13413
rect 395054 -13469 395110 -13413
rect 395178 -13469 395234 -13413
rect 395302 -13469 395358 -13413
rect 395426 -13469 395482 -13413
rect 395550 -13469 395606 -13413
rect 395674 -13469 395730 -13413
rect 395798 -13469 395854 -13413
rect 395922 -13469 395978 -13413
rect 396046 -13469 396102 -13413
rect 396170 -13469 396226 -13413
rect 396294 -13469 396350 -13413
rect 396418 -13469 396474 -13413
rect 396542 -13469 396598 -13413
rect 396666 -13469 396722 -13413
rect 396790 -13469 396846 -13413
rect 396914 -13469 396970 -13413
rect 397038 -13469 397094 -13413
rect 397162 -13469 397218 -13413
rect 397286 -13469 397342 -13413
rect 397410 -13469 397466 -13413
rect 397534 -13469 397590 -13413
rect 397658 -13469 397714 -13413
rect 397782 -13469 397838 -13413
rect 397906 -13469 397962 -13413
rect 398030 -13469 398086 -13413
rect 398154 -13469 398210 -13413
rect 398278 -13469 398334 -13413
rect 398402 -13469 398458 -13413
rect 398526 -13469 398582 -13413
rect 398650 -13469 398706 -13413
rect 398774 -13469 398830 -13413
rect 398898 -13469 398954 -13413
rect 399022 -13469 399078 -13413
rect 399146 -13469 399202 -13413
rect 399270 -13469 399326 -13413
rect 399394 -13469 399450 -13413
rect 399518 -13469 399574 -13413
rect 399642 -13469 399698 -13413
rect 399766 -13469 399822 -13413
rect 399890 -13469 399946 -13413
rect 400014 -13469 400070 -13413
rect 400138 -13469 400194 -13413
rect 400262 -13469 400318 -13413
rect 400386 -13469 400442 -13413
rect 400510 -13469 400566 -13413
rect 400634 -13469 400690 -13413
rect 400758 -13469 400814 -13413
rect 400882 -13469 400938 -13413
rect 401006 -13469 401062 -13413
rect 401130 -13469 401186 -13413
rect 401254 -13469 401310 -13413
rect 387954 -13688 388010 -13632
rect 388078 -13688 388134 -13632
rect 388202 -13688 388258 -13632
rect 388326 -13688 388382 -13632
rect 388450 -13688 388506 -13632
rect 387954 -13812 388010 -13756
rect 388078 -13812 388134 -13756
rect 388202 -13812 388258 -13756
rect 388326 -13812 388382 -13756
rect 388450 -13812 388506 -13756
rect 387954 -13936 388010 -13880
rect 388078 -13936 388134 -13880
rect 388202 -13936 388258 -13880
rect 388326 -13936 388382 -13880
rect 388450 -13936 388506 -13880
rect 387954 -14060 388010 -14004
rect 388078 -14060 388134 -14004
rect 388202 -14060 388258 -14004
rect 388326 -14060 388382 -14004
rect 388450 -14060 388506 -14004
rect 387954 -14184 388010 -14128
rect 388078 -14184 388134 -14128
rect 388202 -14184 388258 -14128
rect 388326 -14184 388382 -14128
rect 388450 -14184 388506 -14128
rect 387954 -14308 388010 -14252
rect 388078 -14308 388134 -14252
rect 388202 -14308 388258 -14252
rect 388326 -14308 388382 -14252
rect 388450 -14308 388506 -14252
rect 387954 -14432 388010 -14376
rect 388078 -14432 388134 -14376
rect 388202 -14432 388258 -14376
rect 388326 -14432 388382 -14376
rect 388450 -14432 388506 -14376
rect 387954 -14556 388010 -14500
rect 388078 -14556 388134 -14500
rect 388202 -14556 388258 -14500
rect 388326 -14556 388382 -14500
rect 388450 -14556 388506 -14500
rect 387954 -14680 388010 -14624
rect 388078 -14680 388134 -14624
rect 388202 -14680 388258 -14624
rect 388326 -14680 388382 -14624
rect 388450 -14680 388506 -14624
rect 387954 -14804 388010 -14748
rect 388078 -14804 388134 -14748
rect 388202 -14804 388258 -14748
rect 388326 -14804 388382 -14748
rect 388450 -14804 388506 -14748
rect 387954 -14928 388010 -14872
rect 388078 -14928 388134 -14872
rect 388202 -14928 388258 -14872
rect 388326 -14928 388382 -14872
rect 388450 -14928 388506 -14872
rect 387954 -15052 388010 -14996
rect 388078 -15052 388134 -14996
rect 388202 -15052 388258 -14996
rect 388326 -15052 388382 -14996
rect 388450 -15052 388506 -14996
rect 387954 -15176 388010 -15120
rect 388078 -15176 388134 -15120
rect 388202 -15176 388258 -15120
rect 388326 -15176 388382 -15120
rect 388450 -15176 388506 -15120
rect 387954 -15300 388010 -15244
rect 388078 -15300 388134 -15244
rect 388202 -15300 388258 -15244
rect 388326 -15300 388382 -15244
rect 388450 -15300 388506 -15244
rect 387954 -15424 388010 -15368
rect 388078 -15424 388134 -15368
rect 388202 -15424 388258 -15368
rect 388326 -15424 388382 -15368
rect 388450 -15424 388506 -15368
rect 387954 -15548 388010 -15492
rect 388078 -15548 388134 -15492
rect 388202 -15548 388258 -15492
rect 388326 -15548 388382 -15492
rect 388450 -15548 388506 -15492
rect 387954 -15672 388010 -15616
rect 388078 -15672 388134 -15616
rect 388202 -15672 388258 -15616
rect 388326 -15672 388382 -15616
rect 388450 -15672 388506 -15616
rect 387954 -15796 388010 -15740
rect 388078 -15796 388134 -15740
rect 388202 -15796 388258 -15740
rect 388326 -15796 388382 -15740
rect 388450 -15796 388506 -15740
rect 387954 -15920 388010 -15864
rect 388078 -15920 388134 -15864
rect 388202 -15920 388258 -15864
rect 388326 -15920 388382 -15864
rect 388450 -15920 388506 -15864
rect 387954 -16044 388010 -15988
rect 388078 -16044 388134 -15988
rect 388202 -16044 388258 -15988
rect 388326 -16044 388382 -15988
rect 388450 -16044 388506 -15988
rect 387954 -16168 388010 -16112
rect 388078 -16168 388134 -16112
rect 388202 -16168 388258 -16112
rect 388326 -16168 388382 -16112
rect 388450 -16168 388506 -16112
rect 387954 -16292 388010 -16236
rect 388078 -16292 388134 -16236
rect 388202 -16292 388258 -16236
rect 388326 -16292 388382 -16236
rect 388450 -16292 388506 -16236
rect 387954 -16416 388010 -16360
rect 388078 -16416 388134 -16360
rect 388202 -16416 388258 -16360
rect 388326 -16416 388382 -16360
rect 388450 -16416 388506 -16360
rect 387954 -16540 388010 -16484
rect 388078 -16540 388134 -16484
rect 388202 -16540 388258 -16484
rect 388326 -16540 388382 -16484
rect 388450 -16540 388506 -16484
rect 387954 -16664 388010 -16608
rect 388078 -16664 388134 -16608
rect 388202 -16664 388258 -16608
rect 388326 -16664 388382 -16608
rect 388450 -16664 388506 -16608
rect 387954 -16788 388010 -16732
rect 388078 -16788 388134 -16732
rect 388202 -16788 388258 -16732
rect 388326 -16788 388382 -16732
rect 388450 -16788 388506 -16732
rect 387954 -16912 388010 -16856
rect 388078 -16912 388134 -16856
rect 388202 -16912 388258 -16856
rect 388326 -16912 388382 -16856
rect 388450 -16912 388506 -16856
rect 387954 -17036 388010 -16980
rect 388078 -17036 388134 -16980
rect 388202 -17036 388258 -16980
rect 388326 -17036 388382 -16980
rect 388450 -17036 388506 -16980
rect 387954 -17160 388010 -17104
rect 388078 -17160 388134 -17104
rect 388202 -17160 388258 -17104
rect 388326 -17160 388382 -17104
rect 388450 -17160 388506 -17104
rect 387954 -17284 388010 -17228
rect 388078 -17284 388134 -17228
rect 388202 -17284 388258 -17228
rect 388326 -17284 388382 -17228
rect 388450 -17284 388506 -17228
rect 387954 -17408 388010 -17352
rect 388078 -17408 388134 -17352
rect 388202 -17408 388258 -17352
rect 388326 -17408 388382 -17352
rect 388450 -17408 388506 -17352
rect 387954 -17532 388010 -17476
rect 388078 -17532 388134 -17476
rect 388202 -17532 388258 -17476
rect 388326 -17532 388382 -17476
rect 388450 -17532 388506 -17476
rect 387954 -17656 388010 -17600
rect 388078 -17656 388134 -17600
rect 388202 -17656 388258 -17600
rect 388326 -17656 388382 -17600
rect 388450 -17656 388506 -17600
rect 387954 -17780 388010 -17724
rect 388078 -17780 388134 -17724
rect 388202 -17780 388258 -17724
rect 388326 -17780 388382 -17724
rect 388450 -17780 388506 -17724
rect 387954 -17904 388010 -17848
rect 388078 -17904 388134 -17848
rect 388202 -17904 388258 -17848
rect 388326 -17904 388382 -17848
rect 388450 -17904 388506 -17848
rect 387954 -18028 388010 -17972
rect 388078 -18028 388134 -17972
rect 388202 -18028 388258 -17972
rect 388326 -18028 388382 -17972
rect 388450 -18028 388506 -17972
rect 387954 -18152 388010 -18096
rect 388078 -18152 388134 -18096
rect 388202 -18152 388258 -18096
rect 388326 -18152 388382 -18096
rect 388450 -18152 388506 -18096
rect 387954 -18276 388010 -18220
rect 388078 -18276 388134 -18220
rect 388202 -18276 388258 -18220
rect 388326 -18276 388382 -18220
rect 388450 -18276 388506 -18220
rect 387954 -18400 388010 -18344
rect 388078 -18400 388134 -18344
rect 388202 -18400 388258 -18344
rect 388326 -18400 388382 -18344
rect 388450 -18400 388506 -18344
rect 387954 -18524 388010 -18468
rect 388078 -18524 388134 -18468
rect 388202 -18524 388258 -18468
rect 388326 -18524 388382 -18468
rect 388450 -18524 388506 -18468
rect 387954 -18648 388010 -18592
rect 388078 -18648 388134 -18592
rect 388202 -18648 388258 -18592
rect 388326 -18648 388382 -18592
rect 388450 -18648 388506 -18592
rect 387954 -18772 388010 -18716
rect 388078 -18772 388134 -18716
rect 388202 -18772 388258 -18716
rect 388326 -18772 388382 -18716
rect 388450 -18772 388506 -18716
rect 387954 -18896 388010 -18840
rect 388078 -18896 388134 -18840
rect 388202 -18896 388258 -18840
rect 388326 -18896 388382 -18840
rect 388450 -18896 388506 -18840
rect 387954 -19020 388010 -18964
rect 388078 -19020 388134 -18964
rect 388202 -19020 388258 -18964
rect 388326 -19020 388382 -18964
rect 388450 -19020 388506 -18964
rect 387954 -19144 388010 -19088
rect 388078 -19144 388134 -19088
rect 388202 -19144 388258 -19088
rect 388326 -19144 388382 -19088
rect 388450 -19144 388506 -19088
rect 387954 -19268 388010 -19212
rect 388078 -19268 388134 -19212
rect 388202 -19268 388258 -19212
rect 388326 -19268 388382 -19212
rect 388450 -19268 388506 -19212
rect 387954 -19392 388010 -19336
rect 388078 -19392 388134 -19336
rect 388202 -19392 388258 -19336
rect 388326 -19392 388382 -19336
rect 388450 -19392 388506 -19336
rect 387954 -19516 388010 -19460
rect 388078 -19516 388134 -19460
rect 388202 -19516 388258 -19460
rect 388326 -19516 388382 -19460
rect 388450 -19516 388506 -19460
rect 387954 -19640 388010 -19584
rect 388078 -19640 388134 -19584
rect 388202 -19640 388258 -19584
rect 388326 -19640 388382 -19584
rect 388450 -19640 388506 -19584
rect 387954 -19764 388010 -19708
rect 388078 -19764 388134 -19708
rect 388202 -19764 388258 -19708
rect 388326 -19764 388382 -19708
rect 388450 -19764 388506 -19708
rect 387954 -19888 388010 -19832
rect 388078 -19888 388134 -19832
rect 388202 -19888 388258 -19832
rect 388326 -19888 388382 -19832
rect 388450 -19888 388506 -19832
rect 387954 -20012 388010 -19956
rect 388078 -20012 388134 -19956
rect 388202 -20012 388258 -19956
rect 388326 -20012 388382 -19956
rect 388450 -20012 388506 -19956
rect 387954 -20136 388010 -20080
rect 388078 -20136 388134 -20080
rect 388202 -20136 388258 -20080
rect 388326 -20136 388382 -20080
rect 388450 -20136 388506 -20080
rect 387954 -20260 388010 -20204
rect 388078 -20260 388134 -20204
rect 388202 -20260 388258 -20204
rect 388326 -20260 388382 -20204
rect 388450 -20260 388506 -20204
rect 387954 -20384 388010 -20328
rect 388078 -20384 388134 -20328
rect 388202 -20384 388258 -20328
rect 388326 -20384 388382 -20328
rect 388450 -20384 388506 -20328
rect 387954 -20508 388010 -20452
rect 388078 -20508 388134 -20452
rect 388202 -20508 388258 -20452
rect 388326 -20508 388382 -20452
rect 388450 -20508 388506 -20452
rect 387954 -20632 388010 -20576
rect 388078 -20632 388134 -20576
rect 388202 -20632 388258 -20576
rect 388326 -20632 388382 -20576
rect 388450 -20632 388506 -20576
rect 387954 -20756 388010 -20700
rect 388078 -20756 388134 -20700
rect 388202 -20756 388258 -20700
rect 388326 -20756 388382 -20700
rect 388450 -20756 388506 -20700
rect 387954 -20880 388010 -20824
rect 388078 -20880 388134 -20824
rect 388202 -20880 388258 -20824
rect 388326 -20880 388382 -20824
rect 388450 -20880 388506 -20824
rect 387954 -21004 388010 -20948
rect 388078 -21004 388134 -20948
rect 388202 -21004 388258 -20948
rect 388326 -21004 388382 -20948
rect 388450 -21004 388506 -20948
rect 387954 -21128 388010 -21072
rect 388078 -21128 388134 -21072
rect 388202 -21128 388258 -21072
rect 388326 -21128 388382 -21072
rect 388450 -21128 388506 -21072
rect 387954 -21252 388010 -21196
rect 388078 -21252 388134 -21196
rect 388202 -21252 388258 -21196
rect 388326 -21252 388382 -21196
rect 388450 -21252 388506 -21196
rect 387954 -21376 388010 -21320
rect 388078 -21376 388134 -21320
rect 388202 -21376 388258 -21320
rect 388326 -21376 388382 -21320
rect 388450 -21376 388506 -21320
rect 387954 -21500 388010 -21444
rect 388078 -21500 388134 -21444
rect 388202 -21500 388258 -21444
rect 388326 -21500 388382 -21444
rect 388450 -21500 388506 -21444
rect 387954 -21624 388010 -21568
rect 388078 -21624 388134 -21568
rect 388202 -21624 388258 -21568
rect 388326 -21624 388382 -21568
rect 388450 -21624 388506 -21568
rect 387954 -21748 388010 -21692
rect 388078 -21748 388134 -21692
rect 388202 -21748 388258 -21692
rect 388326 -21748 388382 -21692
rect 388450 -21748 388506 -21692
rect 387954 -21872 388010 -21816
rect 388078 -21872 388134 -21816
rect 388202 -21872 388258 -21816
rect 388326 -21872 388382 -21816
rect 388450 -21872 388506 -21816
rect 387954 -21996 388010 -21940
rect 388078 -21996 388134 -21940
rect 388202 -21996 388258 -21940
rect 388326 -21996 388382 -21940
rect 388450 -21996 388506 -21940
rect 387954 -22120 388010 -22064
rect 388078 -22120 388134 -22064
rect 388202 -22120 388258 -22064
rect 388326 -22120 388382 -22064
rect 388450 -22120 388506 -22064
rect 387954 -22244 388010 -22188
rect 388078 -22244 388134 -22188
rect 388202 -22244 388258 -22188
rect 388326 -22244 388382 -22188
rect 388450 -22244 388506 -22188
rect 387954 -22368 388010 -22312
rect 388078 -22368 388134 -22312
rect 388202 -22368 388258 -22312
rect 388326 -22368 388382 -22312
rect 388450 -22368 388506 -22312
rect 387954 -22492 388010 -22436
rect 388078 -22492 388134 -22436
rect 388202 -22492 388258 -22436
rect 388326 -22492 388382 -22436
rect 388450 -22492 388506 -22436
rect 387954 -22616 388010 -22560
rect 388078 -22616 388134 -22560
rect 388202 -22616 388258 -22560
rect 388326 -22616 388382 -22560
rect 388450 -22616 388506 -22560
rect 387954 -22740 388010 -22684
rect 388078 -22740 388134 -22684
rect 388202 -22740 388258 -22684
rect 388326 -22740 388382 -22684
rect 388450 -22740 388506 -22684
rect 387954 -22864 388010 -22808
rect 388078 -22864 388134 -22808
rect 388202 -22864 388258 -22808
rect 388326 -22864 388382 -22808
rect 388450 -22864 388506 -22808
rect 387954 -22988 388010 -22932
rect 388078 -22988 388134 -22932
rect 388202 -22988 388258 -22932
rect 388326 -22988 388382 -22932
rect 388450 -22988 388506 -22932
rect 387954 -23112 388010 -23056
rect 388078 -23112 388134 -23056
rect 388202 -23112 388258 -23056
rect 388326 -23112 388382 -23056
rect 388450 -23112 388506 -23056
rect 387954 -23236 388010 -23180
rect 388078 -23236 388134 -23180
rect 388202 -23236 388258 -23180
rect 388326 -23236 388382 -23180
rect 388450 -23236 388506 -23180
rect 387954 -23360 388010 -23304
rect 388078 -23360 388134 -23304
rect 388202 -23360 388258 -23304
rect 388326 -23360 388382 -23304
rect 388450 -23360 388506 -23304
rect 387954 -23484 388010 -23428
rect 388078 -23484 388134 -23428
rect 388202 -23484 388258 -23428
rect 388326 -23484 388382 -23428
rect 388450 -23484 388506 -23428
rect 387954 -23608 388010 -23552
rect 388078 -23608 388134 -23552
rect 388202 -23608 388258 -23552
rect 388326 -23608 388382 -23552
rect 388450 -23608 388506 -23552
rect 387954 -23732 388010 -23676
rect 388078 -23732 388134 -23676
rect 388202 -23732 388258 -23676
rect 388326 -23732 388382 -23676
rect 388450 -23732 388506 -23676
rect 387954 -23856 388010 -23800
rect 388078 -23856 388134 -23800
rect 388202 -23856 388258 -23800
rect 388326 -23856 388382 -23800
rect 388450 -23856 388506 -23800
rect 387954 -23980 388010 -23924
rect 388078 -23980 388134 -23924
rect 388202 -23980 388258 -23924
rect 388326 -23980 388382 -23924
rect 388450 -23980 388506 -23924
rect 387954 -24104 388010 -24048
rect 388078 -24104 388134 -24048
rect 388202 -24104 388258 -24048
rect 388326 -24104 388382 -24048
rect 388450 -24104 388506 -24048
rect 387954 -24228 388010 -24172
rect 388078 -24228 388134 -24172
rect 388202 -24228 388258 -24172
rect 388326 -24228 388382 -24172
rect 388450 -24228 388506 -24172
rect 387954 -24352 388010 -24296
rect 388078 -24352 388134 -24296
rect 388202 -24352 388258 -24296
rect 388326 -24352 388382 -24296
rect 388450 -24352 388506 -24296
rect 387954 -24476 388010 -24420
rect 388078 -24476 388134 -24420
rect 388202 -24476 388258 -24420
rect 388326 -24476 388382 -24420
rect 388450 -24476 388506 -24420
rect 387954 -24600 388010 -24544
rect 388078 -24600 388134 -24544
rect 388202 -24600 388258 -24544
rect 388326 -24600 388382 -24544
rect 388450 -24600 388506 -24544
rect 387954 -24724 388010 -24668
rect 388078 -24724 388134 -24668
rect 388202 -24724 388258 -24668
rect 388326 -24724 388382 -24668
rect 388450 -24724 388506 -24668
rect 387954 -24848 388010 -24792
rect 388078 -24848 388134 -24792
rect 388202 -24848 388258 -24792
rect 388326 -24848 388382 -24792
rect 388450 -24848 388506 -24792
rect 387954 -24972 388010 -24916
rect 388078 -24972 388134 -24916
rect 388202 -24972 388258 -24916
rect 388326 -24972 388382 -24916
rect 388450 -24972 388506 -24916
rect 387954 -25096 388010 -25040
rect 388078 -25096 388134 -25040
rect 388202 -25096 388258 -25040
rect 388326 -25096 388382 -25040
rect 388450 -25096 388506 -25040
rect 387954 -25220 388010 -25164
rect 388078 -25220 388134 -25164
rect 388202 -25220 388258 -25164
rect 388326 -25220 388382 -25164
rect 388450 -25220 388506 -25164
rect 387954 -25344 388010 -25288
rect 388078 -25344 388134 -25288
rect 388202 -25344 388258 -25288
rect 388326 -25344 388382 -25288
rect 388450 -25344 388506 -25288
rect 387954 -25468 388010 -25412
rect 388078 -25468 388134 -25412
rect 388202 -25468 388258 -25412
rect 388326 -25468 388382 -25412
rect 388450 -25468 388506 -25412
rect 388981 -13736 389037 -13680
rect 389123 -13736 389179 -13680
rect 388981 -13878 389037 -13822
rect 389123 -13878 389179 -13822
rect 388981 -14020 389037 -13964
rect 389123 -14020 389179 -13964
rect 388981 -14162 389037 -14106
rect 389123 -14162 389179 -14106
rect 388981 -14304 389037 -14248
rect 389123 -14304 389179 -14248
rect 388981 -14446 389037 -14390
rect 389123 -14446 389179 -14390
rect 388981 -14588 389037 -14532
rect 389123 -14588 389179 -14532
rect 388981 -14730 389037 -14674
rect 389123 -14730 389179 -14674
rect 388981 -14872 389037 -14816
rect 389123 -14872 389179 -14816
rect 388981 -15014 389037 -14958
rect 389123 -15014 389179 -14958
rect 388981 -15156 389037 -15100
rect 389123 -15156 389179 -15100
rect 388981 -15298 389037 -15242
rect 389123 -15298 389179 -15242
rect 388981 -15440 389037 -15384
rect 389123 -15440 389179 -15384
rect 388981 -15582 389037 -15526
rect 389123 -15582 389179 -15526
rect 388981 -15724 389037 -15668
rect 389123 -15724 389179 -15668
rect 388981 -15866 389037 -15810
rect 389123 -15866 389179 -15810
rect 388981 -16008 389037 -15952
rect 389123 -16008 389179 -15952
rect 388981 -16150 389037 -16094
rect 389123 -16150 389179 -16094
rect 388981 -16292 389037 -16236
rect 389123 -16292 389179 -16236
rect 388981 -16434 389037 -16378
rect 389123 -16434 389179 -16378
rect 388981 -16576 389037 -16520
rect 389123 -16576 389179 -16520
rect 388981 -16718 389037 -16662
rect 389123 -16718 389179 -16662
rect 388981 -16860 389037 -16804
rect 389123 -16860 389179 -16804
rect 388981 -17002 389037 -16946
rect 389123 -17002 389179 -16946
rect 388981 -17144 389037 -17088
rect 389123 -17144 389179 -17088
rect 388981 -17286 389037 -17230
rect 389123 -17286 389179 -17230
rect 388981 -17428 389037 -17372
rect 389123 -17428 389179 -17372
rect 388981 -17570 389037 -17514
rect 389123 -17570 389179 -17514
rect 388981 -17712 389037 -17656
rect 389123 -17712 389179 -17656
rect 388981 -17854 389037 -17798
rect 389123 -17854 389179 -17798
rect 388981 -17996 389037 -17940
rect 389123 -17996 389179 -17940
rect 388981 -18138 389037 -18082
rect 389123 -18138 389179 -18082
rect 388981 -18280 389037 -18224
rect 389123 -18280 389179 -18224
rect 388981 -18422 389037 -18366
rect 389123 -18422 389179 -18366
rect 388981 -18564 389037 -18508
rect 389123 -18564 389179 -18508
rect 388981 -18706 389037 -18650
rect 389123 -18706 389179 -18650
rect 388981 -18848 389037 -18792
rect 389123 -18848 389179 -18792
rect 388981 -18990 389037 -18934
rect 389123 -18990 389179 -18934
rect 388981 -19132 389037 -19076
rect 389123 -19132 389179 -19076
rect 388981 -19274 389037 -19218
rect 389123 -19274 389179 -19218
rect 388981 -19416 389037 -19360
rect 389123 -19416 389179 -19360
rect 388981 -19558 389037 -19502
rect 389123 -19558 389179 -19502
rect 388981 -19700 389037 -19644
rect 389123 -19700 389179 -19644
rect 388981 -19842 389037 -19786
rect 389123 -19842 389179 -19786
rect 388981 -19984 389037 -19928
rect 389123 -19984 389179 -19928
rect 388981 -20126 389037 -20070
rect 389123 -20126 389179 -20070
rect 388981 -20268 389037 -20212
rect 389123 -20268 389179 -20212
rect 388981 -20410 389037 -20354
rect 389123 -20410 389179 -20354
rect 388981 -20552 389037 -20496
rect 389123 -20552 389179 -20496
rect 388981 -20694 389037 -20638
rect 389123 -20694 389179 -20638
rect 388981 -20836 389037 -20780
rect 389123 -20836 389179 -20780
rect 388981 -20978 389037 -20922
rect 389123 -20978 389179 -20922
rect 388981 -21120 389037 -21064
rect 389123 -21120 389179 -21064
rect 388981 -21262 389037 -21206
rect 389123 -21262 389179 -21206
rect 388981 -21404 389037 -21348
rect 389123 -21404 389179 -21348
rect 388981 -21546 389037 -21490
rect 389123 -21546 389179 -21490
rect 388981 -21688 389037 -21632
rect 389123 -21688 389179 -21632
rect 388981 -21830 389037 -21774
rect 389123 -21830 389179 -21774
rect 388981 -21972 389037 -21916
rect 389123 -21972 389179 -21916
rect 388981 -22114 389037 -22058
rect 389123 -22114 389179 -22058
rect 388981 -22256 389037 -22200
rect 389123 -22256 389179 -22200
rect 388981 -22398 389037 -22342
rect 389123 -22398 389179 -22342
rect 388981 -22540 389037 -22484
rect 389123 -22540 389179 -22484
rect 388981 -22682 389037 -22626
rect 389123 -22682 389179 -22626
rect 388981 -22824 389037 -22768
rect 389123 -22824 389179 -22768
rect 388981 -22966 389037 -22910
rect 389123 -22966 389179 -22910
rect 388981 -23108 389037 -23052
rect 389123 -23108 389179 -23052
rect 388981 -23250 389037 -23194
rect 389123 -23250 389179 -23194
rect 388981 -23392 389037 -23336
rect 389123 -23392 389179 -23336
rect 388981 -23534 389037 -23478
rect 389123 -23534 389179 -23478
rect 388981 -23676 389037 -23620
rect 389123 -23676 389179 -23620
rect 388981 -23818 389037 -23762
rect 389123 -23818 389179 -23762
rect 388981 -23960 389037 -23904
rect 389123 -23960 389179 -23904
rect 388981 -24102 389037 -24046
rect 389123 -24102 389179 -24046
rect 388981 -24244 389037 -24188
rect 389123 -24244 389179 -24188
rect 388981 -24386 389037 -24330
rect 389123 -24386 389179 -24330
rect 388981 -24528 389037 -24472
rect 389123 -24528 389179 -24472
rect 388981 -24670 389037 -24614
rect 389123 -24670 389179 -24614
rect 388981 -24812 389037 -24756
rect 389123 -24812 389179 -24756
rect 388981 -24954 389037 -24898
rect 389123 -24954 389179 -24898
rect 388981 -25096 389037 -25040
rect 389123 -25096 389179 -25040
rect 388981 -25238 389037 -25182
rect 389123 -25238 389179 -25182
rect 388981 -25380 389037 -25324
rect 389123 -25380 389179 -25324
rect 388981 -25522 389037 -25466
rect 389123 -25522 389179 -25466
rect 389382 -13736 389438 -13680
rect 389524 -13736 389580 -13680
rect 389382 -13878 389438 -13822
rect 389524 -13878 389580 -13822
rect 389382 -14020 389438 -13964
rect 389524 -14020 389580 -13964
rect 389382 -14162 389438 -14106
rect 389524 -14162 389580 -14106
rect 389382 -14304 389438 -14248
rect 389524 -14304 389580 -14248
rect 389382 -14446 389438 -14390
rect 389524 -14446 389580 -14390
rect 389382 -14588 389438 -14532
rect 389524 -14588 389580 -14532
rect 389382 -14730 389438 -14674
rect 389524 -14730 389580 -14674
rect 389382 -14872 389438 -14816
rect 389524 -14872 389580 -14816
rect 389382 -15014 389438 -14958
rect 389524 -15014 389580 -14958
rect 389382 -15156 389438 -15100
rect 389524 -15156 389580 -15100
rect 389382 -15298 389438 -15242
rect 389524 -15298 389580 -15242
rect 389382 -15440 389438 -15384
rect 389524 -15440 389580 -15384
rect 389382 -15582 389438 -15526
rect 389524 -15582 389580 -15526
rect 389382 -15724 389438 -15668
rect 389524 -15724 389580 -15668
rect 389382 -15866 389438 -15810
rect 389524 -15866 389580 -15810
rect 389382 -16008 389438 -15952
rect 389524 -16008 389580 -15952
rect 389382 -16150 389438 -16094
rect 389524 -16150 389580 -16094
rect 389382 -16292 389438 -16236
rect 389524 -16292 389580 -16236
rect 389382 -16434 389438 -16378
rect 389524 -16434 389580 -16378
rect 389382 -16576 389438 -16520
rect 389524 -16576 389580 -16520
rect 389382 -16718 389438 -16662
rect 389524 -16718 389580 -16662
rect 389382 -16860 389438 -16804
rect 389524 -16860 389580 -16804
rect 389382 -17002 389438 -16946
rect 389524 -17002 389580 -16946
rect 389382 -17144 389438 -17088
rect 389524 -17144 389580 -17088
rect 389382 -17286 389438 -17230
rect 389524 -17286 389580 -17230
rect 389382 -17428 389438 -17372
rect 389524 -17428 389580 -17372
rect 389382 -17570 389438 -17514
rect 389524 -17570 389580 -17514
rect 389382 -17712 389438 -17656
rect 389524 -17712 389580 -17656
rect 389382 -17854 389438 -17798
rect 389524 -17854 389580 -17798
rect 389382 -17996 389438 -17940
rect 389524 -17996 389580 -17940
rect 389382 -18138 389438 -18082
rect 389524 -18138 389580 -18082
rect 389382 -18280 389438 -18224
rect 389524 -18280 389580 -18224
rect 389382 -18422 389438 -18366
rect 389524 -18422 389580 -18366
rect 389382 -18564 389438 -18508
rect 389524 -18564 389580 -18508
rect 389382 -18706 389438 -18650
rect 389524 -18706 389580 -18650
rect 389382 -18848 389438 -18792
rect 389524 -18848 389580 -18792
rect 389382 -18990 389438 -18934
rect 389524 -18990 389580 -18934
rect 389382 -19132 389438 -19076
rect 389524 -19132 389580 -19076
rect 389382 -19274 389438 -19218
rect 389524 -19274 389580 -19218
rect 389382 -19416 389438 -19360
rect 389524 -19416 389580 -19360
rect 389382 -19558 389438 -19502
rect 389524 -19558 389580 -19502
rect 389382 -19700 389438 -19644
rect 389524 -19700 389580 -19644
rect 389382 -19842 389438 -19786
rect 389524 -19842 389580 -19786
rect 389382 -19984 389438 -19928
rect 389524 -19984 389580 -19928
rect 389382 -20126 389438 -20070
rect 389524 -20126 389580 -20070
rect 389382 -20268 389438 -20212
rect 389524 -20268 389580 -20212
rect 389382 -20410 389438 -20354
rect 389524 -20410 389580 -20354
rect 389382 -20552 389438 -20496
rect 389524 -20552 389580 -20496
rect 389382 -20694 389438 -20638
rect 389524 -20694 389580 -20638
rect 389382 -20836 389438 -20780
rect 389524 -20836 389580 -20780
rect 389382 -20978 389438 -20922
rect 389524 -20978 389580 -20922
rect 389382 -21120 389438 -21064
rect 389524 -21120 389580 -21064
rect 389382 -21262 389438 -21206
rect 389524 -21262 389580 -21206
rect 389382 -21404 389438 -21348
rect 389524 -21404 389580 -21348
rect 389382 -21546 389438 -21490
rect 389524 -21546 389580 -21490
rect 389382 -21688 389438 -21632
rect 389524 -21688 389580 -21632
rect 389382 -21830 389438 -21774
rect 389524 -21830 389580 -21774
rect 389382 -21972 389438 -21916
rect 389524 -21972 389580 -21916
rect 389382 -22114 389438 -22058
rect 389524 -22114 389580 -22058
rect 389382 -22256 389438 -22200
rect 389524 -22256 389580 -22200
rect 389382 -22398 389438 -22342
rect 389524 -22398 389580 -22342
rect 389382 -22540 389438 -22484
rect 389524 -22540 389580 -22484
rect 389382 -22682 389438 -22626
rect 389524 -22682 389580 -22626
rect 389382 -22824 389438 -22768
rect 389524 -22824 389580 -22768
rect 389382 -22966 389438 -22910
rect 389524 -22966 389580 -22910
rect 389382 -23108 389438 -23052
rect 389524 -23108 389580 -23052
rect 389382 -23250 389438 -23194
rect 389524 -23250 389580 -23194
rect 389382 -23392 389438 -23336
rect 389524 -23392 389580 -23336
rect 389382 -23534 389438 -23478
rect 389524 -23534 389580 -23478
rect 389382 -23676 389438 -23620
rect 389524 -23676 389580 -23620
rect 389382 -23818 389438 -23762
rect 389524 -23818 389580 -23762
rect 389382 -23960 389438 -23904
rect 389524 -23960 389580 -23904
rect 389382 -24102 389438 -24046
rect 389524 -24102 389580 -24046
rect 389382 -24244 389438 -24188
rect 389524 -24244 389580 -24188
rect 389382 -24386 389438 -24330
rect 389524 -24386 389580 -24330
rect 389382 -24528 389438 -24472
rect 389524 -24528 389580 -24472
rect 389382 -24670 389438 -24614
rect 389524 -24670 389580 -24614
rect 389382 -24812 389438 -24756
rect 389524 -24812 389580 -24756
rect 389382 -24954 389438 -24898
rect 389524 -24954 389580 -24898
rect 389382 -25096 389438 -25040
rect 389524 -25096 389580 -25040
rect 389382 -25238 389438 -25182
rect 389524 -25238 389580 -25182
rect 389382 -25380 389438 -25324
rect 389524 -25380 389580 -25324
rect 389382 -25522 389438 -25466
rect 389524 -25522 389580 -25466
rect 389782 -13736 389838 -13680
rect 389924 -13736 389980 -13680
rect 389782 -13878 389838 -13822
rect 389924 -13878 389980 -13822
rect 389782 -14020 389838 -13964
rect 389924 -14020 389980 -13964
rect 389782 -14162 389838 -14106
rect 389924 -14162 389980 -14106
rect 389782 -14304 389838 -14248
rect 389924 -14304 389980 -14248
rect 389782 -14446 389838 -14390
rect 389924 -14446 389980 -14390
rect 389782 -14588 389838 -14532
rect 389924 -14588 389980 -14532
rect 389782 -14730 389838 -14674
rect 389924 -14730 389980 -14674
rect 389782 -14872 389838 -14816
rect 389924 -14872 389980 -14816
rect 389782 -15014 389838 -14958
rect 389924 -15014 389980 -14958
rect 389782 -15156 389838 -15100
rect 389924 -15156 389980 -15100
rect 389782 -15298 389838 -15242
rect 389924 -15298 389980 -15242
rect 389782 -15440 389838 -15384
rect 389924 -15440 389980 -15384
rect 389782 -15582 389838 -15526
rect 389924 -15582 389980 -15526
rect 389782 -15724 389838 -15668
rect 389924 -15724 389980 -15668
rect 389782 -15866 389838 -15810
rect 389924 -15866 389980 -15810
rect 389782 -16008 389838 -15952
rect 389924 -16008 389980 -15952
rect 389782 -16150 389838 -16094
rect 389924 -16150 389980 -16094
rect 389782 -16292 389838 -16236
rect 389924 -16292 389980 -16236
rect 389782 -16434 389838 -16378
rect 389924 -16434 389980 -16378
rect 389782 -16576 389838 -16520
rect 389924 -16576 389980 -16520
rect 389782 -16718 389838 -16662
rect 389924 -16718 389980 -16662
rect 389782 -16860 389838 -16804
rect 389924 -16860 389980 -16804
rect 389782 -17002 389838 -16946
rect 389924 -17002 389980 -16946
rect 389782 -17144 389838 -17088
rect 389924 -17144 389980 -17088
rect 389782 -17286 389838 -17230
rect 389924 -17286 389980 -17230
rect 389782 -17428 389838 -17372
rect 389924 -17428 389980 -17372
rect 389782 -17570 389838 -17514
rect 389924 -17570 389980 -17514
rect 389782 -17712 389838 -17656
rect 389924 -17712 389980 -17656
rect 389782 -17854 389838 -17798
rect 389924 -17854 389980 -17798
rect 389782 -17996 389838 -17940
rect 389924 -17996 389980 -17940
rect 389782 -18138 389838 -18082
rect 389924 -18138 389980 -18082
rect 389782 -18280 389838 -18224
rect 389924 -18280 389980 -18224
rect 389782 -18422 389838 -18366
rect 389924 -18422 389980 -18366
rect 389782 -18564 389838 -18508
rect 389924 -18564 389980 -18508
rect 389782 -18706 389838 -18650
rect 389924 -18706 389980 -18650
rect 389782 -18848 389838 -18792
rect 389924 -18848 389980 -18792
rect 389782 -18990 389838 -18934
rect 389924 -18990 389980 -18934
rect 389782 -19132 389838 -19076
rect 389924 -19132 389980 -19076
rect 389782 -19274 389838 -19218
rect 389924 -19274 389980 -19218
rect 389782 -19416 389838 -19360
rect 389924 -19416 389980 -19360
rect 389782 -19558 389838 -19502
rect 389924 -19558 389980 -19502
rect 389782 -19700 389838 -19644
rect 389924 -19700 389980 -19644
rect 389782 -19842 389838 -19786
rect 389924 -19842 389980 -19786
rect 389782 -19984 389838 -19928
rect 389924 -19984 389980 -19928
rect 389782 -20126 389838 -20070
rect 389924 -20126 389980 -20070
rect 389782 -20268 389838 -20212
rect 389924 -20268 389980 -20212
rect 389782 -20410 389838 -20354
rect 389924 -20410 389980 -20354
rect 389782 -20552 389838 -20496
rect 389924 -20552 389980 -20496
rect 389782 -20694 389838 -20638
rect 389924 -20694 389980 -20638
rect 389782 -20836 389838 -20780
rect 389924 -20836 389980 -20780
rect 389782 -20978 389838 -20922
rect 389924 -20978 389980 -20922
rect 389782 -21120 389838 -21064
rect 389924 -21120 389980 -21064
rect 389782 -21262 389838 -21206
rect 389924 -21262 389980 -21206
rect 389782 -21404 389838 -21348
rect 389924 -21404 389980 -21348
rect 389782 -21546 389838 -21490
rect 389924 -21546 389980 -21490
rect 389782 -21688 389838 -21632
rect 389924 -21688 389980 -21632
rect 389782 -21830 389838 -21774
rect 389924 -21830 389980 -21774
rect 389782 -21972 389838 -21916
rect 389924 -21972 389980 -21916
rect 389782 -22114 389838 -22058
rect 389924 -22114 389980 -22058
rect 389782 -22256 389838 -22200
rect 389924 -22256 389980 -22200
rect 389782 -22398 389838 -22342
rect 389924 -22398 389980 -22342
rect 389782 -22540 389838 -22484
rect 389924 -22540 389980 -22484
rect 389782 -22682 389838 -22626
rect 389924 -22682 389980 -22626
rect 389782 -22824 389838 -22768
rect 389924 -22824 389980 -22768
rect 389782 -22966 389838 -22910
rect 389924 -22966 389980 -22910
rect 389782 -23108 389838 -23052
rect 389924 -23108 389980 -23052
rect 389782 -23250 389838 -23194
rect 389924 -23250 389980 -23194
rect 389782 -23392 389838 -23336
rect 389924 -23392 389980 -23336
rect 389782 -23534 389838 -23478
rect 389924 -23534 389980 -23478
rect 389782 -23676 389838 -23620
rect 389924 -23676 389980 -23620
rect 389782 -23818 389838 -23762
rect 389924 -23818 389980 -23762
rect 389782 -23960 389838 -23904
rect 389924 -23960 389980 -23904
rect 389782 -24102 389838 -24046
rect 389924 -24102 389980 -24046
rect 389782 -24244 389838 -24188
rect 389924 -24244 389980 -24188
rect 389782 -24386 389838 -24330
rect 389924 -24386 389980 -24330
rect 389782 -24528 389838 -24472
rect 389924 -24528 389980 -24472
rect 389782 -24670 389838 -24614
rect 389924 -24670 389980 -24614
rect 389782 -24812 389838 -24756
rect 389924 -24812 389980 -24756
rect 389782 -24954 389838 -24898
rect 389924 -24954 389980 -24898
rect 389782 -25096 389838 -25040
rect 389924 -25096 389980 -25040
rect 389782 -25238 389838 -25182
rect 389924 -25238 389980 -25182
rect 389782 -25380 389838 -25324
rect 389924 -25380 389980 -25324
rect 389782 -25522 389838 -25466
rect 389924 -25522 389980 -25466
rect 390179 -13736 390235 -13680
rect 390321 -13736 390377 -13680
rect 390179 -13878 390235 -13822
rect 390321 -13878 390377 -13822
rect 390179 -14020 390235 -13964
rect 390321 -14020 390377 -13964
rect 390179 -14162 390235 -14106
rect 390321 -14162 390377 -14106
rect 390179 -14304 390235 -14248
rect 390321 -14304 390377 -14248
rect 390179 -14446 390235 -14390
rect 390321 -14446 390377 -14390
rect 390179 -14588 390235 -14532
rect 390321 -14588 390377 -14532
rect 390179 -14730 390235 -14674
rect 390321 -14730 390377 -14674
rect 390179 -14872 390235 -14816
rect 390321 -14872 390377 -14816
rect 390179 -15014 390235 -14958
rect 390321 -15014 390377 -14958
rect 390179 -15156 390235 -15100
rect 390321 -15156 390377 -15100
rect 390179 -15298 390235 -15242
rect 390321 -15298 390377 -15242
rect 390179 -15440 390235 -15384
rect 390321 -15440 390377 -15384
rect 390179 -15582 390235 -15526
rect 390321 -15582 390377 -15526
rect 390179 -15724 390235 -15668
rect 390321 -15724 390377 -15668
rect 390179 -15866 390235 -15810
rect 390321 -15866 390377 -15810
rect 390179 -16008 390235 -15952
rect 390321 -16008 390377 -15952
rect 390179 -16150 390235 -16094
rect 390321 -16150 390377 -16094
rect 390179 -16292 390235 -16236
rect 390321 -16292 390377 -16236
rect 390179 -16434 390235 -16378
rect 390321 -16434 390377 -16378
rect 390179 -16576 390235 -16520
rect 390321 -16576 390377 -16520
rect 390179 -16718 390235 -16662
rect 390321 -16718 390377 -16662
rect 390179 -16860 390235 -16804
rect 390321 -16860 390377 -16804
rect 390179 -17002 390235 -16946
rect 390321 -17002 390377 -16946
rect 390179 -17144 390235 -17088
rect 390321 -17144 390377 -17088
rect 390179 -17286 390235 -17230
rect 390321 -17286 390377 -17230
rect 390179 -17428 390235 -17372
rect 390321 -17428 390377 -17372
rect 390179 -17570 390235 -17514
rect 390321 -17570 390377 -17514
rect 390179 -17712 390235 -17656
rect 390321 -17712 390377 -17656
rect 390179 -17854 390235 -17798
rect 390321 -17854 390377 -17798
rect 390179 -17996 390235 -17940
rect 390321 -17996 390377 -17940
rect 390179 -18138 390235 -18082
rect 390321 -18138 390377 -18082
rect 390179 -18280 390235 -18224
rect 390321 -18280 390377 -18224
rect 390179 -18422 390235 -18366
rect 390321 -18422 390377 -18366
rect 390179 -18564 390235 -18508
rect 390321 -18564 390377 -18508
rect 390179 -18706 390235 -18650
rect 390321 -18706 390377 -18650
rect 390179 -18848 390235 -18792
rect 390321 -18848 390377 -18792
rect 390179 -18990 390235 -18934
rect 390321 -18990 390377 -18934
rect 390179 -19132 390235 -19076
rect 390321 -19132 390377 -19076
rect 390179 -19274 390235 -19218
rect 390321 -19274 390377 -19218
rect 390179 -19416 390235 -19360
rect 390321 -19416 390377 -19360
rect 390179 -19558 390235 -19502
rect 390321 -19558 390377 -19502
rect 390179 -19700 390235 -19644
rect 390321 -19700 390377 -19644
rect 390179 -19842 390235 -19786
rect 390321 -19842 390377 -19786
rect 390179 -19984 390235 -19928
rect 390321 -19984 390377 -19928
rect 390179 -20126 390235 -20070
rect 390321 -20126 390377 -20070
rect 390179 -20268 390235 -20212
rect 390321 -20268 390377 -20212
rect 390179 -20410 390235 -20354
rect 390321 -20410 390377 -20354
rect 390179 -20552 390235 -20496
rect 390321 -20552 390377 -20496
rect 390179 -20694 390235 -20638
rect 390321 -20694 390377 -20638
rect 390179 -20836 390235 -20780
rect 390321 -20836 390377 -20780
rect 390179 -20978 390235 -20922
rect 390321 -20978 390377 -20922
rect 390179 -21120 390235 -21064
rect 390321 -21120 390377 -21064
rect 390179 -21262 390235 -21206
rect 390321 -21262 390377 -21206
rect 390179 -21404 390235 -21348
rect 390321 -21404 390377 -21348
rect 390179 -21546 390235 -21490
rect 390321 -21546 390377 -21490
rect 390179 -21688 390235 -21632
rect 390321 -21688 390377 -21632
rect 390179 -21830 390235 -21774
rect 390321 -21830 390377 -21774
rect 390179 -21972 390235 -21916
rect 390321 -21972 390377 -21916
rect 390179 -22114 390235 -22058
rect 390321 -22114 390377 -22058
rect 390179 -22256 390235 -22200
rect 390321 -22256 390377 -22200
rect 390179 -22398 390235 -22342
rect 390321 -22398 390377 -22342
rect 390179 -22540 390235 -22484
rect 390321 -22540 390377 -22484
rect 390179 -22682 390235 -22626
rect 390321 -22682 390377 -22626
rect 390179 -22824 390235 -22768
rect 390321 -22824 390377 -22768
rect 390179 -22966 390235 -22910
rect 390321 -22966 390377 -22910
rect 390179 -23108 390235 -23052
rect 390321 -23108 390377 -23052
rect 390179 -23250 390235 -23194
rect 390321 -23250 390377 -23194
rect 390179 -23392 390235 -23336
rect 390321 -23392 390377 -23336
rect 390179 -23534 390235 -23478
rect 390321 -23534 390377 -23478
rect 390179 -23676 390235 -23620
rect 390321 -23676 390377 -23620
rect 390179 -23818 390235 -23762
rect 390321 -23818 390377 -23762
rect 390179 -23960 390235 -23904
rect 390321 -23960 390377 -23904
rect 390179 -24102 390235 -24046
rect 390321 -24102 390377 -24046
rect 390179 -24244 390235 -24188
rect 390321 -24244 390377 -24188
rect 390179 -24386 390235 -24330
rect 390321 -24386 390377 -24330
rect 390179 -24528 390235 -24472
rect 390321 -24528 390377 -24472
rect 390179 -24670 390235 -24614
rect 390321 -24670 390377 -24614
rect 390179 -24812 390235 -24756
rect 390321 -24812 390377 -24756
rect 390179 -24954 390235 -24898
rect 390321 -24954 390377 -24898
rect 390179 -25096 390235 -25040
rect 390321 -25096 390377 -25040
rect 390179 -25238 390235 -25182
rect 390321 -25238 390377 -25182
rect 390179 -25380 390235 -25324
rect 390321 -25380 390377 -25324
rect 390179 -25522 390235 -25466
rect 390321 -25522 390377 -25466
rect 390576 -13736 390632 -13680
rect 390718 -13736 390774 -13680
rect 390576 -13878 390632 -13822
rect 390718 -13878 390774 -13822
rect 390576 -14020 390632 -13964
rect 390718 -14020 390774 -13964
rect 390576 -14162 390632 -14106
rect 390718 -14162 390774 -14106
rect 390576 -14304 390632 -14248
rect 390718 -14304 390774 -14248
rect 390576 -14446 390632 -14390
rect 390718 -14446 390774 -14390
rect 390576 -14588 390632 -14532
rect 390718 -14588 390774 -14532
rect 390576 -14730 390632 -14674
rect 390718 -14730 390774 -14674
rect 390576 -14872 390632 -14816
rect 390718 -14872 390774 -14816
rect 390576 -15014 390632 -14958
rect 390718 -15014 390774 -14958
rect 390576 -15156 390632 -15100
rect 390718 -15156 390774 -15100
rect 390576 -15298 390632 -15242
rect 390718 -15298 390774 -15242
rect 390576 -15440 390632 -15384
rect 390718 -15440 390774 -15384
rect 390576 -15582 390632 -15526
rect 390718 -15582 390774 -15526
rect 390576 -15724 390632 -15668
rect 390718 -15724 390774 -15668
rect 390576 -15866 390632 -15810
rect 390718 -15866 390774 -15810
rect 390576 -16008 390632 -15952
rect 390718 -16008 390774 -15952
rect 390576 -16150 390632 -16094
rect 390718 -16150 390774 -16094
rect 390576 -16292 390632 -16236
rect 390718 -16292 390774 -16236
rect 390576 -16434 390632 -16378
rect 390718 -16434 390774 -16378
rect 390576 -16576 390632 -16520
rect 390718 -16576 390774 -16520
rect 390576 -16718 390632 -16662
rect 390718 -16718 390774 -16662
rect 390576 -16860 390632 -16804
rect 390718 -16860 390774 -16804
rect 390576 -17002 390632 -16946
rect 390718 -17002 390774 -16946
rect 390576 -17144 390632 -17088
rect 390718 -17144 390774 -17088
rect 390576 -17286 390632 -17230
rect 390718 -17286 390774 -17230
rect 390576 -17428 390632 -17372
rect 390718 -17428 390774 -17372
rect 390576 -17570 390632 -17514
rect 390718 -17570 390774 -17514
rect 390576 -17712 390632 -17656
rect 390718 -17712 390774 -17656
rect 390576 -17854 390632 -17798
rect 390718 -17854 390774 -17798
rect 390576 -17996 390632 -17940
rect 390718 -17996 390774 -17940
rect 390576 -18138 390632 -18082
rect 390718 -18138 390774 -18082
rect 390576 -18280 390632 -18224
rect 390718 -18280 390774 -18224
rect 390576 -18422 390632 -18366
rect 390718 -18422 390774 -18366
rect 390576 -18564 390632 -18508
rect 390718 -18564 390774 -18508
rect 390576 -18706 390632 -18650
rect 390718 -18706 390774 -18650
rect 390576 -18848 390632 -18792
rect 390718 -18848 390774 -18792
rect 390576 -18990 390632 -18934
rect 390718 -18990 390774 -18934
rect 390576 -19132 390632 -19076
rect 390718 -19132 390774 -19076
rect 390576 -19274 390632 -19218
rect 390718 -19274 390774 -19218
rect 390576 -19416 390632 -19360
rect 390718 -19416 390774 -19360
rect 390576 -19558 390632 -19502
rect 390718 -19558 390774 -19502
rect 390576 -19700 390632 -19644
rect 390718 -19700 390774 -19644
rect 390576 -19842 390632 -19786
rect 390718 -19842 390774 -19786
rect 390576 -19984 390632 -19928
rect 390718 -19984 390774 -19928
rect 390576 -20126 390632 -20070
rect 390718 -20126 390774 -20070
rect 390576 -20268 390632 -20212
rect 390718 -20268 390774 -20212
rect 390576 -20410 390632 -20354
rect 390718 -20410 390774 -20354
rect 390576 -20552 390632 -20496
rect 390718 -20552 390774 -20496
rect 390576 -20694 390632 -20638
rect 390718 -20694 390774 -20638
rect 390576 -20836 390632 -20780
rect 390718 -20836 390774 -20780
rect 390576 -20978 390632 -20922
rect 390718 -20978 390774 -20922
rect 390576 -21120 390632 -21064
rect 390718 -21120 390774 -21064
rect 390576 -21262 390632 -21206
rect 390718 -21262 390774 -21206
rect 390576 -21404 390632 -21348
rect 390718 -21404 390774 -21348
rect 390576 -21546 390632 -21490
rect 390718 -21546 390774 -21490
rect 390576 -21688 390632 -21632
rect 390718 -21688 390774 -21632
rect 390576 -21830 390632 -21774
rect 390718 -21830 390774 -21774
rect 390576 -21972 390632 -21916
rect 390718 -21972 390774 -21916
rect 390576 -22114 390632 -22058
rect 390718 -22114 390774 -22058
rect 390576 -22256 390632 -22200
rect 390718 -22256 390774 -22200
rect 390576 -22398 390632 -22342
rect 390718 -22398 390774 -22342
rect 390576 -22540 390632 -22484
rect 390718 -22540 390774 -22484
rect 390576 -22682 390632 -22626
rect 390718 -22682 390774 -22626
rect 390576 -22824 390632 -22768
rect 390718 -22824 390774 -22768
rect 390576 -22966 390632 -22910
rect 390718 -22966 390774 -22910
rect 390576 -23108 390632 -23052
rect 390718 -23108 390774 -23052
rect 390576 -23250 390632 -23194
rect 390718 -23250 390774 -23194
rect 390576 -23392 390632 -23336
rect 390718 -23392 390774 -23336
rect 390576 -23534 390632 -23478
rect 390718 -23534 390774 -23478
rect 390576 -23676 390632 -23620
rect 390718 -23676 390774 -23620
rect 390576 -23818 390632 -23762
rect 390718 -23818 390774 -23762
rect 390576 -23960 390632 -23904
rect 390718 -23960 390774 -23904
rect 390576 -24102 390632 -24046
rect 390718 -24102 390774 -24046
rect 390576 -24244 390632 -24188
rect 390718 -24244 390774 -24188
rect 390576 -24386 390632 -24330
rect 390718 -24386 390774 -24330
rect 390576 -24528 390632 -24472
rect 390718 -24528 390774 -24472
rect 390576 -24670 390632 -24614
rect 390718 -24670 390774 -24614
rect 390576 -24812 390632 -24756
rect 390718 -24812 390774 -24756
rect 390576 -24954 390632 -24898
rect 390718 -24954 390774 -24898
rect 390576 -25096 390632 -25040
rect 390718 -25096 390774 -25040
rect 390576 -25238 390632 -25182
rect 390718 -25238 390774 -25182
rect 390576 -25380 390632 -25324
rect 390718 -25380 390774 -25324
rect 390576 -25522 390632 -25466
rect 390718 -25522 390774 -25466
rect 390980 -13736 391036 -13680
rect 391122 -13736 391178 -13680
rect 390980 -13878 391036 -13822
rect 391122 -13878 391178 -13822
rect 390980 -14020 391036 -13964
rect 391122 -14020 391178 -13964
rect 390980 -14162 391036 -14106
rect 391122 -14162 391178 -14106
rect 390980 -14304 391036 -14248
rect 391122 -14304 391178 -14248
rect 390980 -14446 391036 -14390
rect 391122 -14446 391178 -14390
rect 390980 -14588 391036 -14532
rect 391122 -14588 391178 -14532
rect 390980 -14730 391036 -14674
rect 391122 -14730 391178 -14674
rect 390980 -14872 391036 -14816
rect 391122 -14872 391178 -14816
rect 390980 -15014 391036 -14958
rect 391122 -15014 391178 -14958
rect 390980 -15156 391036 -15100
rect 391122 -15156 391178 -15100
rect 390980 -15298 391036 -15242
rect 391122 -15298 391178 -15242
rect 390980 -15440 391036 -15384
rect 391122 -15440 391178 -15384
rect 390980 -15582 391036 -15526
rect 391122 -15582 391178 -15526
rect 390980 -15724 391036 -15668
rect 391122 -15724 391178 -15668
rect 390980 -15866 391036 -15810
rect 391122 -15866 391178 -15810
rect 390980 -16008 391036 -15952
rect 391122 -16008 391178 -15952
rect 390980 -16150 391036 -16094
rect 391122 -16150 391178 -16094
rect 390980 -16292 391036 -16236
rect 391122 -16292 391178 -16236
rect 390980 -16434 391036 -16378
rect 391122 -16434 391178 -16378
rect 390980 -16576 391036 -16520
rect 391122 -16576 391178 -16520
rect 390980 -16718 391036 -16662
rect 391122 -16718 391178 -16662
rect 390980 -16860 391036 -16804
rect 391122 -16860 391178 -16804
rect 390980 -17002 391036 -16946
rect 391122 -17002 391178 -16946
rect 390980 -17144 391036 -17088
rect 391122 -17144 391178 -17088
rect 390980 -17286 391036 -17230
rect 391122 -17286 391178 -17230
rect 390980 -17428 391036 -17372
rect 391122 -17428 391178 -17372
rect 390980 -17570 391036 -17514
rect 391122 -17570 391178 -17514
rect 390980 -17712 391036 -17656
rect 391122 -17712 391178 -17656
rect 390980 -17854 391036 -17798
rect 391122 -17854 391178 -17798
rect 390980 -17996 391036 -17940
rect 391122 -17996 391178 -17940
rect 390980 -18138 391036 -18082
rect 391122 -18138 391178 -18082
rect 390980 -18280 391036 -18224
rect 391122 -18280 391178 -18224
rect 390980 -18422 391036 -18366
rect 391122 -18422 391178 -18366
rect 390980 -18564 391036 -18508
rect 391122 -18564 391178 -18508
rect 390980 -18706 391036 -18650
rect 391122 -18706 391178 -18650
rect 390980 -18848 391036 -18792
rect 391122 -18848 391178 -18792
rect 390980 -18990 391036 -18934
rect 391122 -18990 391178 -18934
rect 390980 -19132 391036 -19076
rect 391122 -19132 391178 -19076
rect 390980 -19274 391036 -19218
rect 391122 -19274 391178 -19218
rect 390980 -19416 391036 -19360
rect 391122 -19416 391178 -19360
rect 390980 -19558 391036 -19502
rect 391122 -19558 391178 -19502
rect 390980 -19700 391036 -19644
rect 391122 -19700 391178 -19644
rect 390980 -19842 391036 -19786
rect 391122 -19842 391178 -19786
rect 390980 -19984 391036 -19928
rect 391122 -19984 391178 -19928
rect 390980 -20126 391036 -20070
rect 391122 -20126 391178 -20070
rect 390980 -20268 391036 -20212
rect 391122 -20268 391178 -20212
rect 390980 -20410 391036 -20354
rect 391122 -20410 391178 -20354
rect 390980 -20552 391036 -20496
rect 391122 -20552 391178 -20496
rect 390980 -20694 391036 -20638
rect 391122 -20694 391178 -20638
rect 390980 -20836 391036 -20780
rect 391122 -20836 391178 -20780
rect 390980 -20978 391036 -20922
rect 391122 -20978 391178 -20922
rect 390980 -21120 391036 -21064
rect 391122 -21120 391178 -21064
rect 390980 -21262 391036 -21206
rect 391122 -21262 391178 -21206
rect 390980 -21404 391036 -21348
rect 391122 -21404 391178 -21348
rect 390980 -21546 391036 -21490
rect 391122 -21546 391178 -21490
rect 390980 -21688 391036 -21632
rect 391122 -21688 391178 -21632
rect 390980 -21830 391036 -21774
rect 391122 -21830 391178 -21774
rect 390980 -21972 391036 -21916
rect 391122 -21972 391178 -21916
rect 390980 -22114 391036 -22058
rect 391122 -22114 391178 -22058
rect 390980 -22256 391036 -22200
rect 391122 -22256 391178 -22200
rect 390980 -22398 391036 -22342
rect 391122 -22398 391178 -22342
rect 390980 -22540 391036 -22484
rect 391122 -22540 391178 -22484
rect 390980 -22682 391036 -22626
rect 391122 -22682 391178 -22626
rect 390980 -22824 391036 -22768
rect 391122 -22824 391178 -22768
rect 390980 -22966 391036 -22910
rect 391122 -22966 391178 -22910
rect 390980 -23108 391036 -23052
rect 391122 -23108 391178 -23052
rect 390980 -23250 391036 -23194
rect 391122 -23250 391178 -23194
rect 390980 -23392 391036 -23336
rect 391122 -23392 391178 -23336
rect 390980 -23534 391036 -23478
rect 391122 -23534 391178 -23478
rect 390980 -23676 391036 -23620
rect 391122 -23676 391178 -23620
rect 390980 -23818 391036 -23762
rect 391122 -23818 391178 -23762
rect 390980 -23960 391036 -23904
rect 391122 -23960 391178 -23904
rect 390980 -24102 391036 -24046
rect 391122 -24102 391178 -24046
rect 390980 -24244 391036 -24188
rect 391122 -24244 391178 -24188
rect 390980 -24386 391036 -24330
rect 391122 -24386 391178 -24330
rect 390980 -24528 391036 -24472
rect 391122 -24528 391178 -24472
rect 390980 -24670 391036 -24614
rect 391122 -24670 391178 -24614
rect 390980 -24812 391036 -24756
rect 391122 -24812 391178 -24756
rect 390980 -24954 391036 -24898
rect 391122 -24954 391178 -24898
rect 390980 -25096 391036 -25040
rect 391122 -25096 391178 -25040
rect 390980 -25238 391036 -25182
rect 391122 -25238 391178 -25182
rect 390980 -25380 391036 -25324
rect 391122 -25380 391178 -25324
rect 390980 -25522 391036 -25466
rect 391122 -25522 391178 -25466
rect 391376 -13736 391432 -13680
rect 391518 -13736 391574 -13680
rect 391376 -13878 391432 -13822
rect 391518 -13878 391574 -13822
rect 391376 -14020 391432 -13964
rect 391518 -14020 391574 -13964
rect 391376 -14162 391432 -14106
rect 391518 -14162 391574 -14106
rect 391376 -14304 391432 -14248
rect 391518 -14304 391574 -14248
rect 391376 -14446 391432 -14390
rect 391518 -14446 391574 -14390
rect 391376 -14588 391432 -14532
rect 391518 -14588 391574 -14532
rect 391376 -14730 391432 -14674
rect 391518 -14730 391574 -14674
rect 391376 -14872 391432 -14816
rect 391518 -14872 391574 -14816
rect 391376 -15014 391432 -14958
rect 391518 -15014 391574 -14958
rect 391376 -15156 391432 -15100
rect 391518 -15156 391574 -15100
rect 391376 -15298 391432 -15242
rect 391518 -15298 391574 -15242
rect 391376 -15440 391432 -15384
rect 391518 -15440 391574 -15384
rect 391376 -15582 391432 -15526
rect 391518 -15582 391574 -15526
rect 391376 -15724 391432 -15668
rect 391518 -15724 391574 -15668
rect 391376 -15866 391432 -15810
rect 391518 -15866 391574 -15810
rect 391376 -16008 391432 -15952
rect 391518 -16008 391574 -15952
rect 391376 -16150 391432 -16094
rect 391518 -16150 391574 -16094
rect 391376 -16292 391432 -16236
rect 391518 -16292 391574 -16236
rect 391376 -16434 391432 -16378
rect 391518 -16434 391574 -16378
rect 391376 -16576 391432 -16520
rect 391518 -16576 391574 -16520
rect 391376 -16718 391432 -16662
rect 391518 -16718 391574 -16662
rect 391376 -16860 391432 -16804
rect 391518 -16860 391574 -16804
rect 391376 -17002 391432 -16946
rect 391518 -17002 391574 -16946
rect 391376 -17144 391432 -17088
rect 391518 -17144 391574 -17088
rect 391376 -17286 391432 -17230
rect 391518 -17286 391574 -17230
rect 391376 -17428 391432 -17372
rect 391518 -17428 391574 -17372
rect 391376 -17570 391432 -17514
rect 391518 -17570 391574 -17514
rect 391376 -17712 391432 -17656
rect 391518 -17712 391574 -17656
rect 391376 -17854 391432 -17798
rect 391518 -17854 391574 -17798
rect 391376 -17996 391432 -17940
rect 391518 -17996 391574 -17940
rect 391376 -18138 391432 -18082
rect 391518 -18138 391574 -18082
rect 391376 -18280 391432 -18224
rect 391518 -18280 391574 -18224
rect 391376 -18422 391432 -18366
rect 391518 -18422 391574 -18366
rect 391376 -18564 391432 -18508
rect 391518 -18564 391574 -18508
rect 391376 -18706 391432 -18650
rect 391518 -18706 391574 -18650
rect 391376 -18848 391432 -18792
rect 391518 -18848 391574 -18792
rect 391376 -18990 391432 -18934
rect 391518 -18990 391574 -18934
rect 391376 -19132 391432 -19076
rect 391518 -19132 391574 -19076
rect 391376 -19274 391432 -19218
rect 391518 -19274 391574 -19218
rect 391376 -19416 391432 -19360
rect 391518 -19416 391574 -19360
rect 391376 -19558 391432 -19502
rect 391518 -19558 391574 -19502
rect 391376 -19700 391432 -19644
rect 391518 -19700 391574 -19644
rect 391376 -19842 391432 -19786
rect 391518 -19842 391574 -19786
rect 391376 -19984 391432 -19928
rect 391518 -19984 391574 -19928
rect 391376 -20126 391432 -20070
rect 391518 -20126 391574 -20070
rect 391376 -20268 391432 -20212
rect 391518 -20268 391574 -20212
rect 391376 -20410 391432 -20354
rect 391518 -20410 391574 -20354
rect 391376 -20552 391432 -20496
rect 391518 -20552 391574 -20496
rect 391376 -20694 391432 -20638
rect 391518 -20694 391574 -20638
rect 391376 -20836 391432 -20780
rect 391518 -20836 391574 -20780
rect 391376 -20978 391432 -20922
rect 391518 -20978 391574 -20922
rect 391376 -21120 391432 -21064
rect 391518 -21120 391574 -21064
rect 391376 -21262 391432 -21206
rect 391518 -21262 391574 -21206
rect 391376 -21404 391432 -21348
rect 391518 -21404 391574 -21348
rect 391376 -21546 391432 -21490
rect 391518 -21546 391574 -21490
rect 391376 -21688 391432 -21632
rect 391518 -21688 391574 -21632
rect 391376 -21830 391432 -21774
rect 391518 -21830 391574 -21774
rect 391376 -21972 391432 -21916
rect 391518 -21972 391574 -21916
rect 391376 -22114 391432 -22058
rect 391518 -22114 391574 -22058
rect 391376 -22256 391432 -22200
rect 391518 -22256 391574 -22200
rect 391376 -22398 391432 -22342
rect 391518 -22398 391574 -22342
rect 391376 -22540 391432 -22484
rect 391518 -22540 391574 -22484
rect 391376 -22682 391432 -22626
rect 391518 -22682 391574 -22626
rect 391376 -22824 391432 -22768
rect 391518 -22824 391574 -22768
rect 391376 -22966 391432 -22910
rect 391518 -22966 391574 -22910
rect 391376 -23108 391432 -23052
rect 391518 -23108 391574 -23052
rect 391376 -23250 391432 -23194
rect 391518 -23250 391574 -23194
rect 391376 -23392 391432 -23336
rect 391518 -23392 391574 -23336
rect 391376 -23534 391432 -23478
rect 391518 -23534 391574 -23478
rect 391376 -23676 391432 -23620
rect 391518 -23676 391574 -23620
rect 391376 -23818 391432 -23762
rect 391518 -23818 391574 -23762
rect 391376 -23960 391432 -23904
rect 391518 -23960 391574 -23904
rect 391376 -24102 391432 -24046
rect 391518 -24102 391574 -24046
rect 391376 -24244 391432 -24188
rect 391518 -24244 391574 -24188
rect 391376 -24386 391432 -24330
rect 391518 -24386 391574 -24330
rect 391376 -24528 391432 -24472
rect 391518 -24528 391574 -24472
rect 391376 -24670 391432 -24614
rect 391518 -24670 391574 -24614
rect 391376 -24812 391432 -24756
rect 391518 -24812 391574 -24756
rect 391376 -24954 391432 -24898
rect 391518 -24954 391574 -24898
rect 391376 -25096 391432 -25040
rect 391518 -25096 391574 -25040
rect 391376 -25238 391432 -25182
rect 391518 -25238 391574 -25182
rect 391376 -25380 391432 -25324
rect 391518 -25380 391574 -25324
rect 391376 -25522 391432 -25466
rect 391518 -25522 391574 -25466
rect 391776 -13736 391832 -13680
rect 391918 -13736 391974 -13680
rect 391776 -13878 391832 -13822
rect 391918 -13878 391974 -13822
rect 391776 -14020 391832 -13964
rect 391918 -14020 391974 -13964
rect 391776 -14162 391832 -14106
rect 391918 -14162 391974 -14106
rect 391776 -14304 391832 -14248
rect 391918 -14304 391974 -14248
rect 391776 -14446 391832 -14390
rect 391918 -14446 391974 -14390
rect 391776 -14588 391832 -14532
rect 391918 -14588 391974 -14532
rect 391776 -14730 391832 -14674
rect 391918 -14730 391974 -14674
rect 391776 -14872 391832 -14816
rect 391918 -14872 391974 -14816
rect 391776 -15014 391832 -14958
rect 391918 -15014 391974 -14958
rect 391776 -15156 391832 -15100
rect 391918 -15156 391974 -15100
rect 391776 -15298 391832 -15242
rect 391918 -15298 391974 -15242
rect 391776 -15440 391832 -15384
rect 391918 -15440 391974 -15384
rect 391776 -15582 391832 -15526
rect 391918 -15582 391974 -15526
rect 391776 -15724 391832 -15668
rect 391918 -15724 391974 -15668
rect 391776 -15866 391832 -15810
rect 391918 -15866 391974 -15810
rect 391776 -16008 391832 -15952
rect 391918 -16008 391974 -15952
rect 391776 -16150 391832 -16094
rect 391918 -16150 391974 -16094
rect 391776 -16292 391832 -16236
rect 391918 -16292 391974 -16236
rect 391776 -16434 391832 -16378
rect 391918 -16434 391974 -16378
rect 391776 -16576 391832 -16520
rect 391918 -16576 391974 -16520
rect 391776 -16718 391832 -16662
rect 391918 -16718 391974 -16662
rect 391776 -16860 391832 -16804
rect 391918 -16860 391974 -16804
rect 391776 -17002 391832 -16946
rect 391918 -17002 391974 -16946
rect 391776 -17144 391832 -17088
rect 391918 -17144 391974 -17088
rect 391776 -17286 391832 -17230
rect 391918 -17286 391974 -17230
rect 391776 -17428 391832 -17372
rect 391918 -17428 391974 -17372
rect 391776 -17570 391832 -17514
rect 391918 -17570 391974 -17514
rect 391776 -17712 391832 -17656
rect 391918 -17712 391974 -17656
rect 391776 -17854 391832 -17798
rect 391918 -17854 391974 -17798
rect 391776 -17996 391832 -17940
rect 391918 -17996 391974 -17940
rect 391776 -18138 391832 -18082
rect 391918 -18138 391974 -18082
rect 391776 -18280 391832 -18224
rect 391918 -18280 391974 -18224
rect 391776 -18422 391832 -18366
rect 391918 -18422 391974 -18366
rect 391776 -18564 391832 -18508
rect 391918 -18564 391974 -18508
rect 391776 -18706 391832 -18650
rect 391918 -18706 391974 -18650
rect 391776 -18848 391832 -18792
rect 391918 -18848 391974 -18792
rect 391776 -18990 391832 -18934
rect 391918 -18990 391974 -18934
rect 391776 -19132 391832 -19076
rect 391918 -19132 391974 -19076
rect 391776 -19274 391832 -19218
rect 391918 -19274 391974 -19218
rect 391776 -19416 391832 -19360
rect 391918 -19416 391974 -19360
rect 391776 -19558 391832 -19502
rect 391918 -19558 391974 -19502
rect 391776 -19700 391832 -19644
rect 391918 -19700 391974 -19644
rect 391776 -19842 391832 -19786
rect 391918 -19842 391974 -19786
rect 391776 -19984 391832 -19928
rect 391918 -19984 391974 -19928
rect 391776 -20126 391832 -20070
rect 391918 -20126 391974 -20070
rect 391776 -20268 391832 -20212
rect 391918 -20268 391974 -20212
rect 391776 -20410 391832 -20354
rect 391918 -20410 391974 -20354
rect 391776 -20552 391832 -20496
rect 391918 -20552 391974 -20496
rect 391776 -20694 391832 -20638
rect 391918 -20694 391974 -20638
rect 391776 -20836 391832 -20780
rect 391918 -20836 391974 -20780
rect 391776 -20978 391832 -20922
rect 391918 -20978 391974 -20922
rect 391776 -21120 391832 -21064
rect 391918 -21120 391974 -21064
rect 391776 -21262 391832 -21206
rect 391918 -21262 391974 -21206
rect 391776 -21404 391832 -21348
rect 391918 -21404 391974 -21348
rect 391776 -21546 391832 -21490
rect 391918 -21546 391974 -21490
rect 391776 -21688 391832 -21632
rect 391918 -21688 391974 -21632
rect 391776 -21830 391832 -21774
rect 391918 -21830 391974 -21774
rect 391776 -21972 391832 -21916
rect 391918 -21972 391974 -21916
rect 391776 -22114 391832 -22058
rect 391918 -22114 391974 -22058
rect 391776 -22256 391832 -22200
rect 391918 -22256 391974 -22200
rect 391776 -22398 391832 -22342
rect 391918 -22398 391974 -22342
rect 391776 -22540 391832 -22484
rect 391918 -22540 391974 -22484
rect 391776 -22682 391832 -22626
rect 391918 -22682 391974 -22626
rect 391776 -22824 391832 -22768
rect 391918 -22824 391974 -22768
rect 391776 -22966 391832 -22910
rect 391918 -22966 391974 -22910
rect 391776 -23108 391832 -23052
rect 391918 -23108 391974 -23052
rect 391776 -23250 391832 -23194
rect 391918 -23250 391974 -23194
rect 391776 -23392 391832 -23336
rect 391918 -23392 391974 -23336
rect 391776 -23534 391832 -23478
rect 391918 -23534 391974 -23478
rect 391776 -23676 391832 -23620
rect 391918 -23676 391974 -23620
rect 391776 -23818 391832 -23762
rect 391918 -23818 391974 -23762
rect 391776 -23960 391832 -23904
rect 391918 -23960 391974 -23904
rect 391776 -24102 391832 -24046
rect 391918 -24102 391974 -24046
rect 391776 -24244 391832 -24188
rect 391918 -24244 391974 -24188
rect 391776 -24386 391832 -24330
rect 391918 -24386 391974 -24330
rect 391776 -24528 391832 -24472
rect 391918 -24528 391974 -24472
rect 391776 -24670 391832 -24614
rect 391918 -24670 391974 -24614
rect 391776 -24812 391832 -24756
rect 391918 -24812 391974 -24756
rect 391776 -24954 391832 -24898
rect 391918 -24954 391974 -24898
rect 391776 -25096 391832 -25040
rect 391918 -25096 391974 -25040
rect 391776 -25238 391832 -25182
rect 391918 -25238 391974 -25182
rect 391776 -25380 391832 -25324
rect 391918 -25380 391974 -25324
rect 391776 -25522 391832 -25466
rect 391918 -25522 391974 -25466
rect 392173 -13736 392229 -13680
rect 392315 -13736 392371 -13680
rect 392173 -13878 392229 -13822
rect 392315 -13878 392371 -13822
rect 392173 -14020 392229 -13964
rect 392315 -14020 392371 -13964
rect 392173 -14162 392229 -14106
rect 392315 -14162 392371 -14106
rect 392173 -14304 392229 -14248
rect 392315 -14304 392371 -14248
rect 392173 -14446 392229 -14390
rect 392315 -14446 392371 -14390
rect 392173 -14588 392229 -14532
rect 392315 -14588 392371 -14532
rect 392173 -14730 392229 -14674
rect 392315 -14730 392371 -14674
rect 392173 -14872 392229 -14816
rect 392315 -14872 392371 -14816
rect 392173 -15014 392229 -14958
rect 392315 -15014 392371 -14958
rect 392173 -15156 392229 -15100
rect 392315 -15156 392371 -15100
rect 392173 -15298 392229 -15242
rect 392315 -15298 392371 -15242
rect 392173 -15440 392229 -15384
rect 392315 -15440 392371 -15384
rect 392173 -15582 392229 -15526
rect 392315 -15582 392371 -15526
rect 392173 -15724 392229 -15668
rect 392315 -15724 392371 -15668
rect 392173 -15866 392229 -15810
rect 392315 -15866 392371 -15810
rect 392173 -16008 392229 -15952
rect 392315 -16008 392371 -15952
rect 392173 -16150 392229 -16094
rect 392315 -16150 392371 -16094
rect 392173 -16292 392229 -16236
rect 392315 -16292 392371 -16236
rect 392173 -16434 392229 -16378
rect 392315 -16434 392371 -16378
rect 392173 -16576 392229 -16520
rect 392315 -16576 392371 -16520
rect 392173 -16718 392229 -16662
rect 392315 -16718 392371 -16662
rect 392173 -16860 392229 -16804
rect 392315 -16860 392371 -16804
rect 392173 -17002 392229 -16946
rect 392315 -17002 392371 -16946
rect 392173 -17144 392229 -17088
rect 392315 -17144 392371 -17088
rect 392173 -17286 392229 -17230
rect 392315 -17286 392371 -17230
rect 392173 -17428 392229 -17372
rect 392315 -17428 392371 -17372
rect 392173 -17570 392229 -17514
rect 392315 -17570 392371 -17514
rect 392173 -17712 392229 -17656
rect 392315 -17712 392371 -17656
rect 392173 -17854 392229 -17798
rect 392315 -17854 392371 -17798
rect 392173 -17996 392229 -17940
rect 392315 -17996 392371 -17940
rect 392173 -18138 392229 -18082
rect 392315 -18138 392371 -18082
rect 392173 -18280 392229 -18224
rect 392315 -18280 392371 -18224
rect 392173 -18422 392229 -18366
rect 392315 -18422 392371 -18366
rect 392173 -18564 392229 -18508
rect 392315 -18564 392371 -18508
rect 392173 -18706 392229 -18650
rect 392315 -18706 392371 -18650
rect 392173 -18848 392229 -18792
rect 392315 -18848 392371 -18792
rect 392173 -18990 392229 -18934
rect 392315 -18990 392371 -18934
rect 392173 -19132 392229 -19076
rect 392315 -19132 392371 -19076
rect 392173 -19274 392229 -19218
rect 392315 -19274 392371 -19218
rect 392173 -19416 392229 -19360
rect 392315 -19416 392371 -19360
rect 392173 -19558 392229 -19502
rect 392315 -19558 392371 -19502
rect 392173 -19700 392229 -19644
rect 392315 -19700 392371 -19644
rect 392173 -19842 392229 -19786
rect 392315 -19842 392371 -19786
rect 392173 -19984 392229 -19928
rect 392315 -19984 392371 -19928
rect 392173 -20126 392229 -20070
rect 392315 -20126 392371 -20070
rect 392173 -20268 392229 -20212
rect 392315 -20268 392371 -20212
rect 392173 -20410 392229 -20354
rect 392315 -20410 392371 -20354
rect 392173 -20552 392229 -20496
rect 392315 -20552 392371 -20496
rect 392173 -20694 392229 -20638
rect 392315 -20694 392371 -20638
rect 392173 -20836 392229 -20780
rect 392315 -20836 392371 -20780
rect 392173 -20978 392229 -20922
rect 392315 -20978 392371 -20922
rect 392173 -21120 392229 -21064
rect 392315 -21120 392371 -21064
rect 392173 -21262 392229 -21206
rect 392315 -21262 392371 -21206
rect 392173 -21404 392229 -21348
rect 392315 -21404 392371 -21348
rect 392173 -21546 392229 -21490
rect 392315 -21546 392371 -21490
rect 392173 -21688 392229 -21632
rect 392315 -21688 392371 -21632
rect 392173 -21830 392229 -21774
rect 392315 -21830 392371 -21774
rect 392173 -21972 392229 -21916
rect 392315 -21972 392371 -21916
rect 392173 -22114 392229 -22058
rect 392315 -22114 392371 -22058
rect 392173 -22256 392229 -22200
rect 392315 -22256 392371 -22200
rect 392173 -22398 392229 -22342
rect 392315 -22398 392371 -22342
rect 392173 -22540 392229 -22484
rect 392315 -22540 392371 -22484
rect 392173 -22682 392229 -22626
rect 392315 -22682 392371 -22626
rect 392173 -22824 392229 -22768
rect 392315 -22824 392371 -22768
rect 392173 -22966 392229 -22910
rect 392315 -22966 392371 -22910
rect 392173 -23108 392229 -23052
rect 392315 -23108 392371 -23052
rect 392173 -23250 392229 -23194
rect 392315 -23250 392371 -23194
rect 392173 -23392 392229 -23336
rect 392315 -23392 392371 -23336
rect 392173 -23534 392229 -23478
rect 392315 -23534 392371 -23478
rect 392173 -23676 392229 -23620
rect 392315 -23676 392371 -23620
rect 392173 -23818 392229 -23762
rect 392315 -23818 392371 -23762
rect 392173 -23960 392229 -23904
rect 392315 -23960 392371 -23904
rect 392173 -24102 392229 -24046
rect 392315 -24102 392371 -24046
rect 392173 -24244 392229 -24188
rect 392315 -24244 392371 -24188
rect 392173 -24386 392229 -24330
rect 392315 -24386 392371 -24330
rect 392173 -24528 392229 -24472
rect 392315 -24528 392371 -24472
rect 392173 -24670 392229 -24614
rect 392315 -24670 392371 -24614
rect 392173 -24812 392229 -24756
rect 392315 -24812 392371 -24756
rect 392173 -24954 392229 -24898
rect 392315 -24954 392371 -24898
rect 392173 -25096 392229 -25040
rect 392315 -25096 392371 -25040
rect 392173 -25238 392229 -25182
rect 392315 -25238 392371 -25182
rect 392173 -25380 392229 -25324
rect 392315 -25380 392371 -25324
rect 392173 -25522 392229 -25466
rect 392315 -25522 392371 -25466
rect 392578 -13736 392634 -13680
rect 392720 -13736 392776 -13680
rect 392578 -13878 392634 -13822
rect 392720 -13878 392776 -13822
rect 392578 -14020 392634 -13964
rect 392720 -14020 392776 -13964
rect 392578 -14162 392634 -14106
rect 392720 -14162 392776 -14106
rect 392578 -14304 392634 -14248
rect 392720 -14304 392776 -14248
rect 392578 -14446 392634 -14390
rect 392720 -14446 392776 -14390
rect 392578 -14588 392634 -14532
rect 392720 -14588 392776 -14532
rect 392578 -14730 392634 -14674
rect 392720 -14730 392776 -14674
rect 392578 -14872 392634 -14816
rect 392720 -14872 392776 -14816
rect 392578 -15014 392634 -14958
rect 392720 -15014 392776 -14958
rect 392578 -15156 392634 -15100
rect 392720 -15156 392776 -15100
rect 392578 -15298 392634 -15242
rect 392720 -15298 392776 -15242
rect 392578 -15440 392634 -15384
rect 392720 -15440 392776 -15384
rect 392578 -15582 392634 -15526
rect 392720 -15582 392776 -15526
rect 392578 -15724 392634 -15668
rect 392720 -15724 392776 -15668
rect 392578 -15866 392634 -15810
rect 392720 -15866 392776 -15810
rect 392578 -16008 392634 -15952
rect 392720 -16008 392776 -15952
rect 392578 -16150 392634 -16094
rect 392720 -16150 392776 -16094
rect 392578 -16292 392634 -16236
rect 392720 -16292 392776 -16236
rect 392578 -16434 392634 -16378
rect 392720 -16434 392776 -16378
rect 392578 -16576 392634 -16520
rect 392720 -16576 392776 -16520
rect 392578 -16718 392634 -16662
rect 392720 -16718 392776 -16662
rect 392578 -16860 392634 -16804
rect 392720 -16860 392776 -16804
rect 392578 -17002 392634 -16946
rect 392720 -17002 392776 -16946
rect 392578 -17144 392634 -17088
rect 392720 -17144 392776 -17088
rect 392578 -17286 392634 -17230
rect 392720 -17286 392776 -17230
rect 392578 -17428 392634 -17372
rect 392720 -17428 392776 -17372
rect 392578 -17570 392634 -17514
rect 392720 -17570 392776 -17514
rect 392578 -17712 392634 -17656
rect 392720 -17712 392776 -17656
rect 392578 -17854 392634 -17798
rect 392720 -17854 392776 -17798
rect 392578 -17996 392634 -17940
rect 392720 -17996 392776 -17940
rect 392578 -18138 392634 -18082
rect 392720 -18138 392776 -18082
rect 392578 -18280 392634 -18224
rect 392720 -18280 392776 -18224
rect 392578 -18422 392634 -18366
rect 392720 -18422 392776 -18366
rect 392578 -18564 392634 -18508
rect 392720 -18564 392776 -18508
rect 392578 -18706 392634 -18650
rect 392720 -18706 392776 -18650
rect 392578 -18848 392634 -18792
rect 392720 -18848 392776 -18792
rect 392578 -18990 392634 -18934
rect 392720 -18990 392776 -18934
rect 392578 -19132 392634 -19076
rect 392720 -19132 392776 -19076
rect 392578 -19274 392634 -19218
rect 392720 -19274 392776 -19218
rect 392578 -19416 392634 -19360
rect 392720 -19416 392776 -19360
rect 392578 -19558 392634 -19502
rect 392720 -19558 392776 -19502
rect 392578 -19700 392634 -19644
rect 392720 -19700 392776 -19644
rect 392578 -19842 392634 -19786
rect 392720 -19842 392776 -19786
rect 392578 -19984 392634 -19928
rect 392720 -19984 392776 -19928
rect 392578 -20126 392634 -20070
rect 392720 -20126 392776 -20070
rect 392578 -20268 392634 -20212
rect 392720 -20268 392776 -20212
rect 392578 -20410 392634 -20354
rect 392720 -20410 392776 -20354
rect 392578 -20552 392634 -20496
rect 392720 -20552 392776 -20496
rect 392578 -20694 392634 -20638
rect 392720 -20694 392776 -20638
rect 392578 -20836 392634 -20780
rect 392720 -20836 392776 -20780
rect 392578 -20978 392634 -20922
rect 392720 -20978 392776 -20922
rect 392578 -21120 392634 -21064
rect 392720 -21120 392776 -21064
rect 392578 -21262 392634 -21206
rect 392720 -21262 392776 -21206
rect 392578 -21404 392634 -21348
rect 392720 -21404 392776 -21348
rect 392578 -21546 392634 -21490
rect 392720 -21546 392776 -21490
rect 392578 -21688 392634 -21632
rect 392720 -21688 392776 -21632
rect 392578 -21830 392634 -21774
rect 392720 -21830 392776 -21774
rect 392578 -21972 392634 -21916
rect 392720 -21972 392776 -21916
rect 392578 -22114 392634 -22058
rect 392720 -22114 392776 -22058
rect 392578 -22256 392634 -22200
rect 392720 -22256 392776 -22200
rect 392578 -22398 392634 -22342
rect 392720 -22398 392776 -22342
rect 392578 -22540 392634 -22484
rect 392720 -22540 392776 -22484
rect 392578 -22682 392634 -22626
rect 392720 -22682 392776 -22626
rect 392578 -22824 392634 -22768
rect 392720 -22824 392776 -22768
rect 392578 -22966 392634 -22910
rect 392720 -22966 392776 -22910
rect 392578 -23108 392634 -23052
rect 392720 -23108 392776 -23052
rect 392578 -23250 392634 -23194
rect 392720 -23250 392776 -23194
rect 392578 -23392 392634 -23336
rect 392720 -23392 392776 -23336
rect 392578 -23534 392634 -23478
rect 392720 -23534 392776 -23478
rect 392578 -23676 392634 -23620
rect 392720 -23676 392776 -23620
rect 392578 -23818 392634 -23762
rect 392720 -23818 392776 -23762
rect 392578 -23960 392634 -23904
rect 392720 -23960 392776 -23904
rect 392578 -24102 392634 -24046
rect 392720 -24102 392776 -24046
rect 392578 -24244 392634 -24188
rect 392720 -24244 392776 -24188
rect 392578 -24386 392634 -24330
rect 392720 -24386 392776 -24330
rect 392578 -24528 392634 -24472
rect 392720 -24528 392776 -24472
rect 392578 -24670 392634 -24614
rect 392720 -24670 392776 -24614
rect 392578 -24812 392634 -24756
rect 392720 -24812 392776 -24756
rect 392578 -24954 392634 -24898
rect 392720 -24954 392776 -24898
rect 392578 -25096 392634 -25040
rect 392720 -25096 392776 -25040
rect 392578 -25238 392634 -25182
rect 392720 -25238 392776 -25182
rect 392578 -25380 392634 -25324
rect 392720 -25380 392776 -25324
rect 392578 -25522 392634 -25466
rect 392720 -25522 392776 -25466
rect 392978 -13736 393034 -13680
rect 393120 -13736 393176 -13680
rect 392978 -13878 393034 -13822
rect 393120 -13878 393176 -13822
rect 392978 -14020 393034 -13964
rect 393120 -14020 393176 -13964
rect 392978 -14162 393034 -14106
rect 393120 -14162 393176 -14106
rect 392978 -14304 393034 -14248
rect 393120 -14304 393176 -14248
rect 392978 -14446 393034 -14390
rect 393120 -14446 393176 -14390
rect 392978 -14588 393034 -14532
rect 393120 -14588 393176 -14532
rect 392978 -14730 393034 -14674
rect 393120 -14730 393176 -14674
rect 392978 -14872 393034 -14816
rect 393120 -14872 393176 -14816
rect 392978 -15014 393034 -14958
rect 393120 -15014 393176 -14958
rect 392978 -15156 393034 -15100
rect 393120 -15156 393176 -15100
rect 392978 -15298 393034 -15242
rect 393120 -15298 393176 -15242
rect 392978 -15440 393034 -15384
rect 393120 -15440 393176 -15384
rect 392978 -15582 393034 -15526
rect 393120 -15582 393176 -15526
rect 392978 -15724 393034 -15668
rect 393120 -15724 393176 -15668
rect 392978 -15866 393034 -15810
rect 393120 -15866 393176 -15810
rect 392978 -16008 393034 -15952
rect 393120 -16008 393176 -15952
rect 392978 -16150 393034 -16094
rect 393120 -16150 393176 -16094
rect 392978 -16292 393034 -16236
rect 393120 -16292 393176 -16236
rect 392978 -16434 393034 -16378
rect 393120 -16434 393176 -16378
rect 392978 -16576 393034 -16520
rect 393120 -16576 393176 -16520
rect 392978 -16718 393034 -16662
rect 393120 -16718 393176 -16662
rect 392978 -16860 393034 -16804
rect 393120 -16860 393176 -16804
rect 392978 -17002 393034 -16946
rect 393120 -17002 393176 -16946
rect 392978 -17144 393034 -17088
rect 393120 -17144 393176 -17088
rect 392978 -17286 393034 -17230
rect 393120 -17286 393176 -17230
rect 392978 -17428 393034 -17372
rect 393120 -17428 393176 -17372
rect 392978 -17570 393034 -17514
rect 393120 -17570 393176 -17514
rect 392978 -17712 393034 -17656
rect 393120 -17712 393176 -17656
rect 392978 -17854 393034 -17798
rect 393120 -17854 393176 -17798
rect 392978 -17996 393034 -17940
rect 393120 -17996 393176 -17940
rect 392978 -18138 393034 -18082
rect 393120 -18138 393176 -18082
rect 392978 -18280 393034 -18224
rect 393120 -18280 393176 -18224
rect 392978 -18422 393034 -18366
rect 393120 -18422 393176 -18366
rect 392978 -18564 393034 -18508
rect 393120 -18564 393176 -18508
rect 392978 -18706 393034 -18650
rect 393120 -18706 393176 -18650
rect 392978 -18848 393034 -18792
rect 393120 -18848 393176 -18792
rect 392978 -18990 393034 -18934
rect 393120 -18990 393176 -18934
rect 392978 -19132 393034 -19076
rect 393120 -19132 393176 -19076
rect 392978 -19274 393034 -19218
rect 393120 -19274 393176 -19218
rect 392978 -19416 393034 -19360
rect 393120 -19416 393176 -19360
rect 392978 -19558 393034 -19502
rect 393120 -19558 393176 -19502
rect 392978 -19700 393034 -19644
rect 393120 -19700 393176 -19644
rect 392978 -19842 393034 -19786
rect 393120 -19842 393176 -19786
rect 392978 -19984 393034 -19928
rect 393120 -19984 393176 -19928
rect 392978 -20126 393034 -20070
rect 393120 -20126 393176 -20070
rect 392978 -20268 393034 -20212
rect 393120 -20268 393176 -20212
rect 392978 -20410 393034 -20354
rect 393120 -20410 393176 -20354
rect 392978 -20552 393034 -20496
rect 393120 -20552 393176 -20496
rect 392978 -20694 393034 -20638
rect 393120 -20694 393176 -20638
rect 392978 -20836 393034 -20780
rect 393120 -20836 393176 -20780
rect 392978 -20978 393034 -20922
rect 393120 -20978 393176 -20922
rect 392978 -21120 393034 -21064
rect 393120 -21120 393176 -21064
rect 392978 -21262 393034 -21206
rect 393120 -21262 393176 -21206
rect 392978 -21404 393034 -21348
rect 393120 -21404 393176 -21348
rect 392978 -21546 393034 -21490
rect 393120 -21546 393176 -21490
rect 392978 -21688 393034 -21632
rect 393120 -21688 393176 -21632
rect 392978 -21830 393034 -21774
rect 393120 -21830 393176 -21774
rect 392978 -21972 393034 -21916
rect 393120 -21972 393176 -21916
rect 392978 -22114 393034 -22058
rect 393120 -22114 393176 -22058
rect 392978 -22256 393034 -22200
rect 393120 -22256 393176 -22200
rect 392978 -22398 393034 -22342
rect 393120 -22398 393176 -22342
rect 392978 -22540 393034 -22484
rect 393120 -22540 393176 -22484
rect 392978 -22682 393034 -22626
rect 393120 -22682 393176 -22626
rect 392978 -22824 393034 -22768
rect 393120 -22824 393176 -22768
rect 392978 -22966 393034 -22910
rect 393120 -22966 393176 -22910
rect 392978 -23108 393034 -23052
rect 393120 -23108 393176 -23052
rect 392978 -23250 393034 -23194
rect 393120 -23250 393176 -23194
rect 392978 -23392 393034 -23336
rect 393120 -23392 393176 -23336
rect 392978 -23534 393034 -23478
rect 393120 -23534 393176 -23478
rect 392978 -23676 393034 -23620
rect 393120 -23676 393176 -23620
rect 392978 -23818 393034 -23762
rect 393120 -23818 393176 -23762
rect 392978 -23960 393034 -23904
rect 393120 -23960 393176 -23904
rect 392978 -24102 393034 -24046
rect 393120 -24102 393176 -24046
rect 392978 -24244 393034 -24188
rect 393120 -24244 393176 -24188
rect 392978 -24386 393034 -24330
rect 393120 -24386 393176 -24330
rect 392978 -24528 393034 -24472
rect 393120 -24528 393176 -24472
rect 392978 -24670 393034 -24614
rect 393120 -24670 393176 -24614
rect 392978 -24812 393034 -24756
rect 393120 -24812 393176 -24756
rect 392978 -24954 393034 -24898
rect 393120 -24954 393176 -24898
rect 392978 -25096 393034 -25040
rect 393120 -25096 393176 -25040
rect 392978 -25238 393034 -25182
rect 393120 -25238 393176 -25182
rect 392978 -25380 393034 -25324
rect 393120 -25380 393176 -25324
rect 392978 -25522 393034 -25466
rect 393120 -25522 393176 -25466
rect 393383 -13736 393439 -13680
rect 393525 -13736 393581 -13680
rect 393383 -13878 393439 -13822
rect 393525 -13878 393581 -13822
rect 393383 -14020 393439 -13964
rect 393525 -14020 393581 -13964
rect 393383 -14162 393439 -14106
rect 393525 -14162 393581 -14106
rect 393383 -14304 393439 -14248
rect 393525 -14304 393581 -14248
rect 393383 -14446 393439 -14390
rect 393525 -14446 393581 -14390
rect 393383 -14588 393439 -14532
rect 393525 -14588 393581 -14532
rect 393383 -14730 393439 -14674
rect 393525 -14730 393581 -14674
rect 393383 -14872 393439 -14816
rect 393525 -14872 393581 -14816
rect 393383 -15014 393439 -14958
rect 393525 -15014 393581 -14958
rect 393383 -15156 393439 -15100
rect 393525 -15156 393581 -15100
rect 393383 -15298 393439 -15242
rect 393525 -15298 393581 -15242
rect 393383 -15440 393439 -15384
rect 393525 -15440 393581 -15384
rect 393383 -15582 393439 -15526
rect 393525 -15582 393581 -15526
rect 393383 -15724 393439 -15668
rect 393525 -15724 393581 -15668
rect 393383 -15866 393439 -15810
rect 393525 -15866 393581 -15810
rect 393383 -16008 393439 -15952
rect 393525 -16008 393581 -15952
rect 393383 -16150 393439 -16094
rect 393525 -16150 393581 -16094
rect 393383 -16292 393439 -16236
rect 393525 -16292 393581 -16236
rect 393383 -16434 393439 -16378
rect 393525 -16434 393581 -16378
rect 393383 -16576 393439 -16520
rect 393525 -16576 393581 -16520
rect 393383 -16718 393439 -16662
rect 393525 -16718 393581 -16662
rect 393383 -16860 393439 -16804
rect 393525 -16860 393581 -16804
rect 393383 -17002 393439 -16946
rect 393525 -17002 393581 -16946
rect 393383 -17144 393439 -17088
rect 393525 -17144 393581 -17088
rect 393383 -17286 393439 -17230
rect 393525 -17286 393581 -17230
rect 393383 -17428 393439 -17372
rect 393525 -17428 393581 -17372
rect 393383 -17570 393439 -17514
rect 393525 -17570 393581 -17514
rect 393383 -17712 393439 -17656
rect 393525 -17712 393581 -17656
rect 393383 -17854 393439 -17798
rect 393525 -17854 393581 -17798
rect 393383 -17996 393439 -17940
rect 393525 -17996 393581 -17940
rect 393383 -18138 393439 -18082
rect 393525 -18138 393581 -18082
rect 393383 -18280 393439 -18224
rect 393525 -18280 393581 -18224
rect 393383 -18422 393439 -18366
rect 393525 -18422 393581 -18366
rect 393383 -18564 393439 -18508
rect 393525 -18564 393581 -18508
rect 393383 -18706 393439 -18650
rect 393525 -18706 393581 -18650
rect 393383 -18848 393439 -18792
rect 393525 -18848 393581 -18792
rect 393383 -18990 393439 -18934
rect 393525 -18990 393581 -18934
rect 393383 -19132 393439 -19076
rect 393525 -19132 393581 -19076
rect 393383 -19274 393439 -19218
rect 393525 -19274 393581 -19218
rect 393383 -19416 393439 -19360
rect 393525 -19416 393581 -19360
rect 393383 -19558 393439 -19502
rect 393525 -19558 393581 -19502
rect 393383 -19700 393439 -19644
rect 393525 -19700 393581 -19644
rect 393383 -19842 393439 -19786
rect 393525 -19842 393581 -19786
rect 393383 -19984 393439 -19928
rect 393525 -19984 393581 -19928
rect 393383 -20126 393439 -20070
rect 393525 -20126 393581 -20070
rect 393383 -20268 393439 -20212
rect 393525 -20268 393581 -20212
rect 393383 -20410 393439 -20354
rect 393525 -20410 393581 -20354
rect 393383 -20552 393439 -20496
rect 393525 -20552 393581 -20496
rect 393383 -20694 393439 -20638
rect 393525 -20694 393581 -20638
rect 393383 -20836 393439 -20780
rect 393525 -20836 393581 -20780
rect 393383 -20978 393439 -20922
rect 393525 -20978 393581 -20922
rect 393383 -21120 393439 -21064
rect 393525 -21120 393581 -21064
rect 393383 -21262 393439 -21206
rect 393525 -21262 393581 -21206
rect 393383 -21404 393439 -21348
rect 393525 -21404 393581 -21348
rect 393383 -21546 393439 -21490
rect 393525 -21546 393581 -21490
rect 393383 -21688 393439 -21632
rect 393525 -21688 393581 -21632
rect 393383 -21830 393439 -21774
rect 393525 -21830 393581 -21774
rect 393383 -21972 393439 -21916
rect 393525 -21972 393581 -21916
rect 393383 -22114 393439 -22058
rect 393525 -22114 393581 -22058
rect 393383 -22256 393439 -22200
rect 393525 -22256 393581 -22200
rect 393383 -22398 393439 -22342
rect 393525 -22398 393581 -22342
rect 393383 -22540 393439 -22484
rect 393525 -22540 393581 -22484
rect 393383 -22682 393439 -22626
rect 393525 -22682 393581 -22626
rect 393383 -22824 393439 -22768
rect 393525 -22824 393581 -22768
rect 393383 -22966 393439 -22910
rect 393525 -22966 393581 -22910
rect 393383 -23108 393439 -23052
rect 393525 -23108 393581 -23052
rect 393383 -23250 393439 -23194
rect 393525 -23250 393581 -23194
rect 393383 -23392 393439 -23336
rect 393525 -23392 393581 -23336
rect 393383 -23534 393439 -23478
rect 393525 -23534 393581 -23478
rect 393383 -23676 393439 -23620
rect 393525 -23676 393581 -23620
rect 393383 -23818 393439 -23762
rect 393525 -23818 393581 -23762
rect 393383 -23960 393439 -23904
rect 393525 -23960 393581 -23904
rect 393383 -24102 393439 -24046
rect 393525 -24102 393581 -24046
rect 393383 -24244 393439 -24188
rect 393525 -24244 393581 -24188
rect 393383 -24386 393439 -24330
rect 393525 -24386 393581 -24330
rect 393383 -24528 393439 -24472
rect 393525 -24528 393581 -24472
rect 393383 -24670 393439 -24614
rect 393525 -24670 393581 -24614
rect 393383 -24812 393439 -24756
rect 393525 -24812 393581 -24756
rect 393383 -24954 393439 -24898
rect 393525 -24954 393581 -24898
rect 393383 -25096 393439 -25040
rect 393525 -25096 393581 -25040
rect 393383 -25238 393439 -25182
rect 393525 -25238 393581 -25182
rect 393383 -25380 393439 -25324
rect 393525 -25380 393581 -25324
rect 393383 -25522 393439 -25466
rect 393525 -25522 393581 -25466
rect 393780 -13736 393836 -13680
rect 393922 -13736 393978 -13680
rect 393780 -13878 393836 -13822
rect 393922 -13878 393978 -13822
rect 393780 -14020 393836 -13964
rect 393922 -14020 393978 -13964
rect 393780 -14162 393836 -14106
rect 393922 -14162 393978 -14106
rect 393780 -14304 393836 -14248
rect 393922 -14304 393978 -14248
rect 393780 -14446 393836 -14390
rect 393922 -14446 393978 -14390
rect 393780 -14588 393836 -14532
rect 393922 -14588 393978 -14532
rect 393780 -14730 393836 -14674
rect 393922 -14730 393978 -14674
rect 393780 -14872 393836 -14816
rect 393922 -14872 393978 -14816
rect 393780 -15014 393836 -14958
rect 393922 -15014 393978 -14958
rect 393780 -15156 393836 -15100
rect 393922 -15156 393978 -15100
rect 393780 -15298 393836 -15242
rect 393922 -15298 393978 -15242
rect 393780 -15440 393836 -15384
rect 393922 -15440 393978 -15384
rect 393780 -15582 393836 -15526
rect 393922 -15582 393978 -15526
rect 393780 -15724 393836 -15668
rect 393922 -15724 393978 -15668
rect 393780 -15866 393836 -15810
rect 393922 -15866 393978 -15810
rect 393780 -16008 393836 -15952
rect 393922 -16008 393978 -15952
rect 393780 -16150 393836 -16094
rect 393922 -16150 393978 -16094
rect 393780 -16292 393836 -16236
rect 393922 -16292 393978 -16236
rect 393780 -16434 393836 -16378
rect 393922 -16434 393978 -16378
rect 393780 -16576 393836 -16520
rect 393922 -16576 393978 -16520
rect 393780 -16718 393836 -16662
rect 393922 -16718 393978 -16662
rect 393780 -16860 393836 -16804
rect 393922 -16860 393978 -16804
rect 393780 -17002 393836 -16946
rect 393922 -17002 393978 -16946
rect 393780 -17144 393836 -17088
rect 393922 -17144 393978 -17088
rect 393780 -17286 393836 -17230
rect 393922 -17286 393978 -17230
rect 393780 -17428 393836 -17372
rect 393922 -17428 393978 -17372
rect 393780 -17570 393836 -17514
rect 393922 -17570 393978 -17514
rect 393780 -17712 393836 -17656
rect 393922 -17712 393978 -17656
rect 393780 -17854 393836 -17798
rect 393922 -17854 393978 -17798
rect 393780 -17996 393836 -17940
rect 393922 -17996 393978 -17940
rect 393780 -18138 393836 -18082
rect 393922 -18138 393978 -18082
rect 393780 -18280 393836 -18224
rect 393922 -18280 393978 -18224
rect 393780 -18422 393836 -18366
rect 393922 -18422 393978 -18366
rect 393780 -18564 393836 -18508
rect 393922 -18564 393978 -18508
rect 393780 -18706 393836 -18650
rect 393922 -18706 393978 -18650
rect 393780 -18848 393836 -18792
rect 393922 -18848 393978 -18792
rect 393780 -18990 393836 -18934
rect 393922 -18990 393978 -18934
rect 393780 -19132 393836 -19076
rect 393922 -19132 393978 -19076
rect 393780 -19274 393836 -19218
rect 393922 -19274 393978 -19218
rect 393780 -19416 393836 -19360
rect 393922 -19416 393978 -19360
rect 393780 -19558 393836 -19502
rect 393922 -19558 393978 -19502
rect 393780 -19700 393836 -19644
rect 393922 -19700 393978 -19644
rect 393780 -19842 393836 -19786
rect 393922 -19842 393978 -19786
rect 393780 -19984 393836 -19928
rect 393922 -19984 393978 -19928
rect 393780 -20126 393836 -20070
rect 393922 -20126 393978 -20070
rect 393780 -20268 393836 -20212
rect 393922 -20268 393978 -20212
rect 393780 -20410 393836 -20354
rect 393922 -20410 393978 -20354
rect 393780 -20552 393836 -20496
rect 393922 -20552 393978 -20496
rect 393780 -20694 393836 -20638
rect 393922 -20694 393978 -20638
rect 393780 -20836 393836 -20780
rect 393922 -20836 393978 -20780
rect 393780 -20978 393836 -20922
rect 393922 -20978 393978 -20922
rect 393780 -21120 393836 -21064
rect 393922 -21120 393978 -21064
rect 393780 -21262 393836 -21206
rect 393922 -21262 393978 -21206
rect 393780 -21404 393836 -21348
rect 393922 -21404 393978 -21348
rect 393780 -21546 393836 -21490
rect 393922 -21546 393978 -21490
rect 393780 -21688 393836 -21632
rect 393922 -21688 393978 -21632
rect 393780 -21830 393836 -21774
rect 393922 -21830 393978 -21774
rect 393780 -21972 393836 -21916
rect 393922 -21972 393978 -21916
rect 393780 -22114 393836 -22058
rect 393922 -22114 393978 -22058
rect 393780 -22256 393836 -22200
rect 393922 -22256 393978 -22200
rect 393780 -22398 393836 -22342
rect 393922 -22398 393978 -22342
rect 393780 -22540 393836 -22484
rect 393922 -22540 393978 -22484
rect 393780 -22682 393836 -22626
rect 393922 -22682 393978 -22626
rect 393780 -22824 393836 -22768
rect 393922 -22824 393978 -22768
rect 393780 -22966 393836 -22910
rect 393922 -22966 393978 -22910
rect 393780 -23108 393836 -23052
rect 393922 -23108 393978 -23052
rect 393780 -23250 393836 -23194
rect 393922 -23250 393978 -23194
rect 393780 -23392 393836 -23336
rect 393922 -23392 393978 -23336
rect 393780 -23534 393836 -23478
rect 393922 -23534 393978 -23478
rect 393780 -23676 393836 -23620
rect 393922 -23676 393978 -23620
rect 393780 -23818 393836 -23762
rect 393922 -23818 393978 -23762
rect 393780 -23960 393836 -23904
rect 393922 -23960 393978 -23904
rect 393780 -24102 393836 -24046
rect 393922 -24102 393978 -24046
rect 393780 -24244 393836 -24188
rect 393922 -24244 393978 -24188
rect 393780 -24386 393836 -24330
rect 393922 -24386 393978 -24330
rect 393780 -24528 393836 -24472
rect 393922 -24528 393978 -24472
rect 393780 -24670 393836 -24614
rect 393922 -24670 393978 -24614
rect 393780 -24812 393836 -24756
rect 393922 -24812 393978 -24756
rect 393780 -24954 393836 -24898
rect 393922 -24954 393978 -24898
rect 393780 -25096 393836 -25040
rect 393922 -25096 393978 -25040
rect 393780 -25238 393836 -25182
rect 393922 -25238 393978 -25182
rect 393780 -25380 393836 -25324
rect 393922 -25380 393978 -25324
rect 393780 -25522 393836 -25466
rect 393922 -25522 393978 -25466
rect 394177 -13736 394233 -13680
rect 394319 -13736 394375 -13680
rect 394177 -13878 394233 -13822
rect 394319 -13878 394375 -13822
rect 394177 -14020 394233 -13964
rect 394319 -14020 394375 -13964
rect 394177 -14162 394233 -14106
rect 394319 -14162 394375 -14106
rect 394177 -14304 394233 -14248
rect 394319 -14304 394375 -14248
rect 394177 -14446 394233 -14390
rect 394319 -14446 394375 -14390
rect 394177 -14588 394233 -14532
rect 394319 -14588 394375 -14532
rect 394177 -14730 394233 -14674
rect 394319 -14730 394375 -14674
rect 394177 -14872 394233 -14816
rect 394319 -14872 394375 -14816
rect 394177 -15014 394233 -14958
rect 394319 -15014 394375 -14958
rect 394177 -15156 394233 -15100
rect 394319 -15156 394375 -15100
rect 394177 -15298 394233 -15242
rect 394319 -15298 394375 -15242
rect 394177 -15440 394233 -15384
rect 394319 -15440 394375 -15384
rect 394177 -15582 394233 -15526
rect 394319 -15582 394375 -15526
rect 394177 -15724 394233 -15668
rect 394319 -15724 394375 -15668
rect 394177 -15866 394233 -15810
rect 394319 -15866 394375 -15810
rect 394177 -16008 394233 -15952
rect 394319 -16008 394375 -15952
rect 394177 -16150 394233 -16094
rect 394319 -16150 394375 -16094
rect 394177 -16292 394233 -16236
rect 394319 -16292 394375 -16236
rect 394177 -16434 394233 -16378
rect 394319 -16434 394375 -16378
rect 394177 -16576 394233 -16520
rect 394319 -16576 394375 -16520
rect 394177 -16718 394233 -16662
rect 394319 -16718 394375 -16662
rect 394177 -16860 394233 -16804
rect 394319 -16860 394375 -16804
rect 394177 -17002 394233 -16946
rect 394319 -17002 394375 -16946
rect 394177 -17144 394233 -17088
rect 394319 -17144 394375 -17088
rect 394177 -17286 394233 -17230
rect 394319 -17286 394375 -17230
rect 394177 -17428 394233 -17372
rect 394319 -17428 394375 -17372
rect 394177 -17570 394233 -17514
rect 394319 -17570 394375 -17514
rect 394177 -17712 394233 -17656
rect 394319 -17712 394375 -17656
rect 394177 -17854 394233 -17798
rect 394319 -17854 394375 -17798
rect 394177 -17996 394233 -17940
rect 394319 -17996 394375 -17940
rect 394177 -18138 394233 -18082
rect 394319 -18138 394375 -18082
rect 394177 -18280 394233 -18224
rect 394319 -18280 394375 -18224
rect 394177 -18422 394233 -18366
rect 394319 -18422 394375 -18366
rect 394177 -18564 394233 -18508
rect 394319 -18564 394375 -18508
rect 394177 -18706 394233 -18650
rect 394319 -18706 394375 -18650
rect 394177 -18848 394233 -18792
rect 394319 -18848 394375 -18792
rect 394177 -18990 394233 -18934
rect 394319 -18990 394375 -18934
rect 394177 -19132 394233 -19076
rect 394319 -19132 394375 -19076
rect 394177 -19274 394233 -19218
rect 394319 -19274 394375 -19218
rect 394177 -19416 394233 -19360
rect 394319 -19416 394375 -19360
rect 394177 -19558 394233 -19502
rect 394319 -19558 394375 -19502
rect 394177 -19700 394233 -19644
rect 394319 -19700 394375 -19644
rect 394177 -19842 394233 -19786
rect 394319 -19842 394375 -19786
rect 394177 -19984 394233 -19928
rect 394319 -19984 394375 -19928
rect 394177 -20126 394233 -20070
rect 394319 -20126 394375 -20070
rect 394177 -20268 394233 -20212
rect 394319 -20268 394375 -20212
rect 394177 -20410 394233 -20354
rect 394319 -20410 394375 -20354
rect 394177 -20552 394233 -20496
rect 394319 -20552 394375 -20496
rect 394177 -20694 394233 -20638
rect 394319 -20694 394375 -20638
rect 394177 -20836 394233 -20780
rect 394319 -20836 394375 -20780
rect 394177 -20978 394233 -20922
rect 394319 -20978 394375 -20922
rect 394177 -21120 394233 -21064
rect 394319 -21120 394375 -21064
rect 394177 -21262 394233 -21206
rect 394319 -21262 394375 -21206
rect 394177 -21404 394233 -21348
rect 394319 -21404 394375 -21348
rect 394177 -21546 394233 -21490
rect 394319 -21546 394375 -21490
rect 394177 -21688 394233 -21632
rect 394319 -21688 394375 -21632
rect 394177 -21830 394233 -21774
rect 394319 -21830 394375 -21774
rect 394177 -21972 394233 -21916
rect 394319 -21972 394375 -21916
rect 394177 -22114 394233 -22058
rect 394319 -22114 394375 -22058
rect 394177 -22256 394233 -22200
rect 394319 -22256 394375 -22200
rect 394177 -22398 394233 -22342
rect 394319 -22398 394375 -22342
rect 394177 -22540 394233 -22484
rect 394319 -22540 394375 -22484
rect 394177 -22682 394233 -22626
rect 394319 -22682 394375 -22626
rect 394177 -22824 394233 -22768
rect 394319 -22824 394375 -22768
rect 394177 -22966 394233 -22910
rect 394319 -22966 394375 -22910
rect 394177 -23108 394233 -23052
rect 394319 -23108 394375 -23052
rect 394177 -23250 394233 -23194
rect 394319 -23250 394375 -23194
rect 394177 -23392 394233 -23336
rect 394319 -23392 394375 -23336
rect 394177 -23534 394233 -23478
rect 394319 -23534 394375 -23478
rect 394177 -23676 394233 -23620
rect 394319 -23676 394375 -23620
rect 394177 -23818 394233 -23762
rect 394319 -23818 394375 -23762
rect 394177 -23960 394233 -23904
rect 394319 -23960 394375 -23904
rect 394177 -24102 394233 -24046
rect 394319 -24102 394375 -24046
rect 394177 -24244 394233 -24188
rect 394319 -24244 394375 -24188
rect 394177 -24386 394233 -24330
rect 394319 -24386 394375 -24330
rect 394177 -24528 394233 -24472
rect 394319 -24528 394375 -24472
rect 394177 -24670 394233 -24614
rect 394319 -24670 394375 -24614
rect 394177 -24812 394233 -24756
rect 394319 -24812 394375 -24756
rect 394177 -24954 394233 -24898
rect 394319 -24954 394375 -24898
rect 394177 -25096 394233 -25040
rect 394319 -25096 394375 -25040
rect 394177 -25238 394233 -25182
rect 394319 -25238 394375 -25182
rect 394177 -25380 394233 -25324
rect 394319 -25380 394375 -25324
rect 394177 -25522 394233 -25466
rect 394319 -25522 394375 -25466
rect 394580 -13736 394636 -13680
rect 394722 -13736 394778 -13680
rect 394580 -13878 394636 -13822
rect 394722 -13878 394778 -13822
rect 394580 -14020 394636 -13964
rect 394722 -14020 394778 -13964
rect 394580 -14162 394636 -14106
rect 394722 -14162 394778 -14106
rect 394580 -14304 394636 -14248
rect 394722 -14304 394778 -14248
rect 394580 -14446 394636 -14390
rect 394722 -14446 394778 -14390
rect 394580 -14588 394636 -14532
rect 394722 -14588 394778 -14532
rect 394580 -14730 394636 -14674
rect 394722 -14730 394778 -14674
rect 394580 -14872 394636 -14816
rect 394722 -14872 394778 -14816
rect 394580 -15014 394636 -14958
rect 394722 -15014 394778 -14958
rect 394580 -15156 394636 -15100
rect 394722 -15156 394778 -15100
rect 394580 -15298 394636 -15242
rect 394722 -15298 394778 -15242
rect 394580 -15440 394636 -15384
rect 394722 -15440 394778 -15384
rect 394580 -15582 394636 -15526
rect 394722 -15582 394778 -15526
rect 394580 -15724 394636 -15668
rect 394722 -15724 394778 -15668
rect 394580 -15866 394636 -15810
rect 394722 -15866 394778 -15810
rect 394580 -16008 394636 -15952
rect 394722 -16008 394778 -15952
rect 394580 -16150 394636 -16094
rect 394722 -16150 394778 -16094
rect 394580 -16292 394636 -16236
rect 394722 -16292 394778 -16236
rect 394580 -16434 394636 -16378
rect 394722 -16434 394778 -16378
rect 394580 -16576 394636 -16520
rect 394722 -16576 394778 -16520
rect 394580 -16718 394636 -16662
rect 394722 -16718 394778 -16662
rect 394580 -16860 394636 -16804
rect 394722 -16860 394778 -16804
rect 394580 -17002 394636 -16946
rect 394722 -17002 394778 -16946
rect 394580 -17144 394636 -17088
rect 394722 -17144 394778 -17088
rect 394580 -17286 394636 -17230
rect 394722 -17286 394778 -17230
rect 394580 -17428 394636 -17372
rect 394722 -17428 394778 -17372
rect 394580 -17570 394636 -17514
rect 394722 -17570 394778 -17514
rect 394580 -17712 394636 -17656
rect 394722 -17712 394778 -17656
rect 394580 -17854 394636 -17798
rect 394722 -17854 394778 -17798
rect 394580 -17996 394636 -17940
rect 394722 -17996 394778 -17940
rect 394580 -18138 394636 -18082
rect 394722 -18138 394778 -18082
rect 394580 -18280 394636 -18224
rect 394722 -18280 394778 -18224
rect 394580 -18422 394636 -18366
rect 394722 -18422 394778 -18366
rect 394580 -18564 394636 -18508
rect 394722 -18564 394778 -18508
rect 394580 -18706 394636 -18650
rect 394722 -18706 394778 -18650
rect 394580 -18848 394636 -18792
rect 394722 -18848 394778 -18792
rect 394580 -18990 394636 -18934
rect 394722 -18990 394778 -18934
rect 394580 -19132 394636 -19076
rect 394722 -19132 394778 -19076
rect 394580 -19274 394636 -19218
rect 394722 -19274 394778 -19218
rect 394580 -19416 394636 -19360
rect 394722 -19416 394778 -19360
rect 394580 -19558 394636 -19502
rect 394722 -19558 394778 -19502
rect 394580 -19700 394636 -19644
rect 394722 -19700 394778 -19644
rect 394580 -19842 394636 -19786
rect 394722 -19842 394778 -19786
rect 394580 -19984 394636 -19928
rect 394722 -19984 394778 -19928
rect 394580 -20126 394636 -20070
rect 394722 -20126 394778 -20070
rect 394580 -20268 394636 -20212
rect 394722 -20268 394778 -20212
rect 394580 -20410 394636 -20354
rect 394722 -20410 394778 -20354
rect 394580 -20552 394636 -20496
rect 394722 -20552 394778 -20496
rect 394580 -20694 394636 -20638
rect 394722 -20694 394778 -20638
rect 394580 -20836 394636 -20780
rect 394722 -20836 394778 -20780
rect 394580 -20978 394636 -20922
rect 394722 -20978 394778 -20922
rect 394580 -21120 394636 -21064
rect 394722 -21120 394778 -21064
rect 394580 -21262 394636 -21206
rect 394722 -21262 394778 -21206
rect 394580 -21404 394636 -21348
rect 394722 -21404 394778 -21348
rect 394580 -21546 394636 -21490
rect 394722 -21546 394778 -21490
rect 394580 -21688 394636 -21632
rect 394722 -21688 394778 -21632
rect 394580 -21830 394636 -21774
rect 394722 -21830 394778 -21774
rect 394580 -21972 394636 -21916
rect 394722 -21972 394778 -21916
rect 394580 -22114 394636 -22058
rect 394722 -22114 394778 -22058
rect 394580 -22256 394636 -22200
rect 394722 -22256 394778 -22200
rect 394580 -22398 394636 -22342
rect 394722 -22398 394778 -22342
rect 394580 -22540 394636 -22484
rect 394722 -22540 394778 -22484
rect 394580 -22682 394636 -22626
rect 394722 -22682 394778 -22626
rect 394580 -22824 394636 -22768
rect 394722 -22824 394778 -22768
rect 394580 -22966 394636 -22910
rect 394722 -22966 394778 -22910
rect 394580 -23108 394636 -23052
rect 394722 -23108 394778 -23052
rect 394580 -23250 394636 -23194
rect 394722 -23250 394778 -23194
rect 394580 -23392 394636 -23336
rect 394722 -23392 394778 -23336
rect 394580 -23534 394636 -23478
rect 394722 -23534 394778 -23478
rect 394580 -23676 394636 -23620
rect 394722 -23676 394778 -23620
rect 394580 -23818 394636 -23762
rect 394722 -23818 394778 -23762
rect 394580 -23960 394636 -23904
rect 394722 -23960 394778 -23904
rect 394580 -24102 394636 -24046
rect 394722 -24102 394778 -24046
rect 394580 -24244 394636 -24188
rect 394722 -24244 394778 -24188
rect 394580 -24386 394636 -24330
rect 394722 -24386 394778 -24330
rect 394580 -24528 394636 -24472
rect 394722 -24528 394778 -24472
rect 394580 -24670 394636 -24614
rect 394722 -24670 394778 -24614
rect 394580 -24812 394636 -24756
rect 394722 -24812 394778 -24756
rect 394580 -24954 394636 -24898
rect 394722 -24954 394778 -24898
rect 394580 -25096 394636 -25040
rect 394722 -25096 394778 -25040
rect 394580 -25238 394636 -25182
rect 394722 -25238 394778 -25182
rect 394580 -25380 394636 -25324
rect 394722 -25380 394778 -25324
rect 394580 -25522 394636 -25466
rect 394722 -25522 394778 -25466
rect 394982 -13736 395038 -13680
rect 395124 -13736 395180 -13680
rect 394982 -13878 395038 -13822
rect 395124 -13878 395180 -13822
rect 394982 -14020 395038 -13964
rect 395124 -14020 395180 -13964
rect 394982 -14162 395038 -14106
rect 395124 -14162 395180 -14106
rect 394982 -14304 395038 -14248
rect 395124 -14304 395180 -14248
rect 394982 -14446 395038 -14390
rect 395124 -14446 395180 -14390
rect 394982 -14588 395038 -14532
rect 395124 -14588 395180 -14532
rect 394982 -14730 395038 -14674
rect 395124 -14730 395180 -14674
rect 394982 -14872 395038 -14816
rect 395124 -14872 395180 -14816
rect 394982 -15014 395038 -14958
rect 395124 -15014 395180 -14958
rect 394982 -15156 395038 -15100
rect 395124 -15156 395180 -15100
rect 394982 -15298 395038 -15242
rect 395124 -15298 395180 -15242
rect 394982 -15440 395038 -15384
rect 395124 -15440 395180 -15384
rect 394982 -15582 395038 -15526
rect 395124 -15582 395180 -15526
rect 394982 -15724 395038 -15668
rect 395124 -15724 395180 -15668
rect 394982 -15866 395038 -15810
rect 395124 -15866 395180 -15810
rect 394982 -16008 395038 -15952
rect 395124 -16008 395180 -15952
rect 394982 -16150 395038 -16094
rect 395124 -16150 395180 -16094
rect 394982 -16292 395038 -16236
rect 395124 -16292 395180 -16236
rect 394982 -16434 395038 -16378
rect 395124 -16434 395180 -16378
rect 394982 -16576 395038 -16520
rect 395124 -16576 395180 -16520
rect 394982 -16718 395038 -16662
rect 395124 -16718 395180 -16662
rect 394982 -16860 395038 -16804
rect 395124 -16860 395180 -16804
rect 394982 -17002 395038 -16946
rect 395124 -17002 395180 -16946
rect 394982 -17144 395038 -17088
rect 395124 -17144 395180 -17088
rect 394982 -17286 395038 -17230
rect 395124 -17286 395180 -17230
rect 394982 -17428 395038 -17372
rect 395124 -17428 395180 -17372
rect 394982 -17570 395038 -17514
rect 395124 -17570 395180 -17514
rect 394982 -17712 395038 -17656
rect 395124 -17712 395180 -17656
rect 394982 -17854 395038 -17798
rect 395124 -17854 395180 -17798
rect 394982 -17996 395038 -17940
rect 395124 -17996 395180 -17940
rect 394982 -18138 395038 -18082
rect 395124 -18138 395180 -18082
rect 394982 -18280 395038 -18224
rect 395124 -18280 395180 -18224
rect 394982 -18422 395038 -18366
rect 395124 -18422 395180 -18366
rect 394982 -18564 395038 -18508
rect 395124 -18564 395180 -18508
rect 394982 -18706 395038 -18650
rect 395124 -18706 395180 -18650
rect 394982 -18848 395038 -18792
rect 395124 -18848 395180 -18792
rect 394982 -18990 395038 -18934
rect 395124 -18990 395180 -18934
rect 394982 -19132 395038 -19076
rect 395124 -19132 395180 -19076
rect 394982 -19274 395038 -19218
rect 395124 -19274 395180 -19218
rect 394982 -19416 395038 -19360
rect 395124 -19416 395180 -19360
rect 394982 -19558 395038 -19502
rect 395124 -19558 395180 -19502
rect 394982 -19700 395038 -19644
rect 395124 -19700 395180 -19644
rect 394982 -19842 395038 -19786
rect 395124 -19842 395180 -19786
rect 394982 -19984 395038 -19928
rect 395124 -19984 395180 -19928
rect 394982 -20126 395038 -20070
rect 395124 -20126 395180 -20070
rect 394982 -20268 395038 -20212
rect 395124 -20268 395180 -20212
rect 394982 -20410 395038 -20354
rect 395124 -20410 395180 -20354
rect 394982 -20552 395038 -20496
rect 395124 -20552 395180 -20496
rect 394982 -20694 395038 -20638
rect 395124 -20694 395180 -20638
rect 394982 -20836 395038 -20780
rect 395124 -20836 395180 -20780
rect 394982 -20978 395038 -20922
rect 395124 -20978 395180 -20922
rect 394982 -21120 395038 -21064
rect 395124 -21120 395180 -21064
rect 394982 -21262 395038 -21206
rect 395124 -21262 395180 -21206
rect 394982 -21404 395038 -21348
rect 395124 -21404 395180 -21348
rect 394982 -21546 395038 -21490
rect 395124 -21546 395180 -21490
rect 394982 -21688 395038 -21632
rect 395124 -21688 395180 -21632
rect 394982 -21830 395038 -21774
rect 395124 -21830 395180 -21774
rect 394982 -21972 395038 -21916
rect 395124 -21972 395180 -21916
rect 394982 -22114 395038 -22058
rect 395124 -22114 395180 -22058
rect 394982 -22256 395038 -22200
rect 395124 -22256 395180 -22200
rect 394982 -22398 395038 -22342
rect 395124 -22398 395180 -22342
rect 394982 -22540 395038 -22484
rect 395124 -22540 395180 -22484
rect 394982 -22682 395038 -22626
rect 395124 -22682 395180 -22626
rect 394982 -22824 395038 -22768
rect 395124 -22824 395180 -22768
rect 394982 -22966 395038 -22910
rect 395124 -22966 395180 -22910
rect 394982 -23108 395038 -23052
rect 395124 -23108 395180 -23052
rect 394982 -23250 395038 -23194
rect 395124 -23250 395180 -23194
rect 394982 -23392 395038 -23336
rect 395124 -23392 395180 -23336
rect 394982 -23534 395038 -23478
rect 395124 -23534 395180 -23478
rect 394982 -23676 395038 -23620
rect 395124 -23676 395180 -23620
rect 394982 -23818 395038 -23762
rect 395124 -23818 395180 -23762
rect 394982 -23960 395038 -23904
rect 395124 -23960 395180 -23904
rect 394982 -24102 395038 -24046
rect 395124 -24102 395180 -24046
rect 394982 -24244 395038 -24188
rect 395124 -24244 395180 -24188
rect 394982 -24386 395038 -24330
rect 395124 -24386 395180 -24330
rect 394982 -24528 395038 -24472
rect 395124 -24528 395180 -24472
rect 394982 -24670 395038 -24614
rect 395124 -24670 395180 -24614
rect 394982 -24812 395038 -24756
rect 395124 -24812 395180 -24756
rect 394982 -24954 395038 -24898
rect 395124 -24954 395180 -24898
rect 394982 -25096 395038 -25040
rect 395124 -25096 395180 -25040
rect 394982 -25238 395038 -25182
rect 395124 -25238 395180 -25182
rect 394982 -25380 395038 -25324
rect 395124 -25380 395180 -25324
rect 394982 -25522 395038 -25466
rect 395124 -25522 395180 -25466
rect 395385 -13736 395441 -13680
rect 395527 -13736 395583 -13680
rect 395385 -13878 395441 -13822
rect 395527 -13878 395583 -13822
rect 395385 -14020 395441 -13964
rect 395527 -14020 395583 -13964
rect 395385 -14162 395441 -14106
rect 395527 -14162 395583 -14106
rect 395385 -14304 395441 -14248
rect 395527 -14304 395583 -14248
rect 395385 -14446 395441 -14390
rect 395527 -14446 395583 -14390
rect 395385 -14588 395441 -14532
rect 395527 -14588 395583 -14532
rect 395385 -14730 395441 -14674
rect 395527 -14730 395583 -14674
rect 395385 -14872 395441 -14816
rect 395527 -14872 395583 -14816
rect 395385 -15014 395441 -14958
rect 395527 -15014 395583 -14958
rect 395385 -15156 395441 -15100
rect 395527 -15156 395583 -15100
rect 395385 -15298 395441 -15242
rect 395527 -15298 395583 -15242
rect 395385 -15440 395441 -15384
rect 395527 -15440 395583 -15384
rect 395385 -15582 395441 -15526
rect 395527 -15582 395583 -15526
rect 395385 -15724 395441 -15668
rect 395527 -15724 395583 -15668
rect 395385 -15866 395441 -15810
rect 395527 -15866 395583 -15810
rect 395385 -16008 395441 -15952
rect 395527 -16008 395583 -15952
rect 395385 -16150 395441 -16094
rect 395527 -16150 395583 -16094
rect 395385 -16292 395441 -16236
rect 395527 -16292 395583 -16236
rect 395385 -16434 395441 -16378
rect 395527 -16434 395583 -16378
rect 395385 -16576 395441 -16520
rect 395527 -16576 395583 -16520
rect 395385 -16718 395441 -16662
rect 395527 -16718 395583 -16662
rect 395385 -16860 395441 -16804
rect 395527 -16860 395583 -16804
rect 395385 -17002 395441 -16946
rect 395527 -17002 395583 -16946
rect 395385 -17144 395441 -17088
rect 395527 -17144 395583 -17088
rect 395385 -17286 395441 -17230
rect 395527 -17286 395583 -17230
rect 395385 -17428 395441 -17372
rect 395527 -17428 395583 -17372
rect 395385 -17570 395441 -17514
rect 395527 -17570 395583 -17514
rect 395385 -17712 395441 -17656
rect 395527 -17712 395583 -17656
rect 395385 -17854 395441 -17798
rect 395527 -17854 395583 -17798
rect 395385 -17996 395441 -17940
rect 395527 -17996 395583 -17940
rect 395385 -18138 395441 -18082
rect 395527 -18138 395583 -18082
rect 395385 -18280 395441 -18224
rect 395527 -18280 395583 -18224
rect 395385 -18422 395441 -18366
rect 395527 -18422 395583 -18366
rect 395385 -18564 395441 -18508
rect 395527 -18564 395583 -18508
rect 395385 -18706 395441 -18650
rect 395527 -18706 395583 -18650
rect 395385 -18848 395441 -18792
rect 395527 -18848 395583 -18792
rect 395385 -18990 395441 -18934
rect 395527 -18990 395583 -18934
rect 395385 -19132 395441 -19076
rect 395527 -19132 395583 -19076
rect 395385 -19274 395441 -19218
rect 395527 -19274 395583 -19218
rect 395385 -19416 395441 -19360
rect 395527 -19416 395583 -19360
rect 395385 -19558 395441 -19502
rect 395527 -19558 395583 -19502
rect 395385 -19700 395441 -19644
rect 395527 -19700 395583 -19644
rect 395385 -19842 395441 -19786
rect 395527 -19842 395583 -19786
rect 395385 -19984 395441 -19928
rect 395527 -19984 395583 -19928
rect 395385 -20126 395441 -20070
rect 395527 -20126 395583 -20070
rect 395385 -20268 395441 -20212
rect 395527 -20268 395583 -20212
rect 395385 -20410 395441 -20354
rect 395527 -20410 395583 -20354
rect 395385 -20552 395441 -20496
rect 395527 -20552 395583 -20496
rect 395385 -20694 395441 -20638
rect 395527 -20694 395583 -20638
rect 395385 -20836 395441 -20780
rect 395527 -20836 395583 -20780
rect 395385 -20978 395441 -20922
rect 395527 -20978 395583 -20922
rect 395385 -21120 395441 -21064
rect 395527 -21120 395583 -21064
rect 395385 -21262 395441 -21206
rect 395527 -21262 395583 -21206
rect 395385 -21404 395441 -21348
rect 395527 -21404 395583 -21348
rect 395385 -21546 395441 -21490
rect 395527 -21546 395583 -21490
rect 395385 -21688 395441 -21632
rect 395527 -21688 395583 -21632
rect 395385 -21830 395441 -21774
rect 395527 -21830 395583 -21774
rect 395385 -21972 395441 -21916
rect 395527 -21972 395583 -21916
rect 395385 -22114 395441 -22058
rect 395527 -22114 395583 -22058
rect 395385 -22256 395441 -22200
rect 395527 -22256 395583 -22200
rect 395385 -22398 395441 -22342
rect 395527 -22398 395583 -22342
rect 395385 -22540 395441 -22484
rect 395527 -22540 395583 -22484
rect 395385 -22682 395441 -22626
rect 395527 -22682 395583 -22626
rect 395385 -22824 395441 -22768
rect 395527 -22824 395583 -22768
rect 395385 -22966 395441 -22910
rect 395527 -22966 395583 -22910
rect 395385 -23108 395441 -23052
rect 395527 -23108 395583 -23052
rect 395385 -23250 395441 -23194
rect 395527 -23250 395583 -23194
rect 395385 -23392 395441 -23336
rect 395527 -23392 395583 -23336
rect 395385 -23534 395441 -23478
rect 395527 -23534 395583 -23478
rect 395385 -23676 395441 -23620
rect 395527 -23676 395583 -23620
rect 395385 -23818 395441 -23762
rect 395527 -23818 395583 -23762
rect 395385 -23960 395441 -23904
rect 395527 -23960 395583 -23904
rect 395385 -24102 395441 -24046
rect 395527 -24102 395583 -24046
rect 395385 -24244 395441 -24188
rect 395527 -24244 395583 -24188
rect 395385 -24386 395441 -24330
rect 395527 -24386 395583 -24330
rect 395385 -24528 395441 -24472
rect 395527 -24528 395583 -24472
rect 395385 -24670 395441 -24614
rect 395527 -24670 395583 -24614
rect 395385 -24812 395441 -24756
rect 395527 -24812 395583 -24756
rect 395385 -24954 395441 -24898
rect 395527 -24954 395583 -24898
rect 395385 -25096 395441 -25040
rect 395527 -25096 395583 -25040
rect 395385 -25238 395441 -25182
rect 395527 -25238 395583 -25182
rect 395385 -25380 395441 -25324
rect 395527 -25380 395583 -25324
rect 395385 -25522 395441 -25466
rect 395527 -25522 395583 -25466
rect 395779 -13736 395835 -13680
rect 395921 -13736 395977 -13680
rect 395779 -13878 395835 -13822
rect 395921 -13878 395977 -13822
rect 395779 -14020 395835 -13964
rect 395921 -14020 395977 -13964
rect 395779 -14162 395835 -14106
rect 395921 -14162 395977 -14106
rect 395779 -14304 395835 -14248
rect 395921 -14304 395977 -14248
rect 395779 -14446 395835 -14390
rect 395921 -14446 395977 -14390
rect 395779 -14588 395835 -14532
rect 395921 -14588 395977 -14532
rect 395779 -14730 395835 -14674
rect 395921 -14730 395977 -14674
rect 395779 -14872 395835 -14816
rect 395921 -14872 395977 -14816
rect 395779 -15014 395835 -14958
rect 395921 -15014 395977 -14958
rect 395779 -15156 395835 -15100
rect 395921 -15156 395977 -15100
rect 395779 -15298 395835 -15242
rect 395921 -15298 395977 -15242
rect 395779 -15440 395835 -15384
rect 395921 -15440 395977 -15384
rect 395779 -15582 395835 -15526
rect 395921 -15582 395977 -15526
rect 395779 -15724 395835 -15668
rect 395921 -15724 395977 -15668
rect 395779 -15866 395835 -15810
rect 395921 -15866 395977 -15810
rect 395779 -16008 395835 -15952
rect 395921 -16008 395977 -15952
rect 395779 -16150 395835 -16094
rect 395921 -16150 395977 -16094
rect 395779 -16292 395835 -16236
rect 395921 -16292 395977 -16236
rect 395779 -16434 395835 -16378
rect 395921 -16434 395977 -16378
rect 395779 -16576 395835 -16520
rect 395921 -16576 395977 -16520
rect 395779 -16718 395835 -16662
rect 395921 -16718 395977 -16662
rect 395779 -16860 395835 -16804
rect 395921 -16860 395977 -16804
rect 395779 -17002 395835 -16946
rect 395921 -17002 395977 -16946
rect 395779 -17144 395835 -17088
rect 395921 -17144 395977 -17088
rect 395779 -17286 395835 -17230
rect 395921 -17286 395977 -17230
rect 395779 -17428 395835 -17372
rect 395921 -17428 395977 -17372
rect 395779 -17570 395835 -17514
rect 395921 -17570 395977 -17514
rect 395779 -17712 395835 -17656
rect 395921 -17712 395977 -17656
rect 395779 -17854 395835 -17798
rect 395921 -17854 395977 -17798
rect 395779 -17996 395835 -17940
rect 395921 -17996 395977 -17940
rect 395779 -18138 395835 -18082
rect 395921 -18138 395977 -18082
rect 395779 -18280 395835 -18224
rect 395921 -18280 395977 -18224
rect 395779 -18422 395835 -18366
rect 395921 -18422 395977 -18366
rect 395779 -18564 395835 -18508
rect 395921 -18564 395977 -18508
rect 395779 -18706 395835 -18650
rect 395921 -18706 395977 -18650
rect 395779 -18848 395835 -18792
rect 395921 -18848 395977 -18792
rect 395779 -18990 395835 -18934
rect 395921 -18990 395977 -18934
rect 395779 -19132 395835 -19076
rect 395921 -19132 395977 -19076
rect 395779 -19274 395835 -19218
rect 395921 -19274 395977 -19218
rect 395779 -19416 395835 -19360
rect 395921 -19416 395977 -19360
rect 395779 -19558 395835 -19502
rect 395921 -19558 395977 -19502
rect 395779 -19700 395835 -19644
rect 395921 -19700 395977 -19644
rect 395779 -19842 395835 -19786
rect 395921 -19842 395977 -19786
rect 395779 -19984 395835 -19928
rect 395921 -19984 395977 -19928
rect 395779 -20126 395835 -20070
rect 395921 -20126 395977 -20070
rect 395779 -20268 395835 -20212
rect 395921 -20268 395977 -20212
rect 395779 -20410 395835 -20354
rect 395921 -20410 395977 -20354
rect 395779 -20552 395835 -20496
rect 395921 -20552 395977 -20496
rect 395779 -20694 395835 -20638
rect 395921 -20694 395977 -20638
rect 395779 -20836 395835 -20780
rect 395921 -20836 395977 -20780
rect 395779 -20978 395835 -20922
rect 395921 -20978 395977 -20922
rect 395779 -21120 395835 -21064
rect 395921 -21120 395977 -21064
rect 395779 -21262 395835 -21206
rect 395921 -21262 395977 -21206
rect 395779 -21404 395835 -21348
rect 395921 -21404 395977 -21348
rect 395779 -21546 395835 -21490
rect 395921 -21546 395977 -21490
rect 395779 -21688 395835 -21632
rect 395921 -21688 395977 -21632
rect 395779 -21830 395835 -21774
rect 395921 -21830 395977 -21774
rect 395779 -21972 395835 -21916
rect 395921 -21972 395977 -21916
rect 395779 -22114 395835 -22058
rect 395921 -22114 395977 -22058
rect 395779 -22256 395835 -22200
rect 395921 -22256 395977 -22200
rect 395779 -22398 395835 -22342
rect 395921 -22398 395977 -22342
rect 395779 -22540 395835 -22484
rect 395921 -22540 395977 -22484
rect 395779 -22682 395835 -22626
rect 395921 -22682 395977 -22626
rect 395779 -22824 395835 -22768
rect 395921 -22824 395977 -22768
rect 395779 -22966 395835 -22910
rect 395921 -22966 395977 -22910
rect 395779 -23108 395835 -23052
rect 395921 -23108 395977 -23052
rect 395779 -23250 395835 -23194
rect 395921 -23250 395977 -23194
rect 395779 -23392 395835 -23336
rect 395921 -23392 395977 -23336
rect 395779 -23534 395835 -23478
rect 395921 -23534 395977 -23478
rect 395779 -23676 395835 -23620
rect 395921 -23676 395977 -23620
rect 395779 -23818 395835 -23762
rect 395921 -23818 395977 -23762
rect 395779 -23960 395835 -23904
rect 395921 -23960 395977 -23904
rect 395779 -24102 395835 -24046
rect 395921 -24102 395977 -24046
rect 395779 -24244 395835 -24188
rect 395921 -24244 395977 -24188
rect 395779 -24386 395835 -24330
rect 395921 -24386 395977 -24330
rect 395779 -24528 395835 -24472
rect 395921 -24528 395977 -24472
rect 395779 -24670 395835 -24614
rect 395921 -24670 395977 -24614
rect 395779 -24812 395835 -24756
rect 395921 -24812 395977 -24756
rect 395779 -24954 395835 -24898
rect 395921 -24954 395977 -24898
rect 395779 -25096 395835 -25040
rect 395921 -25096 395977 -25040
rect 395779 -25238 395835 -25182
rect 395921 -25238 395977 -25182
rect 395779 -25380 395835 -25324
rect 395921 -25380 395977 -25324
rect 395779 -25522 395835 -25466
rect 395921 -25522 395977 -25466
rect 396180 -13736 396236 -13680
rect 396322 -13736 396378 -13680
rect 396180 -13878 396236 -13822
rect 396322 -13878 396378 -13822
rect 396180 -14020 396236 -13964
rect 396322 -14020 396378 -13964
rect 396180 -14162 396236 -14106
rect 396322 -14162 396378 -14106
rect 396180 -14304 396236 -14248
rect 396322 -14304 396378 -14248
rect 396180 -14446 396236 -14390
rect 396322 -14446 396378 -14390
rect 396180 -14588 396236 -14532
rect 396322 -14588 396378 -14532
rect 396180 -14730 396236 -14674
rect 396322 -14730 396378 -14674
rect 396180 -14872 396236 -14816
rect 396322 -14872 396378 -14816
rect 396180 -15014 396236 -14958
rect 396322 -15014 396378 -14958
rect 396180 -15156 396236 -15100
rect 396322 -15156 396378 -15100
rect 396180 -15298 396236 -15242
rect 396322 -15298 396378 -15242
rect 396180 -15440 396236 -15384
rect 396322 -15440 396378 -15384
rect 396180 -15582 396236 -15526
rect 396322 -15582 396378 -15526
rect 396180 -15724 396236 -15668
rect 396322 -15724 396378 -15668
rect 396180 -15866 396236 -15810
rect 396322 -15866 396378 -15810
rect 396180 -16008 396236 -15952
rect 396322 -16008 396378 -15952
rect 396180 -16150 396236 -16094
rect 396322 -16150 396378 -16094
rect 396180 -16292 396236 -16236
rect 396322 -16292 396378 -16236
rect 396180 -16434 396236 -16378
rect 396322 -16434 396378 -16378
rect 396180 -16576 396236 -16520
rect 396322 -16576 396378 -16520
rect 396180 -16718 396236 -16662
rect 396322 -16718 396378 -16662
rect 396180 -16860 396236 -16804
rect 396322 -16860 396378 -16804
rect 396180 -17002 396236 -16946
rect 396322 -17002 396378 -16946
rect 396180 -17144 396236 -17088
rect 396322 -17144 396378 -17088
rect 396180 -17286 396236 -17230
rect 396322 -17286 396378 -17230
rect 396180 -17428 396236 -17372
rect 396322 -17428 396378 -17372
rect 396180 -17570 396236 -17514
rect 396322 -17570 396378 -17514
rect 396180 -17712 396236 -17656
rect 396322 -17712 396378 -17656
rect 396180 -17854 396236 -17798
rect 396322 -17854 396378 -17798
rect 396180 -17996 396236 -17940
rect 396322 -17996 396378 -17940
rect 396180 -18138 396236 -18082
rect 396322 -18138 396378 -18082
rect 396180 -18280 396236 -18224
rect 396322 -18280 396378 -18224
rect 396180 -18422 396236 -18366
rect 396322 -18422 396378 -18366
rect 396180 -18564 396236 -18508
rect 396322 -18564 396378 -18508
rect 396180 -18706 396236 -18650
rect 396322 -18706 396378 -18650
rect 396180 -18848 396236 -18792
rect 396322 -18848 396378 -18792
rect 396180 -18990 396236 -18934
rect 396322 -18990 396378 -18934
rect 396180 -19132 396236 -19076
rect 396322 -19132 396378 -19076
rect 396180 -19274 396236 -19218
rect 396322 -19274 396378 -19218
rect 396180 -19416 396236 -19360
rect 396322 -19416 396378 -19360
rect 396180 -19558 396236 -19502
rect 396322 -19558 396378 -19502
rect 396180 -19700 396236 -19644
rect 396322 -19700 396378 -19644
rect 396180 -19842 396236 -19786
rect 396322 -19842 396378 -19786
rect 396180 -19984 396236 -19928
rect 396322 -19984 396378 -19928
rect 396180 -20126 396236 -20070
rect 396322 -20126 396378 -20070
rect 396180 -20268 396236 -20212
rect 396322 -20268 396378 -20212
rect 396180 -20410 396236 -20354
rect 396322 -20410 396378 -20354
rect 396180 -20552 396236 -20496
rect 396322 -20552 396378 -20496
rect 396180 -20694 396236 -20638
rect 396322 -20694 396378 -20638
rect 396180 -20836 396236 -20780
rect 396322 -20836 396378 -20780
rect 396180 -20978 396236 -20922
rect 396322 -20978 396378 -20922
rect 396180 -21120 396236 -21064
rect 396322 -21120 396378 -21064
rect 396180 -21262 396236 -21206
rect 396322 -21262 396378 -21206
rect 396180 -21404 396236 -21348
rect 396322 -21404 396378 -21348
rect 396180 -21546 396236 -21490
rect 396322 -21546 396378 -21490
rect 396180 -21688 396236 -21632
rect 396322 -21688 396378 -21632
rect 396180 -21830 396236 -21774
rect 396322 -21830 396378 -21774
rect 396180 -21972 396236 -21916
rect 396322 -21972 396378 -21916
rect 396180 -22114 396236 -22058
rect 396322 -22114 396378 -22058
rect 396180 -22256 396236 -22200
rect 396322 -22256 396378 -22200
rect 396180 -22398 396236 -22342
rect 396322 -22398 396378 -22342
rect 396180 -22540 396236 -22484
rect 396322 -22540 396378 -22484
rect 396180 -22682 396236 -22626
rect 396322 -22682 396378 -22626
rect 396180 -22824 396236 -22768
rect 396322 -22824 396378 -22768
rect 396180 -22966 396236 -22910
rect 396322 -22966 396378 -22910
rect 396180 -23108 396236 -23052
rect 396322 -23108 396378 -23052
rect 396180 -23250 396236 -23194
rect 396322 -23250 396378 -23194
rect 396180 -23392 396236 -23336
rect 396322 -23392 396378 -23336
rect 396180 -23534 396236 -23478
rect 396322 -23534 396378 -23478
rect 396180 -23676 396236 -23620
rect 396322 -23676 396378 -23620
rect 396180 -23818 396236 -23762
rect 396322 -23818 396378 -23762
rect 396180 -23960 396236 -23904
rect 396322 -23960 396378 -23904
rect 396180 -24102 396236 -24046
rect 396322 -24102 396378 -24046
rect 396180 -24244 396236 -24188
rect 396322 -24244 396378 -24188
rect 396180 -24386 396236 -24330
rect 396322 -24386 396378 -24330
rect 396180 -24528 396236 -24472
rect 396322 -24528 396378 -24472
rect 396180 -24670 396236 -24614
rect 396322 -24670 396378 -24614
rect 396180 -24812 396236 -24756
rect 396322 -24812 396378 -24756
rect 396180 -24954 396236 -24898
rect 396322 -24954 396378 -24898
rect 396180 -25096 396236 -25040
rect 396322 -25096 396378 -25040
rect 396180 -25238 396236 -25182
rect 396322 -25238 396378 -25182
rect 396180 -25380 396236 -25324
rect 396322 -25380 396378 -25324
rect 396180 -25522 396236 -25466
rect 396322 -25522 396378 -25466
rect 396580 -13736 396636 -13680
rect 396722 -13736 396778 -13680
rect 396580 -13878 396636 -13822
rect 396722 -13878 396778 -13822
rect 396580 -14020 396636 -13964
rect 396722 -14020 396778 -13964
rect 396580 -14162 396636 -14106
rect 396722 -14162 396778 -14106
rect 396580 -14304 396636 -14248
rect 396722 -14304 396778 -14248
rect 396580 -14446 396636 -14390
rect 396722 -14446 396778 -14390
rect 396580 -14588 396636 -14532
rect 396722 -14588 396778 -14532
rect 396580 -14730 396636 -14674
rect 396722 -14730 396778 -14674
rect 396580 -14872 396636 -14816
rect 396722 -14872 396778 -14816
rect 396580 -15014 396636 -14958
rect 396722 -15014 396778 -14958
rect 396580 -15156 396636 -15100
rect 396722 -15156 396778 -15100
rect 396580 -15298 396636 -15242
rect 396722 -15298 396778 -15242
rect 396580 -15440 396636 -15384
rect 396722 -15440 396778 -15384
rect 396580 -15582 396636 -15526
rect 396722 -15582 396778 -15526
rect 396580 -15724 396636 -15668
rect 396722 -15724 396778 -15668
rect 396580 -15866 396636 -15810
rect 396722 -15866 396778 -15810
rect 396580 -16008 396636 -15952
rect 396722 -16008 396778 -15952
rect 396580 -16150 396636 -16094
rect 396722 -16150 396778 -16094
rect 396580 -16292 396636 -16236
rect 396722 -16292 396778 -16236
rect 396580 -16434 396636 -16378
rect 396722 -16434 396778 -16378
rect 396580 -16576 396636 -16520
rect 396722 -16576 396778 -16520
rect 396580 -16718 396636 -16662
rect 396722 -16718 396778 -16662
rect 396580 -16860 396636 -16804
rect 396722 -16860 396778 -16804
rect 396580 -17002 396636 -16946
rect 396722 -17002 396778 -16946
rect 396580 -17144 396636 -17088
rect 396722 -17144 396778 -17088
rect 396580 -17286 396636 -17230
rect 396722 -17286 396778 -17230
rect 396580 -17428 396636 -17372
rect 396722 -17428 396778 -17372
rect 396580 -17570 396636 -17514
rect 396722 -17570 396778 -17514
rect 396580 -17712 396636 -17656
rect 396722 -17712 396778 -17656
rect 396580 -17854 396636 -17798
rect 396722 -17854 396778 -17798
rect 396580 -17996 396636 -17940
rect 396722 -17996 396778 -17940
rect 396580 -18138 396636 -18082
rect 396722 -18138 396778 -18082
rect 396580 -18280 396636 -18224
rect 396722 -18280 396778 -18224
rect 396580 -18422 396636 -18366
rect 396722 -18422 396778 -18366
rect 396580 -18564 396636 -18508
rect 396722 -18564 396778 -18508
rect 396580 -18706 396636 -18650
rect 396722 -18706 396778 -18650
rect 396580 -18848 396636 -18792
rect 396722 -18848 396778 -18792
rect 396580 -18990 396636 -18934
rect 396722 -18990 396778 -18934
rect 396580 -19132 396636 -19076
rect 396722 -19132 396778 -19076
rect 396580 -19274 396636 -19218
rect 396722 -19274 396778 -19218
rect 396580 -19416 396636 -19360
rect 396722 -19416 396778 -19360
rect 396580 -19558 396636 -19502
rect 396722 -19558 396778 -19502
rect 396580 -19700 396636 -19644
rect 396722 -19700 396778 -19644
rect 396580 -19842 396636 -19786
rect 396722 -19842 396778 -19786
rect 396580 -19984 396636 -19928
rect 396722 -19984 396778 -19928
rect 396580 -20126 396636 -20070
rect 396722 -20126 396778 -20070
rect 396580 -20268 396636 -20212
rect 396722 -20268 396778 -20212
rect 396580 -20410 396636 -20354
rect 396722 -20410 396778 -20354
rect 396580 -20552 396636 -20496
rect 396722 -20552 396778 -20496
rect 396580 -20694 396636 -20638
rect 396722 -20694 396778 -20638
rect 396580 -20836 396636 -20780
rect 396722 -20836 396778 -20780
rect 396580 -20978 396636 -20922
rect 396722 -20978 396778 -20922
rect 396580 -21120 396636 -21064
rect 396722 -21120 396778 -21064
rect 396580 -21262 396636 -21206
rect 396722 -21262 396778 -21206
rect 396580 -21404 396636 -21348
rect 396722 -21404 396778 -21348
rect 396580 -21546 396636 -21490
rect 396722 -21546 396778 -21490
rect 396580 -21688 396636 -21632
rect 396722 -21688 396778 -21632
rect 396580 -21830 396636 -21774
rect 396722 -21830 396778 -21774
rect 396580 -21972 396636 -21916
rect 396722 -21972 396778 -21916
rect 396580 -22114 396636 -22058
rect 396722 -22114 396778 -22058
rect 396580 -22256 396636 -22200
rect 396722 -22256 396778 -22200
rect 396580 -22398 396636 -22342
rect 396722 -22398 396778 -22342
rect 396580 -22540 396636 -22484
rect 396722 -22540 396778 -22484
rect 396580 -22682 396636 -22626
rect 396722 -22682 396778 -22626
rect 396580 -22824 396636 -22768
rect 396722 -22824 396778 -22768
rect 396580 -22966 396636 -22910
rect 396722 -22966 396778 -22910
rect 396580 -23108 396636 -23052
rect 396722 -23108 396778 -23052
rect 396580 -23250 396636 -23194
rect 396722 -23250 396778 -23194
rect 396580 -23392 396636 -23336
rect 396722 -23392 396778 -23336
rect 396580 -23534 396636 -23478
rect 396722 -23534 396778 -23478
rect 396580 -23676 396636 -23620
rect 396722 -23676 396778 -23620
rect 396580 -23818 396636 -23762
rect 396722 -23818 396778 -23762
rect 396580 -23960 396636 -23904
rect 396722 -23960 396778 -23904
rect 396580 -24102 396636 -24046
rect 396722 -24102 396778 -24046
rect 396580 -24244 396636 -24188
rect 396722 -24244 396778 -24188
rect 396580 -24386 396636 -24330
rect 396722 -24386 396778 -24330
rect 396580 -24528 396636 -24472
rect 396722 -24528 396778 -24472
rect 396580 -24670 396636 -24614
rect 396722 -24670 396778 -24614
rect 396580 -24812 396636 -24756
rect 396722 -24812 396778 -24756
rect 396580 -24954 396636 -24898
rect 396722 -24954 396778 -24898
rect 396580 -25096 396636 -25040
rect 396722 -25096 396778 -25040
rect 396580 -25238 396636 -25182
rect 396722 -25238 396778 -25182
rect 396580 -25380 396636 -25324
rect 396722 -25380 396778 -25324
rect 396580 -25522 396636 -25466
rect 396722 -25522 396778 -25466
rect 396977 -13736 397033 -13680
rect 397119 -13736 397175 -13680
rect 396977 -13878 397033 -13822
rect 397119 -13878 397175 -13822
rect 396977 -14020 397033 -13964
rect 397119 -14020 397175 -13964
rect 396977 -14162 397033 -14106
rect 397119 -14162 397175 -14106
rect 396977 -14304 397033 -14248
rect 397119 -14304 397175 -14248
rect 396977 -14446 397033 -14390
rect 397119 -14446 397175 -14390
rect 396977 -14588 397033 -14532
rect 397119 -14588 397175 -14532
rect 396977 -14730 397033 -14674
rect 397119 -14730 397175 -14674
rect 396977 -14872 397033 -14816
rect 397119 -14872 397175 -14816
rect 396977 -15014 397033 -14958
rect 397119 -15014 397175 -14958
rect 396977 -15156 397033 -15100
rect 397119 -15156 397175 -15100
rect 396977 -15298 397033 -15242
rect 397119 -15298 397175 -15242
rect 396977 -15440 397033 -15384
rect 397119 -15440 397175 -15384
rect 396977 -15582 397033 -15526
rect 397119 -15582 397175 -15526
rect 396977 -15724 397033 -15668
rect 397119 -15724 397175 -15668
rect 396977 -15866 397033 -15810
rect 397119 -15866 397175 -15810
rect 396977 -16008 397033 -15952
rect 397119 -16008 397175 -15952
rect 396977 -16150 397033 -16094
rect 397119 -16150 397175 -16094
rect 396977 -16292 397033 -16236
rect 397119 -16292 397175 -16236
rect 396977 -16434 397033 -16378
rect 397119 -16434 397175 -16378
rect 396977 -16576 397033 -16520
rect 397119 -16576 397175 -16520
rect 396977 -16718 397033 -16662
rect 397119 -16718 397175 -16662
rect 396977 -16860 397033 -16804
rect 397119 -16860 397175 -16804
rect 396977 -17002 397033 -16946
rect 397119 -17002 397175 -16946
rect 396977 -17144 397033 -17088
rect 397119 -17144 397175 -17088
rect 396977 -17286 397033 -17230
rect 397119 -17286 397175 -17230
rect 396977 -17428 397033 -17372
rect 397119 -17428 397175 -17372
rect 396977 -17570 397033 -17514
rect 397119 -17570 397175 -17514
rect 396977 -17712 397033 -17656
rect 397119 -17712 397175 -17656
rect 396977 -17854 397033 -17798
rect 397119 -17854 397175 -17798
rect 396977 -17996 397033 -17940
rect 397119 -17996 397175 -17940
rect 396977 -18138 397033 -18082
rect 397119 -18138 397175 -18082
rect 396977 -18280 397033 -18224
rect 397119 -18280 397175 -18224
rect 396977 -18422 397033 -18366
rect 397119 -18422 397175 -18366
rect 396977 -18564 397033 -18508
rect 397119 -18564 397175 -18508
rect 396977 -18706 397033 -18650
rect 397119 -18706 397175 -18650
rect 396977 -18848 397033 -18792
rect 397119 -18848 397175 -18792
rect 396977 -18990 397033 -18934
rect 397119 -18990 397175 -18934
rect 396977 -19132 397033 -19076
rect 397119 -19132 397175 -19076
rect 396977 -19274 397033 -19218
rect 397119 -19274 397175 -19218
rect 396977 -19416 397033 -19360
rect 397119 -19416 397175 -19360
rect 396977 -19558 397033 -19502
rect 397119 -19558 397175 -19502
rect 396977 -19700 397033 -19644
rect 397119 -19700 397175 -19644
rect 396977 -19842 397033 -19786
rect 397119 -19842 397175 -19786
rect 396977 -19984 397033 -19928
rect 397119 -19984 397175 -19928
rect 396977 -20126 397033 -20070
rect 397119 -20126 397175 -20070
rect 396977 -20268 397033 -20212
rect 397119 -20268 397175 -20212
rect 396977 -20410 397033 -20354
rect 397119 -20410 397175 -20354
rect 396977 -20552 397033 -20496
rect 397119 -20552 397175 -20496
rect 396977 -20694 397033 -20638
rect 397119 -20694 397175 -20638
rect 396977 -20836 397033 -20780
rect 397119 -20836 397175 -20780
rect 396977 -20978 397033 -20922
rect 397119 -20978 397175 -20922
rect 396977 -21120 397033 -21064
rect 397119 -21120 397175 -21064
rect 396977 -21262 397033 -21206
rect 397119 -21262 397175 -21206
rect 396977 -21404 397033 -21348
rect 397119 -21404 397175 -21348
rect 396977 -21546 397033 -21490
rect 397119 -21546 397175 -21490
rect 396977 -21688 397033 -21632
rect 397119 -21688 397175 -21632
rect 396977 -21830 397033 -21774
rect 397119 -21830 397175 -21774
rect 396977 -21972 397033 -21916
rect 397119 -21972 397175 -21916
rect 396977 -22114 397033 -22058
rect 397119 -22114 397175 -22058
rect 396977 -22256 397033 -22200
rect 397119 -22256 397175 -22200
rect 396977 -22398 397033 -22342
rect 397119 -22398 397175 -22342
rect 396977 -22540 397033 -22484
rect 397119 -22540 397175 -22484
rect 396977 -22682 397033 -22626
rect 397119 -22682 397175 -22626
rect 396977 -22824 397033 -22768
rect 397119 -22824 397175 -22768
rect 396977 -22966 397033 -22910
rect 397119 -22966 397175 -22910
rect 396977 -23108 397033 -23052
rect 397119 -23108 397175 -23052
rect 396977 -23250 397033 -23194
rect 397119 -23250 397175 -23194
rect 396977 -23392 397033 -23336
rect 397119 -23392 397175 -23336
rect 396977 -23534 397033 -23478
rect 397119 -23534 397175 -23478
rect 396977 -23676 397033 -23620
rect 397119 -23676 397175 -23620
rect 396977 -23818 397033 -23762
rect 397119 -23818 397175 -23762
rect 396977 -23960 397033 -23904
rect 397119 -23960 397175 -23904
rect 396977 -24102 397033 -24046
rect 397119 -24102 397175 -24046
rect 396977 -24244 397033 -24188
rect 397119 -24244 397175 -24188
rect 396977 -24386 397033 -24330
rect 397119 -24386 397175 -24330
rect 396977 -24528 397033 -24472
rect 397119 -24528 397175 -24472
rect 396977 -24670 397033 -24614
rect 397119 -24670 397175 -24614
rect 396977 -24812 397033 -24756
rect 397119 -24812 397175 -24756
rect 396977 -24954 397033 -24898
rect 397119 -24954 397175 -24898
rect 396977 -25096 397033 -25040
rect 397119 -25096 397175 -25040
rect 396977 -25238 397033 -25182
rect 397119 -25238 397175 -25182
rect 396977 -25380 397033 -25324
rect 397119 -25380 397175 -25324
rect 396977 -25522 397033 -25466
rect 397119 -25522 397175 -25466
rect 397374 -13736 397430 -13680
rect 397516 -13736 397572 -13680
rect 397374 -13878 397430 -13822
rect 397516 -13878 397572 -13822
rect 397374 -14020 397430 -13964
rect 397516 -14020 397572 -13964
rect 397374 -14162 397430 -14106
rect 397516 -14162 397572 -14106
rect 397374 -14304 397430 -14248
rect 397516 -14304 397572 -14248
rect 397374 -14446 397430 -14390
rect 397516 -14446 397572 -14390
rect 397374 -14588 397430 -14532
rect 397516 -14588 397572 -14532
rect 397374 -14730 397430 -14674
rect 397516 -14730 397572 -14674
rect 397374 -14872 397430 -14816
rect 397516 -14872 397572 -14816
rect 397374 -15014 397430 -14958
rect 397516 -15014 397572 -14958
rect 397374 -15156 397430 -15100
rect 397516 -15156 397572 -15100
rect 397374 -15298 397430 -15242
rect 397516 -15298 397572 -15242
rect 397374 -15440 397430 -15384
rect 397516 -15440 397572 -15384
rect 397374 -15582 397430 -15526
rect 397516 -15582 397572 -15526
rect 397374 -15724 397430 -15668
rect 397516 -15724 397572 -15668
rect 397374 -15866 397430 -15810
rect 397516 -15866 397572 -15810
rect 397374 -16008 397430 -15952
rect 397516 -16008 397572 -15952
rect 397374 -16150 397430 -16094
rect 397516 -16150 397572 -16094
rect 397374 -16292 397430 -16236
rect 397516 -16292 397572 -16236
rect 397374 -16434 397430 -16378
rect 397516 -16434 397572 -16378
rect 397374 -16576 397430 -16520
rect 397516 -16576 397572 -16520
rect 397374 -16718 397430 -16662
rect 397516 -16718 397572 -16662
rect 397374 -16860 397430 -16804
rect 397516 -16860 397572 -16804
rect 397374 -17002 397430 -16946
rect 397516 -17002 397572 -16946
rect 397374 -17144 397430 -17088
rect 397516 -17144 397572 -17088
rect 397374 -17286 397430 -17230
rect 397516 -17286 397572 -17230
rect 397374 -17428 397430 -17372
rect 397516 -17428 397572 -17372
rect 397374 -17570 397430 -17514
rect 397516 -17570 397572 -17514
rect 397374 -17712 397430 -17656
rect 397516 -17712 397572 -17656
rect 397374 -17854 397430 -17798
rect 397516 -17854 397572 -17798
rect 397374 -17996 397430 -17940
rect 397516 -17996 397572 -17940
rect 397374 -18138 397430 -18082
rect 397516 -18138 397572 -18082
rect 397374 -18280 397430 -18224
rect 397516 -18280 397572 -18224
rect 397374 -18422 397430 -18366
rect 397516 -18422 397572 -18366
rect 397374 -18564 397430 -18508
rect 397516 -18564 397572 -18508
rect 397374 -18706 397430 -18650
rect 397516 -18706 397572 -18650
rect 397374 -18848 397430 -18792
rect 397516 -18848 397572 -18792
rect 397374 -18990 397430 -18934
rect 397516 -18990 397572 -18934
rect 397374 -19132 397430 -19076
rect 397516 -19132 397572 -19076
rect 397374 -19274 397430 -19218
rect 397516 -19274 397572 -19218
rect 397374 -19416 397430 -19360
rect 397516 -19416 397572 -19360
rect 397374 -19558 397430 -19502
rect 397516 -19558 397572 -19502
rect 397374 -19700 397430 -19644
rect 397516 -19700 397572 -19644
rect 397374 -19842 397430 -19786
rect 397516 -19842 397572 -19786
rect 397374 -19984 397430 -19928
rect 397516 -19984 397572 -19928
rect 397374 -20126 397430 -20070
rect 397516 -20126 397572 -20070
rect 397374 -20268 397430 -20212
rect 397516 -20268 397572 -20212
rect 397374 -20410 397430 -20354
rect 397516 -20410 397572 -20354
rect 397374 -20552 397430 -20496
rect 397516 -20552 397572 -20496
rect 397374 -20694 397430 -20638
rect 397516 -20694 397572 -20638
rect 397374 -20836 397430 -20780
rect 397516 -20836 397572 -20780
rect 397374 -20978 397430 -20922
rect 397516 -20978 397572 -20922
rect 397374 -21120 397430 -21064
rect 397516 -21120 397572 -21064
rect 397374 -21262 397430 -21206
rect 397516 -21262 397572 -21206
rect 397374 -21404 397430 -21348
rect 397516 -21404 397572 -21348
rect 397374 -21546 397430 -21490
rect 397516 -21546 397572 -21490
rect 397374 -21688 397430 -21632
rect 397516 -21688 397572 -21632
rect 397374 -21830 397430 -21774
rect 397516 -21830 397572 -21774
rect 397374 -21972 397430 -21916
rect 397516 -21972 397572 -21916
rect 397374 -22114 397430 -22058
rect 397516 -22114 397572 -22058
rect 397374 -22256 397430 -22200
rect 397516 -22256 397572 -22200
rect 397374 -22398 397430 -22342
rect 397516 -22398 397572 -22342
rect 397374 -22540 397430 -22484
rect 397516 -22540 397572 -22484
rect 397374 -22682 397430 -22626
rect 397516 -22682 397572 -22626
rect 397374 -22824 397430 -22768
rect 397516 -22824 397572 -22768
rect 397374 -22966 397430 -22910
rect 397516 -22966 397572 -22910
rect 397374 -23108 397430 -23052
rect 397516 -23108 397572 -23052
rect 397374 -23250 397430 -23194
rect 397516 -23250 397572 -23194
rect 397374 -23392 397430 -23336
rect 397516 -23392 397572 -23336
rect 397374 -23534 397430 -23478
rect 397516 -23534 397572 -23478
rect 397374 -23676 397430 -23620
rect 397516 -23676 397572 -23620
rect 397374 -23818 397430 -23762
rect 397516 -23818 397572 -23762
rect 397374 -23960 397430 -23904
rect 397516 -23960 397572 -23904
rect 397374 -24102 397430 -24046
rect 397516 -24102 397572 -24046
rect 397374 -24244 397430 -24188
rect 397516 -24244 397572 -24188
rect 397374 -24386 397430 -24330
rect 397516 -24386 397572 -24330
rect 397374 -24528 397430 -24472
rect 397516 -24528 397572 -24472
rect 397374 -24670 397430 -24614
rect 397516 -24670 397572 -24614
rect 397374 -24812 397430 -24756
rect 397516 -24812 397572 -24756
rect 397374 -24954 397430 -24898
rect 397516 -24954 397572 -24898
rect 397374 -25096 397430 -25040
rect 397516 -25096 397572 -25040
rect 397374 -25238 397430 -25182
rect 397516 -25238 397572 -25182
rect 397374 -25380 397430 -25324
rect 397516 -25380 397572 -25324
rect 397374 -25522 397430 -25466
rect 397516 -25522 397572 -25466
rect 397778 -13736 397834 -13680
rect 397920 -13736 397976 -13680
rect 397778 -13878 397834 -13822
rect 397920 -13878 397976 -13822
rect 397778 -14020 397834 -13964
rect 397920 -14020 397976 -13964
rect 397778 -14162 397834 -14106
rect 397920 -14162 397976 -14106
rect 397778 -14304 397834 -14248
rect 397920 -14304 397976 -14248
rect 397778 -14446 397834 -14390
rect 397920 -14446 397976 -14390
rect 397778 -14588 397834 -14532
rect 397920 -14588 397976 -14532
rect 397778 -14730 397834 -14674
rect 397920 -14730 397976 -14674
rect 397778 -14872 397834 -14816
rect 397920 -14872 397976 -14816
rect 397778 -15014 397834 -14958
rect 397920 -15014 397976 -14958
rect 397778 -15156 397834 -15100
rect 397920 -15156 397976 -15100
rect 397778 -15298 397834 -15242
rect 397920 -15298 397976 -15242
rect 397778 -15440 397834 -15384
rect 397920 -15440 397976 -15384
rect 397778 -15582 397834 -15526
rect 397920 -15582 397976 -15526
rect 397778 -15724 397834 -15668
rect 397920 -15724 397976 -15668
rect 397778 -15866 397834 -15810
rect 397920 -15866 397976 -15810
rect 397778 -16008 397834 -15952
rect 397920 -16008 397976 -15952
rect 397778 -16150 397834 -16094
rect 397920 -16150 397976 -16094
rect 397778 -16292 397834 -16236
rect 397920 -16292 397976 -16236
rect 397778 -16434 397834 -16378
rect 397920 -16434 397976 -16378
rect 397778 -16576 397834 -16520
rect 397920 -16576 397976 -16520
rect 397778 -16718 397834 -16662
rect 397920 -16718 397976 -16662
rect 397778 -16860 397834 -16804
rect 397920 -16860 397976 -16804
rect 397778 -17002 397834 -16946
rect 397920 -17002 397976 -16946
rect 397778 -17144 397834 -17088
rect 397920 -17144 397976 -17088
rect 397778 -17286 397834 -17230
rect 397920 -17286 397976 -17230
rect 397778 -17428 397834 -17372
rect 397920 -17428 397976 -17372
rect 397778 -17570 397834 -17514
rect 397920 -17570 397976 -17514
rect 397778 -17712 397834 -17656
rect 397920 -17712 397976 -17656
rect 397778 -17854 397834 -17798
rect 397920 -17854 397976 -17798
rect 397778 -17996 397834 -17940
rect 397920 -17996 397976 -17940
rect 397778 -18138 397834 -18082
rect 397920 -18138 397976 -18082
rect 397778 -18280 397834 -18224
rect 397920 -18280 397976 -18224
rect 397778 -18422 397834 -18366
rect 397920 -18422 397976 -18366
rect 397778 -18564 397834 -18508
rect 397920 -18564 397976 -18508
rect 397778 -18706 397834 -18650
rect 397920 -18706 397976 -18650
rect 397778 -18848 397834 -18792
rect 397920 -18848 397976 -18792
rect 397778 -18990 397834 -18934
rect 397920 -18990 397976 -18934
rect 397778 -19132 397834 -19076
rect 397920 -19132 397976 -19076
rect 397778 -19274 397834 -19218
rect 397920 -19274 397976 -19218
rect 397778 -19416 397834 -19360
rect 397920 -19416 397976 -19360
rect 397778 -19558 397834 -19502
rect 397920 -19558 397976 -19502
rect 397778 -19700 397834 -19644
rect 397920 -19700 397976 -19644
rect 397778 -19842 397834 -19786
rect 397920 -19842 397976 -19786
rect 397778 -19984 397834 -19928
rect 397920 -19984 397976 -19928
rect 397778 -20126 397834 -20070
rect 397920 -20126 397976 -20070
rect 397778 -20268 397834 -20212
rect 397920 -20268 397976 -20212
rect 397778 -20410 397834 -20354
rect 397920 -20410 397976 -20354
rect 397778 -20552 397834 -20496
rect 397920 -20552 397976 -20496
rect 397778 -20694 397834 -20638
rect 397920 -20694 397976 -20638
rect 397778 -20836 397834 -20780
rect 397920 -20836 397976 -20780
rect 397778 -20978 397834 -20922
rect 397920 -20978 397976 -20922
rect 397778 -21120 397834 -21064
rect 397920 -21120 397976 -21064
rect 397778 -21262 397834 -21206
rect 397920 -21262 397976 -21206
rect 397778 -21404 397834 -21348
rect 397920 -21404 397976 -21348
rect 397778 -21546 397834 -21490
rect 397920 -21546 397976 -21490
rect 397778 -21688 397834 -21632
rect 397920 -21688 397976 -21632
rect 397778 -21830 397834 -21774
rect 397920 -21830 397976 -21774
rect 397778 -21972 397834 -21916
rect 397920 -21972 397976 -21916
rect 397778 -22114 397834 -22058
rect 397920 -22114 397976 -22058
rect 397778 -22256 397834 -22200
rect 397920 -22256 397976 -22200
rect 397778 -22398 397834 -22342
rect 397920 -22398 397976 -22342
rect 397778 -22540 397834 -22484
rect 397920 -22540 397976 -22484
rect 397778 -22682 397834 -22626
rect 397920 -22682 397976 -22626
rect 397778 -22824 397834 -22768
rect 397920 -22824 397976 -22768
rect 397778 -22966 397834 -22910
rect 397920 -22966 397976 -22910
rect 397778 -23108 397834 -23052
rect 397920 -23108 397976 -23052
rect 397778 -23250 397834 -23194
rect 397920 -23250 397976 -23194
rect 397778 -23392 397834 -23336
rect 397920 -23392 397976 -23336
rect 397778 -23534 397834 -23478
rect 397920 -23534 397976 -23478
rect 397778 -23676 397834 -23620
rect 397920 -23676 397976 -23620
rect 397778 -23818 397834 -23762
rect 397920 -23818 397976 -23762
rect 397778 -23960 397834 -23904
rect 397920 -23960 397976 -23904
rect 397778 -24102 397834 -24046
rect 397920 -24102 397976 -24046
rect 397778 -24244 397834 -24188
rect 397920 -24244 397976 -24188
rect 397778 -24386 397834 -24330
rect 397920 -24386 397976 -24330
rect 397778 -24528 397834 -24472
rect 397920 -24528 397976 -24472
rect 397778 -24670 397834 -24614
rect 397920 -24670 397976 -24614
rect 397778 -24812 397834 -24756
rect 397920 -24812 397976 -24756
rect 397778 -24954 397834 -24898
rect 397920 -24954 397976 -24898
rect 397778 -25096 397834 -25040
rect 397920 -25096 397976 -25040
rect 397778 -25238 397834 -25182
rect 397920 -25238 397976 -25182
rect 397778 -25380 397834 -25324
rect 397920 -25380 397976 -25324
rect 397778 -25522 397834 -25466
rect 397920 -25522 397976 -25466
rect 398174 -13736 398230 -13680
rect 398316 -13736 398372 -13680
rect 398174 -13878 398230 -13822
rect 398316 -13878 398372 -13822
rect 398174 -14020 398230 -13964
rect 398316 -14020 398372 -13964
rect 398174 -14162 398230 -14106
rect 398316 -14162 398372 -14106
rect 398174 -14304 398230 -14248
rect 398316 -14304 398372 -14248
rect 398174 -14446 398230 -14390
rect 398316 -14446 398372 -14390
rect 398174 -14588 398230 -14532
rect 398316 -14588 398372 -14532
rect 398174 -14730 398230 -14674
rect 398316 -14730 398372 -14674
rect 398174 -14872 398230 -14816
rect 398316 -14872 398372 -14816
rect 398174 -15014 398230 -14958
rect 398316 -15014 398372 -14958
rect 398174 -15156 398230 -15100
rect 398316 -15156 398372 -15100
rect 398174 -15298 398230 -15242
rect 398316 -15298 398372 -15242
rect 398174 -15440 398230 -15384
rect 398316 -15440 398372 -15384
rect 398174 -15582 398230 -15526
rect 398316 -15582 398372 -15526
rect 398174 -15724 398230 -15668
rect 398316 -15724 398372 -15668
rect 398174 -15866 398230 -15810
rect 398316 -15866 398372 -15810
rect 398174 -16008 398230 -15952
rect 398316 -16008 398372 -15952
rect 398174 -16150 398230 -16094
rect 398316 -16150 398372 -16094
rect 398174 -16292 398230 -16236
rect 398316 -16292 398372 -16236
rect 398174 -16434 398230 -16378
rect 398316 -16434 398372 -16378
rect 398174 -16576 398230 -16520
rect 398316 -16576 398372 -16520
rect 398174 -16718 398230 -16662
rect 398316 -16718 398372 -16662
rect 398174 -16860 398230 -16804
rect 398316 -16860 398372 -16804
rect 398174 -17002 398230 -16946
rect 398316 -17002 398372 -16946
rect 398174 -17144 398230 -17088
rect 398316 -17144 398372 -17088
rect 398174 -17286 398230 -17230
rect 398316 -17286 398372 -17230
rect 398174 -17428 398230 -17372
rect 398316 -17428 398372 -17372
rect 398174 -17570 398230 -17514
rect 398316 -17570 398372 -17514
rect 398174 -17712 398230 -17656
rect 398316 -17712 398372 -17656
rect 398174 -17854 398230 -17798
rect 398316 -17854 398372 -17798
rect 398174 -17996 398230 -17940
rect 398316 -17996 398372 -17940
rect 398174 -18138 398230 -18082
rect 398316 -18138 398372 -18082
rect 398174 -18280 398230 -18224
rect 398316 -18280 398372 -18224
rect 398174 -18422 398230 -18366
rect 398316 -18422 398372 -18366
rect 398174 -18564 398230 -18508
rect 398316 -18564 398372 -18508
rect 398174 -18706 398230 -18650
rect 398316 -18706 398372 -18650
rect 398174 -18848 398230 -18792
rect 398316 -18848 398372 -18792
rect 398174 -18990 398230 -18934
rect 398316 -18990 398372 -18934
rect 398174 -19132 398230 -19076
rect 398316 -19132 398372 -19076
rect 398174 -19274 398230 -19218
rect 398316 -19274 398372 -19218
rect 398174 -19416 398230 -19360
rect 398316 -19416 398372 -19360
rect 398174 -19558 398230 -19502
rect 398316 -19558 398372 -19502
rect 398174 -19700 398230 -19644
rect 398316 -19700 398372 -19644
rect 398174 -19842 398230 -19786
rect 398316 -19842 398372 -19786
rect 398174 -19984 398230 -19928
rect 398316 -19984 398372 -19928
rect 398174 -20126 398230 -20070
rect 398316 -20126 398372 -20070
rect 398174 -20268 398230 -20212
rect 398316 -20268 398372 -20212
rect 398174 -20410 398230 -20354
rect 398316 -20410 398372 -20354
rect 398174 -20552 398230 -20496
rect 398316 -20552 398372 -20496
rect 398174 -20694 398230 -20638
rect 398316 -20694 398372 -20638
rect 398174 -20836 398230 -20780
rect 398316 -20836 398372 -20780
rect 398174 -20978 398230 -20922
rect 398316 -20978 398372 -20922
rect 398174 -21120 398230 -21064
rect 398316 -21120 398372 -21064
rect 398174 -21262 398230 -21206
rect 398316 -21262 398372 -21206
rect 398174 -21404 398230 -21348
rect 398316 -21404 398372 -21348
rect 398174 -21546 398230 -21490
rect 398316 -21546 398372 -21490
rect 398174 -21688 398230 -21632
rect 398316 -21688 398372 -21632
rect 398174 -21830 398230 -21774
rect 398316 -21830 398372 -21774
rect 398174 -21972 398230 -21916
rect 398316 -21972 398372 -21916
rect 398174 -22114 398230 -22058
rect 398316 -22114 398372 -22058
rect 398174 -22256 398230 -22200
rect 398316 -22256 398372 -22200
rect 398174 -22398 398230 -22342
rect 398316 -22398 398372 -22342
rect 398174 -22540 398230 -22484
rect 398316 -22540 398372 -22484
rect 398174 -22682 398230 -22626
rect 398316 -22682 398372 -22626
rect 398174 -22824 398230 -22768
rect 398316 -22824 398372 -22768
rect 398174 -22966 398230 -22910
rect 398316 -22966 398372 -22910
rect 398174 -23108 398230 -23052
rect 398316 -23108 398372 -23052
rect 398174 -23250 398230 -23194
rect 398316 -23250 398372 -23194
rect 398174 -23392 398230 -23336
rect 398316 -23392 398372 -23336
rect 398174 -23534 398230 -23478
rect 398316 -23534 398372 -23478
rect 398174 -23676 398230 -23620
rect 398316 -23676 398372 -23620
rect 398174 -23818 398230 -23762
rect 398316 -23818 398372 -23762
rect 398174 -23960 398230 -23904
rect 398316 -23960 398372 -23904
rect 398174 -24102 398230 -24046
rect 398316 -24102 398372 -24046
rect 398174 -24244 398230 -24188
rect 398316 -24244 398372 -24188
rect 398174 -24386 398230 -24330
rect 398316 -24386 398372 -24330
rect 398174 -24528 398230 -24472
rect 398316 -24528 398372 -24472
rect 398174 -24670 398230 -24614
rect 398316 -24670 398372 -24614
rect 398174 -24812 398230 -24756
rect 398316 -24812 398372 -24756
rect 398174 -24954 398230 -24898
rect 398316 -24954 398372 -24898
rect 398174 -25096 398230 -25040
rect 398316 -25096 398372 -25040
rect 398174 -25238 398230 -25182
rect 398316 -25238 398372 -25182
rect 398174 -25380 398230 -25324
rect 398316 -25380 398372 -25324
rect 398174 -25522 398230 -25466
rect 398316 -25522 398372 -25466
rect 398574 -13736 398630 -13680
rect 398716 -13736 398772 -13680
rect 398574 -13878 398630 -13822
rect 398716 -13878 398772 -13822
rect 398574 -14020 398630 -13964
rect 398716 -14020 398772 -13964
rect 398574 -14162 398630 -14106
rect 398716 -14162 398772 -14106
rect 398574 -14304 398630 -14248
rect 398716 -14304 398772 -14248
rect 398574 -14446 398630 -14390
rect 398716 -14446 398772 -14390
rect 398574 -14588 398630 -14532
rect 398716 -14588 398772 -14532
rect 398574 -14730 398630 -14674
rect 398716 -14730 398772 -14674
rect 398574 -14872 398630 -14816
rect 398716 -14872 398772 -14816
rect 398574 -15014 398630 -14958
rect 398716 -15014 398772 -14958
rect 398574 -15156 398630 -15100
rect 398716 -15156 398772 -15100
rect 398574 -15298 398630 -15242
rect 398716 -15298 398772 -15242
rect 398574 -15440 398630 -15384
rect 398716 -15440 398772 -15384
rect 398574 -15582 398630 -15526
rect 398716 -15582 398772 -15526
rect 398574 -15724 398630 -15668
rect 398716 -15724 398772 -15668
rect 398574 -15866 398630 -15810
rect 398716 -15866 398772 -15810
rect 398574 -16008 398630 -15952
rect 398716 -16008 398772 -15952
rect 398574 -16150 398630 -16094
rect 398716 -16150 398772 -16094
rect 398574 -16292 398630 -16236
rect 398716 -16292 398772 -16236
rect 398574 -16434 398630 -16378
rect 398716 -16434 398772 -16378
rect 398574 -16576 398630 -16520
rect 398716 -16576 398772 -16520
rect 398574 -16718 398630 -16662
rect 398716 -16718 398772 -16662
rect 398574 -16860 398630 -16804
rect 398716 -16860 398772 -16804
rect 398574 -17002 398630 -16946
rect 398716 -17002 398772 -16946
rect 398574 -17144 398630 -17088
rect 398716 -17144 398772 -17088
rect 398574 -17286 398630 -17230
rect 398716 -17286 398772 -17230
rect 398574 -17428 398630 -17372
rect 398716 -17428 398772 -17372
rect 398574 -17570 398630 -17514
rect 398716 -17570 398772 -17514
rect 398574 -17712 398630 -17656
rect 398716 -17712 398772 -17656
rect 398574 -17854 398630 -17798
rect 398716 -17854 398772 -17798
rect 398574 -17996 398630 -17940
rect 398716 -17996 398772 -17940
rect 398574 -18138 398630 -18082
rect 398716 -18138 398772 -18082
rect 398574 -18280 398630 -18224
rect 398716 -18280 398772 -18224
rect 398574 -18422 398630 -18366
rect 398716 -18422 398772 -18366
rect 398574 -18564 398630 -18508
rect 398716 -18564 398772 -18508
rect 398574 -18706 398630 -18650
rect 398716 -18706 398772 -18650
rect 398574 -18848 398630 -18792
rect 398716 -18848 398772 -18792
rect 398574 -18990 398630 -18934
rect 398716 -18990 398772 -18934
rect 398574 -19132 398630 -19076
rect 398716 -19132 398772 -19076
rect 398574 -19274 398630 -19218
rect 398716 -19274 398772 -19218
rect 398574 -19416 398630 -19360
rect 398716 -19416 398772 -19360
rect 398574 -19558 398630 -19502
rect 398716 -19558 398772 -19502
rect 398574 -19700 398630 -19644
rect 398716 -19700 398772 -19644
rect 398574 -19842 398630 -19786
rect 398716 -19842 398772 -19786
rect 398574 -19984 398630 -19928
rect 398716 -19984 398772 -19928
rect 398574 -20126 398630 -20070
rect 398716 -20126 398772 -20070
rect 398574 -20268 398630 -20212
rect 398716 -20268 398772 -20212
rect 398574 -20410 398630 -20354
rect 398716 -20410 398772 -20354
rect 398574 -20552 398630 -20496
rect 398716 -20552 398772 -20496
rect 398574 -20694 398630 -20638
rect 398716 -20694 398772 -20638
rect 398574 -20836 398630 -20780
rect 398716 -20836 398772 -20780
rect 398574 -20978 398630 -20922
rect 398716 -20978 398772 -20922
rect 398574 -21120 398630 -21064
rect 398716 -21120 398772 -21064
rect 398574 -21262 398630 -21206
rect 398716 -21262 398772 -21206
rect 398574 -21404 398630 -21348
rect 398716 -21404 398772 -21348
rect 398574 -21546 398630 -21490
rect 398716 -21546 398772 -21490
rect 398574 -21688 398630 -21632
rect 398716 -21688 398772 -21632
rect 398574 -21830 398630 -21774
rect 398716 -21830 398772 -21774
rect 398574 -21972 398630 -21916
rect 398716 -21972 398772 -21916
rect 398574 -22114 398630 -22058
rect 398716 -22114 398772 -22058
rect 398574 -22256 398630 -22200
rect 398716 -22256 398772 -22200
rect 398574 -22398 398630 -22342
rect 398716 -22398 398772 -22342
rect 398574 -22540 398630 -22484
rect 398716 -22540 398772 -22484
rect 398574 -22682 398630 -22626
rect 398716 -22682 398772 -22626
rect 398574 -22824 398630 -22768
rect 398716 -22824 398772 -22768
rect 398574 -22966 398630 -22910
rect 398716 -22966 398772 -22910
rect 398574 -23108 398630 -23052
rect 398716 -23108 398772 -23052
rect 398574 -23250 398630 -23194
rect 398716 -23250 398772 -23194
rect 398574 -23392 398630 -23336
rect 398716 -23392 398772 -23336
rect 398574 -23534 398630 -23478
rect 398716 -23534 398772 -23478
rect 398574 -23676 398630 -23620
rect 398716 -23676 398772 -23620
rect 398574 -23818 398630 -23762
rect 398716 -23818 398772 -23762
rect 398574 -23960 398630 -23904
rect 398716 -23960 398772 -23904
rect 398574 -24102 398630 -24046
rect 398716 -24102 398772 -24046
rect 398574 -24244 398630 -24188
rect 398716 -24244 398772 -24188
rect 398574 -24386 398630 -24330
rect 398716 -24386 398772 -24330
rect 398574 -24528 398630 -24472
rect 398716 -24528 398772 -24472
rect 398574 -24670 398630 -24614
rect 398716 -24670 398772 -24614
rect 398574 -24812 398630 -24756
rect 398716 -24812 398772 -24756
rect 398574 -24954 398630 -24898
rect 398716 -24954 398772 -24898
rect 398574 -25096 398630 -25040
rect 398716 -25096 398772 -25040
rect 398574 -25238 398630 -25182
rect 398716 -25238 398772 -25182
rect 398574 -25380 398630 -25324
rect 398716 -25380 398772 -25324
rect 398574 -25522 398630 -25466
rect 398716 -25522 398772 -25466
rect 398971 -13736 399027 -13680
rect 399113 -13736 399169 -13680
rect 398971 -13878 399027 -13822
rect 399113 -13878 399169 -13822
rect 398971 -14020 399027 -13964
rect 399113 -14020 399169 -13964
rect 398971 -14162 399027 -14106
rect 399113 -14162 399169 -14106
rect 398971 -14304 399027 -14248
rect 399113 -14304 399169 -14248
rect 398971 -14446 399027 -14390
rect 399113 -14446 399169 -14390
rect 398971 -14588 399027 -14532
rect 399113 -14588 399169 -14532
rect 398971 -14730 399027 -14674
rect 399113 -14730 399169 -14674
rect 398971 -14872 399027 -14816
rect 399113 -14872 399169 -14816
rect 398971 -15014 399027 -14958
rect 399113 -15014 399169 -14958
rect 398971 -15156 399027 -15100
rect 399113 -15156 399169 -15100
rect 398971 -15298 399027 -15242
rect 399113 -15298 399169 -15242
rect 398971 -15440 399027 -15384
rect 399113 -15440 399169 -15384
rect 398971 -15582 399027 -15526
rect 399113 -15582 399169 -15526
rect 398971 -15724 399027 -15668
rect 399113 -15724 399169 -15668
rect 398971 -15866 399027 -15810
rect 399113 -15866 399169 -15810
rect 398971 -16008 399027 -15952
rect 399113 -16008 399169 -15952
rect 398971 -16150 399027 -16094
rect 399113 -16150 399169 -16094
rect 398971 -16292 399027 -16236
rect 399113 -16292 399169 -16236
rect 398971 -16434 399027 -16378
rect 399113 -16434 399169 -16378
rect 398971 -16576 399027 -16520
rect 399113 -16576 399169 -16520
rect 398971 -16718 399027 -16662
rect 399113 -16718 399169 -16662
rect 398971 -16860 399027 -16804
rect 399113 -16860 399169 -16804
rect 398971 -17002 399027 -16946
rect 399113 -17002 399169 -16946
rect 398971 -17144 399027 -17088
rect 399113 -17144 399169 -17088
rect 398971 -17286 399027 -17230
rect 399113 -17286 399169 -17230
rect 398971 -17428 399027 -17372
rect 399113 -17428 399169 -17372
rect 398971 -17570 399027 -17514
rect 399113 -17570 399169 -17514
rect 398971 -17712 399027 -17656
rect 399113 -17712 399169 -17656
rect 398971 -17854 399027 -17798
rect 399113 -17854 399169 -17798
rect 398971 -17996 399027 -17940
rect 399113 -17996 399169 -17940
rect 398971 -18138 399027 -18082
rect 399113 -18138 399169 -18082
rect 398971 -18280 399027 -18224
rect 399113 -18280 399169 -18224
rect 398971 -18422 399027 -18366
rect 399113 -18422 399169 -18366
rect 398971 -18564 399027 -18508
rect 399113 -18564 399169 -18508
rect 398971 -18706 399027 -18650
rect 399113 -18706 399169 -18650
rect 398971 -18848 399027 -18792
rect 399113 -18848 399169 -18792
rect 398971 -18990 399027 -18934
rect 399113 -18990 399169 -18934
rect 398971 -19132 399027 -19076
rect 399113 -19132 399169 -19076
rect 398971 -19274 399027 -19218
rect 399113 -19274 399169 -19218
rect 398971 -19416 399027 -19360
rect 399113 -19416 399169 -19360
rect 398971 -19558 399027 -19502
rect 399113 -19558 399169 -19502
rect 398971 -19700 399027 -19644
rect 399113 -19700 399169 -19644
rect 398971 -19842 399027 -19786
rect 399113 -19842 399169 -19786
rect 398971 -19984 399027 -19928
rect 399113 -19984 399169 -19928
rect 398971 -20126 399027 -20070
rect 399113 -20126 399169 -20070
rect 398971 -20268 399027 -20212
rect 399113 -20268 399169 -20212
rect 398971 -20410 399027 -20354
rect 399113 -20410 399169 -20354
rect 398971 -20552 399027 -20496
rect 399113 -20552 399169 -20496
rect 398971 -20694 399027 -20638
rect 399113 -20694 399169 -20638
rect 398971 -20836 399027 -20780
rect 399113 -20836 399169 -20780
rect 398971 -20978 399027 -20922
rect 399113 -20978 399169 -20922
rect 398971 -21120 399027 -21064
rect 399113 -21120 399169 -21064
rect 398971 -21262 399027 -21206
rect 399113 -21262 399169 -21206
rect 398971 -21404 399027 -21348
rect 399113 -21404 399169 -21348
rect 398971 -21546 399027 -21490
rect 399113 -21546 399169 -21490
rect 398971 -21688 399027 -21632
rect 399113 -21688 399169 -21632
rect 398971 -21830 399027 -21774
rect 399113 -21830 399169 -21774
rect 398971 -21972 399027 -21916
rect 399113 -21972 399169 -21916
rect 398971 -22114 399027 -22058
rect 399113 -22114 399169 -22058
rect 398971 -22256 399027 -22200
rect 399113 -22256 399169 -22200
rect 398971 -22398 399027 -22342
rect 399113 -22398 399169 -22342
rect 398971 -22540 399027 -22484
rect 399113 -22540 399169 -22484
rect 398971 -22682 399027 -22626
rect 399113 -22682 399169 -22626
rect 398971 -22824 399027 -22768
rect 399113 -22824 399169 -22768
rect 398971 -22966 399027 -22910
rect 399113 -22966 399169 -22910
rect 398971 -23108 399027 -23052
rect 399113 -23108 399169 -23052
rect 398971 -23250 399027 -23194
rect 399113 -23250 399169 -23194
rect 398971 -23392 399027 -23336
rect 399113 -23392 399169 -23336
rect 398971 -23534 399027 -23478
rect 399113 -23534 399169 -23478
rect 398971 -23676 399027 -23620
rect 399113 -23676 399169 -23620
rect 398971 -23818 399027 -23762
rect 399113 -23818 399169 -23762
rect 398971 -23960 399027 -23904
rect 399113 -23960 399169 -23904
rect 398971 -24102 399027 -24046
rect 399113 -24102 399169 -24046
rect 398971 -24244 399027 -24188
rect 399113 -24244 399169 -24188
rect 398971 -24386 399027 -24330
rect 399113 -24386 399169 -24330
rect 398971 -24528 399027 -24472
rect 399113 -24528 399169 -24472
rect 398971 -24670 399027 -24614
rect 399113 -24670 399169 -24614
rect 398971 -24812 399027 -24756
rect 399113 -24812 399169 -24756
rect 398971 -24954 399027 -24898
rect 399113 -24954 399169 -24898
rect 398971 -25096 399027 -25040
rect 399113 -25096 399169 -25040
rect 398971 -25238 399027 -25182
rect 399113 -25238 399169 -25182
rect 398971 -25380 399027 -25324
rect 399113 -25380 399169 -25324
rect 398971 -25522 399027 -25466
rect 399113 -25522 399169 -25466
rect 399376 -13736 399432 -13680
rect 399518 -13736 399574 -13680
rect 399376 -13878 399432 -13822
rect 399518 -13878 399574 -13822
rect 399376 -14020 399432 -13964
rect 399518 -14020 399574 -13964
rect 399376 -14162 399432 -14106
rect 399518 -14162 399574 -14106
rect 399376 -14304 399432 -14248
rect 399518 -14304 399574 -14248
rect 399376 -14446 399432 -14390
rect 399518 -14446 399574 -14390
rect 399376 -14588 399432 -14532
rect 399518 -14588 399574 -14532
rect 399376 -14730 399432 -14674
rect 399518 -14730 399574 -14674
rect 399376 -14872 399432 -14816
rect 399518 -14872 399574 -14816
rect 399376 -15014 399432 -14958
rect 399518 -15014 399574 -14958
rect 399376 -15156 399432 -15100
rect 399518 -15156 399574 -15100
rect 399376 -15298 399432 -15242
rect 399518 -15298 399574 -15242
rect 399376 -15440 399432 -15384
rect 399518 -15440 399574 -15384
rect 399376 -15582 399432 -15526
rect 399518 -15582 399574 -15526
rect 399376 -15724 399432 -15668
rect 399518 -15724 399574 -15668
rect 399376 -15866 399432 -15810
rect 399518 -15866 399574 -15810
rect 399376 -16008 399432 -15952
rect 399518 -16008 399574 -15952
rect 399376 -16150 399432 -16094
rect 399518 -16150 399574 -16094
rect 399376 -16292 399432 -16236
rect 399518 -16292 399574 -16236
rect 399376 -16434 399432 -16378
rect 399518 -16434 399574 -16378
rect 399376 -16576 399432 -16520
rect 399518 -16576 399574 -16520
rect 399376 -16718 399432 -16662
rect 399518 -16718 399574 -16662
rect 399376 -16860 399432 -16804
rect 399518 -16860 399574 -16804
rect 399376 -17002 399432 -16946
rect 399518 -17002 399574 -16946
rect 399376 -17144 399432 -17088
rect 399518 -17144 399574 -17088
rect 399376 -17286 399432 -17230
rect 399518 -17286 399574 -17230
rect 399376 -17428 399432 -17372
rect 399518 -17428 399574 -17372
rect 399376 -17570 399432 -17514
rect 399518 -17570 399574 -17514
rect 399376 -17712 399432 -17656
rect 399518 -17712 399574 -17656
rect 399376 -17854 399432 -17798
rect 399518 -17854 399574 -17798
rect 399376 -17996 399432 -17940
rect 399518 -17996 399574 -17940
rect 399376 -18138 399432 -18082
rect 399518 -18138 399574 -18082
rect 399376 -18280 399432 -18224
rect 399518 -18280 399574 -18224
rect 399376 -18422 399432 -18366
rect 399518 -18422 399574 -18366
rect 399376 -18564 399432 -18508
rect 399518 -18564 399574 -18508
rect 399376 -18706 399432 -18650
rect 399518 -18706 399574 -18650
rect 399376 -18848 399432 -18792
rect 399518 -18848 399574 -18792
rect 399376 -18990 399432 -18934
rect 399518 -18990 399574 -18934
rect 399376 -19132 399432 -19076
rect 399518 -19132 399574 -19076
rect 399376 -19274 399432 -19218
rect 399518 -19274 399574 -19218
rect 399376 -19416 399432 -19360
rect 399518 -19416 399574 -19360
rect 399376 -19558 399432 -19502
rect 399518 -19558 399574 -19502
rect 399376 -19700 399432 -19644
rect 399518 -19700 399574 -19644
rect 399376 -19842 399432 -19786
rect 399518 -19842 399574 -19786
rect 399376 -19984 399432 -19928
rect 399518 -19984 399574 -19928
rect 399376 -20126 399432 -20070
rect 399518 -20126 399574 -20070
rect 399376 -20268 399432 -20212
rect 399518 -20268 399574 -20212
rect 399376 -20410 399432 -20354
rect 399518 -20410 399574 -20354
rect 399376 -20552 399432 -20496
rect 399518 -20552 399574 -20496
rect 399376 -20694 399432 -20638
rect 399518 -20694 399574 -20638
rect 399376 -20836 399432 -20780
rect 399518 -20836 399574 -20780
rect 399376 -20978 399432 -20922
rect 399518 -20978 399574 -20922
rect 399376 -21120 399432 -21064
rect 399518 -21120 399574 -21064
rect 399376 -21262 399432 -21206
rect 399518 -21262 399574 -21206
rect 399376 -21404 399432 -21348
rect 399518 -21404 399574 -21348
rect 399376 -21546 399432 -21490
rect 399518 -21546 399574 -21490
rect 399376 -21688 399432 -21632
rect 399518 -21688 399574 -21632
rect 399376 -21830 399432 -21774
rect 399518 -21830 399574 -21774
rect 399376 -21972 399432 -21916
rect 399518 -21972 399574 -21916
rect 399376 -22114 399432 -22058
rect 399518 -22114 399574 -22058
rect 399376 -22256 399432 -22200
rect 399518 -22256 399574 -22200
rect 399376 -22398 399432 -22342
rect 399518 -22398 399574 -22342
rect 399376 -22540 399432 -22484
rect 399518 -22540 399574 -22484
rect 399376 -22682 399432 -22626
rect 399518 -22682 399574 -22626
rect 399376 -22824 399432 -22768
rect 399518 -22824 399574 -22768
rect 399376 -22966 399432 -22910
rect 399518 -22966 399574 -22910
rect 399376 -23108 399432 -23052
rect 399518 -23108 399574 -23052
rect 399376 -23250 399432 -23194
rect 399518 -23250 399574 -23194
rect 399376 -23392 399432 -23336
rect 399518 -23392 399574 -23336
rect 399376 -23534 399432 -23478
rect 399518 -23534 399574 -23478
rect 399376 -23676 399432 -23620
rect 399518 -23676 399574 -23620
rect 399376 -23818 399432 -23762
rect 399518 -23818 399574 -23762
rect 399376 -23960 399432 -23904
rect 399518 -23960 399574 -23904
rect 399376 -24102 399432 -24046
rect 399518 -24102 399574 -24046
rect 399376 -24244 399432 -24188
rect 399518 -24244 399574 -24188
rect 399376 -24386 399432 -24330
rect 399518 -24386 399574 -24330
rect 399376 -24528 399432 -24472
rect 399518 -24528 399574 -24472
rect 399376 -24670 399432 -24614
rect 399518 -24670 399574 -24614
rect 399376 -24812 399432 -24756
rect 399518 -24812 399574 -24756
rect 399376 -24954 399432 -24898
rect 399518 -24954 399574 -24898
rect 399376 -25096 399432 -25040
rect 399518 -25096 399574 -25040
rect 399376 -25238 399432 -25182
rect 399518 -25238 399574 -25182
rect 399376 -25380 399432 -25324
rect 399518 -25380 399574 -25324
rect 399376 -25522 399432 -25466
rect 399518 -25522 399574 -25466
rect 399776 -13736 399832 -13680
rect 399918 -13736 399974 -13680
rect 399776 -13878 399832 -13822
rect 399918 -13878 399974 -13822
rect 399776 -14020 399832 -13964
rect 399918 -14020 399974 -13964
rect 399776 -14162 399832 -14106
rect 399918 -14162 399974 -14106
rect 399776 -14304 399832 -14248
rect 399918 -14304 399974 -14248
rect 399776 -14446 399832 -14390
rect 399918 -14446 399974 -14390
rect 399776 -14588 399832 -14532
rect 399918 -14588 399974 -14532
rect 399776 -14730 399832 -14674
rect 399918 -14730 399974 -14674
rect 399776 -14872 399832 -14816
rect 399918 -14872 399974 -14816
rect 399776 -15014 399832 -14958
rect 399918 -15014 399974 -14958
rect 399776 -15156 399832 -15100
rect 399918 -15156 399974 -15100
rect 399776 -15298 399832 -15242
rect 399918 -15298 399974 -15242
rect 399776 -15440 399832 -15384
rect 399918 -15440 399974 -15384
rect 399776 -15582 399832 -15526
rect 399918 -15582 399974 -15526
rect 399776 -15724 399832 -15668
rect 399918 -15724 399974 -15668
rect 399776 -15866 399832 -15810
rect 399918 -15866 399974 -15810
rect 399776 -16008 399832 -15952
rect 399918 -16008 399974 -15952
rect 399776 -16150 399832 -16094
rect 399918 -16150 399974 -16094
rect 399776 -16292 399832 -16236
rect 399918 -16292 399974 -16236
rect 399776 -16434 399832 -16378
rect 399918 -16434 399974 -16378
rect 399776 -16576 399832 -16520
rect 399918 -16576 399974 -16520
rect 399776 -16718 399832 -16662
rect 399918 -16718 399974 -16662
rect 399776 -16860 399832 -16804
rect 399918 -16860 399974 -16804
rect 399776 -17002 399832 -16946
rect 399918 -17002 399974 -16946
rect 399776 -17144 399832 -17088
rect 399918 -17144 399974 -17088
rect 399776 -17286 399832 -17230
rect 399918 -17286 399974 -17230
rect 399776 -17428 399832 -17372
rect 399918 -17428 399974 -17372
rect 399776 -17570 399832 -17514
rect 399918 -17570 399974 -17514
rect 399776 -17712 399832 -17656
rect 399918 -17712 399974 -17656
rect 399776 -17854 399832 -17798
rect 399918 -17854 399974 -17798
rect 399776 -17996 399832 -17940
rect 399918 -17996 399974 -17940
rect 399776 -18138 399832 -18082
rect 399918 -18138 399974 -18082
rect 399776 -18280 399832 -18224
rect 399918 -18280 399974 -18224
rect 399776 -18422 399832 -18366
rect 399918 -18422 399974 -18366
rect 399776 -18564 399832 -18508
rect 399918 -18564 399974 -18508
rect 399776 -18706 399832 -18650
rect 399918 -18706 399974 -18650
rect 399776 -18848 399832 -18792
rect 399918 -18848 399974 -18792
rect 399776 -18990 399832 -18934
rect 399918 -18990 399974 -18934
rect 399776 -19132 399832 -19076
rect 399918 -19132 399974 -19076
rect 399776 -19274 399832 -19218
rect 399918 -19274 399974 -19218
rect 399776 -19416 399832 -19360
rect 399918 -19416 399974 -19360
rect 399776 -19558 399832 -19502
rect 399918 -19558 399974 -19502
rect 399776 -19700 399832 -19644
rect 399918 -19700 399974 -19644
rect 399776 -19842 399832 -19786
rect 399918 -19842 399974 -19786
rect 399776 -19984 399832 -19928
rect 399918 -19984 399974 -19928
rect 399776 -20126 399832 -20070
rect 399918 -20126 399974 -20070
rect 399776 -20268 399832 -20212
rect 399918 -20268 399974 -20212
rect 399776 -20410 399832 -20354
rect 399918 -20410 399974 -20354
rect 399776 -20552 399832 -20496
rect 399918 -20552 399974 -20496
rect 399776 -20694 399832 -20638
rect 399918 -20694 399974 -20638
rect 399776 -20836 399832 -20780
rect 399918 -20836 399974 -20780
rect 399776 -20978 399832 -20922
rect 399918 -20978 399974 -20922
rect 399776 -21120 399832 -21064
rect 399918 -21120 399974 -21064
rect 399776 -21262 399832 -21206
rect 399918 -21262 399974 -21206
rect 399776 -21404 399832 -21348
rect 399918 -21404 399974 -21348
rect 399776 -21546 399832 -21490
rect 399918 -21546 399974 -21490
rect 399776 -21688 399832 -21632
rect 399918 -21688 399974 -21632
rect 399776 -21830 399832 -21774
rect 399918 -21830 399974 -21774
rect 399776 -21972 399832 -21916
rect 399918 -21972 399974 -21916
rect 399776 -22114 399832 -22058
rect 399918 -22114 399974 -22058
rect 399776 -22256 399832 -22200
rect 399918 -22256 399974 -22200
rect 399776 -22398 399832 -22342
rect 399918 -22398 399974 -22342
rect 399776 -22540 399832 -22484
rect 399918 -22540 399974 -22484
rect 399776 -22682 399832 -22626
rect 399918 -22682 399974 -22626
rect 399776 -22824 399832 -22768
rect 399918 -22824 399974 -22768
rect 399776 -22966 399832 -22910
rect 399918 -22966 399974 -22910
rect 399776 -23108 399832 -23052
rect 399918 -23108 399974 -23052
rect 399776 -23250 399832 -23194
rect 399918 -23250 399974 -23194
rect 399776 -23392 399832 -23336
rect 399918 -23392 399974 -23336
rect 399776 -23534 399832 -23478
rect 399918 -23534 399974 -23478
rect 399776 -23676 399832 -23620
rect 399918 -23676 399974 -23620
rect 399776 -23818 399832 -23762
rect 399918 -23818 399974 -23762
rect 399776 -23960 399832 -23904
rect 399918 -23960 399974 -23904
rect 399776 -24102 399832 -24046
rect 399918 -24102 399974 -24046
rect 399776 -24244 399832 -24188
rect 399918 -24244 399974 -24188
rect 399776 -24386 399832 -24330
rect 399918 -24386 399974 -24330
rect 399776 -24528 399832 -24472
rect 399918 -24528 399974 -24472
rect 399776 -24670 399832 -24614
rect 399918 -24670 399974 -24614
rect 399776 -24812 399832 -24756
rect 399918 -24812 399974 -24756
rect 399776 -24954 399832 -24898
rect 399918 -24954 399974 -24898
rect 399776 -25096 399832 -25040
rect 399918 -25096 399974 -25040
rect 399776 -25238 399832 -25182
rect 399918 -25238 399974 -25182
rect 399776 -25380 399832 -25324
rect 399918 -25380 399974 -25324
rect 399776 -25522 399832 -25466
rect 399918 -25522 399974 -25466
rect 400181 -13736 400237 -13680
rect 400323 -13736 400379 -13680
rect 400181 -13878 400237 -13822
rect 400323 -13878 400379 -13822
rect 400181 -14020 400237 -13964
rect 400323 -14020 400379 -13964
rect 400181 -14162 400237 -14106
rect 400323 -14162 400379 -14106
rect 400181 -14304 400237 -14248
rect 400323 -14304 400379 -14248
rect 400181 -14446 400237 -14390
rect 400323 -14446 400379 -14390
rect 400181 -14588 400237 -14532
rect 400323 -14588 400379 -14532
rect 400181 -14730 400237 -14674
rect 400323 -14730 400379 -14674
rect 400181 -14872 400237 -14816
rect 400323 -14872 400379 -14816
rect 400181 -15014 400237 -14958
rect 400323 -15014 400379 -14958
rect 400181 -15156 400237 -15100
rect 400323 -15156 400379 -15100
rect 400181 -15298 400237 -15242
rect 400323 -15298 400379 -15242
rect 400181 -15440 400237 -15384
rect 400323 -15440 400379 -15384
rect 400181 -15582 400237 -15526
rect 400323 -15582 400379 -15526
rect 400181 -15724 400237 -15668
rect 400323 -15724 400379 -15668
rect 400181 -15866 400237 -15810
rect 400323 -15866 400379 -15810
rect 400181 -16008 400237 -15952
rect 400323 -16008 400379 -15952
rect 400181 -16150 400237 -16094
rect 400323 -16150 400379 -16094
rect 400181 -16292 400237 -16236
rect 400323 -16292 400379 -16236
rect 400181 -16434 400237 -16378
rect 400323 -16434 400379 -16378
rect 400181 -16576 400237 -16520
rect 400323 -16576 400379 -16520
rect 400181 -16718 400237 -16662
rect 400323 -16718 400379 -16662
rect 400181 -16860 400237 -16804
rect 400323 -16860 400379 -16804
rect 400181 -17002 400237 -16946
rect 400323 -17002 400379 -16946
rect 400181 -17144 400237 -17088
rect 400323 -17144 400379 -17088
rect 400181 -17286 400237 -17230
rect 400323 -17286 400379 -17230
rect 400181 -17428 400237 -17372
rect 400323 -17428 400379 -17372
rect 400181 -17570 400237 -17514
rect 400323 -17570 400379 -17514
rect 400181 -17712 400237 -17656
rect 400323 -17712 400379 -17656
rect 400181 -17854 400237 -17798
rect 400323 -17854 400379 -17798
rect 400181 -17996 400237 -17940
rect 400323 -17996 400379 -17940
rect 400181 -18138 400237 -18082
rect 400323 -18138 400379 -18082
rect 400181 -18280 400237 -18224
rect 400323 -18280 400379 -18224
rect 400181 -18422 400237 -18366
rect 400323 -18422 400379 -18366
rect 400181 -18564 400237 -18508
rect 400323 -18564 400379 -18508
rect 400181 -18706 400237 -18650
rect 400323 -18706 400379 -18650
rect 400181 -18848 400237 -18792
rect 400323 -18848 400379 -18792
rect 400181 -18990 400237 -18934
rect 400323 -18990 400379 -18934
rect 400181 -19132 400237 -19076
rect 400323 -19132 400379 -19076
rect 400181 -19274 400237 -19218
rect 400323 -19274 400379 -19218
rect 400181 -19416 400237 -19360
rect 400323 -19416 400379 -19360
rect 400181 -19558 400237 -19502
rect 400323 -19558 400379 -19502
rect 400181 -19700 400237 -19644
rect 400323 -19700 400379 -19644
rect 400181 -19842 400237 -19786
rect 400323 -19842 400379 -19786
rect 400181 -19984 400237 -19928
rect 400323 -19984 400379 -19928
rect 400181 -20126 400237 -20070
rect 400323 -20126 400379 -20070
rect 400181 -20268 400237 -20212
rect 400323 -20268 400379 -20212
rect 400181 -20410 400237 -20354
rect 400323 -20410 400379 -20354
rect 400181 -20552 400237 -20496
rect 400323 -20552 400379 -20496
rect 400181 -20694 400237 -20638
rect 400323 -20694 400379 -20638
rect 400181 -20836 400237 -20780
rect 400323 -20836 400379 -20780
rect 400181 -20978 400237 -20922
rect 400323 -20978 400379 -20922
rect 400181 -21120 400237 -21064
rect 400323 -21120 400379 -21064
rect 400181 -21262 400237 -21206
rect 400323 -21262 400379 -21206
rect 400181 -21404 400237 -21348
rect 400323 -21404 400379 -21348
rect 400181 -21546 400237 -21490
rect 400323 -21546 400379 -21490
rect 400181 -21688 400237 -21632
rect 400323 -21688 400379 -21632
rect 400181 -21830 400237 -21774
rect 400323 -21830 400379 -21774
rect 400181 -21972 400237 -21916
rect 400323 -21972 400379 -21916
rect 400181 -22114 400237 -22058
rect 400323 -22114 400379 -22058
rect 400181 -22256 400237 -22200
rect 400323 -22256 400379 -22200
rect 400181 -22398 400237 -22342
rect 400323 -22398 400379 -22342
rect 400181 -22540 400237 -22484
rect 400323 -22540 400379 -22484
rect 400181 -22682 400237 -22626
rect 400323 -22682 400379 -22626
rect 400181 -22824 400237 -22768
rect 400323 -22824 400379 -22768
rect 400181 -22966 400237 -22910
rect 400323 -22966 400379 -22910
rect 400181 -23108 400237 -23052
rect 400323 -23108 400379 -23052
rect 400181 -23250 400237 -23194
rect 400323 -23250 400379 -23194
rect 400181 -23392 400237 -23336
rect 400323 -23392 400379 -23336
rect 400181 -23534 400237 -23478
rect 400323 -23534 400379 -23478
rect 400181 -23676 400237 -23620
rect 400323 -23676 400379 -23620
rect 400181 -23818 400237 -23762
rect 400323 -23818 400379 -23762
rect 400181 -23960 400237 -23904
rect 400323 -23960 400379 -23904
rect 400181 -24102 400237 -24046
rect 400323 -24102 400379 -24046
rect 400181 -24244 400237 -24188
rect 400323 -24244 400379 -24188
rect 400181 -24386 400237 -24330
rect 400323 -24386 400379 -24330
rect 400181 -24528 400237 -24472
rect 400323 -24528 400379 -24472
rect 400181 -24670 400237 -24614
rect 400323 -24670 400379 -24614
rect 400181 -24812 400237 -24756
rect 400323 -24812 400379 -24756
rect 400181 -24954 400237 -24898
rect 400323 -24954 400379 -24898
rect 400181 -25096 400237 -25040
rect 400323 -25096 400379 -25040
rect 400181 -25238 400237 -25182
rect 400323 -25238 400379 -25182
rect 400181 -25380 400237 -25324
rect 400323 -25380 400379 -25324
rect 400181 -25522 400237 -25466
rect 400323 -25522 400379 -25466
rect 400766 -13688 400822 -13632
rect 400890 -13688 400946 -13632
rect 401014 -13688 401070 -13632
rect 401138 -13688 401194 -13632
rect 401262 -13688 401318 -13632
rect 400766 -13812 400822 -13756
rect 400890 -13812 400946 -13756
rect 401014 -13812 401070 -13756
rect 401138 -13812 401194 -13756
rect 401262 -13812 401318 -13756
rect 400766 -13936 400822 -13880
rect 400890 -13936 400946 -13880
rect 401014 -13936 401070 -13880
rect 401138 -13936 401194 -13880
rect 401262 -13936 401318 -13880
rect 400766 -14060 400822 -14004
rect 400890 -14060 400946 -14004
rect 401014 -14060 401070 -14004
rect 401138 -14060 401194 -14004
rect 401262 -14060 401318 -14004
rect 400766 -14184 400822 -14128
rect 400890 -14184 400946 -14128
rect 401014 -14184 401070 -14128
rect 401138 -14184 401194 -14128
rect 401262 -14184 401318 -14128
rect 400766 -14308 400822 -14252
rect 400890 -14308 400946 -14252
rect 401014 -14308 401070 -14252
rect 401138 -14308 401194 -14252
rect 401262 -14308 401318 -14252
rect 400766 -14432 400822 -14376
rect 400890 -14432 400946 -14376
rect 401014 -14432 401070 -14376
rect 401138 -14432 401194 -14376
rect 401262 -14432 401318 -14376
rect 400766 -14556 400822 -14500
rect 400890 -14556 400946 -14500
rect 401014 -14556 401070 -14500
rect 401138 -14556 401194 -14500
rect 401262 -14556 401318 -14500
rect 400766 -14680 400822 -14624
rect 400890 -14680 400946 -14624
rect 401014 -14680 401070 -14624
rect 401138 -14680 401194 -14624
rect 401262 -14680 401318 -14624
rect 400766 -14804 400822 -14748
rect 400890 -14804 400946 -14748
rect 401014 -14804 401070 -14748
rect 401138 -14804 401194 -14748
rect 401262 -14804 401318 -14748
rect 400766 -14928 400822 -14872
rect 400890 -14928 400946 -14872
rect 401014 -14928 401070 -14872
rect 401138 -14928 401194 -14872
rect 401262 -14928 401318 -14872
rect 400766 -15052 400822 -14996
rect 400890 -15052 400946 -14996
rect 401014 -15052 401070 -14996
rect 401138 -15052 401194 -14996
rect 401262 -15052 401318 -14996
rect 400766 -15176 400822 -15120
rect 400890 -15176 400946 -15120
rect 401014 -15176 401070 -15120
rect 401138 -15176 401194 -15120
rect 401262 -15176 401318 -15120
rect 400766 -15300 400822 -15244
rect 400890 -15300 400946 -15244
rect 401014 -15300 401070 -15244
rect 401138 -15300 401194 -15244
rect 401262 -15300 401318 -15244
rect 400766 -15424 400822 -15368
rect 400890 -15424 400946 -15368
rect 401014 -15424 401070 -15368
rect 401138 -15424 401194 -15368
rect 401262 -15424 401318 -15368
rect 400766 -15548 400822 -15492
rect 400890 -15548 400946 -15492
rect 401014 -15548 401070 -15492
rect 401138 -15548 401194 -15492
rect 401262 -15548 401318 -15492
rect 400766 -15672 400822 -15616
rect 400890 -15672 400946 -15616
rect 401014 -15672 401070 -15616
rect 401138 -15672 401194 -15616
rect 401262 -15672 401318 -15616
rect 400766 -15796 400822 -15740
rect 400890 -15796 400946 -15740
rect 401014 -15796 401070 -15740
rect 401138 -15796 401194 -15740
rect 401262 -15796 401318 -15740
rect 400766 -15920 400822 -15864
rect 400890 -15920 400946 -15864
rect 401014 -15920 401070 -15864
rect 401138 -15920 401194 -15864
rect 401262 -15920 401318 -15864
rect 400766 -16044 400822 -15988
rect 400890 -16044 400946 -15988
rect 401014 -16044 401070 -15988
rect 401138 -16044 401194 -15988
rect 401262 -16044 401318 -15988
rect 400766 -16168 400822 -16112
rect 400890 -16168 400946 -16112
rect 401014 -16168 401070 -16112
rect 401138 -16168 401194 -16112
rect 401262 -16168 401318 -16112
rect 400766 -16292 400822 -16236
rect 400890 -16292 400946 -16236
rect 401014 -16292 401070 -16236
rect 401138 -16292 401194 -16236
rect 401262 -16292 401318 -16236
rect 400766 -16416 400822 -16360
rect 400890 -16416 400946 -16360
rect 401014 -16416 401070 -16360
rect 401138 -16416 401194 -16360
rect 401262 -16416 401318 -16360
rect 400766 -16540 400822 -16484
rect 400890 -16540 400946 -16484
rect 401014 -16540 401070 -16484
rect 401138 -16540 401194 -16484
rect 401262 -16540 401318 -16484
rect 400766 -16664 400822 -16608
rect 400890 -16664 400946 -16608
rect 401014 -16664 401070 -16608
rect 401138 -16664 401194 -16608
rect 401262 -16664 401318 -16608
rect 400766 -16788 400822 -16732
rect 400890 -16788 400946 -16732
rect 401014 -16788 401070 -16732
rect 401138 -16788 401194 -16732
rect 401262 -16788 401318 -16732
rect 400766 -16912 400822 -16856
rect 400890 -16912 400946 -16856
rect 401014 -16912 401070 -16856
rect 401138 -16912 401194 -16856
rect 401262 -16912 401318 -16856
rect 400766 -17036 400822 -16980
rect 400890 -17036 400946 -16980
rect 401014 -17036 401070 -16980
rect 401138 -17036 401194 -16980
rect 401262 -17036 401318 -16980
rect 400766 -17160 400822 -17104
rect 400890 -17160 400946 -17104
rect 401014 -17160 401070 -17104
rect 401138 -17160 401194 -17104
rect 401262 -17160 401318 -17104
rect 400766 -17284 400822 -17228
rect 400890 -17284 400946 -17228
rect 401014 -17284 401070 -17228
rect 401138 -17284 401194 -17228
rect 401262 -17284 401318 -17228
rect 400766 -17408 400822 -17352
rect 400890 -17408 400946 -17352
rect 401014 -17408 401070 -17352
rect 401138 -17408 401194 -17352
rect 401262 -17408 401318 -17352
rect 400766 -17532 400822 -17476
rect 400890 -17532 400946 -17476
rect 401014 -17532 401070 -17476
rect 401138 -17532 401194 -17476
rect 401262 -17532 401318 -17476
rect 400766 -17656 400822 -17600
rect 400890 -17656 400946 -17600
rect 401014 -17656 401070 -17600
rect 401138 -17656 401194 -17600
rect 401262 -17656 401318 -17600
rect 400766 -17780 400822 -17724
rect 400890 -17780 400946 -17724
rect 401014 -17780 401070 -17724
rect 401138 -17780 401194 -17724
rect 401262 -17780 401318 -17724
rect 400766 -17904 400822 -17848
rect 400890 -17904 400946 -17848
rect 401014 -17904 401070 -17848
rect 401138 -17904 401194 -17848
rect 401262 -17904 401318 -17848
rect 400766 -18028 400822 -17972
rect 400890 -18028 400946 -17972
rect 401014 -18028 401070 -17972
rect 401138 -18028 401194 -17972
rect 401262 -18028 401318 -17972
rect 400766 -18152 400822 -18096
rect 400890 -18152 400946 -18096
rect 401014 -18152 401070 -18096
rect 401138 -18152 401194 -18096
rect 401262 -18152 401318 -18096
rect 400766 -18276 400822 -18220
rect 400890 -18276 400946 -18220
rect 401014 -18276 401070 -18220
rect 401138 -18276 401194 -18220
rect 401262 -18276 401318 -18220
rect 400766 -18400 400822 -18344
rect 400890 -18400 400946 -18344
rect 401014 -18400 401070 -18344
rect 401138 -18400 401194 -18344
rect 401262 -18400 401318 -18344
rect 400766 -18524 400822 -18468
rect 400890 -18524 400946 -18468
rect 401014 -18524 401070 -18468
rect 401138 -18524 401194 -18468
rect 401262 -18524 401318 -18468
rect 400766 -18648 400822 -18592
rect 400890 -18648 400946 -18592
rect 401014 -18648 401070 -18592
rect 401138 -18648 401194 -18592
rect 401262 -18648 401318 -18592
rect 400766 -18772 400822 -18716
rect 400890 -18772 400946 -18716
rect 401014 -18772 401070 -18716
rect 401138 -18772 401194 -18716
rect 401262 -18772 401318 -18716
rect 400766 -18896 400822 -18840
rect 400890 -18896 400946 -18840
rect 401014 -18896 401070 -18840
rect 401138 -18896 401194 -18840
rect 401262 -18896 401318 -18840
rect 400766 -19020 400822 -18964
rect 400890 -19020 400946 -18964
rect 401014 -19020 401070 -18964
rect 401138 -19020 401194 -18964
rect 401262 -19020 401318 -18964
rect 400766 -19144 400822 -19088
rect 400890 -19144 400946 -19088
rect 401014 -19144 401070 -19088
rect 401138 -19144 401194 -19088
rect 401262 -19144 401318 -19088
rect 400766 -19268 400822 -19212
rect 400890 -19268 400946 -19212
rect 401014 -19268 401070 -19212
rect 401138 -19268 401194 -19212
rect 401262 -19268 401318 -19212
rect 400766 -19392 400822 -19336
rect 400890 -19392 400946 -19336
rect 401014 -19392 401070 -19336
rect 401138 -19392 401194 -19336
rect 401262 -19392 401318 -19336
rect 400766 -19516 400822 -19460
rect 400890 -19516 400946 -19460
rect 401014 -19516 401070 -19460
rect 401138 -19516 401194 -19460
rect 401262 -19516 401318 -19460
rect 400766 -19640 400822 -19584
rect 400890 -19640 400946 -19584
rect 401014 -19640 401070 -19584
rect 401138 -19640 401194 -19584
rect 401262 -19640 401318 -19584
rect 400766 -19764 400822 -19708
rect 400890 -19764 400946 -19708
rect 401014 -19764 401070 -19708
rect 401138 -19764 401194 -19708
rect 401262 -19764 401318 -19708
rect 400766 -19888 400822 -19832
rect 400890 -19888 400946 -19832
rect 401014 -19888 401070 -19832
rect 401138 -19888 401194 -19832
rect 401262 -19888 401318 -19832
rect 400766 -20012 400822 -19956
rect 400890 -20012 400946 -19956
rect 401014 -20012 401070 -19956
rect 401138 -20012 401194 -19956
rect 401262 -20012 401318 -19956
rect 400766 -20136 400822 -20080
rect 400890 -20136 400946 -20080
rect 401014 -20136 401070 -20080
rect 401138 -20136 401194 -20080
rect 401262 -20136 401318 -20080
rect 400766 -20260 400822 -20204
rect 400890 -20260 400946 -20204
rect 401014 -20260 401070 -20204
rect 401138 -20260 401194 -20204
rect 401262 -20260 401318 -20204
rect 400766 -20384 400822 -20328
rect 400890 -20384 400946 -20328
rect 401014 -20384 401070 -20328
rect 401138 -20384 401194 -20328
rect 401262 -20384 401318 -20328
rect 400766 -20508 400822 -20452
rect 400890 -20508 400946 -20452
rect 401014 -20508 401070 -20452
rect 401138 -20508 401194 -20452
rect 401262 -20508 401318 -20452
rect 400766 -20632 400822 -20576
rect 400890 -20632 400946 -20576
rect 401014 -20632 401070 -20576
rect 401138 -20632 401194 -20576
rect 401262 -20632 401318 -20576
rect 400766 -20756 400822 -20700
rect 400890 -20756 400946 -20700
rect 401014 -20756 401070 -20700
rect 401138 -20756 401194 -20700
rect 401262 -20756 401318 -20700
rect 400766 -20880 400822 -20824
rect 400890 -20880 400946 -20824
rect 401014 -20880 401070 -20824
rect 401138 -20880 401194 -20824
rect 401262 -20880 401318 -20824
rect 400766 -21004 400822 -20948
rect 400890 -21004 400946 -20948
rect 401014 -21004 401070 -20948
rect 401138 -21004 401194 -20948
rect 401262 -21004 401318 -20948
rect 400766 -21128 400822 -21072
rect 400890 -21128 400946 -21072
rect 401014 -21128 401070 -21072
rect 401138 -21128 401194 -21072
rect 401262 -21128 401318 -21072
rect 400766 -21252 400822 -21196
rect 400890 -21252 400946 -21196
rect 401014 -21252 401070 -21196
rect 401138 -21252 401194 -21196
rect 401262 -21252 401318 -21196
rect 400766 -21376 400822 -21320
rect 400890 -21376 400946 -21320
rect 401014 -21376 401070 -21320
rect 401138 -21376 401194 -21320
rect 401262 -21376 401318 -21320
rect 400766 -21500 400822 -21444
rect 400890 -21500 400946 -21444
rect 401014 -21500 401070 -21444
rect 401138 -21500 401194 -21444
rect 401262 -21500 401318 -21444
rect 400766 -21624 400822 -21568
rect 400890 -21624 400946 -21568
rect 401014 -21624 401070 -21568
rect 401138 -21624 401194 -21568
rect 401262 -21624 401318 -21568
rect 400766 -21748 400822 -21692
rect 400890 -21748 400946 -21692
rect 401014 -21748 401070 -21692
rect 401138 -21748 401194 -21692
rect 401262 -21748 401318 -21692
rect 400766 -21872 400822 -21816
rect 400890 -21872 400946 -21816
rect 401014 -21872 401070 -21816
rect 401138 -21872 401194 -21816
rect 401262 -21872 401318 -21816
rect 400766 -21996 400822 -21940
rect 400890 -21996 400946 -21940
rect 401014 -21996 401070 -21940
rect 401138 -21996 401194 -21940
rect 401262 -21996 401318 -21940
rect 400766 -22120 400822 -22064
rect 400890 -22120 400946 -22064
rect 401014 -22120 401070 -22064
rect 401138 -22120 401194 -22064
rect 401262 -22120 401318 -22064
rect 400766 -22244 400822 -22188
rect 400890 -22244 400946 -22188
rect 401014 -22244 401070 -22188
rect 401138 -22244 401194 -22188
rect 401262 -22244 401318 -22188
rect 400766 -22368 400822 -22312
rect 400890 -22368 400946 -22312
rect 401014 -22368 401070 -22312
rect 401138 -22368 401194 -22312
rect 401262 -22368 401318 -22312
rect 400766 -22492 400822 -22436
rect 400890 -22492 400946 -22436
rect 401014 -22492 401070 -22436
rect 401138 -22492 401194 -22436
rect 401262 -22492 401318 -22436
rect 400766 -22616 400822 -22560
rect 400890 -22616 400946 -22560
rect 401014 -22616 401070 -22560
rect 401138 -22616 401194 -22560
rect 401262 -22616 401318 -22560
rect 400766 -22740 400822 -22684
rect 400890 -22740 400946 -22684
rect 401014 -22740 401070 -22684
rect 401138 -22740 401194 -22684
rect 401262 -22740 401318 -22684
rect 400766 -22864 400822 -22808
rect 400890 -22864 400946 -22808
rect 401014 -22864 401070 -22808
rect 401138 -22864 401194 -22808
rect 401262 -22864 401318 -22808
rect 400766 -22988 400822 -22932
rect 400890 -22988 400946 -22932
rect 401014 -22988 401070 -22932
rect 401138 -22988 401194 -22932
rect 401262 -22988 401318 -22932
rect 400766 -23112 400822 -23056
rect 400890 -23112 400946 -23056
rect 401014 -23112 401070 -23056
rect 401138 -23112 401194 -23056
rect 401262 -23112 401318 -23056
rect 400766 -23236 400822 -23180
rect 400890 -23236 400946 -23180
rect 401014 -23236 401070 -23180
rect 401138 -23236 401194 -23180
rect 401262 -23236 401318 -23180
rect 400766 -23360 400822 -23304
rect 400890 -23360 400946 -23304
rect 401014 -23360 401070 -23304
rect 401138 -23360 401194 -23304
rect 401262 -23360 401318 -23304
rect 400766 -23484 400822 -23428
rect 400890 -23484 400946 -23428
rect 401014 -23484 401070 -23428
rect 401138 -23484 401194 -23428
rect 401262 -23484 401318 -23428
rect 400766 -23608 400822 -23552
rect 400890 -23608 400946 -23552
rect 401014 -23608 401070 -23552
rect 401138 -23608 401194 -23552
rect 401262 -23608 401318 -23552
rect 400766 -23732 400822 -23676
rect 400890 -23732 400946 -23676
rect 401014 -23732 401070 -23676
rect 401138 -23732 401194 -23676
rect 401262 -23732 401318 -23676
rect 400766 -23856 400822 -23800
rect 400890 -23856 400946 -23800
rect 401014 -23856 401070 -23800
rect 401138 -23856 401194 -23800
rect 401262 -23856 401318 -23800
rect 400766 -23980 400822 -23924
rect 400890 -23980 400946 -23924
rect 401014 -23980 401070 -23924
rect 401138 -23980 401194 -23924
rect 401262 -23980 401318 -23924
rect 400766 -24104 400822 -24048
rect 400890 -24104 400946 -24048
rect 401014 -24104 401070 -24048
rect 401138 -24104 401194 -24048
rect 401262 -24104 401318 -24048
rect 400766 -24228 400822 -24172
rect 400890 -24228 400946 -24172
rect 401014 -24228 401070 -24172
rect 401138 -24228 401194 -24172
rect 401262 -24228 401318 -24172
rect 400766 -24352 400822 -24296
rect 400890 -24352 400946 -24296
rect 401014 -24352 401070 -24296
rect 401138 -24352 401194 -24296
rect 401262 -24352 401318 -24296
rect 400766 -24476 400822 -24420
rect 400890 -24476 400946 -24420
rect 401014 -24476 401070 -24420
rect 401138 -24476 401194 -24420
rect 401262 -24476 401318 -24420
rect 400766 -24600 400822 -24544
rect 400890 -24600 400946 -24544
rect 401014 -24600 401070 -24544
rect 401138 -24600 401194 -24544
rect 401262 -24600 401318 -24544
rect 400766 -24724 400822 -24668
rect 400890 -24724 400946 -24668
rect 401014 -24724 401070 -24668
rect 401138 -24724 401194 -24668
rect 401262 -24724 401318 -24668
rect 400766 -24848 400822 -24792
rect 400890 -24848 400946 -24792
rect 401014 -24848 401070 -24792
rect 401138 -24848 401194 -24792
rect 401262 -24848 401318 -24792
rect 400766 -24972 400822 -24916
rect 400890 -24972 400946 -24916
rect 401014 -24972 401070 -24916
rect 401138 -24972 401194 -24916
rect 401262 -24972 401318 -24916
rect 400766 -25096 400822 -25040
rect 400890 -25096 400946 -25040
rect 401014 -25096 401070 -25040
rect 401138 -25096 401194 -25040
rect 401262 -25096 401318 -25040
rect 400766 -25220 400822 -25164
rect 400890 -25220 400946 -25164
rect 401014 -25220 401070 -25164
rect 401138 -25220 401194 -25164
rect 401262 -25220 401318 -25164
rect 400766 -25344 400822 -25288
rect 400890 -25344 400946 -25288
rect 401014 -25344 401070 -25288
rect 401138 -25344 401194 -25288
rect 401262 -25344 401318 -25288
rect 400766 -25468 400822 -25412
rect 400890 -25468 400946 -25412
rect 401014 -25468 401070 -25412
rect 401138 -25468 401194 -25412
rect 401262 -25468 401318 -25412
rect 387954 -25592 388010 -25536
rect 388078 -25592 388134 -25536
rect 388202 -25592 388258 -25536
rect 388326 -25592 388382 -25536
rect 388450 -25592 388506 -25536
rect 400766 -25592 400822 -25536
rect 400890 -25592 400946 -25536
rect 401014 -25592 401070 -25536
rect 401138 -25592 401194 -25536
rect 401262 -25592 401318 -25536
rect 387954 -25716 388010 -25660
rect 388078 -25716 388134 -25660
rect 388202 -25716 388258 -25660
rect 388326 -25716 388382 -25660
rect 388450 -25716 388506 -25660
rect 388655 -25744 388711 -25688
rect 388797 -25744 388853 -25688
rect 388939 -25744 388995 -25688
rect 389081 -25744 389137 -25688
rect 389223 -25744 389279 -25688
rect 389365 -25744 389421 -25688
rect 389507 -25744 389563 -25688
rect 389649 -25744 389705 -25688
rect 389791 -25744 389847 -25688
rect 389933 -25744 389989 -25688
rect 390075 -25744 390131 -25688
rect 390217 -25744 390273 -25688
rect 390359 -25744 390415 -25688
rect 390501 -25744 390557 -25688
rect 390643 -25744 390699 -25688
rect 390785 -25744 390841 -25688
rect 390927 -25744 390983 -25688
rect 391069 -25744 391125 -25688
rect 391211 -25744 391267 -25688
rect 391353 -25744 391409 -25688
rect 391495 -25744 391551 -25688
rect 391637 -25744 391693 -25688
rect 391779 -25744 391835 -25688
rect 391921 -25744 391977 -25688
rect 392063 -25744 392119 -25688
rect 392205 -25744 392261 -25688
rect 392347 -25744 392403 -25688
rect 392489 -25744 392545 -25688
rect 392631 -25744 392687 -25688
rect 392773 -25744 392829 -25688
rect 392915 -25744 392971 -25688
rect 393057 -25744 393113 -25688
rect 393199 -25744 393255 -25688
rect 393341 -25744 393397 -25688
rect 393483 -25744 393539 -25688
rect 393625 -25744 393681 -25688
rect 393767 -25744 393823 -25688
rect 393909 -25744 393965 -25688
rect 394051 -25744 394107 -25688
rect 394193 -25744 394249 -25688
rect 394335 -25744 394391 -25688
rect 394477 -25744 394533 -25688
rect 394619 -25744 394675 -25688
rect 394761 -25744 394817 -25688
rect 394903 -25744 394959 -25688
rect 395045 -25744 395101 -25688
rect 395187 -25744 395243 -25688
rect 395329 -25744 395385 -25688
rect 395471 -25744 395527 -25688
rect 395613 -25744 395669 -25688
rect 395755 -25744 395811 -25688
rect 395897 -25744 395953 -25688
rect 396039 -25744 396095 -25688
rect 396181 -25744 396237 -25688
rect 396323 -25744 396379 -25688
rect 396465 -25744 396521 -25688
rect 396607 -25744 396663 -25688
rect 396749 -25744 396805 -25688
rect 396891 -25744 396947 -25688
rect 397033 -25744 397089 -25688
rect 397175 -25744 397231 -25688
rect 397317 -25744 397373 -25688
rect 397459 -25744 397515 -25688
rect 397601 -25744 397657 -25688
rect 397743 -25744 397799 -25688
rect 397885 -25744 397941 -25688
rect 398027 -25744 398083 -25688
rect 398169 -25744 398225 -25688
rect 398311 -25744 398367 -25688
rect 398453 -25744 398509 -25688
rect 398595 -25744 398651 -25688
rect 398737 -25744 398793 -25688
rect 398879 -25744 398935 -25688
rect 399021 -25744 399077 -25688
rect 399163 -25744 399219 -25688
rect 399305 -25744 399361 -25688
rect 399447 -25744 399503 -25688
rect 399589 -25744 399645 -25688
rect 399731 -25744 399787 -25688
rect 399873 -25744 399929 -25688
rect 400015 -25744 400071 -25688
rect 400157 -25744 400213 -25688
rect 400299 -25744 400355 -25688
rect 400441 -25744 400497 -25688
rect 400583 -25744 400639 -25688
rect 400766 -25716 400822 -25660
rect 400890 -25716 400946 -25660
rect 401014 -25716 401070 -25660
rect 401138 -25716 401194 -25660
rect 401262 -25716 401318 -25660
rect 387954 -25840 388010 -25784
rect 388078 -25840 388134 -25784
rect 388202 -25840 388258 -25784
rect 388326 -25840 388382 -25784
rect 388450 -25840 388506 -25784
rect 388655 -25886 388711 -25830
rect 388797 -25886 388853 -25830
rect 388939 -25886 388995 -25830
rect 389081 -25886 389137 -25830
rect 389223 -25886 389279 -25830
rect 389365 -25886 389421 -25830
rect 389507 -25886 389563 -25830
rect 389649 -25886 389705 -25830
rect 389791 -25886 389847 -25830
rect 389933 -25886 389989 -25830
rect 390075 -25886 390131 -25830
rect 390217 -25886 390273 -25830
rect 390359 -25886 390415 -25830
rect 390501 -25886 390557 -25830
rect 390643 -25886 390699 -25830
rect 390785 -25886 390841 -25830
rect 390927 -25886 390983 -25830
rect 391069 -25886 391125 -25830
rect 391211 -25886 391267 -25830
rect 391353 -25886 391409 -25830
rect 391495 -25886 391551 -25830
rect 391637 -25886 391693 -25830
rect 391779 -25886 391835 -25830
rect 391921 -25886 391977 -25830
rect 392063 -25886 392119 -25830
rect 392205 -25886 392261 -25830
rect 392347 -25886 392403 -25830
rect 392489 -25886 392545 -25830
rect 392631 -25886 392687 -25830
rect 392773 -25886 392829 -25830
rect 392915 -25886 392971 -25830
rect 393057 -25886 393113 -25830
rect 393199 -25886 393255 -25830
rect 393341 -25886 393397 -25830
rect 393483 -25886 393539 -25830
rect 393625 -25886 393681 -25830
rect 393767 -25886 393823 -25830
rect 393909 -25886 393965 -25830
rect 394051 -25886 394107 -25830
rect 394193 -25886 394249 -25830
rect 394335 -25886 394391 -25830
rect 394477 -25886 394533 -25830
rect 394619 -25886 394675 -25830
rect 394761 -25886 394817 -25830
rect 394903 -25886 394959 -25830
rect 395045 -25886 395101 -25830
rect 395187 -25886 395243 -25830
rect 395329 -25886 395385 -25830
rect 395471 -25886 395527 -25830
rect 395613 -25886 395669 -25830
rect 395755 -25886 395811 -25830
rect 395897 -25886 395953 -25830
rect 396039 -25886 396095 -25830
rect 396181 -25886 396237 -25830
rect 396323 -25886 396379 -25830
rect 396465 -25886 396521 -25830
rect 396607 -25886 396663 -25830
rect 396749 -25886 396805 -25830
rect 396891 -25886 396947 -25830
rect 397033 -25886 397089 -25830
rect 397175 -25886 397231 -25830
rect 397317 -25886 397373 -25830
rect 397459 -25886 397515 -25830
rect 397601 -25886 397657 -25830
rect 397743 -25886 397799 -25830
rect 397885 -25886 397941 -25830
rect 398027 -25886 398083 -25830
rect 398169 -25886 398225 -25830
rect 398311 -25886 398367 -25830
rect 398453 -25886 398509 -25830
rect 398595 -25886 398651 -25830
rect 398737 -25886 398793 -25830
rect 398879 -25886 398935 -25830
rect 399021 -25886 399077 -25830
rect 399163 -25886 399219 -25830
rect 399305 -25886 399361 -25830
rect 399447 -25886 399503 -25830
rect 399589 -25886 399645 -25830
rect 399731 -25886 399787 -25830
rect 399873 -25886 399929 -25830
rect 400015 -25886 400071 -25830
rect 400157 -25886 400213 -25830
rect 400299 -25886 400355 -25830
rect 400441 -25886 400497 -25830
rect 400583 -25886 400639 -25830
rect 400766 -25840 400822 -25784
rect 400890 -25840 400946 -25784
rect 401014 -25840 401070 -25784
rect 401138 -25840 401194 -25784
rect 401262 -25840 401318 -25784
<< metal5 >>
rect 387840 -13041 401440 -12925
rect 387840 -13097 387986 -13041
rect 388042 -13097 388110 -13041
rect 388166 -13097 388234 -13041
rect 388290 -13097 388358 -13041
rect 388414 -13097 388482 -13041
rect 388538 -13097 388606 -13041
rect 388662 -13097 388730 -13041
rect 388786 -13097 388854 -13041
rect 388910 -13097 388978 -13041
rect 389034 -13097 389102 -13041
rect 389158 -13097 389226 -13041
rect 389282 -13097 389350 -13041
rect 389406 -13097 389474 -13041
rect 389530 -13097 389598 -13041
rect 389654 -13097 389722 -13041
rect 389778 -13097 389846 -13041
rect 389902 -13097 389970 -13041
rect 390026 -13097 390094 -13041
rect 390150 -13097 390218 -13041
rect 390274 -13097 390342 -13041
rect 390398 -13097 390466 -13041
rect 390522 -13097 390590 -13041
rect 390646 -13097 390714 -13041
rect 390770 -13097 390838 -13041
rect 390894 -13097 390962 -13041
rect 391018 -13097 391086 -13041
rect 391142 -13097 391210 -13041
rect 391266 -13097 391334 -13041
rect 391390 -13097 391458 -13041
rect 391514 -13097 391582 -13041
rect 391638 -13097 391706 -13041
rect 391762 -13097 391830 -13041
rect 391886 -13097 391954 -13041
rect 392010 -13097 392078 -13041
rect 392134 -13097 392202 -13041
rect 392258 -13097 392326 -13041
rect 392382 -13097 392450 -13041
rect 392506 -13097 392574 -13041
rect 392630 -13097 392698 -13041
rect 392754 -13097 392822 -13041
rect 392878 -13097 392946 -13041
rect 393002 -13097 393070 -13041
rect 393126 -13097 393194 -13041
rect 393250 -13097 393318 -13041
rect 393374 -13097 393442 -13041
rect 393498 -13097 393566 -13041
rect 393622 -13097 393690 -13041
rect 393746 -13097 393814 -13041
rect 393870 -13097 393938 -13041
rect 393994 -13097 394062 -13041
rect 394118 -13097 394186 -13041
rect 394242 -13097 394310 -13041
rect 394366 -13097 394434 -13041
rect 394490 -13097 394558 -13041
rect 394614 -13097 394682 -13041
rect 394738 -13097 394806 -13041
rect 394862 -13097 394930 -13041
rect 394986 -13097 395054 -13041
rect 395110 -13097 395178 -13041
rect 395234 -13097 395302 -13041
rect 395358 -13097 395426 -13041
rect 395482 -13097 395550 -13041
rect 395606 -13097 395674 -13041
rect 395730 -13097 395798 -13041
rect 395854 -13097 395922 -13041
rect 395978 -13097 396046 -13041
rect 396102 -13097 396170 -13041
rect 396226 -13097 396294 -13041
rect 396350 -13097 396418 -13041
rect 396474 -13097 396542 -13041
rect 396598 -13097 396666 -13041
rect 396722 -13097 396790 -13041
rect 396846 -13097 396914 -13041
rect 396970 -13097 397038 -13041
rect 397094 -13097 397162 -13041
rect 397218 -13097 397286 -13041
rect 397342 -13097 397410 -13041
rect 397466 -13097 397534 -13041
rect 397590 -13097 397658 -13041
rect 397714 -13097 397782 -13041
rect 397838 -13097 397906 -13041
rect 397962 -13097 398030 -13041
rect 398086 -13097 398154 -13041
rect 398210 -13097 398278 -13041
rect 398334 -13097 398402 -13041
rect 398458 -13097 398526 -13041
rect 398582 -13097 398650 -13041
rect 398706 -13097 398774 -13041
rect 398830 -13097 398898 -13041
rect 398954 -13097 399022 -13041
rect 399078 -13097 399146 -13041
rect 399202 -13097 399270 -13041
rect 399326 -13097 399394 -13041
rect 399450 -13097 399518 -13041
rect 399574 -13097 399642 -13041
rect 399698 -13097 399766 -13041
rect 399822 -13097 399890 -13041
rect 399946 -13097 400014 -13041
rect 400070 -13097 400138 -13041
rect 400194 -13097 400262 -13041
rect 400318 -13097 400386 -13041
rect 400442 -13097 400510 -13041
rect 400566 -13097 400634 -13041
rect 400690 -13097 400758 -13041
rect 400814 -13097 400882 -13041
rect 400938 -13097 401006 -13041
rect 401062 -13097 401130 -13041
rect 401186 -13097 401254 -13041
rect 401310 -13097 401440 -13041
rect 387840 -13165 401440 -13097
rect 387840 -13221 387986 -13165
rect 388042 -13221 388110 -13165
rect 388166 -13221 388234 -13165
rect 388290 -13221 388358 -13165
rect 388414 -13221 388482 -13165
rect 388538 -13221 388606 -13165
rect 388662 -13221 388730 -13165
rect 388786 -13221 388854 -13165
rect 388910 -13221 388978 -13165
rect 389034 -13221 389102 -13165
rect 389158 -13221 389226 -13165
rect 389282 -13221 389350 -13165
rect 389406 -13221 389474 -13165
rect 389530 -13221 389598 -13165
rect 389654 -13221 389722 -13165
rect 389778 -13221 389846 -13165
rect 389902 -13221 389970 -13165
rect 390026 -13221 390094 -13165
rect 390150 -13221 390218 -13165
rect 390274 -13221 390342 -13165
rect 390398 -13221 390466 -13165
rect 390522 -13221 390590 -13165
rect 390646 -13221 390714 -13165
rect 390770 -13221 390838 -13165
rect 390894 -13221 390962 -13165
rect 391018 -13221 391086 -13165
rect 391142 -13221 391210 -13165
rect 391266 -13221 391334 -13165
rect 391390 -13221 391458 -13165
rect 391514 -13221 391582 -13165
rect 391638 -13221 391706 -13165
rect 391762 -13221 391830 -13165
rect 391886 -13221 391954 -13165
rect 392010 -13221 392078 -13165
rect 392134 -13221 392202 -13165
rect 392258 -13221 392326 -13165
rect 392382 -13221 392450 -13165
rect 392506 -13221 392574 -13165
rect 392630 -13221 392698 -13165
rect 392754 -13221 392822 -13165
rect 392878 -13221 392946 -13165
rect 393002 -13221 393070 -13165
rect 393126 -13221 393194 -13165
rect 393250 -13221 393318 -13165
rect 393374 -13221 393442 -13165
rect 393498 -13221 393566 -13165
rect 393622 -13221 393690 -13165
rect 393746 -13221 393814 -13165
rect 393870 -13221 393938 -13165
rect 393994 -13221 394062 -13165
rect 394118 -13221 394186 -13165
rect 394242 -13221 394310 -13165
rect 394366 -13221 394434 -13165
rect 394490 -13221 394558 -13165
rect 394614 -13221 394682 -13165
rect 394738 -13221 394806 -13165
rect 394862 -13221 394930 -13165
rect 394986 -13221 395054 -13165
rect 395110 -13221 395178 -13165
rect 395234 -13221 395302 -13165
rect 395358 -13221 395426 -13165
rect 395482 -13221 395550 -13165
rect 395606 -13221 395674 -13165
rect 395730 -13221 395798 -13165
rect 395854 -13221 395922 -13165
rect 395978 -13221 396046 -13165
rect 396102 -13221 396170 -13165
rect 396226 -13221 396294 -13165
rect 396350 -13221 396418 -13165
rect 396474 -13221 396542 -13165
rect 396598 -13221 396666 -13165
rect 396722 -13221 396790 -13165
rect 396846 -13221 396914 -13165
rect 396970 -13221 397038 -13165
rect 397094 -13221 397162 -13165
rect 397218 -13221 397286 -13165
rect 397342 -13221 397410 -13165
rect 397466 -13221 397534 -13165
rect 397590 -13221 397658 -13165
rect 397714 -13221 397782 -13165
rect 397838 -13221 397906 -13165
rect 397962 -13221 398030 -13165
rect 398086 -13221 398154 -13165
rect 398210 -13221 398278 -13165
rect 398334 -13221 398402 -13165
rect 398458 -13221 398526 -13165
rect 398582 -13221 398650 -13165
rect 398706 -13221 398774 -13165
rect 398830 -13221 398898 -13165
rect 398954 -13221 399022 -13165
rect 399078 -13221 399146 -13165
rect 399202 -13221 399270 -13165
rect 399326 -13221 399394 -13165
rect 399450 -13221 399518 -13165
rect 399574 -13221 399642 -13165
rect 399698 -13221 399766 -13165
rect 399822 -13221 399890 -13165
rect 399946 -13221 400014 -13165
rect 400070 -13221 400138 -13165
rect 400194 -13221 400262 -13165
rect 400318 -13221 400386 -13165
rect 400442 -13221 400510 -13165
rect 400566 -13221 400634 -13165
rect 400690 -13221 400758 -13165
rect 400814 -13221 400882 -13165
rect 400938 -13221 401006 -13165
rect 401062 -13221 401130 -13165
rect 401186 -13221 401254 -13165
rect 401310 -13221 401440 -13165
rect 387840 -13289 401440 -13221
rect 387840 -13345 387986 -13289
rect 388042 -13345 388110 -13289
rect 388166 -13345 388234 -13289
rect 388290 -13345 388358 -13289
rect 388414 -13345 388482 -13289
rect 388538 -13345 388606 -13289
rect 388662 -13345 388730 -13289
rect 388786 -13345 388854 -13289
rect 388910 -13345 388978 -13289
rect 389034 -13345 389102 -13289
rect 389158 -13345 389226 -13289
rect 389282 -13345 389350 -13289
rect 389406 -13345 389474 -13289
rect 389530 -13345 389598 -13289
rect 389654 -13345 389722 -13289
rect 389778 -13345 389846 -13289
rect 389902 -13345 389970 -13289
rect 390026 -13345 390094 -13289
rect 390150 -13345 390218 -13289
rect 390274 -13345 390342 -13289
rect 390398 -13345 390466 -13289
rect 390522 -13345 390590 -13289
rect 390646 -13345 390714 -13289
rect 390770 -13345 390838 -13289
rect 390894 -13345 390962 -13289
rect 391018 -13345 391086 -13289
rect 391142 -13345 391210 -13289
rect 391266 -13345 391334 -13289
rect 391390 -13345 391458 -13289
rect 391514 -13345 391582 -13289
rect 391638 -13345 391706 -13289
rect 391762 -13345 391830 -13289
rect 391886 -13345 391954 -13289
rect 392010 -13345 392078 -13289
rect 392134 -13345 392202 -13289
rect 392258 -13345 392326 -13289
rect 392382 -13345 392450 -13289
rect 392506 -13345 392574 -13289
rect 392630 -13345 392698 -13289
rect 392754 -13345 392822 -13289
rect 392878 -13345 392946 -13289
rect 393002 -13345 393070 -13289
rect 393126 -13345 393194 -13289
rect 393250 -13345 393318 -13289
rect 393374 -13345 393442 -13289
rect 393498 -13345 393566 -13289
rect 393622 -13345 393690 -13289
rect 393746 -13345 393814 -13289
rect 393870 -13345 393938 -13289
rect 393994 -13345 394062 -13289
rect 394118 -13345 394186 -13289
rect 394242 -13345 394310 -13289
rect 394366 -13345 394434 -13289
rect 394490 -13345 394558 -13289
rect 394614 -13345 394682 -13289
rect 394738 -13345 394806 -13289
rect 394862 -13345 394930 -13289
rect 394986 -13345 395054 -13289
rect 395110 -13345 395178 -13289
rect 395234 -13345 395302 -13289
rect 395358 -13345 395426 -13289
rect 395482 -13345 395550 -13289
rect 395606 -13345 395674 -13289
rect 395730 -13345 395798 -13289
rect 395854 -13345 395922 -13289
rect 395978 -13345 396046 -13289
rect 396102 -13345 396170 -13289
rect 396226 -13345 396294 -13289
rect 396350 -13345 396418 -13289
rect 396474 -13345 396542 -13289
rect 396598 -13345 396666 -13289
rect 396722 -13345 396790 -13289
rect 396846 -13345 396914 -13289
rect 396970 -13345 397038 -13289
rect 397094 -13345 397162 -13289
rect 397218 -13345 397286 -13289
rect 397342 -13345 397410 -13289
rect 397466 -13345 397534 -13289
rect 397590 -13345 397658 -13289
rect 397714 -13345 397782 -13289
rect 397838 -13345 397906 -13289
rect 397962 -13345 398030 -13289
rect 398086 -13345 398154 -13289
rect 398210 -13345 398278 -13289
rect 398334 -13345 398402 -13289
rect 398458 -13345 398526 -13289
rect 398582 -13345 398650 -13289
rect 398706 -13345 398774 -13289
rect 398830 -13345 398898 -13289
rect 398954 -13345 399022 -13289
rect 399078 -13345 399146 -13289
rect 399202 -13345 399270 -13289
rect 399326 -13345 399394 -13289
rect 399450 -13345 399518 -13289
rect 399574 -13345 399642 -13289
rect 399698 -13345 399766 -13289
rect 399822 -13345 399890 -13289
rect 399946 -13345 400014 -13289
rect 400070 -13345 400138 -13289
rect 400194 -13345 400262 -13289
rect 400318 -13345 400386 -13289
rect 400442 -13345 400510 -13289
rect 400566 -13345 400634 -13289
rect 400690 -13345 400758 -13289
rect 400814 -13345 400882 -13289
rect 400938 -13345 401006 -13289
rect 401062 -13345 401130 -13289
rect 401186 -13345 401254 -13289
rect 401310 -13345 401440 -13289
rect 387840 -13413 401440 -13345
rect 387840 -13469 387986 -13413
rect 388042 -13469 388110 -13413
rect 388166 -13469 388234 -13413
rect 388290 -13469 388358 -13413
rect 388414 -13469 388482 -13413
rect 388538 -13469 388606 -13413
rect 388662 -13469 388730 -13413
rect 388786 -13469 388854 -13413
rect 388910 -13469 388978 -13413
rect 389034 -13469 389102 -13413
rect 389158 -13469 389226 -13413
rect 389282 -13469 389350 -13413
rect 389406 -13469 389474 -13413
rect 389530 -13469 389598 -13413
rect 389654 -13469 389722 -13413
rect 389778 -13469 389846 -13413
rect 389902 -13469 389970 -13413
rect 390026 -13469 390094 -13413
rect 390150 -13469 390218 -13413
rect 390274 -13469 390342 -13413
rect 390398 -13469 390466 -13413
rect 390522 -13469 390590 -13413
rect 390646 -13469 390714 -13413
rect 390770 -13469 390838 -13413
rect 390894 -13469 390962 -13413
rect 391018 -13469 391086 -13413
rect 391142 -13469 391210 -13413
rect 391266 -13469 391334 -13413
rect 391390 -13469 391458 -13413
rect 391514 -13469 391582 -13413
rect 391638 -13469 391706 -13413
rect 391762 -13469 391830 -13413
rect 391886 -13469 391954 -13413
rect 392010 -13469 392078 -13413
rect 392134 -13469 392202 -13413
rect 392258 -13469 392326 -13413
rect 392382 -13469 392450 -13413
rect 392506 -13469 392574 -13413
rect 392630 -13469 392698 -13413
rect 392754 -13469 392822 -13413
rect 392878 -13469 392946 -13413
rect 393002 -13469 393070 -13413
rect 393126 -13469 393194 -13413
rect 393250 -13469 393318 -13413
rect 393374 -13469 393442 -13413
rect 393498 -13469 393566 -13413
rect 393622 -13469 393690 -13413
rect 393746 -13469 393814 -13413
rect 393870 -13469 393938 -13413
rect 393994 -13469 394062 -13413
rect 394118 -13469 394186 -13413
rect 394242 -13469 394310 -13413
rect 394366 -13469 394434 -13413
rect 394490 -13469 394558 -13413
rect 394614 -13469 394682 -13413
rect 394738 -13469 394806 -13413
rect 394862 -13469 394930 -13413
rect 394986 -13469 395054 -13413
rect 395110 -13469 395178 -13413
rect 395234 -13469 395302 -13413
rect 395358 -13469 395426 -13413
rect 395482 -13469 395550 -13413
rect 395606 -13469 395674 -13413
rect 395730 -13469 395798 -13413
rect 395854 -13469 395922 -13413
rect 395978 -13469 396046 -13413
rect 396102 -13469 396170 -13413
rect 396226 -13469 396294 -13413
rect 396350 -13469 396418 -13413
rect 396474 -13469 396542 -13413
rect 396598 -13469 396666 -13413
rect 396722 -13469 396790 -13413
rect 396846 -13469 396914 -13413
rect 396970 -13469 397038 -13413
rect 397094 -13469 397162 -13413
rect 397218 -13469 397286 -13413
rect 397342 -13469 397410 -13413
rect 397466 -13469 397534 -13413
rect 397590 -13469 397658 -13413
rect 397714 -13469 397782 -13413
rect 397838 -13469 397906 -13413
rect 397962 -13469 398030 -13413
rect 398086 -13469 398154 -13413
rect 398210 -13469 398278 -13413
rect 398334 -13469 398402 -13413
rect 398458 -13469 398526 -13413
rect 398582 -13469 398650 -13413
rect 398706 -13469 398774 -13413
rect 398830 -13469 398898 -13413
rect 398954 -13469 399022 -13413
rect 399078 -13469 399146 -13413
rect 399202 -13469 399270 -13413
rect 399326 -13469 399394 -13413
rect 399450 -13469 399518 -13413
rect 399574 -13469 399642 -13413
rect 399698 -13469 399766 -13413
rect 399822 -13469 399890 -13413
rect 399946 -13469 400014 -13413
rect 400070 -13469 400138 -13413
rect 400194 -13469 400262 -13413
rect 400318 -13469 400386 -13413
rect 400442 -13469 400510 -13413
rect 400566 -13469 400634 -13413
rect 400690 -13469 400758 -13413
rect 400814 -13469 400882 -13413
rect 400938 -13469 401006 -13413
rect 401062 -13469 401130 -13413
rect 401186 -13469 401254 -13413
rect 401310 -13469 401440 -13413
rect 387840 -13590 401440 -13469
rect 387840 -13632 402640 -13590
rect 387840 -13688 387954 -13632
rect 388010 -13688 388078 -13632
rect 388134 -13688 388202 -13632
rect 388258 -13688 388326 -13632
rect 388382 -13688 388450 -13632
rect 388506 -13680 400766 -13632
rect 388506 -13688 388981 -13680
rect 387840 -13736 388981 -13688
rect 389037 -13736 389123 -13680
rect 389179 -13736 389382 -13680
rect 389438 -13736 389524 -13680
rect 389580 -13736 389782 -13680
rect 389838 -13736 389924 -13680
rect 389980 -13736 390179 -13680
rect 390235 -13736 390321 -13680
rect 390377 -13736 390576 -13680
rect 390632 -13736 390718 -13680
rect 390774 -13736 390980 -13680
rect 391036 -13736 391122 -13680
rect 391178 -13736 391376 -13680
rect 391432 -13736 391518 -13680
rect 391574 -13736 391776 -13680
rect 391832 -13736 391918 -13680
rect 391974 -13736 392173 -13680
rect 392229 -13736 392315 -13680
rect 392371 -13736 392578 -13680
rect 392634 -13736 392720 -13680
rect 392776 -13736 392978 -13680
rect 393034 -13736 393120 -13680
rect 393176 -13736 393383 -13680
rect 393439 -13736 393525 -13680
rect 393581 -13736 393780 -13680
rect 393836 -13736 393922 -13680
rect 393978 -13736 394177 -13680
rect 394233 -13736 394319 -13680
rect 394375 -13736 394580 -13680
rect 394636 -13736 394722 -13680
rect 394778 -13736 394982 -13680
rect 395038 -13736 395124 -13680
rect 395180 -13736 395385 -13680
rect 395441 -13736 395527 -13680
rect 395583 -13736 395779 -13680
rect 395835 -13736 395921 -13680
rect 395977 -13736 396180 -13680
rect 396236 -13736 396322 -13680
rect 396378 -13736 396580 -13680
rect 396636 -13736 396722 -13680
rect 396778 -13736 396977 -13680
rect 397033 -13736 397119 -13680
rect 397175 -13736 397374 -13680
rect 397430 -13736 397516 -13680
rect 397572 -13736 397778 -13680
rect 397834 -13736 397920 -13680
rect 397976 -13736 398174 -13680
rect 398230 -13736 398316 -13680
rect 398372 -13736 398574 -13680
rect 398630 -13736 398716 -13680
rect 398772 -13736 398971 -13680
rect 399027 -13736 399113 -13680
rect 399169 -13736 399376 -13680
rect 399432 -13736 399518 -13680
rect 399574 -13736 399776 -13680
rect 399832 -13736 399918 -13680
rect 399974 -13736 400181 -13680
rect 400237 -13736 400323 -13680
rect 400379 -13688 400766 -13680
rect 400822 -13688 400890 -13632
rect 400946 -13688 401014 -13632
rect 401070 -13688 401138 -13632
rect 401194 -13688 401262 -13632
rect 401318 -13688 402640 -13632
rect 400379 -13736 402640 -13688
rect 387840 -13756 402640 -13736
rect 387840 -13812 387954 -13756
rect 388010 -13812 388078 -13756
rect 388134 -13812 388202 -13756
rect 388258 -13812 388326 -13756
rect 388382 -13812 388450 -13756
rect 388506 -13812 400766 -13756
rect 400822 -13812 400890 -13756
rect 400946 -13812 401014 -13756
rect 401070 -13812 401138 -13756
rect 401194 -13812 401262 -13756
rect 401318 -13812 402640 -13756
rect 387840 -13822 402640 -13812
rect 387840 -13878 388981 -13822
rect 389037 -13878 389123 -13822
rect 389179 -13878 389382 -13822
rect 389438 -13878 389524 -13822
rect 389580 -13878 389782 -13822
rect 389838 -13878 389924 -13822
rect 389980 -13878 390179 -13822
rect 390235 -13878 390321 -13822
rect 390377 -13878 390576 -13822
rect 390632 -13878 390718 -13822
rect 390774 -13878 390980 -13822
rect 391036 -13878 391122 -13822
rect 391178 -13878 391376 -13822
rect 391432 -13878 391518 -13822
rect 391574 -13878 391776 -13822
rect 391832 -13878 391918 -13822
rect 391974 -13878 392173 -13822
rect 392229 -13878 392315 -13822
rect 392371 -13878 392578 -13822
rect 392634 -13878 392720 -13822
rect 392776 -13878 392978 -13822
rect 393034 -13878 393120 -13822
rect 393176 -13878 393383 -13822
rect 393439 -13878 393525 -13822
rect 393581 -13878 393780 -13822
rect 393836 -13878 393922 -13822
rect 393978 -13878 394177 -13822
rect 394233 -13878 394319 -13822
rect 394375 -13878 394580 -13822
rect 394636 -13878 394722 -13822
rect 394778 -13878 394982 -13822
rect 395038 -13878 395124 -13822
rect 395180 -13878 395385 -13822
rect 395441 -13878 395527 -13822
rect 395583 -13878 395779 -13822
rect 395835 -13878 395921 -13822
rect 395977 -13878 396180 -13822
rect 396236 -13878 396322 -13822
rect 396378 -13878 396580 -13822
rect 396636 -13878 396722 -13822
rect 396778 -13878 396977 -13822
rect 397033 -13878 397119 -13822
rect 397175 -13878 397374 -13822
rect 397430 -13878 397516 -13822
rect 397572 -13878 397778 -13822
rect 397834 -13878 397920 -13822
rect 397976 -13878 398174 -13822
rect 398230 -13878 398316 -13822
rect 398372 -13878 398574 -13822
rect 398630 -13878 398716 -13822
rect 398772 -13878 398971 -13822
rect 399027 -13878 399113 -13822
rect 399169 -13878 399376 -13822
rect 399432 -13878 399518 -13822
rect 399574 -13878 399776 -13822
rect 399832 -13878 399918 -13822
rect 399974 -13878 400181 -13822
rect 400237 -13878 400323 -13822
rect 400379 -13878 402640 -13822
rect 387840 -13880 402640 -13878
rect 387840 -13936 387954 -13880
rect 388010 -13936 388078 -13880
rect 388134 -13936 388202 -13880
rect 388258 -13936 388326 -13880
rect 388382 -13936 388450 -13880
rect 388506 -13936 400766 -13880
rect 400822 -13936 400890 -13880
rect 400946 -13936 401014 -13880
rect 401070 -13936 401138 -13880
rect 401194 -13936 401262 -13880
rect 401318 -13936 402640 -13880
rect 387840 -13964 402640 -13936
rect 387840 -14004 388981 -13964
rect 387840 -14060 387954 -14004
rect 388010 -14060 388078 -14004
rect 388134 -14060 388202 -14004
rect 388258 -14060 388326 -14004
rect 388382 -14060 388450 -14004
rect 388506 -14020 388981 -14004
rect 389037 -14020 389123 -13964
rect 389179 -14020 389382 -13964
rect 389438 -14020 389524 -13964
rect 389580 -14020 389782 -13964
rect 389838 -14020 389924 -13964
rect 389980 -14020 390179 -13964
rect 390235 -14020 390321 -13964
rect 390377 -14020 390576 -13964
rect 390632 -14020 390718 -13964
rect 390774 -14020 390980 -13964
rect 391036 -14020 391122 -13964
rect 391178 -14020 391376 -13964
rect 391432 -14020 391518 -13964
rect 391574 -14020 391776 -13964
rect 391832 -14020 391918 -13964
rect 391974 -14020 392173 -13964
rect 392229 -14020 392315 -13964
rect 392371 -14020 392578 -13964
rect 392634 -14020 392720 -13964
rect 392776 -14020 392978 -13964
rect 393034 -14020 393120 -13964
rect 393176 -14020 393383 -13964
rect 393439 -14020 393525 -13964
rect 393581 -14020 393780 -13964
rect 393836 -14020 393922 -13964
rect 393978 -14020 394177 -13964
rect 394233 -14020 394319 -13964
rect 394375 -14020 394580 -13964
rect 394636 -14020 394722 -13964
rect 394778 -14020 394982 -13964
rect 395038 -14020 395124 -13964
rect 395180 -14020 395385 -13964
rect 395441 -14020 395527 -13964
rect 395583 -14020 395779 -13964
rect 395835 -14020 395921 -13964
rect 395977 -14020 396180 -13964
rect 396236 -14020 396322 -13964
rect 396378 -14020 396580 -13964
rect 396636 -14020 396722 -13964
rect 396778 -14020 396977 -13964
rect 397033 -14020 397119 -13964
rect 397175 -14020 397374 -13964
rect 397430 -14020 397516 -13964
rect 397572 -14020 397778 -13964
rect 397834 -14020 397920 -13964
rect 397976 -14020 398174 -13964
rect 398230 -14020 398316 -13964
rect 398372 -14020 398574 -13964
rect 398630 -14020 398716 -13964
rect 398772 -14020 398971 -13964
rect 399027 -14020 399113 -13964
rect 399169 -14020 399376 -13964
rect 399432 -14020 399518 -13964
rect 399574 -14020 399776 -13964
rect 399832 -14020 399918 -13964
rect 399974 -14020 400181 -13964
rect 400237 -14020 400323 -13964
rect 400379 -14004 402640 -13964
rect 400379 -14020 400766 -14004
rect 388506 -14060 400766 -14020
rect 400822 -14060 400890 -14004
rect 400946 -14060 401014 -14004
rect 401070 -14060 401138 -14004
rect 401194 -14060 401262 -14004
rect 401318 -14060 402640 -14004
rect 387840 -14106 402640 -14060
rect 387840 -14128 388981 -14106
rect 387840 -14184 387954 -14128
rect 388010 -14184 388078 -14128
rect 388134 -14184 388202 -14128
rect 388258 -14184 388326 -14128
rect 388382 -14184 388450 -14128
rect 388506 -14162 388981 -14128
rect 389037 -14162 389123 -14106
rect 389179 -14162 389382 -14106
rect 389438 -14162 389524 -14106
rect 389580 -14162 389782 -14106
rect 389838 -14162 389924 -14106
rect 389980 -14162 390179 -14106
rect 390235 -14162 390321 -14106
rect 390377 -14162 390576 -14106
rect 390632 -14162 390718 -14106
rect 390774 -14162 390980 -14106
rect 391036 -14162 391122 -14106
rect 391178 -14162 391376 -14106
rect 391432 -14162 391518 -14106
rect 391574 -14162 391776 -14106
rect 391832 -14162 391918 -14106
rect 391974 -14162 392173 -14106
rect 392229 -14162 392315 -14106
rect 392371 -14162 392578 -14106
rect 392634 -14162 392720 -14106
rect 392776 -14162 392978 -14106
rect 393034 -14162 393120 -14106
rect 393176 -14162 393383 -14106
rect 393439 -14162 393525 -14106
rect 393581 -14162 393780 -14106
rect 393836 -14162 393922 -14106
rect 393978 -14162 394177 -14106
rect 394233 -14162 394319 -14106
rect 394375 -14162 394580 -14106
rect 394636 -14162 394722 -14106
rect 394778 -14162 394982 -14106
rect 395038 -14162 395124 -14106
rect 395180 -14162 395385 -14106
rect 395441 -14162 395527 -14106
rect 395583 -14162 395779 -14106
rect 395835 -14162 395921 -14106
rect 395977 -14162 396180 -14106
rect 396236 -14162 396322 -14106
rect 396378 -14162 396580 -14106
rect 396636 -14162 396722 -14106
rect 396778 -14162 396977 -14106
rect 397033 -14162 397119 -14106
rect 397175 -14162 397374 -14106
rect 397430 -14162 397516 -14106
rect 397572 -14162 397778 -14106
rect 397834 -14162 397920 -14106
rect 397976 -14162 398174 -14106
rect 398230 -14162 398316 -14106
rect 398372 -14162 398574 -14106
rect 398630 -14162 398716 -14106
rect 398772 -14162 398971 -14106
rect 399027 -14162 399113 -14106
rect 399169 -14162 399376 -14106
rect 399432 -14162 399518 -14106
rect 399574 -14162 399776 -14106
rect 399832 -14162 399918 -14106
rect 399974 -14162 400181 -14106
rect 400237 -14162 400323 -14106
rect 400379 -14128 402640 -14106
rect 400379 -14162 400766 -14128
rect 388506 -14184 400766 -14162
rect 400822 -14184 400890 -14128
rect 400946 -14184 401014 -14128
rect 401070 -14184 401138 -14128
rect 401194 -14184 401262 -14128
rect 401318 -14184 402640 -14128
rect 387840 -14248 402640 -14184
rect 387840 -14252 388981 -14248
rect 387840 -14308 387954 -14252
rect 388010 -14308 388078 -14252
rect 388134 -14308 388202 -14252
rect 388258 -14308 388326 -14252
rect 388382 -14308 388450 -14252
rect 388506 -14304 388981 -14252
rect 389037 -14304 389123 -14248
rect 389179 -14304 389382 -14248
rect 389438 -14304 389524 -14248
rect 389580 -14304 389782 -14248
rect 389838 -14304 389924 -14248
rect 389980 -14304 390179 -14248
rect 390235 -14304 390321 -14248
rect 390377 -14304 390576 -14248
rect 390632 -14304 390718 -14248
rect 390774 -14304 390980 -14248
rect 391036 -14304 391122 -14248
rect 391178 -14304 391376 -14248
rect 391432 -14304 391518 -14248
rect 391574 -14304 391776 -14248
rect 391832 -14304 391918 -14248
rect 391974 -14304 392173 -14248
rect 392229 -14304 392315 -14248
rect 392371 -14304 392578 -14248
rect 392634 -14304 392720 -14248
rect 392776 -14304 392978 -14248
rect 393034 -14304 393120 -14248
rect 393176 -14304 393383 -14248
rect 393439 -14304 393525 -14248
rect 393581 -14304 393780 -14248
rect 393836 -14304 393922 -14248
rect 393978 -14304 394177 -14248
rect 394233 -14304 394319 -14248
rect 394375 -14304 394580 -14248
rect 394636 -14304 394722 -14248
rect 394778 -14304 394982 -14248
rect 395038 -14304 395124 -14248
rect 395180 -14304 395385 -14248
rect 395441 -14304 395527 -14248
rect 395583 -14304 395779 -14248
rect 395835 -14304 395921 -14248
rect 395977 -14304 396180 -14248
rect 396236 -14304 396322 -14248
rect 396378 -14304 396580 -14248
rect 396636 -14304 396722 -14248
rect 396778 -14304 396977 -14248
rect 397033 -14304 397119 -14248
rect 397175 -14304 397374 -14248
rect 397430 -14304 397516 -14248
rect 397572 -14304 397778 -14248
rect 397834 -14304 397920 -14248
rect 397976 -14304 398174 -14248
rect 398230 -14304 398316 -14248
rect 398372 -14304 398574 -14248
rect 398630 -14304 398716 -14248
rect 398772 -14304 398971 -14248
rect 399027 -14304 399113 -14248
rect 399169 -14304 399376 -14248
rect 399432 -14304 399518 -14248
rect 399574 -14304 399776 -14248
rect 399832 -14304 399918 -14248
rect 399974 -14304 400181 -14248
rect 400237 -14304 400323 -14248
rect 400379 -14252 402640 -14248
rect 400379 -14304 400766 -14252
rect 388506 -14308 400766 -14304
rect 400822 -14308 400890 -14252
rect 400946 -14308 401014 -14252
rect 401070 -14308 401138 -14252
rect 401194 -14308 401262 -14252
rect 401318 -14308 402640 -14252
rect 387840 -14376 402640 -14308
rect 387840 -14432 387954 -14376
rect 388010 -14432 388078 -14376
rect 388134 -14432 388202 -14376
rect 388258 -14432 388326 -14376
rect 388382 -14432 388450 -14376
rect 388506 -14390 400766 -14376
rect 388506 -14432 388981 -14390
rect 387840 -14446 388981 -14432
rect 389037 -14446 389123 -14390
rect 389179 -14446 389382 -14390
rect 389438 -14446 389524 -14390
rect 389580 -14446 389782 -14390
rect 389838 -14446 389924 -14390
rect 389980 -14446 390179 -14390
rect 390235 -14446 390321 -14390
rect 390377 -14446 390576 -14390
rect 390632 -14446 390718 -14390
rect 390774 -14446 390980 -14390
rect 391036 -14446 391122 -14390
rect 391178 -14446 391376 -14390
rect 391432 -14446 391518 -14390
rect 391574 -14446 391776 -14390
rect 391832 -14446 391918 -14390
rect 391974 -14446 392173 -14390
rect 392229 -14446 392315 -14390
rect 392371 -14446 392578 -14390
rect 392634 -14446 392720 -14390
rect 392776 -14446 392978 -14390
rect 393034 -14446 393120 -14390
rect 393176 -14446 393383 -14390
rect 393439 -14446 393525 -14390
rect 393581 -14446 393780 -14390
rect 393836 -14446 393922 -14390
rect 393978 -14446 394177 -14390
rect 394233 -14446 394319 -14390
rect 394375 -14446 394580 -14390
rect 394636 -14446 394722 -14390
rect 394778 -14446 394982 -14390
rect 395038 -14446 395124 -14390
rect 395180 -14446 395385 -14390
rect 395441 -14446 395527 -14390
rect 395583 -14446 395779 -14390
rect 395835 -14446 395921 -14390
rect 395977 -14446 396180 -14390
rect 396236 -14446 396322 -14390
rect 396378 -14446 396580 -14390
rect 396636 -14446 396722 -14390
rect 396778 -14446 396977 -14390
rect 397033 -14446 397119 -14390
rect 397175 -14446 397374 -14390
rect 397430 -14446 397516 -14390
rect 397572 -14446 397778 -14390
rect 397834 -14446 397920 -14390
rect 397976 -14446 398174 -14390
rect 398230 -14446 398316 -14390
rect 398372 -14446 398574 -14390
rect 398630 -14446 398716 -14390
rect 398772 -14446 398971 -14390
rect 399027 -14446 399113 -14390
rect 399169 -14446 399376 -14390
rect 399432 -14446 399518 -14390
rect 399574 -14446 399776 -14390
rect 399832 -14446 399918 -14390
rect 399974 -14446 400181 -14390
rect 400237 -14446 400323 -14390
rect 400379 -14432 400766 -14390
rect 400822 -14432 400890 -14376
rect 400946 -14432 401014 -14376
rect 401070 -14432 401138 -14376
rect 401194 -14432 401262 -14376
rect 401318 -14432 402640 -14376
rect 400379 -14446 402640 -14432
rect 387840 -14500 402640 -14446
rect 387840 -14556 387954 -14500
rect 388010 -14556 388078 -14500
rect 388134 -14556 388202 -14500
rect 388258 -14556 388326 -14500
rect 388382 -14556 388450 -14500
rect 388506 -14532 400766 -14500
rect 388506 -14556 388981 -14532
rect 387840 -14588 388981 -14556
rect 389037 -14588 389123 -14532
rect 389179 -14588 389382 -14532
rect 389438 -14588 389524 -14532
rect 389580 -14588 389782 -14532
rect 389838 -14588 389924 -14532
rect 389980 -14588 390179 -14532
rect 390235 -14588 390321 -14532
rect 390377 -14588 390576 -14532
rect 390632 -14588 390718 -14532
rect 390774 -14588 390980 -14532
rect 391036 -14588 391122 -14532
rect 391178 -14588 391376 -14532
rect 391432 -14588 391518 -14532
rect 391574 -14588 391776 -14532
rect 391832 -14588 391918 -14532
rect 391974 -14588 392173 -14532
rect 392229 -14588 392315 -14532
rect 392371 -14588 392578 -14532
rect 392634 -14588 392720 -14532
rect 392776 -14588 392978 -14532
rect 393034 -14588 393120 -14532
rect 393176 -14588 393383 -14532
rect 393439 -14588 393525 -14532
rect 393581 -14588 393780 -14532
rect 393836 -14588 393922 -14532
rect 393978 -14588 394177 -14532
rect 394233 -14588 394319 -14532
rect 394375 -14588 394580 -14532
rect 394636 -14588 394722 -14532
rect 394778 -14588 394982 -14532
rect 395038 -14588 395124 -14532
rect 395180 -14588 395385 -14532
rect 395441 -14588 395527 -14532
rect 395583 -14588 395779 -14532
rect 395835 -14588 395921 -14532
rect 395977 -14588 396180 -14532
rect 396236 -14588 396322 -14532
rect 396378 -14588 396580 -14532
rect 396636 -14588 396722 -14532
rect 396778 -14588 396977 -14532
rect 397033 -14588 397119 -14532
rect 397175 -14588 397374 -14532
rect 397430 -14588 397516 -14532
rect 397572 -14588 397778 -14532
rect 397834 -14588 397920 -14532
rect 397976 -14588 398174 -14532
rect 398230 -14588 398316 -14532
rect 398372 -14588 398574 -14532
rect 398630 -14588 398716 -14532
rect 398772 -14588 398971 -14532
rect 399027 -14588 399113 -14532
rect 399169 -14588 399376 -14532
rect 399432 -14588 399518 -14532
rect 399574 -14588 399776 -14532
rect 399832 -14588 399918 -14532
rect 399974 -14588 400181 -14532
rect 400237 -14588 400323 -14532
rect 400379 -14556 400766 -14532
rect 400822 -14556 400890 -14500
rect 400946 -14556 401014 -14500
rect 401070 -14556 401138 -14500
rect 401194 -14556 401262 -14500
rect 401318 -14556 402640 -14500
rect 400379 -14588 402640 -14556
rect 387840 -14624 402640 -14588
rect 387840 -14680 387954 -14624
rect 388010 -14680 388078 -14624
rect 388134 -14680 388202 -14624
rect 388258 -14680 388326 -14624
rect 388382 -14680 388450 -14624
rect 388506 -14674 400766 -14624
rect 388506 -14680 388981 -14674
rect 387840 -14730 388981 -14680
rect 389037 -14730 389123 -14674
rect 389179 -14730 389382 -14674
rect 389438 -14730 389524 -14674
rect 389580 -14730 389782 -14674
rect 389838 -14730 389924 -14674
rect 389980 -14730 390179 -14674
rect 390235 -14730 390321 -14674
rect 390377 -14730 390576 -14674
rect 390632 -14730 390718 -14674
rect 390774 -14730 390980 -14674
rect 391036 -14730 391122 -14674
rect 391178 -14730 391376 -14674
rect 391432 -14730 391518 -14674
rect 391574 -14730 391776 -14674
rect 391832 -14730 391918 -14674
rect 391974 -14730 392173 -14674
rect 392229 -14730 392315 -14674
rect 392371 -14730 392578 -14674
rect 392634 -14730 392720 -14674
rect 392776 -14730 392978 -14674
rect 393034 -14730 393120 -14674
rect 393176 -14730 393383 -14674
rect 393439 -14730 393525 -14674
rect 393581 -14730 393780 -14674
rect 393836 -14730 393922 -14674
rect 393978 -14730 394177 -14674
rect 394233 -14730 394319 -14674
rect 394375 -14730 394580 -14674
rect 394636 -14730 394722 -14674
rect 394778 -14730 394982 -14674
rect 395038 -14730 395124 -14674
rect 395180 -14730 395385 -14674
rect 395441 -14730 395527 -14674
rect 395583 -14730 395779 -14674
rect 395835 -14730 395921 -14674
rect 395977 -14730 396180 -14674
rect 396236 -14730 396322 -14674
rect 396378 -14730 396580 -14674
rect 396636 -14730 396722 -14674
rect 396778 -14730 396977 -14674
rect 397033 -14730 397119 -14674
rect 397175 -14730 397374 -14674
rect 397430 -14730 397516 -14674
rect 397572 -14730 397778 -14674
rect 397834 -14730 397920 -14674
rect 397976 -14730 398174 -14674
rect 398230 -14730 398316 -14674
rect 398372 -14730 398574 -14674
rect 398630 -14730 398716 -14674
rect 398772 -14730 398971 -14674
rect 399027 -14730 399113 -14674
rect 399169 -14730 399376 -14674
rect 399432 -14730 399518 -14674
rect 399574 -14730 399776 -14674
rect 399832 -14730 399918 -14674
rect 399974 -14730 400181 -14674
rect 400237 -14730 400323 -14674
rect 400379 -14680 400766 -14674
rect 400822 -14680 400890 -14624
rect 400946 -14680 401014 -14624
rect 401070 -14680 401138 -14624
rect 401194 -14680 401262 -14624
rect 401318 -14680 402640 -14624
rect 400379 -14730 402640 -14680
rect 387840 -14748 402640 -14730
rect 387840 -14804 387954 -14748
rect 388010 -14804 388078 -14748
rect 388134 -14804 388202 -14748
rect 388258 -14804 388326 -14748
rect 388382 -14804 388450 -14748
rect 388506 -14804 400766 -14748
rect 400822 -14804 400890 -14748
rect 400946 -14804 401014 -14748
rect 401070 -14804 401138 -14748
rect 401194 -14804 401262 -14748
rect 401318 -14804 402640 -14748
rect 387840 -14816 402640 -14804
rect 387840 -14872 388981 -14816
rect 389037 -14872 389123 -14816
rect 389179 -14872 389382 -14816
rect 389438 -14872 389524 -14816
rect 389580 -14872 389782 -14816
rect 389838 -14872 389924 -14816
rect 389980 -14872 390179 -14816
rect 390235 -14872 390321 -14816
rect 390377 -14872 390576 -14816
rect 390632 -14872 390718 -14816
rect 390774 -14872 390980 -14816
rect 391036 -14872 391122 -14816
rect 391178 -14872 391376 -14816
rect 391432 -14872 391518 -14816
rect 391574 -14872 391776 -14816
rect 391832 -14872 391918 -14816
rect 391974 -14872 392173 -14816
rect 392229 -14872 392315 -14816
rect 392371 -14872 392578 -14816
rect 392634 -14872 392720 -14816
rect 392776 -14872 392978 -14816
rect 393034 -14872 393120 -14816
rect 393176 -14872 393383 -14816
rect 393439 -14872 393525 -14816
rect 393581 -14872 393780 -14816
rect 393836 -14872 393922 -14816
rect 393978 -14872 394177 -14816
rect 394233 -14872 394319 -14816
rect 394375 -14872 394580 -14816
rect 394636 -14872 394722 -14816
rect 394778 -14872 394982 -14816
rect 395038 -14872 395124 -14816
rect 395180 -14872 395385 -14816
rect 395441 -14872 395527 -14816
rect 395583 -14872 395779 -14816
rect 395835 -14872 395921 -14816
rect 395977 -14872 396180 -14816
rect 396236 -14872 396322 -14816
rect 396378 -14872 396580 -14816
rect 396636 -14872 396722 -14816
rect 396778 -14872 396977 -14816
rect 397033 -14872 397119 -14816
rect 397175 -14872 397374 -14816
rect 397430 -14872 397516 -14816
rect 397572 -14872 397778 -14816
rect 397834 -14872 397920 -14816
rect 397976 -14872 398174 -14816
rect 398230 -14872 398316 -14816
rect 398372 -14872 398574 -14816
rect 398630 -14872 398716 -14816
rect 398772 -14872 398971 -14816
rect 399027 -14872 399113 -14816
rect 399169 -14872 399376 -14816
rect 399432 -14872 399518 -14816
rect 399574 -14872 399776 -14816
rect 399832 -14872 399918 -14816
rect 399974 -14872 400181 -14816
rect 400237 -14872 400323 -14816
rect 400379 -14872 402640 -14816
rect 387840 -14928 387954 -14872
rect 388010 -14928 388078 -14872
rect 388134 -14928 388202 -14872
rect 388258 -14928 388326 -14872
rect 388382 -14928 388450 -14872
rect 388506 -14928 400766 -14872
rect 400822 -14928 400890 -14872
rect 400946 -14928 401014 -14872
rect 401070 -14928 401138 -14872
rect 401194 -14928 401262 -14872
rect 401318 -14928 402640 -14872
rect 387840 -14958 402640 -14928
rect 387840 -14996 388981 -14958
rect 387840 -15052 387954 -14996
rect 388010 -15052 388078 -14996
rect 388134 -15052 388202 -14996
rect 388258 -15052 388326 -14996
rect 388382 -15052 388450 -14996
rect 388506 -15014 388981 -14996
rect 389037 -15014 389123 -14958
rect 389179 -15014 389382 -14958
rect 389438 -15014 389524 -14958
rect 389580 -15014 389782 -14958
rect 389838 -15014 389924 -14958
rect 389980 -15014 390179 -14958
rect 390235 -15014 390321 -14958
rect 390377 -15014 390576 -14958
rect 390632 -15014 390718 -14958
rect 390774 -15014 390980 -14958
rect 391036 -15014 391122 -14958
rect 391178 -15014 391376 -14958
rect 391432 -15014 391518 -14958
rect 391574 -15014 391776 -14958
rect 391832 -15014 391918 -14958
rect 391974 -15014 392173 -14958
rect 392229 -15014 392315 -14958
rect 392371 -15014 392578 -14958
rect 392634 -15014 392720 -14958
rect 392776 -15014 392978 -14958
rect 393034 -15014 393120 -14958
rect 393176 -15014 393383 -14958
rect 393439 -15014 393525 -14958
rect 393581 -15014 393780 -14958
rect 393836 -15014 393922 -14958
rect 393978 -15014 394177 -14958
rect 394233 -15014 394319 -14958
rect 394375 -15014 394580 -14958
rect 394636 -15014 394722 -14958
rect 394778 -15014 394982 -14958
rect 395038 -15014 395124 -14958
rect 395180 -15014 395385 -14958
rect 395441 -15014 395527 -14958
rect 395583 -15014 395779 -14958
rect 395835 -15014 395921 -14958
rect 395977 -15014 396180 -14958
rect 396236 -15014 396322 -14958
rect 396378 -15014 396580 -14958
rect 396636 -15014 396722 -14958
rect 396778 -15014 396977 -14958
rect 397033 -15014 397119 -14958
rect 397175 -15014 397374 -14958
rect 397430 -15014 397516 -14958
rect 397572 -15014 397778 -14958
rect 397834 -15014 397920 -14958
rect 397976 -15014 398174 -14958
rect 398230 -15014 398316 -14958
rect 398372 -15014 398574 -14958
rect 398630 -15014 398716 -14958
rect 398772 -15014 398971 -14958
rect 399027 -15014 399113 -14958
rect 399169 -15014 399376 -14958
rect 399432 -15014 399518 -14958
rect 399574 -15014 399776 -14958
rect 399832 -15014 399918 -14958
rect 399974 -15014 400181 -14958
rect 400237 -15014 400323 -14958
rect 400379 -14996 402640 -14958
rect 400379 -15014 400766 -14996
rect 388506 -15052 400766 -15014
rect 400822 -15052 400890 -14996
rect 400946 -15052 401014 -14996
rect 401070 -15052 401138 -14996
rect 401194 -15052 401262 -14996
rect 401318 -15052 402640 -14996
rect 387840 -15100 402640 -15052
rect 387840 -15120 388981 -15100
rect 387840 -15176 387954 -15120
rect 388010 -15176 388078 -15120
rect 388134 -15176 388202 -15120
rect 388258 -15176 388326 -15120
rect 388382 -15176 388450 -15120
rect 388506 -15156 388981 -15120
rect 389037 -15156 389123 -15100
rect 389179 -15156 389382 -15100
rect 389438 -15156 389524 -15100
rect 389580 -15156 389782 -15100
rect 389838 -15156 389924 -15100
rect 389980 -15156 390179 -15100
rect 390235 -15156 390321 -15100
rect 390377 -15156 390576 -15100
rect 390632 -15156 390718 -15100
rect 390774 -15156 390980 -15100
rect 391036 -15156 391122 -15100
rect 391178 -15156 391376 -15100
rect 391432 -15156 391518 -15100
rect 391574 -15156 391776 -15100
rect 391832 -15156 391918 -15100
rect 391974 -15156 392173 -15100
rect 392229 -15156 392315 -15100
rect 392371 -15156 392578 -15100
rect 392634 -15156 392720 -15100
rect 392776 -15156 392978 -15100
rect 393034 -15156 393120 -15100
rect 393176 -15156 393383 -15100
rect 393439 -15156 393525 -15100
rect 393581 -15156 393780 -15100
rect 393836 -15156 393922 -15100
rect 393978 -15156 394177 -15100
rect 394233 -15156 394319 -15100
rect 394375 -15156 394580 -15100
rect 394636 -15156 394722 -15100
rect 394778 -15156 394982 -15100
rect 395038 -15156 395124 -15100
rect 395180 -15156 395385 -15100
rect 395441 -15156 395527 -15100
rect 395583 -15156 395779 -15100
rect 395835 -15156 395921 -15100
rect 395977 -15156 396180 -15100
rect 396236 -15156 396322 -15100
rect 396378 -15156 396580 -15100
rect 396636 -15156 396722 -15100
rect 396778 -15156 396977 -15100
rect 397033 -15156 397119 -15100
rect 397175 -15156 397374 -15100
rect 397430 -15156 397516 -15100
rect 397572 -15156 397778 -15100
rect 397834 -15156 397920 -15100
rect 397976 -15156 398174 -15100
rect 398230 -15156 398316 -15100
rect 398372 -15156 398574 -15100
rect 398630 -15156 398716 -15100
rect 398772 -15156 398971 -15100
rect 399027 -15156 399113 -15100
rect 399169 -15156 399376 -15100
rect 399432 -15156 399518 -15100
rect 399574 -15156 399776 -15100
rect 399832 -15156 399918 -15100
rect 399974 -15156 400181 -15100
rect 400237 -15156 400323 -15100
rect 400379 -15120 402640 -15100
rect 400379 -15156 400766 -15120
rect 388506 -15176 400766 -15156
rect 400822 -15176 400890 -15120
rect 400946 -15176 401014 -15120
rect 401070 -15176 401138 -15120
rect 401194 -15176 401262 -15120
rect 401318 -15176 402640 -15120
rect 387840 -15242 402640 -15176
rect 387840 -15244 388981 -15242
rect 387840 -15300 387954 -15244
rect 388010 -15300 388078 -15244
rect 388134 -15300 388202 -15244
rect 388258 -15300 388326 -15244
rect 388382 -15300 388450 -15244
rect 388506 -15298 388981 -15244
rect 389037 -15298 389123 -15242
rect 389179 -15298 389382 -15242
rect 389438 -15298 389524 -15242
rect 389580 -15298 389782 -15242
rect 389838 -15298 389924 -15242
rect 389980 -15298 390179 -15242
rect 390235 -15298 390321 -15242
rect 390377 -15298 390576 -15242
rect 390632 -15298 390718 -15242
rect 390774 -15298 390980 -15242
rect 391036 -15298 391122 -15242
rect 391178 -15298 391376 -15242
rect 391432 -15298 391518 -15242
rect 391574 -15298 391776 -15242
rect 391832 -15298 391918 -15242
rect 391974 -15298 392173 -15242
rect 392229 -15298 392315 -15242
rect 392371 -15298 392578 -15242
rect 392634 -15298 392720 -15242
rect 392776 -15298 392978 -15242
rect 393034 -15298 393120 -15242
rect 393176 -15298 393383 -15242
rect 393439 -15298 393525 -15242
rect 393581 -15298 393780 -15242
rect 393836 -15298 393922 -15242
rect 393978 -15298 394177 -15242
rect 394233 -15298 394319 -15242
rect 394375 -15298 394580 -15242
rect 394636 -15298 394722 -15242
rect 394778 -15298 394982 -15242
rect 395038 -15298 395124 -15242
rect 395180 -15298 395385 -15242
rect 395441 -15298 395527 -15242
rect 395583 -15298 395779 -15242
rect 395835 -15298 395921 -15242
rect 395977 -15298 396180 -15242
rect 396236 -15298 396322 -15242
rect 396378 -15298 396580 -15242
rect 396636 -15298 396722 -15242
rect 396778 -15298 396977 -15242
rect 397033 -15298 397119 -15242
rect 397175 -15298 397374 -15242
rect 397430 -15298 397516 -15242
rect 397572 -15298 397778 -15242
rect 397834 -15298 397920 -15242
rect 397976 -15298 398174 -15242
rect 398230 -15298 398316 -15242
rect 398372 -15298 398574 -15242
rect 398630 -15298 398716 -15242
rect 398772 -15298 398971 -15242
rect 399027 -15298 399113 -15242
rect 399169 -15298 399376 -15242
rect 399432 -15298 399518 -15242
rect 399574 -15298 399776 -15242
rect 399832 -15298 399918 -15242
rect 399974 -15298 400181 -15242
rect 400237 -15298 400323 -15242
rect 400379 -15244 402640 -15242
rect 400379 -15298 400766 -15244
rect 388506 -15300 400766 -15298
rect 400822 -15300 400890 -15244
rect 400946 -15300 401014 -15244
rect 401070 -15300 401138 -15244
rect 401194 -15300 401262 -15244
rect 401318 -15300 402640 -15244
rect 387840 -15368 402640 -15300
rect 387840 -15424 387954 -15368
rect 388010 -15424 388078 -15368
rect 388134 -15424 388202 -15368
rect 388258 -15424 388326 -15368
rect 388382 -15424 388450 -15368
rect 388506 -15384 400766 -15368
rect 388506 -15424 388981 -15384
rect 387840 -15440 388981 -15424
rect 389037 -15440 389123 -15384
rect 389179 -15440 389382 -15384
rect 389438 -15440 389524 -15384
rect 389580 -15440 389782 -15384
rect 389838 -15440 389924 -15384
rect 389980 -15440 390179 -15384
rect 390235 -15440 390321 -15384
rect 390377 -15440 390576 -15384
rect 390632 -15440 390718 -15384
rect 390774 -15440 390980 -15384
rect 391036 -15440 391122 -15384
rect 391178 -15440 391376 -15384
rect 391432 -15440 391518 -15384
rect 391574 -15440 391776 -15384
rect 391832 -15440 391918 -15384
rect 391974 -15440 392173 -15384
rect 392229 -15440 392315 -15384
rect 392371 -15440 392578 -15384
rect 392634 -15440 392720 -15384
rect 392776 -15440 392978 -15384
rect 393034 -15440 393120 -15384
rect 393176 -15440 393383 -15384
rect 393439 -15440 393525 -15384
rect 393581 -15440 393780 -15384
rect 393836 -15440 393922 -15384
rect 393978 -15440 394177 -15384
rect 394233 -15440 394319 -15384
rect 394375 -15440 394580 -15384
rect 394636 -15440 394722 -15384
rect 394778 -15440 394982 -15384
rect 395038 -15440 395124 -15384
rect 395180 -15440 395385 -15384
rect 395441 -15440 395527 -15384
rect 395583 -15440 395779 -15384
rect 395835 -15440 395921 -15384
rect 395977 -15440 396180 -15384
rect 396236 -15440 396322 -15384
rect 396378 -15440 396580 -15384
rect 396636 -15440 396722 -15384
rect 396778 -15440 396977 -15384
rect 397033 -15440 397119 -15384
rect 397175 -15440 397374 -15384
rect 397430 -15440 397516 -15384
rect 397572 -15440 397778 -15384
rect 397834 -15440 397920 -15384
rect 397976 -15440 398174 -15384
rect 398230 -15440 398316 -15384
rect 398372 -15440 398574 -15384
rect 398630 -15440 398716 -15384
rect 398772 -15440 398971 -15384
rect 399027 -15440 399113 -15384
rect 399169 -15440 399376 -15384
rect 399432 -15440 399518 -15384
rect 399574 -15440 399776 -15384
rect 399832 -15440 399918 -15384
rect 399974 -15440 400181 -15384
rect 400237 -15440 400323 -15384
rect 400379 -15424 400766 -15384
rect 400822 -15424 400890 -15368
rect 400946 -15424 401014 -15368
rect 401070 -15424 401138 -15368
rect 401194 -15424 401262 -15368
rect 401318 -15424 402640 -15368
rect 400379 -15440 402640 -15424
rect 387840 -15492 402640 -15440
rect 387840 -15548 387954 -15492
rect 388010 -15548 388078 -15492
rect 388134 -15548 388202 -15492
rect 388258 -15548 388326 -15492
rect 388382 -15548 388450 -15492
rect 388506 -15526 400766 -15492
rect 388506 -15548 388981 -15526
rect 387840 -15582 388981 -15548
rect 389037 -15582 389123 -15526
rect 389179 -15582 389382 -15526
rect 389438 -15582 389524 -15526
rect 389580 -15582 389782 -15526
rect 389838 -15582 389924 -15526
rect 389980 -15582 390179 -15526
rect 390235 -15582 390321 -15526
rect 390377 -15582 390576 -15526
rect 390632 -15582 390718 -15526
rect 390774 -15582 390980 -15526
rect 391036 -15582 391122 -15526
rect 391178 -15582 391376 -15526
rect 391432 -15582 391518 -15526
rect 391574 -15582 391776 -15526
rect 391832 -15582 391918 -15526
rect 391974 -15582 392173 -15526
rect 392229 -15582 392315 -15526
rect 392371 -15582 392578 -15526
rect 392634 -15582 392720 -15526
rect 392776 -15582 392978 -15526
rect 393034 -15582 393120 -15526
rect 393176 -15582 393383 -15526
rect 393439 -15582 393525 -15526
rect 393581 -15582 393780 -15526
rect 393836 -15582 393922 -15526
rect 393978 -15582 394177 -15526
rect 394233 -15582 394319 -15526
rect 394375 -15582 394580 -15526
rect 394636 -15582 394722 -15526
rect 394778 -15582 394982 -15526
rect 395038 -15582 395124 -15526
rect 395180 -15582 395385 -15526
rect 395441 -15582 395527 -15526
rect 395583 -15582 395779 -15526
rect 395835 -15582 395921 -15526
rect 395977 -15582 396180 -15526
rect 396236 -15582 396322 -15526
rect 396378 -15582 396580 -15526
rect 396636 -15582 396722 -15526
rect 396778 -15582 396977 -15526
rect 397033 -15582 397119 -15526
rect 397175 -15582 397374 -15526
rect 397430 -15582 397516 -15526
rect 397572 -15582 397778 -15526
rect 397834 -15582 397920 -15526
rect 397976 -15582 398174 -15526
rect 398230 -15582 398316 -15526
rect 398372 -15582 398574 -15526
rect 398630 -15582 398716 -15526
rect 398772 -15582 398971 -15526
rect 399027 -15582 399113 -15526
rect 399169 -15582 399376 -15526
rect 399432 -15582 399518 -15526
rect 399574 -15582 399776 -15526
rect 399832 -15582 399918 -15526
rect 399974 -15582 400181 -15526
rect 400237 -15582 400323 -15526
rect 400379 -15548 400766 -15526
rect 400822 -15548 400890 -15492
rect 400946 -15548 401014 -15492
rect 401070 -15548 401138 -15492
rect 401194 -15548 401262 -15492
rect 401318 -15548 402640 -15492
rect 400379 -15582 402640 -15548
rect 387840 -15616 402640 -15582
rect 387840 -15672 387954 -15616
rect 388010 -15672 388078 -15616
rect 388134 -15672 388202 -15616
rect 388258 -15672 388326 -15616
rect 388382 -15672 388450 -15616
rect 388506 -15668 400766 -15616
rect 388506 -15672 388981 -15668
rect 387840 -15724 388981 -15672
rect 389037 -15724 389123 -15668
rect 389179 -15724 389382 -15668
rect 389438 -15724 389524 -15668
rect 389580 -15724 389782 -15668
rect 389838 -15724 389924 -15668
rect 389980 -15724 390179 -15668
rect 390235 -15724 390321 -15668
rect 390377 -15724 390576 -15668
rect 390632 -15724 390718 -15668
rect 390774 -15724 390980 -15668
rect 391036 -15724 391122 -15668
rect 391178 -15724 391376 -15668
rect 391432 -15724 391518 -15668
rect 391574 -15724 391776 -15668
rect 391832 -15724 391918 -15668
rect 391974 -15724 392173 -15668
rect 392229 -15724 392315 -15668
rect 392371 -15724 392578 -15668
rect 392634 -15724 392720 -15668
rect 392776 -15724 392978 -15668
rect 393034 -15724 393120 -15668
rect 393176 -15724 393383 -15668
rect 393439 -15724 393525 -15668
rect 393581 -15724 393780 -15668
rect 393836 -15724 393922 -15668
rect 393978 -15724 394177 -15668
rect 394233 -15724 394319 -15668
rect 394375 -15724 394580 -15668
rect 394636 -15724 394722 -15668
rect 394778 -15724 394982 -15668
rect 395038 -15724 395124 -15668
rect 395180 -15724 395385 -15668
rect 395441 -15724 395527 -15668
rect 395583 -15724 395779 -15668
rect 395835 -15724 395921 -15668
rect 395977 -15724 396180 -15668
rect 396236 -15724 396322 -15668
rect 396378 -15724 396580 -15668
rect 396636 -15724 396722 -15668
rect 396778 -15724 396977 -15668
rect 397033 -15724 397119 -15668
rect 397175 -15724 397374 -15668
rect 397430 -15724 397516 -15668
rect 397572 -15724 397778 -15668
rect 397834 -15724 397920 -15668
rect 397976 -15724 398174 -15668
rect 398230 -15724 398316 -15668
rect 398372 -15724 398574 -15668
rect 398630 -15724 398716 -15668
rect 398772 -15724 398971 -15668
rect 399027 -15724 399113 -15668
rect 399169 -15724 399376 -15668
rect 399432 -15724 399518 -15668
rect 399574 -15724 399776 -15668
rect 399832 -15724 399918 -15668
rect 399974 -15724 400181 -15668
rect 400237 -15724 400323 -15668
rect 400379 -15672 400766 -15668
rect 400822 -15672 400890 -15616
rect 400946 -15672 401014 -15616
rect 401070 -15672 401138 -15616
rect 401194 -15672 401262 -15616
rect 401318 -15672 402640 -15616
rect 400379 -15724 402640 -15672
rect 387840 -15740 402640 -15724
rect 387840 -15796 387954 -15740
rect 388010 -15796 388078 -15740
rect 388134 -15796 388202 -15740
rect 388258 -15796 388326 -15740
rect 388382 -15796 388450 -15740
rect 388506 -15796 400766 -15740
rect 400822 -15796 400890 -15740
rect 400946 -15796 401014 -15740
rect 401070 -15796 401138 -15740
rect 401194 -15796 401262 -15740
rect 401318 -15796 402640 -15740
rect 387840 -15810 402640 -15796
rect 387840 -15864 388981 -15810
rect 387840 -15920 387954 -15864
rect 388010 -15920 388078 -15864
rect 388134 -15920 388202 -15864
rect 388258 -15920 388326 -15864
rect 388382 -15920 388450 -15864
rect 388506 -15866 388981 -15864
rect 389037 -15866 389123 -15810
rect 389179 -15866 389382 -15810
rect 389438 -15866 389524 -15810
rect 389580 -15866 389782 -15810
rect 389838 -15866 389924 -15810
rect 389980 -15866 390179 -15810
rect 390235 -15866 390321 -15810
rect 390377 -15866 390576 -15810
rect 390632 -15866 390718 -15810
rect 390774 -15866 390980 -15810
rect 391036 -15866 391122 -15810
rect 391178 -15866 391376 -15810
rect 391432 -15866 391518 -15810
rect 391574 -15866 391776 -15810
rect 391832 -15866 391918 -15810
rect 391974 -15866 392173 -15810
rect 392229 -15866 392315 -15810
rect 392371 -15866 392578 -15810
rect 392634 -15866 392720 -15810
rect 392776 -15866 392978 -15810
rect 393034 -15866 393120 -15810
rect 393176 -15866 393383 -15810
rect 393439 -15866 393525 -15810
rect 393581 -15866 393780 -15810
rect 393836 -15866 393922 -15810
rect 393978 -15866 394177 -15810
rect 394233 -15866 394319 -15810
rect 394375 -15866 394580 -15810
rect 394636 -15866 394722 -15810
rect 394778 -15866 394982 -15810
rect 395038 -15866 395124 -15810
rect 395180 -15866 395385 -15810
rect 395441 -15866 395527 -15810
rect 395583 -15866 395779 -15810
rect 395835 -15866 395921 -15810
rect 395977 -15866 396180 -15810
rect 396236 -15866 396322 -15810
rect 396378 -15866 396580 -15810
rect 396636 -15866 396722 -15810
rect 396778 -15866 396977 -15810
rect 397033 -15866 397119 -15810
rect 397175 -15866 397374 -15810
rect 397430 -15866 397516 -15810
rect 397572 -15866 397778 -15810
rect 397834 -15866 397920 -15810
rect 397976 -15866 398174 -15810
rect 398230 -15866 398316 -15810
rect 398372 -15866 398574 -15810
rect 398630 -15866 398716 -15810
rect 398772 -15866 398971 -15810
rect 399027 -15866 399113 -15810
rect 399169 -15866 399376 -15810
rect 399432 -15866 399518 -15810
rect 399574 -15866 399776 -15810
rect 399832 -15866 399918 -15810
rect 399974 -15866 400181 -15810
rect 400237 -15866 400323 -15810
rect 400379 -15864 402640 -15810
rect 400379 -15866 400766 -15864
rect 388506 -15920 400766 -15866
rect 400822 -15920 400890 -15864
rect 400946 -15920 401014 -15864
rect 401070 -15920 401138 -15864
rect 401194 -15920 401262 -15864
rect 401318 -15920 402640 -15864
rect 387840 -15952 402640 -15920
rect 387840 -15988 388981 -15952
rect 387840 -16044 387954 -15988
rect 388010 -16044 388078 -15988
rect 388134 -16044 388202 -15988
rect 388258 -16044 388326 -15988
rect 388382 -16044 388450 -15988
rect 388506 -16008 388981 -15988
rect 389037 -16008 389123 -15952
rect 389179 -16008 389382 -15952
rect 389438 -16008 389524 -15952
rect 389580 -16008 389782 -15952
rect 389838 -16008 389924 -15952
rect 389980 -16008 390179 -15952
rect 390235 -16008 390321 -15952
rect 390377 -16008 390576 -15952
rect 390632 -16008 390718 -15952
rect 390774 -16008 390980 -15952
rect 391036 -16008 391122 -15952
rect 391178 -16008 391376 -15952
rect 391432 -16008 391518 -15952
rect 391574 -16008 391776 -15952
rect 391832 -16008 391918 -15952
rect 391974 -16008 392173 -15952
rect 392229 -16008 392315 -15952
rect 392371 -16008 392578 -15952
rect 392634 -16008 392720 -15952
rect 392776 -16008 392978 -15952
rect 393034 -16008 393120 -15952
rect 393176 -16008 393383 -15952
rect 393439 -16008 393525 -15952
rect 393581 -16008 393780 -15952
rect 393836 -16008 393922 -15952
rect 393978 -16008 394177 -15952
rect 394233 -16008 394319 -15952
rect 394375 -16008 394580 -15952
rect 394636 -16008 394722 -15952
rect 394778 -16008 394982 -15952
rect 395038 -16008 395124 -15952
rect 395180 -16008 395385 -15952
rect 395441 -16008 395527 -15952
rect 395583 -16008 395779 -15952
rect 395835 -16008 395921 -15952
rect 395977 -16008 396180 -15952
rect 396236 -16008 396322 -15952
rect 396378 -16008 396580 -15952
rect 396636 -16008 396722 -15952
rect 396778 -16008 396977 -15952
rect 397033 -16008 397119 -15952
rect 397175 -16008 397374 -15952
rect 397430 -16008 397516 -15952
rect 397572 -16008 397778 -15952
rect 397834 -16008 397920 -15952
rect 397976 -16008 398174 -15952
rect 398230 -16008 398316 -15952
rect 398372 -16008 398574 -15952
rect 398630 -16008 398716 -15952
rect 398772 -16008 398971 -15952
rect 399027 -16008 399113 -15952
rect 399169 -16008 399376 -15952
rect 399432 -16008 399518 -15952
rect 399574 -16008 399776 -15952
rect 399832 -16008 399918 -15952
rect 399974 -16008 400181 -15952
rect 400237 -16008 400323 -15952
rect 400379 -15988 402640 -15952
rect 400379 -16008 400766 -15988
rect 388506 -16044 400766 -16008
rect 400822 -16044 400890 -15988
rect 400946 -16044 401014 -15988
rect 401070 -16044 401138 -15988
rect 401194 -16044 401262 -15988
rect 401318 -16044 402640 -15988
rect 387840 -16094 402640 -16044
rect 387840 -16112 388981 -16094
rect 387840 -16168 387954 -16112
rect 388010 -16168 388078 -16112
rect 388134 -16168 388202 -16112
rect 388258 -16168 388326 -16112
rect 388382 -16168 388450 -16112
rect 388506 -16150 388981 -16112
rect 389037 -16150 389123 -16094
rect 389179 -16150 389382 -16094
rect 389438 -16150 389524 -16094
rect 389580 -16150 389782 -16094
rect 389838 -16150 389924 -16094
rect 389980 -16150 390179 -16094
rect 390235 -16150 390321 -16094
rect 390377 -16150 390576 -16094
rect 390632 -16150 390718 -16094
rect 390774 -16150 390980 -16094
rect 391036 -16150 391122 -16094
rect 391178 -16150 391376 -16094
rect 391432 -16150 391518 -16094
rect 391574 -16150 391776 -16094
rect 391832 -16150 391918 -16094
rect 391974 -16150 392173 -16094
rect 392229 -16150 392315 -16094
rect 392371 -16150 392578 -16094
rect 392634 -16150 392720 -16094
rect 392776 -16150 392978 -16094
rect 393034 -16150 393120 -16094
rect 393176 -16150 393383 -16094
rect 393439 -16150 393525 -16094
rect 393581 -16150 393780 -16094
rect 393836 -16150 393922 -16094
rect 393978 -16150 394177 -16094
rect 394233 -16150 394319 -16094
rect 394375 -16150 394580 -16094
rect 394636 -16150 394722 -16094
rect 394778 -16150 394982 -16094
rect 395038 -16150 395124 -16094
rect 395180 -16150 395385 -16094
rect 395441 -16150 395527 -16094
rect 395583 -16150 395779 -16094
rect 395835 -16150 395921 -16094
rect 395977 -16150 396180 -16094
rect 396236 -16150 396322 -16094
rect 396378 -16150 396580 -16094
rect 396636 -16150 396722 -16094
rect 396778 -16150 396977 -16094
rect 397033 -16150 397119 -16094
rect 397175 -16150 397374 -16094
rect 397430 -16150 397516 -16094
rect 397572 -16150 397778 -16094
rect 397834 -16150 397920 -16094
rect 397976 -16150 398174 -16094
rect 398230 -16150 398316 -16094
rect 398372 -16150 398574 -16094
rect 398630 -16150 398716 -16094
rect 398772 -16150 398971 -16094
rect 399027 -16150 399113 -16094
rect 399169 -16150 399376 -16094
rect 399432 -16150 399518 -16094
rect 399574 -16150 399776 -16094
rect 399832 -16150 399918 -16094
rect 399974 -16150 400181 -16094
rect 400237 -16150 400323 -16094
rect 400379 -16112 402640 -16094
rect 400379 -16150 400766 -16112
rect 388506 -16168 400766 -16150
rect 400822 -16168 400890 -16112
rect 400946 -16168 401014 -16112
rect 401070 -16168 401138 -16112
rect 401194 -16168 401262 -16112
rect 401318 -16168 402640 -16112
rect 387840 -16236 402640 -16168
rect 387840 -16292 387954 -16236
rect 388010 -16292 388078 -16236
rect 388134 -16292 388202 -16236
rect 388258 -16292 388326 -16236
rect 388382 -16292 388450 -16236
rect 388506 -16292 388981 -16236
rect 389037 -16292 389123 -16236
rect 389179 -16292 389382 -16236
rect 389438 -16292 389524 -16236
rect 389580 -16292 389782 -16236
rect 389838 -16292 389924 -16236
rect 389980 -16292 390179 -16236
rect 390235 -16292 390321 -16236
rect 390377 -16292 390576 -16236
rect 390632 -16292 390718 -16236
rect 390774 -16292 390980 -16236
rect 391036 -16292 391122 -16236
rect 391178 -16292 391376 -16236
rect 391432 -16292 391518 -16236
rect 391574 -16292 391776 -16236
rect 391832 -16292 391918 -16236
rect 391974 -16292 392173 -16236
rect 392229 -16292 392315 -16236
rect 392371 -16292 392578 -16236
rect 392634 -16292 392720 -16236
rect 392776 -16292 392978 -16236
rect 393034 -16292 393120 -16236
rect 393176 -16292 393383 -16236
rect 393439 -16292 393525 -16236
rect 393581 -16292 393780 -16236
rect 393836 -16292 393922 -16236
rect 393978 -16292 394177 -16236
rect 394233 -16292 394319 -16236
rect 394375 -16292 394580 -16236
rect 394636 -16292 394722 -16236
rect 394778 -16292 394982 -16236
rect 395038 -16292 395124 -16236
rect 395180 -16292 395385 -16236
rect 395441 -16292 395527 -16236
rect 395583 -16292 395779 -16236
rect 395835 -16292 395921 -16236
rect 395977 -16292 396180 -16236
rect 396236 -16292 396322 -16236
rect 396378 -16292 396580 -16236
rect 396636 -16292 396722 -16236
rect 396778 -16292 396977 -16236
rect 397033 -16292 397119 -16236
rect 397175 -16292 397374 -16236
rect 397430 -16292 397516 -16236
rect 397572 -16292 397778 -16236
rect 397834 -16292 397920 -16236
rect 397976 -16292 398174 -16236
rect 398230 -16292 398316 -16236
rect 398372 -16292 398574 -16236
rect 398630 -16292 398716 -16236
rect 398772 -16292 398971 -16236
rect 399027 -16292 399113 -16236
rect 399169 -16292 399376 -16236
rect 399432 -16292 399518 -16236
rect 399574 -16292 399776 -16236
rect 399832 -16292 399918 -16236
rect 399974 -16292 400181 -16236
rect 400237 -16292 400323 -16236
rect 400379 -16292 400766 -16236
rect 400822 -16292 400890 -16236
rect 400946 -16292 401014 -16236
rect 401070 -16292 401138 -16236
rect 401194 -16292 401262 -16236
rect 401318 -16292 402640 -16236
rect 387840 -16360 402640 -16292
rect 387840 -16416 387954 -16360
rect 388010 -16416 388078 -16360
rect 388134 -16416 388202 -16360
rect 388258 -16416 388326 -16360
rect 388382 -16416 388450 -16360
rect 388506 -16378 400766 -16360
rect 388506 -16416 388981 -16378
rect 387840 -16434 388981 -16416
rect 389037 -16434 389123 -16378
rect 389179 -16434 389382 -16378
rect 389438 -16434 389524 -16378
rect 389580 -16434 389782 -16378
rect 389838 -16434 389924 -16378
rect 389980 -16434 390179 -16378
rect 390235 -16434 390321 -16378
rect 390377 -16434 390576 -16378
rect 390632 -16434 390718 -16378
rect 390774 -16434 390980 -16378
rect 391036 -16434 391122 -16378
rect 391178 -16434 391376 -16378
rect 391432 -16434 391518 -16378
rect 391574 -16434 391776 -16378
rect 391832 -16434 391918 -16378
rect 391974 -16434 392173 -16378
rect 392229 -16434 392315 -16378
rect 392371 -16434 392578 -16378
rect 392634 -16434 392720 -16378
rect 392776 -16434 392978 -16378
rect 393034 -16434 393120 -16378
rect 393176 -16434 393383 -16378
rect 393439 -16434 393525 -16378
rect 393581 -16434 393780 -16378
rect 393836 -16434 393922 -16378
rect 393978 -16434 394177 -16378
rect 394233 -16434 394319 -16378
rect 394375 -16434 394580 -16378
rect 394636 -16434 394722 -16378
rect 394778 -16434 394982 -16378
rect 395038 -16434 395124 -16378
rect 395180 -16434 395385 -16378
rect 395441 -16434 395527 -16378
rect 395583 -16434 395779 -16378
rect 395835 -16434 395921 -16378
rect 395977 -16434 396180 -16378
rect 396236 -16434 396322 -16378
rect 396378 -16434 396580 -16378
rect 396636 -16434 396722 -16378
rect 396778 -16434 396977 -16378
rect 397033 -16434 397119 -16378
rect 397175 -16434 397374 -16378
rect 397430 -16434 397516 -16378
rect 397572 -16434 397778 -16378
rect 397834 -16434 397920 -16378
rect 397976 -16434 398174 -16378
rect 398230 -16434 398316 -16378
rect 398372 -16434 398574 -16378
rect 398630 -16434 398716 -16378
rect 398772 -16434 398971 -16378
rect 399027 -16434 399113 -16378
rect 399169 -16434 399376 -16378
rect 399432 -16434 399518 -16378
rect 399574 -16434 399776 -16378
rect 399832 -16434 399918 -16378
rect 399974 -16434 400181 -16378
rect 400237 -16434 400323 -16378
rect 400379 -16416 400766 -16378
rect 400822 -16416 400890 -16360
rect 400946 -16416 401014 -16360
rect 401070 -16416 401138 -16360
rect 401194 -16416 401262 -16360
rect 401318 -16416 402640 -16360
rect 400379 -16434 402640 -16416
rect 387840 -16484 402640 -16434
rect 387840 -16540 387954 -16484
rect 388010 -16540 388078 -16484
rect 388134 -16540 388202 -16484
rect 388258 -16540 388326 -16484
rect 388382 -16540 388450 -16484
rect 388506 -16520 400766 -16484
rect 388506 -16540 388981 -16520
rect 387840 -16576 388981 -16540
rect 389037 -16576 389123 -16520
rect 389179 -16576 389382 -16520
rect 389438 -16576 389524 -16520
rect 389580 -16576 389782 -16520
rect 389838 -16576 389924 -16520
rect 389980 -16576 390179 -16520
rect 390235 -16576 390321 -16520
rect 390377 -16576 390576 -16520
rect 390632 -16576 390718 -16520
rect 390774 -16576 390980 -16520
rect 391036 -16576 391122 -16520
rect 391178 -16576 391376 -16520
rect 391432 -16576 391518 -16520
rect 391574 -16576 391776 -16520
rect 391832 -16576 391918 -16520
rect 391974 -16576 392173 -16520
rect 392229 -16576 392315 -16520
rect 392371 -16576 392578 -16520
rect 392634 -16576 392720 -16520
rect 392776 -16576 392978 -16520
rect 393034 -16576 393120 -16520
rect 393176 -16576 393383 -16520
rect 393439 -16576 393525 -16520
rect 393581 -16576 393780 -16520
rect 393836 -16576 393922 -16520
rect 393978 -16576 394177 -16520
rect 394233 -16576 394319 -16520
rect 394375 -16576 394580 -16520
rect 394636 -16576 394722 -16520
rect 394778 -16576 394982 -16520
rect 395038 -16576 395124 -16520
rect 395180 -16576 395385 -16520
rect 395441 -16576 395527 -16520
rect 395583 -16576 395779 -16520
rect 395835 -16576 395921 -16520
rect 395977 -16576 396180 -16520
rect 396236 -16576 396322 -16520
rect 396378 -16576 396580 -16520
rect 396636 -16576 396722 -16520
rect 396778 -16576 396977 -16520
rect 397033 -16576 397119 -16520
rect 397175 -16576 397374 -16520
rect 397430 -16576 397516 -16520
rect 397572 -16576 397778 -16520
rect 397834 -16576 397920 -16520
rect 397976 -16576 398174 -16520
rect 398230 -16576 398316 -16520
rect 398372 -16576 398574 -16520
rect 398630 -16576 398716 -16520
rect 398772 -16576 398971 -16520
rect 399027 -16576 399113 -16520
rect 399169 -16576 399376 -16520
rect 399432 -16576 399518 -16520
rect 399574 -16576 399776 -16520
rect 399832 -16576 399918 -16520
rect 399974 -16576 400181 -16520
rect 400237 -16576 400323 -16520
rect 400379 -16540 400766 -16520
rect 400822 -16540 400890 -16484
rect 400946 -16540 401014 -16484
rect 401070 -16540 401138 -16484
rect 401194 -16540 401262 -16484
rect 401318 -16540 402640 -16484
rect 400379 -16576 402640 -16540
rect 387840 -16608 402640 -16576
rect 387840 -16664 387954 -16608
rect 388010 -16664 388078 -16608
rect 388134 -16664 388202 -16608
rect 388258 -16664 388326 -16608
rect 388382 -16664 388450 -16608
rect 388506 -16662 400766 -16608
rect 388506 -16664 388981 -16662
rect 387840 -16718 388981 -16664
rect 389037 -16718 389123 -16662
rect 389179 -16718 389382 -16662
rect 389438 -16718 389524 -16662
rect 389580 -16718 389782 -16662
rect 389838 -16718 389924 -16662
rect 389980 -16718 390179 -16662
rect 390235 -16718 390321 -16662
rect 390377 -16718 390576 -16662
rect 390632 -16718 390718 -16662
rect 390774 -16718 390980 -16662
rect 391036 -16718 391122 -16662
rect 391178 -16718 391376 -16662
rect 391432 -16718 391518 -16662
rect 391574 -16718 391776 -16662
rect 391832 -16718 391918 -16662
rect 391974 -16718 392173 -16662
rect 392229 -16718 392315 -16662
rect 392371 -16718 392578 -16662
rect 392634 -16718 392720 -16662
rect 392776 -16718 392978 -16662
rect 393034 -16718 393120 -16662
rect 393176 -16718 393383 -16662
rect 393439 -16718 393525 -16662
rect 393581 -16718 393780 -16662
rect 393836 -16718 393922 -16662
rect 393978 -16718 394177 -16662
rect 394233 -16718 394319 -16662
rect 394375 -16718 394580 -16662
rect 394636 -16718 394722 -16662
rect 394778 -16718 394982 -16662
rect 395038 -16718 395124 -16662
rect 395180 -16718 395385 -16662
rect 395441 -16718 395527 -16662
rect 395583 -16718 395779 -16662
rect 395835 -16718 395921 -16662
rect 395977 -16718 396180 -16662
rect 396236 -16718 396322 -16662
rect 396378 -16718 396580 -16662
rect 396636 -16718 396722 -16662
rect 396778 -16718 396977 -16662
rect 397033 -16718 397119 -16662
rect 397175 -16718 397374 -16662
rect 397430 -16718 397516 -16662
rect 397572 -16718 397778 -16662
rect 397834 -16718 397920 -16662
rect 397976 -16718 398174 -16662
rect 398230 -16718 398316 -16662
rect 398372 -16718 398574 -16662
rect 398630 -16718 398716 -16662
rect 398772 -16718 398971 -16662
rect 399027 -16718 399113 -16662
rect 399169 -16718 399376 -16662
rect 399432 -16718 399518 -16662
rect 399574 -16718 399776 -16662
rect 399832 -16718 399918 -16662
rect 399974 -16718 400181 -16662
rect 400237 -16718 400323 -16662
rect 400379 -16664 400766 -16662
rect 400822 -16664 400890 -16608
rect 400946 -16664 401014 -16608
rect 401070 -16664 401138 -16608
rect 401194 -16664 401262 -16608
rect 401318 -16664 402640 -16608
rect 400379 -16718 402640 -16664
rect 387840 -16732 402640 -16718
rect 387840 -16788 387954 -16732
rect 388010 -16788 388078 -16732
rect 388134 -16788 388202 -16732
rect 388258 -16788 388326 -16732
rect 388382 -16788 388450 -16732
rect 388506 -16788 400766 -16732
rect 400822 -16788 400890 -16732
rect 400946 -16788 401014 -16732
rect 401070 -16788 401138 -16732
rect 401194 -16788 401262 -16732
rect 401318 -16788 402640 -16732
rect 387840 -16804 402640 -16788
rect 387840 -16856 388981 -16804
rect 387840 -16912 387954 -16856
rect 388010 -16912 388078 -16856
rect 388134 -16912 388202 -16856
rect 388258 -16912 388326 -16856
rect 388382 -16912 388450 -16856
rect 388506 -16860 388981 -16856
rect 389037 -16860 389123 -16804
rect 389179 -16860 389382 -16804
rect 389438 -16860 389524 -16804
rect 389580 -16860 389782 -16804
rect 389838 -16860 389924 -16804
rect 389980 -16860 390179 -16804
rect 390235 -16860 390321 -16804
rect 390377 -16860 390576 -16804
rect 390632 -16860 390718 -16804
rect 390774 -16860 390980 -16804
rect 391036 -16860 391122 -16804
rect 391178 -16860 391376 -16804
rect 391432 -16860 391518 -16804
rect 391574 -16860 391776 -16804
rect 391832 -16860 391918 -16804
rect 391974 -16860 392173 -16804
rect 392229 -16860 392315 -16804
rect 392371 -16860 392578 -16804
rect 392634 -16860 392720 -16804
rect 392776 -16860 392978 -16804
rect 393034 -16860 393120 -16804
rect 393176 -16860 393383 -16804
rect 393439 -16860 393525 -16804
rect 393581 -16860 393780 -16804
rect 393836 -16860 393922 -16804
rect 393978 -16860 394177 -16804
rect 394233 -16860 394319 -16804
rect 394375 -16860 394580 -16804
rect 394636 -16860 394722 -16804
rect 394778 -16860 394982 -16804
rect 395038 -16860 395124 -16804
rect 395180 -16860 395385 -16804
rect 395441 -16860 395527 -16804
rect 395583 -16860 395779 -16804
rect 395835 -16860 395921 -16804
rect 395977 -16860 396180 -16804
rect 396236 -16860 396322 -16804
rect 396378 -16860 396580 -16804
rect 396636 -16860 396722 -16804
rect 396778 -16860 396977 -16804
rect 397033 -16860 397119 -16804
rect 397175 -16860 397374 -16804
rect 397430 -16860 397516 -16804
rect 397572 -16860 397778 -16804
rect 397834 -16860 397920 -16804
rect 397976 -16860 398174 -16804
rect 398230 -16860 398316 -16804
rect 398372 -16860 398574 -16804
rect 398630 -16860 398716 -16804
rect 398772 -16860 398971 -16804
rect 399027 -16860 399113 -16804
rect 399169 -16860 399376 -16804
rect 399432 -16860 399518 -16804
rect 399574 -16860 399776 -16804
rect 399832 -16860 399918 -16804
rect 399974 -16860 400181 -16804
rect 400237 -16860 400323 -16804
rect 400379 -16856 402640 -16804
rect 400379 -16860 400766 -16856
rect 388506 -16912 400766 -16860
rect 400822 -16912 400890 -16856
rect 400946 -16912 401014 -16856
rect 401070 -16912 401138 -16856
rect 401194 -16912 401262 -16856
rect 401318 -16912 402640 -16856
rect 387840 -16946 402640 -16912
rect 387840 -16980 388981 -16946
rect 387840 -17036 387954 -16980
rect 388010 -17036 388078 -16980
rect 388134 -17036 388202 -16980
rect 388258 -17036 388326 -16980
rect 388382 -17036 388450 -16980
rect 388506 -17002 388981 -16980
rect 389037 -17002 389123 -16946
rect 389179 -17002 389382 -16946
rect 389438 -17002 389524 -16946
rect 389580 -17002 389782 -16946
rect 389838 -17002 389924 -16946
rect 389980 -17002 390179 -16946
rect 390235 -17002 390321 -16946
rect 390377 -17002 390576 -16946
rect 390632 -17002 390718 -16946
rect 390774 -17002 390980 -16946
rect 391036 -17002 391122 -16946
rect 391178 -17002 391376 -16946
rect 391432 -17002 391518 -16946
rect 391574 -17002 391776 -16946
rect 391832 -17002 391918 -16946
rect 391974 -17002 392173 -16946
rect 392229 -17002 392315 -16946
rect 392371 -17002 392578 -16946
rect 392634 -17002 392720 -16946
rect 392776 -17002 392978 -16946
rect 393034 -17002 393120 -16946
rect 393176 -17002 393383 -16946
rect 393439 -17002 393525 -16946
rect 393581 -17002 393780 -16946
rect 393836 -17002 393922 -16946
rect 393978 -17002 394177 -16946
rect 394233 -17002 394319 -16946
rect 394375 -17002 394580 -16946
rect 394636 -17002 394722 -16946
rect 394778 -17002 394982 -16946
rect 395038 -17002 395124 -16946
rect 395180 -17002 395385 -16946
rect 395441 -17002 395527 -16946
rect 395583 -17002 395779 -16946
rect 395835 -17002 395921 -16946
rect 395977 -17002 396180 -16946
rect 396236 -17002 396322 -16946
rect 396378 -17002 396580 -16946
rect 396636 -17002 396722 -16946
rect 396778 -17002 396977 -16946
rect 397033 -17002 397119 -16946
rect 397175 -17002 397374 -16946
rect 397430 -17002 397516 -16946
rect 397572 -17002 397778 -16946
rect 397834 -17002 397920 -16946
rect 397976 -17002 398174 -16946
rect 398230 -17002 398316 -16946
rect 398372 -17002 398574 -16946
rect 398630 -17002 398716 -16946
rect 398772 -17002 398971 -16946
rect 399027 -17002 399113 -16946
rect 399169 -17002 399376 -16946
rect 399432 -17002 399518 -16946
rect 399574 -17002 399776 -16946
rect 399832 -17002 399918 -16946
rect 399974 -17002 400181 -16946
rect 400237 -17002 400323 -16946
rect 400379 -16980 402640 -16946
rect 400379 -17002 400766 -16980
rect 388506 -17036 400766 -17002
rect 400822 -17036 400890 -16980
rect 400946 -17036 401014 -16980
rect 401070 -17036 401138 -16980
rect 401194 -17036 401262 -16980
rect 401318 -17036 402640 -16980
rect 387840 -17088 402640 -17036
rect 387840 -17104 388981 -17088
rect 387840 -17160 387954 -17104
rect 388010 -17160 388078 -17104
rect 388134 -17160 388202 -17104
rect 388258 -17160 388326 -17104
rect 388382 -17160 388450 -17104
rect 388506 -17144 388981 -17104
rect 389037 -17144 389123 -17088
rect 389179 -17144 389382 -17088
rect 389438 -17144 389524 -17088
rect 389580 -17144 389782 -17088
rect 389838 -17144 389924 -17088
rect 389980 -17144 390179 -17088
rect 390235 -17144 390321 -17088
rect 390377 -17144 390576 -17088
rect 390632 -17144 390718 -17088
rect 390774 -17144 390980 -17088
rect 391036 -17144 391122 -17088
rect 391178 -17144 391376 -17088
rect 391432 -17144 391518 -17088
rect 391574 -17144 391776 -17088
rect 391832 -17144 391918 -17088
rect 391974 -17144 392173 -17088
rect 392229 -17144 392315 -17088
rect 392371 -17144 392578 -17088
rect 392634 -17144 392720 -17088
rect 392776 -17144 392978 -17088
rect 393034 -17144 393120 -17088
rect 393176 -17144 393383 -17088
rect 393439 -17144 393525 -17088
rect 393581 -17144 393780 -17088
rect 393836 -17144 393922 -17088
rect 393978 -17144 394177 -17088
rect 394233 -17144 394319 -17088
rect 394375 -17144 394580 -17088
rect 394636 -17144 394722 -17088
rect 394778 -17144 394982 -17088
rect 395038 -17144 395124 -17088
rect 395180 -17144 395385 -17088
rect 395441 -17144 395527 -17088
rect 395583 -17144 395779 -17088
rect 395835 -17144 395921 -17088
rect 395977 -17144 396180 -17088
rect 396236 -17144 396322 -17088
rect 396378 -17144 396580 -17088
rect 396636 -17144 396722 -17088
rect 396778 -17144 396977 -17088
rect 397033 -17144 397119 -17088
rect 397175 -17144 397374 -17088
rect 397430 -17144 397516 -17088
rect 397572 -17144 397778 -17088
rect 397834 -17144 397920 -17088
rect 397976 -17144 398174 -17088
rect 398230 -17144 398316 -17088
rect 398372 -17144 398574 -17088
rect 398630 -17144 398716 -17088
rect 398772 -17144 398971 -17088
rect 399027 -17144 399113 -17088
rect 399169 -17144 399376 -17088
rect 399432 -17144 399518 -17088
rect 399574 -17144 399776 -17088
rect 399832 -17144 399918 -17088
rect 399974 -17144 400181 -17088
rect 400237 -17144 400323 -17088
rect 400379 -17104 402640 -17088
rect 400379 -17144 400766 -17104
rect 388506 -17160 400766 -17144
rect 400822 -17160 400890 -17104
rect 400946 -17160 401014 -17104
rect 401070 -17160 401138 -17104
rect 401194 -17160 401262 -17104
rect 401318 -17160 402640 -17104
rect 387840 -17228 402640 -17160
rect 387840 -17284 387954 -17228
rect 388010 -17284 388078 -17228
rect 388134 -17284 388202 -17228
rect 388258 -17284 388326 -17228
rect 388382 -17284 388450 -17228
rect 388506 -17230 400766 -17228
rect 388506 -17284 388981 -17230
rect 387840 -17286 388981 -17284
rect 389037 -17286 389123 -17230
rect 389179 -17286 389382 -17230
rect 389438 -17286 389524 -17230
rect 389580 -17286 389782 -17230
rect 389838 -17286 389924 -17230
rect 389980 -17286 390179 -17230
rect 390235 -17286 390321 -17230
rect 390377 -17286 390576 -17230
rect 390632 -17286 390718 -17230
rect 390774 -17286 390980 -17230
rect 391036 -17286 391122 -17230
rect 391178 -17286 391376 -17230
rect 391432 -17286 391518 -17230
rect 391574 -17286 391776 -17230
rect 391832 -17286 391918 -17230
rect 391974 -17286 392173 -17230
rect 392229 -17286 392315 -17230
rect 392371 -17286 392578 -17230
rect 392634 -17286 392720 -17230
rect 392776 -17286 392978 -17230
rect 393034 -17286 393120 -17230
rect 393176 -17286 393383 -17230
rect 393439 -17286 393525 -17230
rect 393581 -17286 393780 -17230
rect 393836 -17286 393922 -17230
rect 393978 -17286 394177 -17230
rect 394233 -17286 394319 -17230
rect 394375 -17286 394580 -17230
rect 394636 -17286 394722 -17230
rect 394778 -17286 394982 -17230
rect 395038 -17286 395124 -17230
rect 395180 -17286 395385 -17230
rect 395441 -17286 395527 -17230
rect 395583 -17286 395779 -17230
rect 395835 -17286 395921 -17230
rect 395977 -17286 396180 -17230
rect 396236 -17286 396322 -17230
rect 396378 -17286 396580 -17230
rect 396636 -17286 396722 -17230
rect 396778 -17286 396977 -17230
rect 397033 -17286 397119 -17230
rect 397175 -17286 397374 -17230
rect 397430 -17286 397516 -17230
rect 397572 -17286 397778 -17230
rect 397834 -17286 397920 -17230
rect 397976 -17286 398174 -17230
rect 398230 -17286 398316 -17230
rect 398372 -17286 398574 -17230
rect 398630 -17286 398716 -17230
rect 398772 -17286 398971 -17230
rect 399027 -17286 399113 -17230
rect 399169 -17286 399376 -17230
rect 399432 -17286 399518 -17230
rect 399574 -17286 399776 -17230
rect 399832 -17286 399918 -17230
rect 399974 -17286 400181 -17230
rect 400237 -17286 400323 -17230
rect 400379 -17284 400766 -17230
rect 400822 -17284 400890 -17228
rect 400946 -17284 401014 -17228
rect 401070 -17284 401138 -17228
rect 401194 -17284 401262 -17228
rect 401318 -17284 402640 -17228
rect 400379 -17286 402640 -17284
rect 387840 -17352 402640 -17286
rect 387840 -17408 387954 -17352
rect 388010 -17408 388078 -17352
rect 388134 -17408 388202 -17352
rect 388258 -17408 388326 -17352
rect 388382 -17408 388450 -17352
rect 388506 -17372 400766 -17352
rect 388506 -17408 388981 -17372
rect 387840 -17428 388981 -17408
rect 389037 -17428 389123 -17372
rect 389179 -17428 389382 -17372
rect 389438 -17428 389524 -17372
rect 389580 -17428 389782 -17372
rect 389838 -17428 389924 -17372
rect 389980 -17428 390179 -17372
rect 390235 -17428 390321 -17372
rect 390377 -17428 390576 -17372
rect 390632 -17428 390718 -17372
rect 390774 -17428 390980 -17372
rect 391036 -17428 391122 -17372
rect 391178 -17428 391376 -17372
rect 391432 -17428 391518 -17372
rect 391574 -17428 391776 -17372
rect 391832 -17428 391918 -17372
rect 391974 -17428 392173 -17372
rect 392229 -17428 392315 -17372
rect 392371 -17428 392578 -17372
rect 392634 -17428 392720 -17372
rect 392776 -17428 392978 -17372
rect 393034 -17428 393120 -17372
rect 393176 -17428 393383 -17372
rect 393439 -17428 393525 -17372
rect 393581 -17428 393780 -17372
rect 393836 -17428 393922 -17372
rect 393978 -17428 394177 -17372
rect 394233 -17428 394319 -17372
rect 394375 -17428 394580 -17372
rect 394636 -17428 394722 -17372
rect 394778 -17428 394982 -17372
rect 395038 -17428 395124 -17372
rect 395180 -17428 395385 -17372
rect 395441 -17428 395527 -17372
rect 395583 -17428 395779 -17372
rect 395835 -17428 395921 -17372
rect 395977 -17428 396180 -17372
rect 396236 -17428 396322 -17372
rect 396378 -17428 396580 -17372
rect 396636 -17428 396722 -17372
rect 396778 -17428 396977 -17372
rect 397033 -17428 397119 -17372
rect 397175 -17428 397374 -17372
rect 397430 -17428 397516 -17372
rect 397572 -17428 397778 -17372
rect 397834 -17428 397920 -17372
rect 397976 -17428 398174 -17372
rect 398230 -17428 398316 -17372
rect 398372 -17428 398574 -17372
rect 398630 -17428 398716 -17372
rect 398772 -17428 398971 -17372
rect 399027 -17428 399113 -17372
rect 399169 -17428 399376 -17372
rect 399432 -17428 399518 -17372
rect 399574 -17428 399776 -17372
rect 399832 -17428 399918 -17372
rect 399974 -17428 400181 -17372
rect 400237 -17428 400323 -17372
rect 400379 -17408 400766 -17372
rect 400822 -17408 400890 -17352
rect 400946 -17408 401014 -17352
rect 401070 -17408 401138 -17352
rect 401194 -17408 401262 -17352
rect 401318 -17408 402640 -17352
rect 400379 -17428 402640 -17408
rect 387840 -17476 402640 -17428
rect 387840 -17532 387954 -17476
rect 388010 -17532 388078 -17476
rect 388134 -17532 388202 -17476
rect 388258 -17532 388326 -17476
rect 388382 -17532 388450 -17476
rect 388506 -17514 400766 -17476
rect 388506 -17532 388981 -17514
rect 387840 -17570 388981 -17532
rect 389037 -17570 389123 -17514
rect 389179 -17570 389382 -17514
rect 389438 -17570 389524 -17514
rect 389580 -17570 389782 -17514
rect 389838 -17570 389924 -17514
rect 389980 -17570 390179 -17514
rect 390235 -17570 390321 -17514
rect 390377 -17570 390576 -17514
rect 390632 -17570 390718 -17514
rect 390774 -17570 390980 -17514
rect 391036 -17570 391122 -17514
rect 391178 -17570 391376 -17514
rect 391432 -17570 391518 -17514
rect 391574 -17570 391776 -17514
rect 391832 -17570 391918 -17514
rect 391974 -17570 392173 -17514
rect 392229 -17570 392315 -17514
rect 392371 -17570 392578 -17514
rect 392634 -17570 392720 -17514
rect 392776 -17570 392978 -17514
rect 393034 -17570 393120 -17514
rect 393176 -17570 393383 -17514
rect 393439 -17570 393525 -17514
rect 393581 -17570 393780 -17514
rect 393836 -17570 393922 -17514
rect 393978 -17570 394177 -17514
rect 394233 -17570 394319 -17514
rect 394375 -17570 394580 -17514
rect 394636 -17570 394722 -17514
rect 394778 -17570 394982 -17514
rect 395038 -17570 395124 -17514
rect 395180 -17570 395385 -17514
rect 395441 -17570 395527 -17514
rect 395583 -17570 395779 -17514
rect 395835 -17570 395921 -17514
rect 395977 -17570 396180 -17514
rect 396236 -17570 396322 -17514
rect 396378 -17570 396580 -17514
rect 396636 -17570 396722 -17514
rect 396778 -17570 396977 -17514
rect 397033 -17570 397119 -17514
rect 397175 -17570 397374 -17514
rect 397430 -17570 397516 -17514
rect 397572 -17570 397778 -17514
rect 397834 -17570 397920 -17514
rect 397976 -17570 398174 -17514
rect 398230 -17570 398316 -17514
rect 398372 -17570 398574 -17514
rect 398630 -17570 398716 -17514
rect 398772 -17570 398971 -17514
rect 399027 -17570 399113 -17514
rect 399169 -17570 399376 -17514
rect 399432 -17570 399518 -17514
rect 399574 -17570 399776 -17514
rect 399832 -17570 399918 -17514
rect 399974 -17570 400181 -17514
rect 400237 -17570 400323 -17514
rect 400379 -17532 400766 -17514
rect 400822 -17532 400890 -17476
rect 400946 -17532 401014 -17476
rect 401070 -17532 401138 -17476
rect 401194 -17532 401262 -17476
rect 401318 -17532 402640 -17476
rect 400379 -17570 402640 -17532
rect 387840 -17600 402640 -17570
rect 387840 -17656 387954 -17600
rect 388010 -17656 388078 -17600
rect 388134 -17656 388202 -17600
rect 388258 -17656 388326 -17600
rect 388382 -17656 388450 -17600
rect 388506 -17656 400766 -17600
rect 400822 -17656 400890 -17600
rect 400946 -17656 401014 -17600
rect 401070 -17656 401138 -17600
rect 401194 -17656 401262 -17600
rect 401318 -17656 402640 -17600
rect 387840 -17712 388981 -17656
rect 389037 -17712 389123 -17656
rect 389179 -17712 389382 -17656
rect 389438 -17712 389524 -17656
rect 389580 -17712 389782 -17656
rect 389838 -17712 389924 -17656
rect 389980 -17712 390179 -17656
rect 390235 -17712 390321 -17656
rect 390377 -17712 390576 -17656
rect 390632 -17712 390718 -17656
rect 390774 -17712 390980 -17656
rect 391036 -17712 391122 -17656
rect 391178 -17712 391376 -17656
rect 391432 -17712 391518 -17656
rect 391574 -17712 391776 -17656
rect 391832 -17712 391918 -17656
rect 391974 -17712 392173 -17656
rect 392229 -17712 392315 -17656
rect 392371 -17712 392578 -17656
rect 392634 -17712 392720 -17656
rect 392776 -17712 392978 -17656
rect 393034 -17712 393120 -17656
rect 393176 -17712 393383 -17656
rect 393439 -17712 393525 -17656
rect 393581 -17712 393780 -17656
rect 393836 -17712 393922 -17656
rect 393978 -17712 394177 -17656
rect 394233 -17712 394319 -17656
rect 394375 -17712 394580 -17656
rect 394636 -17712 394722 -17656
rect 394778 -17712 394982 -17656
rect 395038 -17712 395124 -17656
rect 395180 -17712 395385 -17656
rect 395441 -17712 395527 -17656
rect 395583 -17712 395779 -17656
rect 395835 -17712 395921 -17656
rect 395977 -17712 396180 -17656
rect 396236 -17712 396322 -17656
rect 396378 -17712 396580 -17656
rect 396636 -17712 396722 -17656
rect 396778 -17712 396977 -17656
rect 397033 -17712 397119 -17656
rect 397175 -17712 397374 -17656
rect 397430 -17712 397516 -17656
rect 397572 -17712 397778 -17656
rect 397834 -17712 397920 -17656
rect 397976 -17712 398174 -17656
rect 398230 -17712 398316 -17656
rect 398372 -17712 398574 -17656
rect 398630 -17712 398716 -17656
rect 398772 -17712 398971 -17656
rect 399027 -17712 399113 -17656
rect 399169 -17712 399376 -17656
rect 399432 -17712 399518 -17656
rect 399574 -17712 399776 -17656
rect 399832 -17712 399918 -17656
rect 399974 -17712 400181 -17656
rect 400237 -17712 400323 -17656
rect 400379 -17712 402640 -17656
rect 387840 -17724 402640 -17712
rect 387840 -17780 387954 -17724
rect 388010 -17780 388078 -17724
rect 388134 -17780 388202 -17724
rect 388258 -17780 388326 -17724
rect 388382 -17780 388450 -17724
rect 388506 -17780 400766 -17724
rect 400822 -17780 400890 -17724
rect 400946 -17780 401014 -17724
rect 401070 -17780 401138 -17724
rect 401194 -17780 401262 -17724
rect 401318 -17780 402640 -17724
rect 387840 -17798 402640 -17780
rect 387840 -17848 388981 -17798
rect 387840 -17904 387954 -17848
rect 388010 -17904 388078 -17848
rect 388134 -17904 388202 -17848
rect 388258 -17904 388326 -17848
rect 388382 -17904 388450 -17848
rect 388506 -17854 388981 -17848
rect 389037 -17854 389123 -17798
rect 389179 -17854 389382 -17798
rect 389438 -17854 389524 -17798
rect 389580 -17854 389782 -17798
rect 389838 -17854 389924 -17798
rect 389980 -17854 390179 -17798
rect 390235 -17854 390321 -17798
rect 390377 -17854 390576 -17798
rect 390632 -17854 390718 -17798
rect 390774 -17854 390980 -17798
rect 391036 -17854 391122 -17798
rect 391178 -17854 391376 -17798
rect 391432 -17854 391518 -17798
rect 391574 -17854 391776 -17798
rect 391832 -17854 391918 -17798
rect 391974 -17854 392173 -17798
rect 392229 -17854 392315 -17798
rect 392371 -17854 392578 -17798
rect 392634 -17854 392720 -17798
rect 392776 -17854 392978 -17798
rect 393034 -17854 393120 -17798
rect 393176 -17854 393383 -17798
rect 393439 -17854 393525 -17798
rect 393581 -17854 393780 -17798
rect 393836 -17854 393922 -17798
rect 393978 -17854 394177 -17798
rect 394233 -17854 394319 -17798
rect 394375 -17854 394580 -17798
rect 394636 -17854 394722 -17798
rect 394778 -17854 394982 -17798
rect 395038 -17854 395124 -17798
rect 395180 -17854 395385 -17798
rect 395441 -17854 395527 -17798
rect 395583 -17854 395779 -17798
rect 395835 -17854 395921 -17798
rect 395977 -17854 396180 -17798
rect 396236 -17854 396322 -17798
rect 396378 -17854 396580 -17798
rect 396636 -17854 396722 -17798
rect 396778 -17854 396977 -17798
rect 397033 -17854 397119 -17798
rect 397175 -17854 397374 -17798
rect 397430 -17854 397516 -17798
rect 397572 -17854 397778 -17798
rect 397834 -17854 397920 -17798
rect 397976 -17854 398174 -17798
rect 398230 -17854 398316 -17798
rect 398372 -17854 398574 -17798
rect 398630 -17854 398716 -17798
rect 398772 -17854 398971 -17798
rect 399027 -17854 399113 -17798
rect 399169 -17854 399376 -17798
rect 399432 -17854 399518 -17798
rect 399574 -17854 399776 -17798
rect 399832 -17854 399918 -17798
rect 399974 -17854 400181 -17798
rect 400237 -17854 400323 -17798
rect 400379 -17848 402640 -17798
rect 400379 -17854 400766 -17848
rect 388506 -17904 400766 -17854
rect 400822 -17904 400890 -17848
rect 400946 -17904 401014 -17848
rect 401070 -17904 401138 -17848
rect 401194 -17904 401262 -17848
rect 401318 -17904 402640 -17848
rect 387840 -17940 402640 -17904
rect 387840 -17972 388981 -17940
rect 387840 -18028 387954 -17972
rect 388010 -18028 388078 -17972
rect 388134 -18028 388202 -17972
rect 388258 -18028 388326 -17972
rect 388382 -18028 388450 -17972
rect 388506 -17996 388981 -17972
rect 389037 -17996 389123 -17940
rect 389179 -17996 389382 -17940
rect 389438 -17996 389524 -17940
rect 389580 -17996 389782 -17940
rect 389838 -17996 389924 -17940
rect 389980 -17996 390179 -17940
rect 390235 -17996 390321 -17940
rect 390377 -17996 390576 -17940
rect 390632 -17996 390718 -17940
rect 390774 -17996 390980 -17940
rect 391036 -17996 391122 -17940
rect 391178 -17996 391376 -17940
rect 391432 -17996 391518 -17940
rect 391574 -17996 391776 -17940
rect 391832 -17996 391918 -17940
rect 391974 -17996 392173 -17940
rect 392229 -17996 392315 -17940
rect 392371 -17996 392578 -17940
rect 392634 -17996 392720 -17940
rect 392776 -17996 392978 -17940
rect 393034 -17996 393120 -17940
rect 393176 -17996 393383 -17940
rect 393439 -17996 393525 -17940
rect 393581 -17996 393780 -17940
rect 393836 -17996 393922 -17940
rect 393978 -17996 394177 -17940
rect 394233 -17996 394319 -17940
rect 394375 -17996 394580 -17940
rect 394636 -17996 394722 -17940
rect 394778 -17996 394982 -17940
rect 395038 -17996 395124 -17940
rect 395180 -17996 395385 -17940
rect 395441 -17996 395527 -17940
rect 395583 -17996 395779 -17940
rect 395835 -17996 395921 -17940
rect 395977 -17996 396180 -17940
rect 396236 -17996 396322 -17940
rect 396378 -17996 396580 -17940
rect 396636 -17996 396722 -17940
rect 396778 -17996 396977 -17940
rect 397033 -17996 397119 -17940
rect 397175 -17996 397374 -17940
rect 397430 -17996 397516 -17940
rect 397572 -17996 397778 -17940
rect 397834 -17996 397920 -17940
rect 397976 -17996 398174 -17940
rect 398230 -17996 398316 -17940
rect 398372 -17996 398574 -17940
rect 398630 -17996 398716 -17940
rect 398772 -17996 398971 -17940
rect 399027 -17996 399113 -17940
rect 399169 -17996 399376 -17940
rect 399432 -17996 399518 -17940
rect 399574 -17996 399776 -17940
rect 399832 -17996 399918 -17940
rect 399974 -17996 400181 -17940
rect 400237 -17996 400323 -17940
rect 400379 -17972 402640 -17940
rect 400379 -17996 400766 -17972
rect 388506 -18028 400766 -17996
rect 400822 -18028 400890 -17972
rect 400946 -18028 401014 -17972
rect 401070 -18028 401138 -17972
rect 401194 -18028 401262 -17972
rect 401318 -18028 402640 -17972
rect 387840 -18082 402640 -18028
rect 387840 -18096 388981 -18082
rect 387840 -18152 387954 -18096
rect 388010 -18152 388078 -18096
rect 388134 -18152 388202 -18096
rect 388258 -18152 388326 -18096
rect 388382 -18152 388450 -18096
rect 388506 -18138 388981 -18096
rect 389037 -18138 389123 -18082
rect 389179 -18138 389382 -18082
rect 389438 -18138 389524 -18082
rect 389580 -18138 389782 -18082
rect 389838 -18138 389924 -18082
rect 389980 -18138 390179 -18082
rect 390235 -18138 390321 -18082
rect 390377 -18138 390576 -18082
rect 390632 -18138 390718 -18082
rect 390774 -18138 390980 -18082
rect 391036 -18138 391122 -18082
rect 391178 -18138 391376 -18082
rect 391432 -18138 391518 -18082
rect 391574 -18138 391776 -18082
rect 391832 -18138 391918 -18082
rect 391974 -18138 392173 -18082
rect 392229 -18138 392315 -18082
rect 392371 -18138 392578 -18082
rect 392634 -18138 392720 -18082
rect 392776 -18138 392978 -18082
rect 393034 -18138 393120 -18082
rect 393176 -18138 393383 -18082
rect 393439 -18138 393525 -18082
rect 393581 -18138 393780 -18082
rect 393836 -18138 393922 -18082
rect 393978 -18138 394177 -18082
rect 394233 -18138 394319 -18082
rect 394375 -18138 394580 -18082
rect 394636 -18138 394722 -18082
rect 394778 -18138 394982 -18082
rect 395038 -18138 395124 -18082
rect 395180 -18138 395385 -18082
rect 395441 -18138 395527 -18082
rect 395583 -18138 395779 -18082
rect 395835 -18138 395921 -18082
rect 395977 -18138 396180 -18082
rect 396236 -18138 396322 -18082
rect 396378 -18138 396580 -18082
rect 396636 -18138 396722 -18082
rect 396778 -18138 396977 -18082
rect 397033 -18138 397119 -18082
rect 397175 -18138 397374 -18082
rect 397430 -18138 397516 -18082
rect 397572 -18138 397778 -18082
rect 397834 -18138 397920 -18082
rect 397976 -18138 398174 -18082
rect 398230 -18138 398316 -18082
rect 398372 -18138 398574 -18082
rect 398630 -18138 398716 -18082
rect 398772 -18138 398971 -18082
rect 399027 -18138 399113 -18082
rect 399169 -18138 399376 -18082
rect 399432 -18138 399518 -18082
rect 399574 -18138 399776 -18082
rect 399832 -18138 399918 -18082
rect 399974 -18138 400181 -18082
rect 400237 -18138 400323 -18082
rect 400379 -18096 402640 -18082
rect 400379 -18138 400766 -18096
rect 388506 -18152 400766 -18138
rect 400822 -18152 400890 -18096
rect 400946 -18152 401014 -18096
rect 401070 -18152 401138 -18096
rect 401194 -18152 401262 -18096
rect 401318 -18152 402640 -18096
rect 387840 -18220 402640 -18152
rect 387840 -18276 387954 -18220
rect 388010 -18276 388078 -18220
rect 388134 -18276 388202 -18220
rect 388258 -18276 388326 -18220
rect 388382 -18276 388450 -18220
rect 388506 -18224 400766 -18220
rect 388506 -18276 388981 -18224
rect 387840 -18280 388981 -18276
rect 389037 -18280 389123 -18224
rect 389179 -18280 389382 -18224
rect 389438 -18280 389524 -18224
rect 389580 -18280 389782 -18224
rect 389838 -18280 389924 -18224
rect 389980 -18280 390179 -18224
rect 390235 -18280 390321 -18224
rect 390377 -18280 390576 -18224
rect 390632 -18280 390718 -18224
rect 390774 -18280 390980 -18224
rect 391036 -18280 391122 -18224
rect 391178 -18280 391376 -18224
rect 391432 -18280 391518 -18224
rect 391574 -18280 391776 -18224
rect 391832 -18280 391918 -18224
rect 391974 -18280 392173 -18224
rect 392229 -18280 392315 -18224
rect 392371 -18280 392578 -18224
rect 392634 -18280 392720 -18224
rect 392776 -18280 392978 -18224
rect 393034 -18280 393120 -18224
rect 393176 -18280 393383 -18224
rect 393439 -18280 393525 -18224
rect 393581 -18280 393780 -18224
rect 393836 -18280 393922 -18224
rect 393978 -18280 394177 -18224
rect 394233 -18280 394319 -18224
rect 394375 -18280 394580 -18224
rect 394636 -18280 394722 -18224
rect 394778 -18280 394982 -18224
rect 395038 -18280 395124 -18224
rect 395180 -18280 395385 -18224
rect 395441 -18280 395527 -18224
rect 395583 -18280 395779 -18224
rect 395835 -18280 395921 -18224
rect 395977 -18280 396180 -18224
rect 396236 -18280 396322 -18224
rect 396378 -18280 396580 -18224
rect 396636 -18280 396722 -18224
rect 396778 -18280 396977 -18224
rect 397033 -18280 397119 -18224
rect 397175 -18280 397374 -18224
rect 397430 -18280 397516 -18224
rect 397572 -18280 397778 -18224
rect 397834 -18280 397920 -18224
rect 397976 -18280 398174 -18224
rect 398230 -18280 398316 -18224
rect 398372 -18280 398574 -18224
rect 398630 -18280 398716 -18224
rect 398772 -18280 398971 -18224
rect 399027 -18280 399113 -18224
rect 399169 -18280 399376 -18224
rect 399432 -18280 399518 -18224
rect 399574 -18280 399776 -18224
rect 399832 -18280 399918 -18224
rect 399974 -18280 400181 -18224
rect 400237 -18280 400323 -18224
rect 400379 -18276 400766 -18224
rect 400822 -18276 400890 -18220
rect 400946 -18276 401014 -18220
rect 401070 -18276 401138 -18220
rect 401194 -18276 401262 -18220
rect 401318 -18276 402640 -18220
rect 400379 -18280 402640 -18276
rect 387840 -18344 402640 -18280
rect 387840 -18400 387954 -18344
rect 388010 -18400 388078 -18344
rect 388134 -18400 388202 -18344
rect 388258 -18400 388326 -18344
rect 388382 -18400 388450 -18344
rect 388506 -18366 400766 -18344
rect 388506 -18400 388981 -18366
rect 387840 -18422 388981 -18400
rect 389037 -18422 389123 -18366
rect 389179 -18422 389382 -18366
rect 389438 -18422 389524 -18366
rect 389580 -18422 389782 -18366
rect 389838 -18422 389924 -18366
rect 389980 -18422 390179 -18366
rect 390235 -18422 390321 -18366
rect 390377 -18422 390576 -18366
rect 390632 -18422 390718 -18366
rect 390774 -18422 390980 -18366
rect 391036 -18422 391122 -18366
rect 391178 -18422 391376 -18366
rect 391432 -18422 391518 -18366
rect 391574 -18422 391776 -18366
rect 391832 -18422 391918 -18366
rect 391974 -18422 392173 -18366
rect 392229 -18422 392315 -18366
rect 392371 -18422 392578 -18366
rect 392634 -18422 392720 -18366
rect 392776 -18422 392978 -18366
rect 393034 -18422 393120 -18366
rect 393176 -18422 393383 -18366
rect 393439 -18422 393525 -18366
rect 393581 -18422 393780 -18366
rect 393836 -18422 393922 -18366
rect 393978 -18422 394177 -18366
rect 394233 -18422 394319 -18366
rect 394375 -18422 394580 -18366
rect 394636 -18422 394722 -18366
rect 394778 -18422 394982 -18366
rect 395038 -18422 395124 -18366
rect 395180 -18422 395385 -18366
rect 395441 -18422 395527 -18366
rect 395583 -18422 395779 -18366
rect 395835 -18422 395921 -18366
rect 395977 -18422 396180 -18366
rect 396236 -18422 396322 -18366
rect 396378 -18422 396580 -18366
rect 396636 -18422 396722 -18366
rect 396778 -18422 396977 -18366
rect 397033 -18422 397119 -18366
rect 397175 -18422 397374 -18366
rect 397430 -18422 397516 -18366
rect 397572 -18422 397778 -18366
rect 397834 -18422 397920 -18366
rect 397976 -18422 398174 -18366
rect 398230 -18422 398316 -18366
rect 398372 -18422 398574 -18366
rect 398630 -18422 398716 -18366
rect 398772 -18422 398971 -18366
rect 399027 -18422 399113 -18366
rect 399169 -18422 399376 -18366
rect 399432 -18422 399518 -18366
rect 399574 -18422 399776 -18366
rect 399832 -18422 399918 -18366
rect 399974 -18422 400181 -18366
rect 400237 -18422 400323 -18366
rect 400379 -18400 400766 -18366
rect 400822 -18400 400890 -18344
rect 400946 -18400 401014 -18344
rect 401070 -18400 401138 -18344
rect 401194 -18400 401262 -18344
rect 401318 -18400 402640 -18344
rect 400379 -18422 402640 -18400
rect 387840 -18468 402640 -18422
rect 387840 -18524 387954 -18468
rect 388010 -18524 388078 -18468
rect 388134 -18524 388202 -18468
rect 388258 -18524 388326 -18468
rect 388382 -18524 388450 -18468
rect 388506 -18508 400766 -18468
rect 388506 -18524 388981 -18508
rect 387840 -18564 388981 -18524
rect 389037 -18564 389123 -18508
rect 389179 -18564 389382 -18508
rect 389438 -18564 389524 -18508
rect 389580 -18564 389782 -18508
rect 389838 -18564 389924 -18508
rect 389980 -18564 390179 -18508
rect 390235 -18564 390321 -18508
rect 390377 -18564 390576 -18508
rect 390632 -18564 390718 -18508
rect 390774 -18564 390980 -18508
rect 391036 -18564 391122 -18508
rect 391178 -18564 391376 -18508
rect 391432 -18564 391518 -18508
rect 391574 -18564 391776 -18508
rect 391832 -18564 391918 -18508
rect 391974 -18564 392173 -18508
rect 392229 -18564 392315 -18508
rect 392371 -18564 392578 -18508
rect 392634 -18564 392720 -18508
rect 392776 -18564 392978 -18508
rect 393034 -18564 393120 -18508
rect 393176 -18564 393383 -18508
rect 393439 -18564 393525 -18508
rect 393581 -18564 393780 -18508
rect 393836 -18564 393922 -18508
rect 393978 -18564 394177 -18508
rect 394233 -18564 394319 -18508
rect 394375 -18564 394580 -18508
rect 394636 -18564 394722 -18508
rect 394778 -18564 394982 -18508
rect 395038 -18564 395124 -18508
rect 395180 -18564 395385 -18508
rect 395441 -18564 395527 -18508
rect 395583 -18564 395779 -18508
rect 395835 -18564 395921 -18508
rect 395977 -18564 396180 -18508
rect 396236 -18564 396322 -18508
rect 396378 -18564 396580 -18508
rect 396636 -18564 396722 -18508
rect 396778 -18564 396977 -18508
rect 397033 -18564 397119 -18508
rect 397175 -18564 397374 -18508
rect 397430 -18564 397516 -18508
rect 397572 -18564 397778 -18508
rect 397834 -18564 397920 -18508
rect 397976 -18564 398174 -18508
rect 398230 -18564 398316 -18508
rect 398372 -18564 398574 -18508
rect 398630 -18564 398716 -18508
rect 398772 -18564 398971 -18508
rect 399027 -18564 399113 -18508
rect 399169 -18564 399376 -18508
rect 399432 -18564 399518 -18508
rect 399574 -18564 399776 -18508
rect 399832 -18564 399918 -18508
rect 399974 -18564 400181 -18508
rect 400237 -18564 400323 -18508
rect 400379 -18524 400766 -18508
rect 400822 -18524 400890 -18468
rect 400946 -18524 401014 -18468
rect 401070 -18524 401138 -18468
rect 401194 -18524 401262 -18468
rect 401318 -18524 402640 -18468
rect 400379 -18564 402640 -18524
rect 387840 -18592 402640 -18564
rect 387840 -18648 387954 -18592
rect 388010 -18648 388078 -18592
rect 388134 -18648 388202 -18592
rect 388258 -18648 388326 -18592
rect 388382 -18648 388450 -18592
rect 388506 -18648 400766 -18592
rect 400822 -18648 400890 -18592
rect 400946 -18648 401014 -18592
rect 401070 -18648 401138 -18592
rect 401194 -18648 401262 -18592
rect 401318 -18648 402640 -18592
rect 387840 -18650 402640 -18648
rect 387840 -18706 388981 -18650
rect 389037 -18706 389123 -18650
rect 389179 -18706 389382 -18650
rect 389438 -18706 389524 -18650
rect 389580 -18706 389782 -18650
rect 389838 -18706 389924 -18650
rect 389980 -18706 390179 -18650
rect 390235 -18706 390321 -18650
rect 390377 -18706 390576 -18650
rect 390632 -18706 390718 -18650
rect 390774 -18706 390980 -18650
rect 391036 -18706 391122 -18650
rect 391178 -18706 391376 -18650
rect 391432 -18706 391518 -18650
rect 391574 -18706 391776 -18650
rect 391832 -18706 391918 -18650
rect 391974 -18706 392173 -18650
rect 392229 -18706 392315 -18650
rect 392371 -18706 392578 -18650
rect 392634 -18706 392720 -18650
rect 392776 -18706 392978 -18650
rect 393034 -18706 393120 -18650
rect 393176 -18706 393383 -18650
rect 393439 -18706 393525 -18650
rect 393581 -18706 393780 -18650
rect 393836 -18706 393922 -18650
rect 393978 -18706 394177 -18650
rect 394233 -18706 394319 -18650
rect 394375 -18706 394580 -18650
rect 394636 -18706 394722 -18650
rect 394778 -18706 394982 -18650
rect 395038 -18706 395124 -18650
rect 395180 -18706 395385 -18650
rect 395441 -18706 395527 -18650
rect 395583 -18706 395779 -18650
rect 395835 -18706 395921 -18650
rect 395977 -18706 396180 -18650
rect 396236 -18706 396322 -18650
rect 396378 -18706 396580 -18650
rect 396636 -18706 396722 -18650
rect 396778 -18706 396977 -18650
rect 397033 -18706 397119 -18650
rect 397175 -18706 397374 -18650
rect 397430 -18706 397516 -18650
rect 397572 -18706 397778 -18650
rect 397834 -18706 397920 -18650
rect 397976 -18706 398174 -18650
rect 398230 -18706 398316 -18650
rect 398372 -18706 398574 -18650
rect 398630 -18706 398716 -18650
rect 398772 -18706 398971 -18650
rect 399027 -18706 399113 -18650
rect 399169 -18706 399376 -18650
rect 399432 -18706 399518 -18650
rect 399574 -18706 399776 -18650
rect 399832 -18706 399918 -18650
rect 399974 -18706 400181 -18650
rect 400237 -18706 400323 -18650
rect 400379 -18706 402640 -18650
rect 387840 -18716 402640 -18706
rect 387840 -18772 387954 -18716
rect 388010 -18772 388078 -18716
rect 388134 -18772 388202 -18716
rect 388258 -18772 388326 -18716
rect 388382 -18772 388450 -18716
rect 388506 -18772 400766 -18716
rect 400822 -18772 400890 -18716
rect 400946 -18772 401014 -18716
rect 401070 -18772 401138 -18716
rect 401194 -18772 401262 -18716
rect 401318 -18772 402640 -18716
rect 387840 -18792 402640 -18772
rect 387840 -18840 388981 -18792
rect 387840 -18896 387954 -18840
rect 388010 -18896 388078 -18840
rect 388134 -18896 388202 -18840
rect 388258 -18896 388326 -18840
rect 388382 -18896 388450 -18840
rect 388506 -18848 388981 -18840
rect 389037 -18848 389123 -18792
rect 389179 -18848 389382 -18792
rect 389438 -18848 389524 -18792
rect 389580 -18848 389782 -18792
rect 389838 -18848 389924 -18792
rect 389980 -18848 390179 -18792
rect 390235 -18848 390321 -18792
rect 390377 -18848 390576 -18792
rect 390632 -18848 390718 -18792
rect 390774 -18848 390980 -18792
rect 391036 -18848 391122 -18792
rect 391178 -18848 391376 -18792
rect 391432 -18848 391518 -18792
rect 391574 -18848 391776 -18792
rect 391832 -18848 391918 -18792
rect 391974 -18848 392173 -18792
rect 392229 -18848 392315 -18792
rect 392371 -18848 392578 -18792
rect 392634 -18848 392720 -18792
rect 392776 -18848 392978 -18792
rect 393034 -18848 393120 -18792
rect 393176 -18848 393383 -18792
rect 393439 -18848 393525 -18792
rect 393581 -18848 393780 -18792
rect 393836 -18848 393922 -18792
rect 393978 -18848 394177 -18792
rect 394233 -18848 394319 -18792
rect 394375 -18848 394580 -18792
rect 394636 -18848 394722 -18792
rect 394778 -18848 394982 -18792
rect 395038 -18848 395124 -18792
rect 395180 -18848 395385 -18792
rect 395441 -18848 395527 -18792
rect 395583 -18848 395779 -18792
rect 395835 -18848 395921 -18792
rect 395977 -18848 396180 -18792
rect 396236 -18848 396322 -18792
rect 396378 -18848 396580 -18792
rect 396636 -18848 396722 -18792
rect 396778 -18848 396977 -18792
rect 397033 -18848 397119 -18792
rect 397175 -18848 397374 -18792
rect 397430 -18848 397516 -18792
rect 397572 -18848 397778 -18792
rect 397834 -18848 397920 -18792
rect 397976 -18848 398174 -18792
rect 398230 -18848 398316 -18792
rect 398372 -18848 398574 -18792
rect 398630 -18848 398716 -18792
rect 398772 -18848 398971 -18792
rect 399027 -18848 399113 -18792
rect 399169 -18848 399376 -18792
rect 399432 -18848 399518 -18792
rect 399574 -18848 399776 -18792
rect 399832 -18848 399918 -18792
rect 399974 -18848 400181 -18792
rect 400237 -18848 400323 -18792
rect 400379 -18840 402640 -18792
rect 400379 -18848 400766 -18840
rect 388506 -18896 400766 -18848
rect 400822 -18896 400890 -18840
rect 400946 -18896 401014 -18840
rect 401070 -18896 401138 -18840
rect 401194 -18896 401262 -18840
rect 401318 -18896 402640 -18840
rect 387840 -18934 402640 -18896
rect 387840 -18964 388981 -18934
rect 387840 -19020 387954 -18964
rect 388010 -19020 388078 -18964
rect 388134 -19020 388202 -18964
rect 388258 -19020 388326 -18964
rect 388382 -19020 388450 -18964
rect 388506 -18990 388981 -18964
rect 389037 -18990 389123 -18934
rect 389179 -18990 389382 -18934
rect 389438 -18990 389524 -18934
rect 389580 -18990 389782 -18934
rect 389838 -18990 389924 -18934
rect 389980 -18990 390179 -18934
rect 390235 -18990 390321 -18934
rect 390377 -18990 390576 -18934
rect 390632 -18990 390718 -18934
rect 390774 -18990 390980 -18934
rect 391036 -18990 391122 -18934
rect 391178 -18990 391376 -18934
rect 391432 -18990 391518 -18934
rect 391574 -18990 391776 -18934
rect 391832 -18990 391918 -18934
rect 391974 -18990 392173 -18934
rect 392229 -18990 392315 -18934
rect 392371 -18990 392578 -18934
rect 392634 -18990 392720 -18934
rect 392776 -18990 392978 -18934
rect 393034 -18990 393120 -18934
rect 393176 -18990 393383 -18934
rect 393439 -18990 393525 -18934
rect 393581 -18990 393780 -18934
rect 393836 -18990 393922 -18934
rect 393978 -18990 394177 -18934
rect 394233 -18990 394319 -18934
rect 394375 -18990 394580 -18934
rect 394636 -18990 394722 -18934
rect 394778 -18990 394982 -18934
rect 395038 -18990 395124 -18934
rect 395180 -18990 395385 -18934
rect 395441 -18990 395527 -18934
rect 395583 -18990 395779 -18934
rect 395835 -18990 395921 -18934
rect 395977 -18990 396180 -18934
rect 396236 -18990 396322 -18934
rect 396378 -18990 396580 -18934
rect 396636 -18990 396722 -18934
rect 396778 -18990 396977 -18934
rect 397033 -18990 397119 -18934
rect 397175 -18990 397374 -18934
rect 397430 -18990 397516 -18934
rect 397572 -18990 397778 -18934
rect 397834 -18990 397920 -18934
rect 397976 -18990 398174 -18934
rect 398230 -18990 398316 -18934
rect 398372 -18990 398574 -18934
rect 398630 -18990 398716 -18934
rect 398772 -18990 398971 -18934
rect 399027 -18990 399113 -18934
rect 399169 -18990 399376 -18934
rect 399432 -18990 399518 -18934
rect 399574 -18990 399776 -18934
rect 399832 -18990 399918 -18934
rect 399974 -18990 400181 -18934
rect 400237 -18990 400323 -18934
rect 400379 -18964 402640 -18934
rect 400379 -18990 400766 -18964
rect 388506 -19020 400766 -18990
rect 400822 -19020 400890 -18964
rect 400946 -19020 401014 -18964
rect 401070 -19020 401138 -18964
rect 401194 -19020 401262 -18964
rect 401318 -19020 402640 -18964
rect 387840 -19076 402640 -19020
rect 387840 -19088 388981 -19076
rect 387840 -19144 387954 -19088
rect 388010 -19144 388078 -19088
rect 388134 -19144 388202 -19088
rect 388258 -19144 388326 -19088
rect 388382 -19144 388450 -19088
rect 388506 -19132 388981 -19088
rect 389037 -19132 389123 -19076
rect 389179 -19132 389382 -19076
rect 389438 -19132 389524 -19076
rect 389580 -19132 389782 -19076
rect 389838 -19132 389924 -19076
rect 389980 -19132 390179 -19076
rect 390235 -19132 390321 -19076
rect 390377 -19132 390576 -19076
rect 390632 -19132 390718 -19076
rect 390774 -19132 390980 -19076
rect 391036 -19132 391122 -19076
rect 391178 -19132 391376 -19076
rect 391432 -19132 391518 -19076
rect 391574 -19132 391776 -19076
rect 391832 -19132 391918 -19076
rect 391974 -19132 392173 -19076
rect 392229 -19132 392315 -19076
rect 392371 -19132 392578 -19076
rect 392634 -19132 392720 -19076
rect 392776 -19132 392978 -19076
rect 393034 -19132 393120 -19076
rect 393176 -19132 393383 -19076
rect 393439 -19132 393525 -19076
rect 393581 -19132 393780 -19076
rect 393836 -19132 393922 -19076
rect 393978 -19132 394177 -19076
rect 394233 -19132 394319 -19076
rect 394375 -19132 394580 -19076
rect 394636 -19132 394722 -19076
rect 394778 -19132 394982 -19076
rect 395038 -19132 395124 -19076
rect 395180 -19132 395385 -19076
rect 395441 -19132 395527 -19076
rect 395583 -19132 395779 -19076
rect 395835 -19132 395921 -19076
rect 395977 -19132 396180 -19076
rect 396236 -19132 396322 -19076
rect 396378 -19132 396580 -19076
rect 396636 -19132 396722 -19076
rect 396778 -19132 396977 -19076
rect 397033 -19132 397119 -19076
rect 397175 -19132 397374 -19076
rect 397430 -19132 397516 -19076
rect 397572 -19132 397778 -19076
rect 397834 -19132 397920 -19076
rect 397976 -19132 398174 -19076
rect 398230 -19132 398316 -19076
rect 398372 -19132 398574 -19076
rect 398630 -19132 398716 -19076
rect 398772 -19132 398971 -19076
rect 399027 -19132 399113 -19076
rect 399169 -19132 399376 -19076
rect 399432 -19132 399518 -19076
rect 399574 -19132 399776 -19076
rect 399832 -19132 399918 -19076
rect 399974 -19132 400181 -19076
rect 400237 -19132 400323 -19076
rect 400379 -19088 402640 -19076
rect 400379 -19132 400766 -19088
rect 388506 -19144 400766 -19132
rect 400822 -19144 400890 -19088
rect 400946 -19144 401014 -19088
rect 401070 -19144 401138 -19088
rect 401194 -19144 401262 -19088
rect 401318 -19144 402640 -19088
rect 387840 -19212 402640 -19144
rect 387840 -19268 387954 -19212
rect 388010 -19268 388078 -19212
rect 388134 -19268 388202 -19212
rect 388258 -19268 388326 -19212
rect 388382 -19268 388450 -19212
rect 388506 -19218 400766 -19212
rect 388506 -19268 388981 -19218
rect 387840 -19274 388981 -19268
rect 389037 -19274 389123 -19218
rect 389179 -19274 389382 -19218
rect 389438 -19274 389524 -19218
rect 389580 -19274 389782 -19218
rect 389838 -19274 389924 -19218
rect 389980 -19274 390179 -19218
rect 390235 -19274 390321 -19218
rect 390377 -19274 390576 -19218
rect 390632 -19274 390718 -19218
rect 390774 -19274 390980 -19218
rect 391036 -19274 391122 -19218
rect 391178 -19274 391376 -19218
rect 391432 -19274 391518 -19218
rect 391574 -19274 391776 -19218
rect 391832 -19274 391918 -19218
rect 391974 -19274 392173 -19218
rect 392229 -19274 392315 -19218
rect 392371 -19274 392578 -19218
rect 392634 -19274 392720 -19218
rect 392776 -19274 392978 -19218
rect 393034 -19274 393120 -19218
rect 393176 -19274 393383 -19218
rect 393439 -19274 393525 -19218
rect 393581 -19274 393780 -19218
rect 393836 -19274 393922 -19218
rect 393978 -19274 394177 -19218
rect 394233 -19274 394319 -19218
rect 394375 -19274 394580 -19218
rect 394636 -19274 394722 -19218
rect 394778 -19274 394982 -19218
rect 395038 -19274 395124 -19218
rect 395180 -19274 395385 -19218
rect 395441 -19274 395527 -19218
rect 395583 -19274 395779 -19218
rect 395835 -19274 395921 -19218
rect 395977 -19274 396180 -19218
rect 396236 -19274 396322 -19218
rect 396378 -19274 396580 -19218
rect 396636 -19274 396722 -19218
rect 396778 -19274 396977 -19218
rect 397033 -19274 397119 -19218
rect 397175 -19274 397374 -19218
rect 397430 -19274 397516 -19218
rect 397572 -19274 397778 -19218
rect 397834 -19274 397920 -19218
rect 397976 -19274 398174 -19218
rect 398230 -19274 398316 -19218
rect 398372 -19274 398574 -19218
rect 398630 -19274 398716 -19218
rect 398772 -19274 398971 -19218
rect 399027 -19274 399113 -19218
rect 399169 -19274 399376 -19218
rect 399432 -19274 399518 -19218
rect 399574 -19274 399776 -19218
rect 399832 -19274 399918 -19218
rect 399974 -19274 400181 -19218
rect 400237 -19274 400323 -19218
rect 400379 -19268 400766 -19218
rect 400822 -19268 400890 -19212
rect 400946 -19268 401014 -19212
rect 401070 -19268 401138 -19212
rect 401194 -19268 401262 -19212
rect 401318 -19268 402640 -19212
rect 400379 -19274 402640 -19268
rect 387840 -19336 402640 -19274
rect 387840 -19392 387954 -19336
rect 388010 -19392 388078 -19336
rect 388134 -19392 388202 -19336
rect 388258 -19392 388326 -19336
rect 388382 -19392 388450 -19336
rect 388506 -19360 400766 -19336
rect 388506 -19392 388981 -19360
rect 387840 -19416 388981 -19392
rect 389037 -19416 389123 -19360
rect 389179 -19416 389382 -19360
rect 389438 -19416 389524 -19360
rect 389580 -19416 389782 -19360
rect 389838 -19416 389924 -19360
rect 389980 -19416 390179 -19360
rect 390235 -19416 390321 -19360
rect 390377 -19416 390576 -19360
rect 390632 -19416 390718 -19360
rect 390774 -19416 390980 -19360
rect 391036 -19416 391122 -19360
rect 391178 -19416 391376 -19360
rect 391432 -19416 391518 -19360
rect 391574 -19416 391776 -19360
rect 391832 -19416 391918 -19360
rect 391974 -19416 392173 -19360
rect 392229 -19416 392315 -19360
rect 392371 -19416 392578 -19360
rect 392634 -19416 392720 -19360
rect 392776 -19416 392978 -19360
rect 393034 -19416 393120 -19360
rect 393176 -19416 393383 -19360
rect 393439 -19416 393525 -19360
rect 393581 -19416 393780 -19360
rect 393836 -19416 393922 -19360
rect 393978 -19416 394177 -19360
rect 394233 -19416 394319 -19360
rect 394375 -19416 394580 -19360
rect 394636 -19416 394722 -19360
rect 394778 -19416 394982 -19360
rect 395038 -19416 395124 -19360
rect 395180 -19416 395385 -19360
rect 395441 -19416 395527 -19360
rect 395583 -19416 395779 -19360
rect 395835 -19416 395921 -19360
rect 395977 -19416 396180 -19360
rect 396236 -19416 396322 -19360
rect 396378 -19416 396580 -19360
rect 396636 -19416 396722 -19360
rect 396778 -19416 396977 -19360
rect 397033 -19416 397119 -19360
rect 397175 -19416 397374 -19360
rect 397430 -19416 397516 -19360
rect 397572 -19416 397778 -19360
rect 397834 -19416 397920 -19360
rect 397976 -19416 398174 -19360
rect 398230 -19416 398316 -19360
rect 398372 -19416 398574 -19360
rect 398630 -19416 398716 -19360
rect 398772 -19416 398971 -19360
rect 399027 -19416 399113 -19360
rect 399169 -19416 399376 -19360
rect 399432 -19416 399518 -19360
rect 399574 -19416 399776 -19360
rect 399832 -19416 399918 -19360
rect 399974 -19416 400181 -19360
rect 400237 -19416 400323 -19360
rect 400379 -19392 400766 -19360
rect 400822 -19392 400890 -19336
rect 400946 -19392 401014 -19336
rect 401070 -19392 401138 -19336
rect 401194 -19392 401262 -19336
rect 401318 -19392 402640 -19336
rect 400379 -19416 402640 -19392
rect 387840 -19460 402640 -19416
rect 387840 -19516 387954 -19460
rect 388010 -19516 388078 -19460
rect 388134 -19516 388202 -19460
rect 388258 -19516 388326 -19460
rect 388382 -19516 388450 -19460
rect 388506 -19502 400766 -19460
rect 388506 -19516 388981 -19502
rect 387840 -19558 388981 -19516
rect 389037 -19558 389123 -19502
rect 389179 -19558 389382 -19502
rect 389438 -19558 389524 -19502
rect 389580 -19558 389782 -19502
rect 389838 -19558 389924 -19502
rect 389980 -19558 390179 -19502
rect 390235 -19558 390321 -19502
rect 390377 -19558 390576 -19502
rect 390632 -19558 390718 -19502
rect 390774 -19558 390980 -19502
rect 391036 -19558 391122 -19502
rect 391178 -19558 391376 -19502
rect 391432 -19558 391518 -19502
rect 391574 -19558 391776 -19502
rect 391832 -19558 391918 -19502
rect 391974 -19558 392173 -19502
rect 392229 -19558 392315 -19502
rect 392371 -19558 392578 -19502
rect 392634 -19558 392720 -19502
rect 392776 -19558 392978 -19502
rect 393034 -19558 393120 -19502
rect 393176 -19558 393383 -19502
rect 393439 -19558 393525 -19502
rect 393581 -19558 393780 -19502
rect 393836 -19558 393922 -19502
rect 393978 -19558 394177 -19502
rect 394233 -19558 394319 -19502
rect 394375 -19558 394580 -19502
rect 394636 -19558 394722 -19502
rect 394778 -19558 394982 -19502
rect 395038 -19558 395124 -19502
rect 395180 -19558 395385 -19502
rect 395441 -19558 395527 -19502
rect 395583 -19558 395779 -19502
rect 395835 -19558 395921 -19502
rect 395977 -19558 396180 -19502
rect 396236 -19558 396322 -19502
rect 396378 -19558 396580 -19502
rect 396636 -19558 396722 -19502
rect 396778 -19558 396977 -19502
rect 397033 -19558 397119 -19502
rect 397175 -19558 397374 -19502
rect 397430 -19558 397516 -19502
rect 397572 -19558 397778 -19502
rect 397834 -19558 397920 -19502
rect 397976 -19558 398174 -19502
rect 398230 -19558 398316 -19502
rect 398372 -19558 398574 -19502
rect 398630 -19558 398716 -19502
rect 398772 -19558 398971 -19502
rect 399027 -19558 399113 -19502
rect 399169 -19558 399376 -19502
rect 399432 -19558 399518 -19502
rect 399574 -19558 399776 -19502
rect 399832 -19558 399918 -19502
rect 399974 -19558 400181 -19502
rect 400237 -19558 400323 -19502
rect 400379 -19516 400766 -19502
rect 400822 -19516 400890 -19460
rect 400946 -19516 401014 -19460
rect 401070 -19516 401138 -19460
rect 401194 -19516 401262 -19460
rect 401318 -19516 402640 -19460
rect 400379 -19558 402640 -19516
rect 387840 -19584 402640 -19558
rect 387840 -19640 387954 -19584
rect 388010 -19640 388078 -19584
rect 388134 -19640 388202 -19584
rect 388258 -19640 388326 -19584
rect 388382 -19640 388450 -19584
rect 388506 -19640 400766 -19584
rect 400822 -19640 400890 -19584
rect 400946 -19640 401014 -19584
rect 401070 -19640 401138 -19584
rect 401194 -19640 401262 -19584
rect 401318 -19640 402640 -19584
rect 387840 -19644 402640 -19640
rect 387840 -19700 388981 -19644
rect 389037 -19700 389123 -19644
rect 389179 -19700 389382 -19644
rect 389438 -19700 389524 -19644
rect 389580 -19700 389782 -19644
rect 389838 -19700 389924 -19644
rect 389980 -19700 390179 -19644
rect 390235 -19700 390321 -19644
rect 390377 -19700 390576 -19644
rect 390632 -19700 390718 -19644
rect 390774 -19700 390980 -19644
rect 391036 -19700 391122 -19644
rect 391178 -19700 391376 -19644
rect 391432 -19700 391518 -19644
rect 391574 -19700 391776 -19644
rect 391832 -19700 391918 -19644
rect 391974 -19700 392173 -19644
rect 392229 -19700 392315 -19644
rect 392371 -19700 392578 -19644
rect 392634 -19700 392720 -19644
rect 392776 -19700 392978 -19644
rect 393034 -19700 393120 -19644
rect 393176 -19700 393383 -19644
rect 393439 -19700 393525 -19644
rect 393581 -19700 393780 -19644
rect 393836 -19700 393922 -19644
rect 393978 -19700 394177 -19644
rect 394233 -19700 394319 -19644
rect 394375 -19700 394580 -19644
rect 394636 -19700 394722 -19644
rect 394778 -19700 394982 -19644
rect 395038 -19700 395124 -19644
rect 395180 -19700 395385 -19644
rect 395441 -19700 395527 -19644
rect 395583 -19700 395779 -19644
rect 395835 -19700 395921 -19644
rect 395977 -19700 396180 -19644
rect 396236 -19700 396322 -19644
rect 396378 -19700 396580 -19644
rect 396636 -19700 396722 -19644
rect 396778 -19700 396977 -19644
rect 397033 -19700 397119 -19644
rect 397175 -19700 397374 -19644
rect 397430 -19700 397516 -19644
rect 397572 -19700 397778 -19644
rect 397834 -19700 397920 -19644
rect 397976 -19700 398174 -19644
rect 398230 -19700 398316 -19644
rect 398372 -19700 398574 -19644
rect 398630 -19700 398716 -19644
rect 398772 -19700 398971 -19644
rect 399027 -19700 399113 -19644
rect 399169 -19700 399376 -19644
rect 399432 -19700 399518 -19644
rect 399574 -19700 399776 -19644
rect 399832 -19700 399918 -19644
rect 399974 -19700 400181 -19644
rect 400237 -19700 400323 -19644
rect 400379 -19700 402640 -19644
rect 387840 -19708 402640 -19700
rect 387840 -19764 387954 -19708
rect 388010 -19764 388078 -19708
rect 388134 -19764 388202 -19708
rect 388258 -19764 388326 -19708
rect 388382 -19764 388450 -19708
rect 388506 -19764 400766 -19708
rect 400822 -19764 400890 -19708
rect 400946 -19764 401014 -19708
rect 401070 -19764 401138 -19708
rect 401194 -19764 401262 -19708
rect 401318 -19764 402640 -19708
rect 387840 -19786 402640 -19764
rect 387840 -19832 388981 -19786
rect 387840 -19888 387954 -19832
rect 388010 -19888 388078 -19832
rect 388134 -19888 388202 -19832
rect 388258 -19888 388326 -19832
rect 388382 -19888 388450 -19832
rect 388506 -19842 388981 -19832
rect 389037 -19842 389123 -19786
rect 389179 -19842 389382 -19786
rect 389438 -19842 389524 -19786
rect 389580 -19842 389782 -19786
rect 389838 -19842 389924 -19786
rect 389980 -19842 390179 -19786
rect 390235 -19842 390321 -19786
rect 390377 -19842 390576 -19786
rect 390632 -19842 390718 -19786
rect 390774 -19842 390980 -19786
rect 391036 -19842 391122 -19786
rect 391178 -19842 391376 -19786
rect 391432 -19842 391518 -19786
rect 391574 -19842 391776 -19786
rect 391832 -19842 391918 -19786
rect 391974 -19842 392173 -19786
rect 392229 -19842 392315 -19786
rect 392371 -19842 392578 -19786
rect 392634 -19842 392720 -19786
rect 392776 -19842 392978 -19786
rect 393034 -19842 393120 -19786
rect 393176 -19842 393383 -19786
rect 393439 -19842 393525 -19786
rect 393581 -19842 393780 -19786
rect 393836 -19842 393922 -19786
rect 393978 -19842 394177 -19786
rect 394233 -19842 394319 -19786
rect 394375 -19842 394580 -19786
rect 394636 -19842 394722 -19786
rect 394778 -19842 394982 -19786
rect 395038 -19842 395124 -19786
rect 395180 -19842 395385 -19786
rect 395441 -19842 395527 -19786
rect 395583 -19842 395779 -19786
rect 395835 -19842 395921 -19786
rect 395977 -19842 396180 -19786
rect 396236 -19842 396322 -19786
rect 396378 -19842 396580 -19786
rect 396636 -19842 396722 -19786
rect 396778 -19842 396977 -19786
rect 397033 -19842 397119 -19786
rect 397175 -19842 397374 -19786
rect 397430 -19842 397516 -19786
rect 397572 -19842 397778 -19786
rect 397834 -19842 397920 -19786
rect 397976 -19842 398174 -19786
rect 398230 -19842 398316 -19786
rect 398372 -19842 398574 -19786
rect 398630 -19842 398716 -19786
rect 398772 -19842 398971 -19786
rect 399027 -19842 399113 -19786
rect 399169 -19842 399376 -19786
rect 399432 -19842 399518 -19786
rect 399574 -19842 399776 -19786
rect 399832 -19842 399918 -19786
rect 399974 -19842 400181 -19786
rect 400237 -19842 400323 -19786
rect 400379 -19832 402640 -19786
rect 400379 -19842 400766 -19832
rect 388506 -19888 400766 -19842
rect 400822 -19888 400890 -19832
rect 400946 -19888 401014 -19832
rect 401070 -19888 401138 -19832
rect 401194 -19888 401262 -19832
rect 401318 -19888 402640 -19832
rect 387840 -19928 402640 -19888
rect 387840 -19956 388981 -19928
rect 387840 -20012 387954 -19956
rect 388010 -20012 388078 -19956
rect 388134 -20012 388202 -19956
rect 388258 -20012 388326 -19956
rect 388382 -20012 388450 -19956
rect 388506 -19984 388981 -19956
rect 389037 -19984 389123 -19928
rect 389179 -19984 389382 -19928
rect 389438 -19984 389524 -19928
rect 389580 -19984 389782 -19928
rect 389838 -19984 389924 -19928
rect 389980 -19984 390179 -19928
rect 390235 -19984 390321 -19928
rect 390377 -19984 390576 -19928
rect 390632 -19984 390718 -19928
rect 390774 -19984 390980 -19928
rect 391036 -19984 391122 -19928
rect 391178 -19984 391376 -19928
rect 391432 -19984 391518 -19928
rect 391574 -19984 391776 -19928
rect 391832 -19984 391918 -19928
rect 391974 -19984 392173 -19928
rect 392229 -19984 392315 -19928
rect 392371 -19984 392578 -19928
rect 392634 -19984 392720 -19928
rect 392776 -19984 392978 -19928
rect 393034 -19984 393120 -19928
rect 393176 -19984 393383 -19928
rect 393439 -19984 393525 -19928
rect 393581 -19984 393780 -19928
rect 393836 -19984 393922 -19928
rect 393978 -19984 394177 -19928
rect 394233 -19984 394319 -19928
rect 394375 -19984 394580 -19928
rect 394636 -19984 394722 -19928
rect 394778 -19984 394982 -19928
rect 395038 -19984 395124 -19928
rect 395180 -19984 395385 -19928
rect 395441 -19984 395527 -19928
rect 395583 -19984 395779 -19928
rect 395835 -19984 395921 -19928
rect 395977 -19984 396180 -19928
rect 396236 -19984 396322 -19928
rect 396378 -19984 396580 -19928
rect 396636 -19984 396722 -19928
rect 396778 -19984 396977 -19928
rect 397033 -19984 397119 -19928
rect 397175 -19984 397374 -19928
rect 397430 -19984 397516 -19928
rect 397572 -19984 397778 -19928
rect 397834 -19984 397920 -19928
rect 397976 -19984 398174 -19928
rect 398230 -19984 398316 -19928
rect 398372 -19984 398574 -19928
rect 398630 -19984 398716 -19928
rect 398772 -19984 398971 -19928
rect 399027 -19984 399113 -19928
rect 399169 -19984 399376 -19928
rect 399432 -19984 399518 -19928
rect 399574 -19984 399776 -19928
rect 399832 -19984 399918 -19928
rect 399974 -19984 400181 -19928
rect 400237 -19984 400323 -19928
rect 400379 -19956 402640 -19928
rect 400379 -19984 400766 -19956
rect 388506 -20012 400766 -19984
rect 400822 -20012 400890 -19956
rect 400946 -20012 401014 -19956
rect 401070 -20012 401138 -19956
rect 401194 -20012 401262 -19956
rect 401318 -20012 402640 -19956
rect 387840 -20070 402640 -20012
rect 387840 -20080 388981 -20070
rect 387840 -20136 387954 -20080
rect 388010 -20136 388078 -20080
rect 388134 -20136 388202 -20080
rect 388258 -20136 388326 -20080
rect 388382 -20136 388450 -20080
rect 388506 -20126 388981 -20080
rect 389037 -20126 389123 -20070
rect 389179 -20126 389382 -20070
rect 389438 -20126 389524 -20070
rect 389580 -20126 389782 -20070
rect 389838 -20126 389924 -20070
rect 389980 -20126 390179 -20070
rect 390235 -20126 390321 -20070
rect 390377 -20126 390576 -20070
rect 390632 -20126 390718 -20070
rect 390774 -20126 390980 -20070
rect 391036 -20126 391122 -20070
rect 391178 -20126 391376 -20070
rect 391432 -20126 391518 -20070
rect 391574 -20126 391776 -20070
rect 391832 -20126 391918 -20070
rect 391974 -20126 392173 -20070
rect 392229 -20126 392315 -20070
rect 392371 -20126 392578 -20070
rect 392634 -20126 392720 -20070
rect 392776 -20126 392978 -20070
rect 393034 -20126 393120 -20070
rect 393176 -20126 393383 -20070
rect 393439 -20126 393525 -20070
rect 393581 -20126 393780 -20070
rect 393836 -20126 393922 -20070
rect 393978 -20126 394177 -20070
rect 394233 -20126 394319 -20070
rect 394375 -20126 394580 -20070
rect 394636 -20126 394722 -20070
rect 394778 -20126 394982 -20070
rect 395038 -20126 395124 -20070
rect 395180 -20126 395385 -20070
rect 395441 -20126 395527 -20070
rect 395583 -20126 395779 -20070
rect 395835 -20126 395921 -20070
rect 395977 -20126 396180 -20070
rect 396236 -20126 396322 -20070
rect 396378 -20126 396580 -20070
rect 396636 -20126 396722 -20070
rect 396778 -20126 396977 -20070
rect 397033 -20126 397119 -20070
rect 397175 -20126 397374 -20070
rect 397430 -20126 397516 -20070
rect 397572 -20126 397778 -20070
rect 397834 -20126 397920 -20070
rect 397976 -20126 398174 -20070
rect 398230 -20126 398316 -20070
rect 398372 -20126 398574 -20070
rect 398630 -20126 398716 -20070
rect 398772 -20126 398971 -20070
rect 399027 -20126 399113 -20070
rect 399169 -20126 399376 -20070
rect 399432 -20126 399518 -20070
rect 399574 -20126 399776 -20070
rect 399832 -20126 399918 -20070
rect 399974 -20126 400181 -20070
rect 400237 -20126 400323 -20070
rect 400379 -20080 402640 -20070
rect 400379 -20126 400766 -20080
rect 388506 -20136 400766 -20126
rect 400822 -20136 400890 -20080
rect 400946 -20136 401014 -20080
rect 401070 -20136 401138 -20080
rect 401194 -20136 401262 -20080
rect 401318 -20136 402640 -20080
rect 387840 -20204 402640 -20136
rect 387840 -20260 387954 -20204
rect 388010 -20260 388078 -20204
rect 388134 -20260 388202 -20204
rect 388258 -20260 388326 -20204
rect 388382 -20260 388450 -20204
rect 388506 -20212 400766 -20204
rect 388506 -20260 388981 -20212
rect 387840 -20268 388981 -20260
rect 389037 -20268 389123 -20212
rect 389179 -20268 389382 -20212
rect 389438 -20268 389524 -20212
rect 389580 -20268 389782 -20212
rect 389838 -20268 389924 -20212
rect 389980 -20268 390179 -20212
rect 390235 -20268 390321 -20212
rect 390377 -20268 390576 -20212
rect 390632 -20268 390718 -20212
rect 390774 -20268 390980 -20212
rect 391036 -20268 391122 -20212
rect 391178 -20268 391376 -20212
rect 391432 -20268 391518 -20212
rect 391574 -20268 391776 -20212
rect 391832 -20268 391918 -20212
rect 391974 -20268 392173 -20212
rect 392229 -20268 392315 -20212
rect 392371 -20268 392578 -20212
rect 392634 -20268 392720 -20212
rect 392776 -20268 392978 -20212
rect 393034 -20268 393120 -20212
rect 393176 -20268 393383 -20212
rect 393439 -20268 393525 -20212
rect 393581 -20268 393780 -20212
rect 393836 -20268 393922 -20212
rect 393978 -20268 394177 -20212
rect 394233 -20268 394319 -20212
rect 394375 -20268 394580 -20212
rect 394636 -20268 394722 -20212
rect 394778 -20268 394982 -20212
rect 395038 -20268 395124 -20212
rect 395180 -20268 395385 -20212
rect 395441 -20268 395527 -20212
rect 395583 -20268 395779 -20212
rect 395835 -20268 395921 -20212
rect 395977 -20268 396180 -20212
rect 396236 -20268 396322 -20212
rect 396378 -20268 396580 -20212
rect 396636 -20268 396722 -20212
rect 396778 -20268 396977 -20212
rect 397033 -20268 397119 -20212
rect 397175 -20268 397374 -20212
rect 397430 -20268 397516 -20212
rect 397572 -20268 397778 -20212
rect 397834 -20268 397920 -20212
rect 397976 -20268 398174 -20212
rect 398230 -20268 398316 -20212
rect 398372 -20268 398574 -20212
rect 398630 -20268 398716 -20212
rect 398772 -20268 398971 -20212
rect 399027 -20268 399113 -20212
rect 399169 -20268 399376 -20212
rect 399432 -20268 399518 -20212
rect 399574 -20268 399776 -20212
rect 399832 -20268 399918 -20212
rect 399974 -20268 400181 -20212
rect 400237 -20268 400323 -20212
rect 400379 -20260 400766 -20212
rect 400822 -20260 400890 -20204
rect 400946 -20260 401014 -20204
rect 401070 -20260 401138 -20204
rect 401194 -20260 401262 -20204
rect 401318 -20260 402640 -20204
rect 400379 -20268 402640 -20260
rect 387840 -20328 402640 -20268
rect 387840 -20384 387954 -20328
rect 388010 -20384 388078 -20328
rect 388134 -20384 388202 -20328
rect 388258 -20384 388326 -20328
rect 388382 -20384 388450 -20328
rect 388506 -20354 400766 -20328
rect 388506 -20384 388981 -20354
rect 387840 -20410 388981 -20384
rect 389037 -20410 389123 -20354
rect 389179 -20410 389382 -20354
rect 389438 -20410 389524 -20354
rect 389580 -20410 389782 -20354
rect 389838 -20410 389924 -20354
rect 389980 -20410 390179 -20354
rect 390235 -20410 390321 -20354
rect 390377 -20410 390576 -20354
rect 390632 -20410 390718 -20354
rect 390774 -20410 390980 -20354
rect 391036 -20410 391122 -20354
rect 391178 -20410 391376 -20354
rect 391432 -20410 391518 -20354
rect 391574 -20410 391776 -20354
rect 391832 -20410 391918 -20354
rect 391974 -20410 392173 -20354
rect 392229 -20410 392315 -20354
rect 392371 -20410 392578 -20354
rect 392634 -20410 392720 -20354
rect 392776 -20410 392978 -20354
rect 393034 -20410 393120 -20354
rect 393176 -20410 393383 -20354
rect 393439 -20410 393525 -20354
rect 393581 -20410 393780 -20354
rect 393836 -20410 393922 -20354
rect 393978 -20410 394177 -20354
rect 394233 -20410 394319 -20354
rect 394375 -20410 394580 -20354
rect 394636 -20410 394722 -20354
rect 394778 -20410 394982 -20354
rect 395038 -20410 395124 -20354
rect 395180 -20410 395385 -20354
rect 395441 -20410 395527 -20354
rect 395583 -20410 395779 -20354
rect 395835 -20410 395921 -20354
rect 395977 -20410 396180 -20354
rect 396236 -20410 396322 -20354
rect 396378 -20410 396580 -20354
rect 396636 -20410 396722 -20354
rect 396778 -20410 396977 -20354
rect 397033 -20410 397119 -20354
rect 397175 -20410 397374 -20354
rect 397430 -20410 397516 -20354
rect 397572 -20410 397778 -20354
rect 397834 -20410 397920 -20354
rect 397976 -20410 398174 -20354
rect 398230 -20410 398316 -20354
rect 398372 -20410 398574 -20354
rect 398630 -20410 398716 -20354
rect 398772 -20410 398971 -20354
rect 399027 -20410 399113 -20354
rect 399169 -20410 399376 -20354
rect 399432 -20410 399518 -20354
rect 399574 -20410 399776 -20354
rect 399832 -20410 399918 -20354
rect 399974 -20410 400181 -20354
rect 400237 -20410 400323 -20354
rect 400379 -20384 400766 -20354
rect 400822 -20384 400890 -20328
rect 400946 -20384 401014 -20328
rect 401070 -20384 401138 -20328
rect 401194 -20384 401262 -20328
rect 401318 -20384 402640 -20328
rect 400379 -20410 402640 -20384
rect 387840 -20452 402640 -20410
rect 387840 -20508 387954 -20452
rect 388010 -20508 388078 -20452
rect 388134 -20508 388202 -20452
rect 388258 -20508 388326 -20452
rect 388382 -20508 388450 -20452
rect 388506 -20496 400766 -20452
rect 388506 -20508 388981 -20496
rect 387840 -20552 388981 -20508
rect 389037 -20552 389123 -20496
rect 389179 -20552 389382 -20496
rect 389438 -20552 389524 -20496
rect 389580 -20552 389782 -20496
rect 389838 -20552 389924 -20496
rect 389980 -20552 390179 -20496
rect 390235 -20552 390321 -20496
rect 390377 -20552 390576 -20496
rect 390632 -20552 390718 -20496
rect 390774 -20552 390980 -20496
rect 391036 -20552 391122 -20496
rect 391178 -20552 391376 -20496
rect 391432 -20552 391518 -20496
rect 391574 -20552 391776 -20496
rect 391832 -20552 391918 -20496
rect 391974 -20552 392173 -20496
rect 392229 -20552 392315 -20496
rect 392371 -20552 392578 -20496
rect 392634 -20552 392720 -20496
rect 392776 -20552 392978 -20496
rect 393034 -20552 393120 -20496
rect 393176 -20552 393383 -20496
rect 393439 -20552 393525 -20496
rect 393581 -20552 393780 -20496
rect 393836 -20552 393922 -20496
rect 393978 -20552 394177 -20496
rect 394233 -20552 394319 -20496
rect 394375 -20552 394580 -20496
rect 394636 -20552 394722 -20496
rect 394778 -20552 394982 -20496
rect 395038 -20552 395124 -20496
rect 395180 -20552 395385 -20496
rect 395441 -20552 395527 -20496
rect 395583 -20552 395779 -20496
rect 395835 -20552 395921 -20496
rect 395977 -20552 396180 -20496
rect 396236 -20552 396322 -20496
rect 396378 -20552 396580 -20496
rect 396636 -20552 396722 -20496
rect 396778 -20552 396977 -20496
rect 397033 -20552 397119 -20496
rect 397175 -20552 397374 -20496
rect 397430 -20552 397516 -20496
rect 397572 -20552 397778 -20496
rect 397834 -20552 397920 -20496
rect 397976 -20552 398174 -20496
rect 398230 -20552 398316 -20496
rect 398372 -20552 398574 -20496
rect 398630 -20552 398716 -20496
rect 398772 -20552 398971 -20496
rect 399027 -20552 399113 -20496
rect 399169 -20552 399376 -20496
rect 399432 -20552 399518 -20496
rect 399574 -20552 399776 -20496
rect 399832 -20552 399918 -20496
rect 399974 -20552 400181 -20496
rect 400237 -20552 400323 -20496
rect 400379 -20508 400766 -20496
rect 400822 -20508 400890 -20452
rect 400946 -20508 401014 -20452
rect 401070 -20508 401138 -20452
rect 401194 -20508 401262 -20452
rect 401318 -20508 402640 -20452
rect 400379 -20552 402640 -20508
rect 387840 -20576 402640 -20552
rect 387840 -20632 387954 -20576
rect 388010 -20632 388078 -20576
rect 388134 -20632 388202 -20576
rect 388258 -20632 388326 -20576
rect 388382 -20632 388450 -20576
rect 388506 -20632 400766 -20576
rect 400822 -20632 400890 -20576
rect 400946 -20632 401014 -20576
rect 401070 -20632 401138 -20576
rect 401194 -20632 401262 -20576
rect 401318 -20632 402640 -20576
rect 387840 -20638 402640 -20632
rect 387840 -20694 388981 -20638
rect 389037 -20694 389123 -20638
rect 389179 -20694 389382 -20638
rect 389438 -20694 389524 -20638
rect 389580 -20694 389782 -20638
rect 389838 -20694 389924 -20638
rect 389980 -20694 390179 -20638
rect 390235 -20694 390321 -20638
rect 390377 -20694 390576 -20638
rect 390632 -20694 390718 -20638
rect 390774 -20694 390980 -20638
rect 391036 -20694 391122 -20638
rect 391178 -20694 391376 -20638
rect 391432 -20694 391518 -20638
rect 391574 -20694 391776 -20638
rect 391832 -20694 391918 -20638
rect 391974 -20694 392173 -20638
rect 392229 -20694 392315 -20638
rect 392371 -20694 392578 -20638
rect 392634 -20694 392720 -20638
rect 392776 -20694 392978 -20638
rect 393034 -20694 393120 -20638
rect 393176 -20694 393383 -20638
rect 393439 -20694 393525 -20638
rect 393581 -20694 393780 -20638
rect 393836 -20694 393922 -20638
rect 393978 -20694 394177 -20638
rect 394233 -20694 394319 -20638
rect 394375 -20694 394580 -20638
rect 394636 -20694 394722 -20638
rect 394778 -20694 394982 -20638
rect 395038 -20694 395124 -20638
rect 395180 -20694 395385 -20638
rect 395441 -20694 395527 -20638
rect 395583 -20694 395779 -20638
rect 395835 -20694 395921 -20638
rect 395977 -20694 396180 -20638
rect 396236 -20694 396322 -20638
rect 396378 -20694 396580 -20638
rect 396636 -20694 396722 -20638
rect 396778 -20694 396977 -20638
rect 397033 -20694 397119 -20638
rect 397175 -20694 397374 -20638
rect 397430 -20694 397516 -20638
rect 397572 -20694 397778 -20638
rect 397834 -20694 397920 -20638
rect 397976 -20694 398174 -20638
rect 398230 -20694 398316 -20638
rect 398372 -20694 398574 -20638
rect 398630 -20694 398716 -20638
rect 398772 -20694 398971 -20638
rect 399027 -20694 399113 -20638
rect 399169 -20694 399376 -20638
rect 399432 -20694 399518 -20638
rect 399574 -20694 399776 -20638
rect 399832 -20694 399918 -20638
rect 399974 -20694 400181 -20638
rect 400237 -20694 400323 -20638
rect 400379 -20694 402640 -20638
rect 387840 -20700 402640 -20694
rect 387840 -20756 387954 -20700
rect 388010 -20756 388078 -20700
rect 388134 -20756 388202 -20700
rect 388258 -20756 388326 -20700
rect 388382 -20756 388450 -20700
rect 388506 -20756 400766 -20700
rect 400822 -20756 400890 -20700
rect 400946 -20756 401014 -20700
rect 401070 -20756 401138 -20700
rect 401194 -20756 401262 -20700
rect 401318 -20756 402640 -20700
rect 387840 -20780 402640 -20756
rect 387840 -20824 388981 -20780
rect 387840 -20880 387954 -20824
rect 388010 -20880 388078 -20824
rect 388134 -20880 388202 -20824
rect 388258 -20880 388326 -20824
rect 388382 -20880 388450 -20824
rect 388506 -20836 388981 -20824
rect 389037 -20836 389123 -20780
rect 389179 -20836 389382 -20780
rect 389438 -20836 389524 -20780
rect 389580 -20836 389782 -20780
rect 389838 -20836 389924 -20780
rect 389980 -20836 390179 -20780
rect 390235 -20836 390321 -20780
rect 390377 -20836 390576 -20780
rect 390632 -20836 390718 -20780
rect 390774 -20836 390980 -20780
rect 391036 -20836 391122 -20780
rect 391178 -20836 391376 -20780
rect 391432 -20836 391518 -20780
rect 391574 -20836 391776 -20780
rect 391832 -20836 391918 -20780
rect 391974 -20836 392173 -20780
rect 392229 -20836 392315 -20780
rect 392371 -20836 392578 -20780
rect 392634 -20836 392720 -20780
rect 392776 -20836 392978 -20780
rect 393034 -20836 393120 -20780
rect 393176 -20836 393383 -20780
rect 393439 -20836 393525 -20780
rect 393581 -20836 393780 -20780
rect 393836 -20836 393922 -20780
rect 393978 -20836 394177 -20780
rect 394233 -20836 394319 -20780
rect 394375 -20836 394580 -20780
rect 394636 -20836 394722 -20780
rect 394778 -20836 394982 -20780
rect 395038 -20836 395124 -20780
rect 395180 -20836 395385 -20780
rect 395441 -20836 395527 -20780
rect 395583 -20836 395779 -20780
rect 395835 -20836 395921 -20780
rect 395977 -20836 396180 -20780
rect 396236 -20836 396322 -20780
rect 396378 -20836 396580 -20780
rect 396636 -20836 396722 -20780
rect 396778 -20836 396977 -20780
rect 397033 -20836 397119 -20780
rect 397175 -20836 397374 -20780
rect 397430 -20836 397516 -20780
rect 397572 -20836 397778 -20780
rect 397834 -20836 397920 -20780
rect 397976 -20836 398174 -20780
rect 398230 -20836 398316 -20780
rect 398372 -20836 398574 -20780
rect 398630 -20836 398716 -20780
rect 398772 -20836 398971 -20780
rect 399027 -20836 399113 -20780
rect 399169 -20836 399376 -20780
rect 399432 -20836 399518 -20780
rect 399574 -20836 399776 -20780
rect 399832 -20836 399918 -20780
rect 399974 -20836 400181 -20780
rect 400237 -20836 400323 -20780
rect 400379 -20824 402640 -20780
rect 400379 -20836 400766 -20824
rect 388506 -20880 400766 -20836
rect 400822 -20880 400890 -20824
rect 400946 -20880 401014 -20824
rect 401070 -20880 401138 -20824
rect 401194 -20880 401262 -20824
rect 401318 -20880 402640 -20824
rect 387840 -20922 402640 -20880
rect 387840 -20948 388981 -20922
rect 387840 -21004 387954 -20948
rect 388010 -21004 388078 -20948
rect 388134 -21004 388202 -20948
rect 388258 -21004 388326 -20948
rect 388382 -21004 388450 -20948
rect 388506 -20978 388981 -20948
rect 389037 -20978 389123 -20922
rect 389179 -20978 389382 -20922
rect 389438 -20978 389524 -20922
rect 389580 -20978 389782 -20922
rect 389838 -20978 389924 -20922
rect 389980 -20978 390179 -20922
rect 390235 -20978 390321 -20922
rect 390377 -20978 390576 -20922
rect 390632 -20978 390718 -20922
rect 390774 -20978 390980 -20922
rect 391036 -20978 391122 -20922
rect 391178 -20978 391376 -20922
rect 391432 -20978 391518 -20922
rect 391574 -20978 391776 -20922
rect 391832 -20978 391918 -20922
rect 391974 -20978 392173 -20922
rect 392229 -20978 392315 -20922
rect 392371 -20978 392578 -20922
rect 392634 -20978 392720 -20922
rect 392776 -20978 392978 -20922
rect 393034 -20978 393120 -20922
rect 393176 -20978 393383 -20922
rect 393439 -20978 393525 -20922
rect 393581 -20978 393780 -20922
rect 393836 -20978 393922 -20922
rect 393978 -20978 394177 -20922
rect 394233 -20978 394319 -20922
rect 394375 -20978 394580 -20922
rect 394636 -20978 394722 -20922
rect 394778 -20978 394982 -20922
rect 395038 -20978 395124 -20922
rect 395180 -20978 395385 -20922
rect 395441 -20978 395527 -20922
rect 395583 -20978 395779 -20922
rect 395835 -20978 395921 -20922
rect 395977 -20978 396180 -20922
rect 396236 -20978 396322 -20922
rect 396378 -20978 396580 -20922
rect 396636 -20978 396722 -20922
rect 396778 -20978 396977 -20922
rect 397033 -20978 397119 -20922
rect 397175 -20978 397374 -20922
rect 397430 -20978 397516 -20922
rect 397572 -20978 397778 -20922
rect 397834 -20978 397920 -20922
rect 397976 -20978 398174 -20922
rect 398230 -20978 398316 -20922
rect 398372 -20978 398574 -20922
rect 398630 -20978 398716 -20922
rect 398772 -20978 398971 -20922
rect 399027 -20978 399113 -20922
rect 399169 -20978 399376 -20922
rect 399432 -20978 399518 -20922
rect 399574 -20978 399776 -20922
rect 399832 -20978 399918 -20922
rect 399974 -20978 400181 -20922
rect 400237 -20978 400323 -20922
rect 400379 -20948 402640 -20922
rect 400379 -20978 400766 -20948
rect 388506 -21004 400766 -20978
rect 400822 -21004 400890 -20948
rect 400946 -21004 401014 -20948
rect 401070 -21004 401138 -20948
rect 401194 -21004 401262 -20948
rect 401318 -21004 402640 -20948
rect 387840 -21064 402640 -21004
rect 387840 -21072 388981 -21064
rect 387840 -21128 387954 -21072
rect 388010 -21128 388078 -21072
rect 388134 -21128 388202 -21072
rect 388258 -21128 388326 -21072
rect 388382 -21128 388450 -21072
rect 388506 -21120 388981 -21072
rect 389037 -21120 389123 -21064
rect 389179 -21120 389382 -21064
rect 389438 -21120 389524 -21064
rect 389580 -21120 389782 -21064
rect 389838 -21120 389924 -21064
rect 389980 -21120 390179 -21064
rect 390235 -21120 390321 -21064
rect 390377 -21120 390576 -21064
rect 390632 -21120 390718 -21064
rect 390774 -21120 390980 -21064
rect 391036 -21120 391122 -21064
rect 391178 -21120 391376 -21064
rect 391432 -21120 391518 -21064
rect 391574 -21120 391776 -21064
rect 391832 -21120 391918 -21064
rect 391974 -21120 392173 -21064
rect 392229 -21120 392315 -21064
rect 392371 -21120 392578 -21064
rect 392634 -21120 392720 -21064
rect 392776 -21120 392978 -21064
rect 393034 -21120 393120 -21064
rect 393176 -21120 393383 -21064
rect 393439 -21120 393525 -21064
rect 393581 -21120 393780 -21064
rect 393836 -21120 393922 -21064
rect 393978 -21120 394177 -21064
rect 394233 -21120 394319 -21064
rect 394375 -21120 394580 -21064
rect 394636 -21120 394722 -21064
rect 394778 -21120 394982 -21064
rect 395038 -21120 395124 -21064
rect 395180 -21120 395385 -21064
rect 395441 -21120 395527 -21064
rect 395583 -21120 395779 -21064
rect 395835 -21120 395921 -21064
rect 395977 -21120 396180 -21064
rect 396236 -21120 396322 -21064
rect 396378 -21120 396580 -21064
rect 396636 -21120 396722 -21064
rect 396778 -21120 396977 -21064
rect 397033 -21120 397119 -21064
rect 397175 -21120 397374 -21064
rect 397430 -21120 397516 -21064
rect 397572 -21120 397778 -21064
rect 397834 -21120 397920 -21064
rect 397976 -21120 398174 -21064
rect 398230 -21120 398316 -21064
rect 398372 -21120 398574 -21064
rect 398630 -21120 398716 -21064
rect 398772 -21120 398971 -21064
rect 399027 -21120 399113 -21064
rect 399169 -21120 399376 -21064
rect 399432 -21120 399518 -21064
rect 399574 -21120 399776 -21064
rect 399832 -21120 399918 -21064
rect 399974 -21120 400181 -21064
rect 400237 -21120 400323 -21064
rect 400379 -21072 402640 -21064
rect 400379 -21120 400766 -21072
rect 388506 -21128 400766 -21120
rect 400822 -21128 400890 -21072
rect 400946 -21128 401014 -21072
rect 401070 -21128 401138 -21072
rect 401194 -21128 401262 -21072
rect 401318 -21128 402640 -21072
rect 387840 -21196 402640 -21128
rect 387840 -21252 387954 -21196
rect 388010 -21252 388078 -21196
rect 388134 -21252 388202 -21196
rect 388258 -21252 388326 -21196
rect 388382 -21252 388450 -21196
rect 388506 -21206 400766 -21196
rect 388506 -21252 388981 -21206
rect 387840 -21262 388981 -21252
rect 389037 -21262 389123 -21206
rect 389179 -21262 389382 -21206
rect 389438 -21262 389524 -21206
rect 389580 -21262 389782 -21206
rect 389838 -21262 389924 -21206
rect 389980 -21262 390179 -21206
rect 390235 -21262 390321 -21206
rect 390377 -21262 390576 -21206
rect 390632 -21262 390718 -21206
rect 390774 -21262 390980 -21206
rect 391036 -21262 391122 -21206
rect 391178 -21262 391376 -21206
rect 391432 -21262 391518 -21206
rect 391574 -21262 391776 -21206
rect 391832 -21262 391918 -21206
rect 391974 -21262 392173 -21206
rect 392229 -21262 392315 -21206
rect 392371 -21262 392578 -21206
rect 392634 -21262 392720 -21206
rect 392776 -21262 392978 -21206
rect 393034 -21262 393120 -21206
rect 393176 -21262 393383 -21206
rect 393439 -21262 393525 -21206
rect 393581 -21262 393780 -21206
rect 393836 -21262 393922 -21206
rect 393978 -21262 394177 -21206
rect 394233 -21262 394319 -21206
rect 394375 -21262 394580 -21206
rect 394636 -21262 394722 -21206
rect 394778 -21262 394982 -21206
rect 395038 -21262 395124 -21206
rect 395180 -21262 395385 -21206
rect 395441 -21262 395527 -21206
rect 395583 -21262 395779 -21206
rect 395835 -21262 395921 -21206
rect 395977 -21262 396180 -21206
rect 396236 -21262 396322 -21206
rect 396378 -21262 396580 -21206
rect 396636 -21262 396722 -21206
rect 396778 -21262 396977 -21206
rect 397033 -21262 397119 -21206
rect 397175 -21262 397374 -21206
rect 397430 -21262 397516 -21206
rect 397572 -21262 397778 -21206
rect 397834 -21262 397920 -21206
rect 397976 -21262 398174 -21206
rect 398230 -21262 398316 -21206
rect 398372 -21262 398574 -21206
rect 398630 -21262 398716 -21206
rect 398772 -21262 398971 -21206
rect 399027 -21262 399113 -21206
rect 399169 -21262 399376 -21206
rect 399432 -21262 399518 -21206
rect 399574 -21262 399776 -21206
rect 399832 -21262 399918 -21206
rect 399974 -21262 400181 -21206
rect 400237 -21262 400323 -21206
rect 400379 -21252 400766 -21206
rect 400822 -21252 400890 -21196
rect 400946 -21252 401014 -21196
rect 401070 -21252 401138 -21196
rect 401194 -21252 401262 -21196
rect 401318 -21252 402640 -21196
rect 400379 -21262 402640 -21252
rect 387840 -21320 402640 -21262
rect 387840 -21376 387954 -21320
rect 388010 -21376 388078 -21320
rect 388134 -21376 388202 -21320
rect 388258 -21376 388326 -21320
rect 388382 -21376 388450 -21320
rect 388506 -21348 400766 -21320
rect 388506 -21376 388981 -21348
rect 387840 -21404 388981 -21376
rect 389037 -21404 389123 -21348
rect 389179 -21404 389382 -21348
rect 389438 -21404 389524 -21348
rect 389580 -21404 389782 -21348
rect 389838 -21404 389924 -21348
rect 389980 -21404 390179 -21348
rect 390235 -21404 390321 -21348
rect 390377 -21404 390576 -21348
rect 390632 -21404 390718 -21348
rect 390774 -21404 390980 -21348
rect 391036 -21404 391122 -21348
rect 391178 -21404 391376 -21348
rect 391432 -21404 391518 -21348
rect 391574 -21404 391776 -21348
rect 391832 -21404 391918 -21348
rect 391974 -21404 392173 -21348
rect 392229 -21404 392315 -21348
rect 392371 -21404 392578 -21348
rect 392634 -21404 392720 -21348
rect 392776 -21404 392978 -21348
rect 393034 -21404 393120 -21348
rect 393176 -21404 393383 -21348
rect 393439 -21404 393525 -21348
rect 393581 -21404 393780 -21348
rect 393836 -21404 393922 -21348
rect 393978 -21404 394177 -21348
rect 394233 -21404 394319 -21348
rect 394375 -21404 394580 -21348
rect 394636 -21404 394722 -21348
rect 394778 -21404 394982 -21348
rect 395038 -21404 395124 -21348
rect 395180 -21404 395385 -21348
rect 395441 -21404 395527 -21348
rect 395583 -21404 395779 -21348
rect 395835 -21404 395921 -21348
rect 395977 -21404 396180 -21348
rect 396236 -21404 396322 -21348
rect 396378 -21404 396580 -21348
rect 396636 -21404 396722 -21348
rect 396778 -21404 396977 -21348
rect 397033 -21404 397119 -21348
rect 397175 -21404 397374 -21348
rect 397430 -21404 397516 -21348
rect 397572 -21404 397778 -21348
rect 397834 -21404 397920 -21348
rect 397976 -21404 398174 -21348
rect 398230 -21404 398316 -21348
rect 398372 -21404 398574 -21348
rect 398630 -21404 398716 -21348
rect 398772 -21404 398971 -21348
rect 399027 -21404 399113 -21348
rect 399169 -21404 399376 -21348
rect 399432 -21404 399518 -21348
rect 399574 -21404 399776 -21348
rect 399832 -21404 399918 -21348
rect 399974 -21404 400181 -21348
rect 400237 -21404 400323 -21348
rect 400379 -21376 400766 -21348
rect 400822 -21376 400890 -21320
rect 400946 -21376 401014 -21320
rect 401070 -21376 401138 -21320
rect 401194 -21376 401262 -21320
rect 401318 -21376 402640 -21320
rect 400379 -21404 402640 -21376
rect 387840 -21444 402640 -21404
rect 387840 -21500 387954 -21444
rect 388010 -21500 388078 -21444
rect 388134 -21500 388202 -21444
rect 388258 -21500 388326 -21444
rect 388382 -21500 388450 -21444
rect 388506 -21490 400766 -21444
rect 388506 -21500 388981 -21490
rect 387840 -21546 388981 -21500
rect 389037 -21546 389123 -21490
rect 389179 -21546 389382 -21490
rect 389438 -21546 389524 -21490
rect 389580 -21546 389782 -21490
rect 389838 -21546 389924 -21490
rect 389980 -21546 390179 -21490
rect 390235 -21546 390321 -21490
rect 390377 -21546 390576 -21490
rect 390632 -21546 390718 -21490
rect 390774 -21546 390980 -21490
rect 391036 -21546 391122 -21490
rect 391178 -21546 391376 -21490
rect 391432 -21546 391518 -21490
rect 391574 -21546 391776 -21490
rect 391832 -21546 391918 -21490
rect 391974 -21546 392173 -21490
rect 392229 -21546 392315 -21490
rect 392371 -21546 392578 -21490
rect 392634 -21546 392720 -21490
rect 392776 -21546 392978 -21490
rect 393034 -21546 393120 -21490
rect 393176 -21546 393383 -21490
rect 393439 -21546 393525 -21490
rect 393581 -21546 393780 -21490
rect 393836 -21546 393922 -21490
rect 393978 -21546 394177 -21490
rect 394233 -21546 394319 -21490
rect 394375 -21546 394580 -21490
rect 394636 -21546 394722 -21490
rect 394778 -21546 394982 -21490
rect 395038 -21546 395124 -21490
rect 395180 -21546 395385 -21490
rect 395441 -21546 395527 -21490
rect 395583 -21546 395779 -21490
rect 395835 -21546 395921 -21490
rect 395977 -21546 396180 -21490
rect 396236 -21546 396322 -21490
rect 396378 -21546 396580 -21490
rect 396636 -21546 396722 -21490
rect 396778 -21546 396977 -21490
rect 397033 -21546 397119 -21490
rect 397175 -21546 397374 -21490
rect 397430 -21546 397516 -21490
rect 397572 -21546 397778 -21490
rect 397834 -21546 397920 -21490
rect 397976 -21546 398174 -21490
rect 398230 -21546 398316 -21490
rect 398372 -21546 398574 -21490
rect 398630 -21546 398716 -21490
rect 398772 -21546 398971 -21490
rect 399027 -21546 399113 -21490
rect 399169 -21546 399376 -21490
rect 399432 -21546 399518 -21490
rect 399574 -21546 399776 -21490
rect 399832 -21546 399918 -21490
rect 399974 -21546 400181 -21490
rect 400237 -21546 400323 -21490
rect 400379 -21500 400766 -21490
rect 400822 -21500 400890 -21444
rect 400946 -21500 401014 -21444
rect 401070 -21500 401138 -21444
rect 401194 -21500 401262 -21444
rect 401318 -21500 402640 -21444
rect 400379 -21546 402640 -21500
rect 387840 -21568 402640 -21546
rect 387840 -21624 387954 -21568
rect 388010 -21624 388078 -21568
rect 388134 -21624 388202 -21568
rect 388258 -21624 388326 -21568
rect 388382 -21624 388450 -21568
rect 388506 -21624 400766 -21568
rect 400822 -21624 400890 -21568
rect 400946 -21624 401014 -21568
rect 401070 -21624 401138 -21568
rect 401194 -21624 401262 -21568
rect 401318 -21624 402640 -21568
rect 387840 -21632 402640 -21624
rect 387840 -21688 388981 -21632
rect 389037 -21688 389123 -21632
rect 389179 -21688 389382 -21632
rect 389438 -21688 389524 -21632
rect 389580 -21688 389782 -21632
rect 389838 -21688 389924 -21632
rect 389980 -21688 390179 -21632
rect 390235 -21688 390321 -21632
rect 390377 -21688 390576 -21632
rect 390632 -21688 390718 -21632
rect 390774 -21688 390980 -21632
rect 391036 -21688 391122 -21632
rect 391178 -21688 391376 -21632
rect 391432 -21688 391518 -21632
rect 391574 -21688 391776 -21632
rect 391832 -21688 391918 -21632
rect 391974 -21688 392173 -21632
rect 392229 -21688 392315 -21632
rect 392371 -21688 392578 -21632
rect 392634 -21688 392720 -21632
rect 392776 -21688 392978 -21632
rect 393034 -21688 393120 -21632
rect 393176 -21688 393383 -21632
rect 393439 -21688 393525 -21632
rect 393581 -21688 393780 -21632
rect 393836 -21688 393922 -21632
rect 393978 -21688 394177 -21632
rect 394233 -21688 394319 -21632
rect 394375 -21688 394580 -21632
rect 394636 -21688 394722 -21632
rect 394778 -21688 394982 -21632
rect 395038 -21688 395124 -21632
rect 395180 -21688 395385 -21632
rect 395441 -21688 395527 -21632
rect 395583 -21688 395779 -21632
rect 395835 -21688 395921 -21632
rect 395977 -21688 396180 -21632
rect 396236 -21688 396322 -21632
rect 396378 -21688 396580 -21632
rect 396636 -21688 396722 -21632
rect 396778 -21688 396977 -21632
rect 397033 -21688 397119 -21632
rect 397175 -21688 397374 -21632
rect 397430 -21688 397516 -21632
rect 397572 -21688 397778 -21632
rect 397834 -21688 397920 -21632
rect 397976 -21688 398174 -21632
rect 398230 -21688 398316 -21632
rect 398372 -21688 398574 -21632
rect 398630 -21688 398716 -21632
rect 398772 -21688 398971 -21632
rect 399027 -21688 399113 -21632
rect 399169 -21688 399376 -21632
rect 399432 -21688 399518 -21632
rect 399574 -21688 399776 -21632
rect 399832 -21688 399918 -21632
rect 399974 -21688 400181 -21632
rect 400237 -21688 400323 -21632
rect 400379 -21688 402640 -21632
rect 387840 -21692 402640 -21688
rect 387840 -21748 387954 -21692
rect 388010 -21748 388078 -21692
rect 388134 -21748 388202 -21692
rect 388258 -21748 388326 -21692
rect 388382 -21748 388450 -21692
rect 388506 -21748 400766 -21692
rect 400822 -21748 400890 -21692
rect 400946 -21748 401014 -21692
rect 401070 -21748 401138 -21692
rect 401194 -21748 401262 -21692
rect 401318 -21748 402640 -21692
rect 387840 -21774 402640 -21748
rect 387840 -21816 388981 -21774
rect 387840 -21872 387954 -21816
rect 388010 -21872 388078 -21816
rect 388134 -21872 388202 -21816
rect 388258 -21872 388326 -21816
rect 388382 -21872 388450 -21816
rect 388506 -21830 388981 -21816
rect 389037 -21830 389123 -21774
rect 389179 -21830 389382 -21774
rect 389438 -21830 389524 -21774
rect 389580 -21830 389782 -21774
rect 389838 -21830 389924 -21774
rect 389980 -21830 390179 -21774
rect 390235 -21830 390321 -21774
rect 390377 -21830 390576 -21774
rect 390632 -21830 390718 -21774
rect 390774 -21830 390980 -21774
rect 391036 -21830 391122 -21774
rect 391178 -21830 391376 -21774
rect 391432 -21830 391518 -21774
rect 391574 -21830 391776 -21774
rect 391832 -21830 391918 -21774
rect 391974 -21830 392173 -21774
rect 392229 -21830 392315 -21774
rect 392371 -21830 392578 -21774
rect 392634 -21830 392720 -21774
rect 392776 -21830 392978 -21774
rect 393034 -21830 393120 -21774
rect 393176 -21830 393383 -21774
rect 393439 -21830 393525 -21774
rect 393581 -21830 393780 -21774
rect 393836 -21830 393922 -21774
rect 393978 -21830 394177 -21774
rect 394233 -21830 394319 -21774
rect 394375 -21830 394580 -21774
rect 394636 -21830 394722 -21774
rect 394778 -21830 394982 -21774
rect 395038 -21830 395124 -21774
rect 395180 -21830 395385 -21774
rect 395441 -21830 395527 -21774
rect 395583 -21830 395779 -21774
rect 395835 -21830 395921 -21774
rect 395977 -21830 396180 -21774
rect 396236 -21830 396322 -21774
rect 396378 -21830 396580 -21774
rect 396636 -21830 396722 -21774
rect 396778 -21830 396977 -21774
rect 397033 -21830 397119 -21774
rect 397175 -21830 397374 -21774
rect 397430 -21830 397516 -21774
rect 397572 -21830 397778 -21774
rect 397834 -21830 397920 -21774
rect 397976 -21830 398174 -21774
rect 398230 -21830 398316 -21774
rect 398372 -21830 398574 -21774
rect 398630 -21830 398716 -21774
rect 398772 -21830 398971 -21774
rect 399027 -21830 399113 -21774
rect 399169 -21830 399376 -21774
rect 399432 -21830 399518 -21774
rect 399574 -21830 399776 -21774
rect 399832 -21830 399918 -21774
rect 399974 -21830 400181 -21774
rect 400237 -21830 400323 -21774
rect 400379 -21816 402640 -21774
rect 400379 -21830 400766 -21816
rect 388506 -21872 400766 -21830
rect 400822 -21872 400890 -21816
rect 400946 -21872 401014 -21816
rect 401070 -21872 401138 -21816
rect 401194 -21872 401262 -21816
rect 401318 -21872 402640 -21816
rect 387840 -21916 402640 -21872
rect 387840 -21940 388981 -21916
rect 387840 -21996 387954 -21940
rect 388010 -21996 388078 -21940
rect 388134 -21996 388202 -21940
rect 388258 -21996 388326 -21940
rect 388382 -21996 388450 -21940
rect 388506 -21972 388981 -21940
rect 389037 -21972 389123 -21916
rect 389179 -21972 389382 -21916
rect 389438 -21972 389524 -21916
rect 389580 -21972 389782 -21916
rect 389838 -21972 389924 -21916
rect 389980 -21972 390179 -21916
rect 390235 -21972 390321 -21916
rect 390377 -21972 390576 -21916
rect 390632 -21972 390718 -21916
rect 390774 -21972 390980 -21916
rect 391036 -21972 391122 -21916
rect 391178 -21972 391376 -21916
rect 391432 -21972 391518 -21916
rect 391574 -21972 391776 -21916
rect 391832 -21972 391918 -21916
rect 391974 -21972 392173 -21916
rect 392229 -21972 392315 -21916
rect 392371 -21972 392578 -21916
rect 392634 -21972 392720 -21916
rect 392776 -21972 392978 -21916
rect 393034 -21972 393120 -21916
rect 393176 -21972 393383 -21916
rect 393439 -21972 393525 -21916
rect 393581 -21972 393780 -21916
rect 393836 -21972 393922 -21916
rect 393978 -21972 394177 -21916
rect 394233 -21972 394319 -21916
rect 394375 -21972 394580 -21916
rect 394636 -21972 394722 -21916
rect 394778 -21972 394982 -21916
rect 395038 -21972 395124 -21916
rect 395180 -21972 395385 -21916
rect 395441 -21972 395527 -21916
rect 395583 -21972 395779 -21916
rect 395835 -21972 395921 -21916
rect 395977 -21972 396180 -21916
rect 396236 -21972 396322 -21916
rect 396378 -21972 396580 -21916
rect 396636 -21972 396722 -21916
rect 396778 -21972 396977 -21916
rect 397033 -21972 397119 -21916
rect 397175 -21972 397374 -21916
rect 397430 -21972 397516 -21916
rect 397572 -21972 397778 -21916
rect 397834 -21972 397920 -21916
rect 397976 -21972 398174 -21916
rect 398230 -21972 398316 -21916
rect 398372 -21972 398574 -21916
rect 398630 -21972 398716 -21916
rect 398772 -21972 398971 -21916
rect 399027 -21972 399113 -21916
rect 399169 -21972 399376 -21916
rect 399432 -21972 399518 -21916
rect 399574 -21972 399776 -21916
rect 399832 -21972 399918 -21916
rect 399974 -21972 400181 -21916
rect 400237 -21972 400323 -21916
rect 400379 -21940 402640 -21916
rect 400379 -21972 400766 -21940
rect 388506 -21996 400766 -21972
rect 400822 -21996 400890 -21940
rect 400946 -21996 401014 -21940
rect 401070 -21996 401138 -21940
rect 401194 -21996 401262 -21940
rect 401318 -21996 402640 -21940
rect 387840 -22058 402640 -21996
rect 387840 -22064 388981 -22058
rect 387840 -22120 387954 -22064
rect 388010 -22120 388078 -22064
rect 388134 -22120 388202 -22064
rect 388258 -22120 388326 -22064
rect 388382 -22120 388450 -22064
rect 388506 -22114 388981 -22064
rect 389037 -22114 389123 -22058
rect 389179 -22114 389382 -22058
rect 389438 -22114 389524 -22058
rect 389580 -22114 389782 -22058
rect 389838 -22114 389924 -22058
rect 389980 -22114 390179 -22058
rect 390235 -22114 390321 -22058
rect 390377 -22114 390576 -22058
rect 390632 -22114 390718 -22058
rect 390774 -22114 390980 -22058
rect 391036 -22114 391122 -22058
rect 391178 -22114 391376 -22058
rect 391432 -22114 391518 -22058
rect 391574 -22114 391776 -22058
rect 391832 -22114 391918 -22058
rect 391974 -22114 392173 -22058
rect 392229 -22114 392315 -22058
rect 392371 -22114 392578 -22058
rect 392634 -22114 392720 -22058
rect 392776 -22114 392978 -22058
rect 393034 -22114 393120 -22058
rect 393176 -22114 393383 -22058
rect 393439 -22114 393525 -22058
rect 393581 -22114 393780 -22058
rect 393836 -22114 393922 -22058
rect 393978 -22114 394177 -22058
rect 394233 -22114 394319 -22058
rect 394375 -22114 394580 -22058
rect 394636 -22114 394722 -22058
rect 394778 -22114 394982 -22058
rect 395038 -22114 395124 -22058
rect 395180 -22114 395385 -22058
rect 395441 -22114 395527 -22058
rect 395583 -22114 395779 -22058
rect 395835 -22114 395921 -22058
rect 395977 -22114 396180 -22058
rect 396236 -22114 396322 -22058
rect 396378 -22114 396580 -22058
rect 396636 -22114 396722 -22058
rect 396778 -22114 396977 -22058
rect 397033 -22114 397119 -22058
rect 397175 -22114 397374 -22058
rect 397430 -22114 397516 -22058
rect 397572 -22114 397778 -22058
rect 397834 -22114 397920 -22058
rect 397976 -22114 398174 -22058
rect 398230 -22114 398316 -22058
rect 398372 -22114 398574 -22058
rect 398630 -22114 398716 -22058
rect 398772 -22114 398971 -22058
rect 399027 -22114 399113 -22058
rect 399169 -22114 399376 -22058
rect 399432 -22114 399518 -22058
rect 399574 -22114 399776 -22058
rect 399832 -22114 399918 -22058
rect 399974 -22114 400181 -22058
rect 400237 -22114 400323 -22058
rect 400379 -22064 402640 -22058
rect 400379 -22114 400766 -22064
rect 388506 -22120 400766 -22114
rect 400822 -22120 400890 -22064
rect 400946 -22120 401014 -22064
rect 401070 -22120 401138 -22064
rect 401194 -22120 401262 -22064
rect 401318 -22120 402640 -22064
rect 387840 -22188 402640 -22120
rect 387840 -22244 387954 -22188
rect 388010 -22244 388078 -22188
rect 388134 -22244 388202 -22188
rect 388258 -22244 388326 -22188
rect 388382 -22244 388450 -22188
rect 388506 -22200 400766 -22188
rect 388506 -22244 388981 -22200
rect 387840 -22256 388981 -22244
rect 389037 -22256 389123 -22200
rect 389179 -22256 389382 -22200
rect 389438 -22256 389524 -22200
rect 389580 -22256 389782 -22200
rect 389838 -22256 389924 -22200
rect 389980 -22256 390179 -22200
rect 390235 -22256 390321 -22200
rect 390377 -22256 390576 -22200
rect 390632 -22256 390718 -22200
rect 390774 -22256 390980 -22200
rect 391036 -22256 391122 -22200
rect 391178 -22256 391376 -22200
rect 391432 -22256 391518 -22200
rect 391574 -22256 391776 -22200
rect 391832 -22256 391918 -22200
rect 391974 -22256 392173 -22200
rect 392229 -22256 392315 -22200
rect 392371 -22256 392578 -22200
rect 392634 -22256 392720 -22200
rect 392776 -22256 392978 -22200
rect 393034 -22256 393120 -22200
rect 393176 -22256 393383 -22200
rect 393439 -22256 393525 -22200
rect 393581 -22256 393780 -22200
rect 393836 -22256 393922 -22200
rect 393978 -22256 394177 -22200
rect 394233 -22256 394319 -22200
rect 394375 -22256 394580 -22200
rect 394636 -22256 394722 -22200
rect 394778 -22256 394982 -22200
rect 395038 -22256 395124 -22200
rect 395180 -22256 395385 -22200
rect 395441 -22256 395527 -22200
rect 395583 -22256 395779 -22200
rect 395835 -22256 395921 -22200
rect 395977 -22256 396180 -22200
rect 396236 -22256 396322 -22200
rect 396378 -22256 396580 -22200
rect 396636 -22256 396722 -22200
rect 396778 -22256 396977 -22200
rect 397033 -22256 397119 -22200
rect 397175 -22256 397374 -22200
rect 397430 -22256 397516 -22200
rect 397572 -22256 397778 -22200
rect 397834 -22256 397920 -22200
rect 397976 -22256 398174 -22200
rect 398230 -22256 398316 -22200
rect 398372 -22256 398574 -22200
rect 398630 -22256 398716 -22200
rect 398772 -22256 398971 -22200
rect 399027 -22256 399113 -22200
rect 399169 -22256 399376 -22200
rect 399432 -22256 399518 -22200
rect 399574 -22256 399776 -22200
rect 399832 -22256 399918 -22200
rect 399974 -22256 400181 -22200
rect 400237 -22256 400323 -22200
rect 400379 -22244 400766 -22200
rect 400822 -22244 400890 -22188
rect 400946 -22244 401014 -22188
rect 401070 -22244 401138 -22188
rect 401194 -22244 401262 -22188
rect 401318 -22244 402640 -22188
rect 400379 -22256 402640 -22244
rect 387840 -22312 402640 -22256
rect 387840 -22368 387954 -22312
rect 388010 -22368 388078 -22312
rect 388134 -22368 388202 -22312
rect 388258 -22368 388326 -22312
rect 388382 -22368 388450 -22312
rect 388506 -22342 400766 -22312
rect 388506 -22368 388981 -22342
rect 387840 -22398 388981 -22368
rect 389037 -22398 389123 -22342
rect 389179 -22398 389382 -22342
rect 389438 -22398 389524 -22342
rect 389580 -22398 389782 -22342
rect 389838 -22398 389924 -22342
rect 389980 -22398 390179 -22342
rect 390235 -22398 390321 -22342
rect 390377 -22398 390576 -22342
rect 390632 -22398 390718 -22342
rect 390774 -22398 390980 -22342
rect 391036 -22398 391122 -22342
rect 391178 -22398 391376 -22342
rect 391432 -22398 391518 -22342
rect 391574 -22398 391776 -22342
rect 391832 -22398 391918 -22342
rect 391974 -22398 392173 -22342
rect 392229 -22398 392315 -22342
rect 392371 -22398 392578 -22342
rect 392634 -22398 392720 -22342
rect 392776 -22398 392978 -22342
rect 393034 -22398 393120 -22342
rect 393176 -22398 393383 -22342
rect 393439 -22398 393525 -22342
rect 393581 -22398 393780 -22342
rect 393836 -22398 393922 -22342
rect 393978 -22398 394177 -22342
rect 394233 -22398 394319 -22342
rect 394375 -22398 394580 -22342
rect 394636 -22398 394722 -22342
rect 394778 -22398 394982 -22342
rect 395038 -22398 395124 -22342
rect 395180 -22398 395385 -22342
rect 395441 -22398 395527 -22342
rect 395583 -22398 395779 -22342
rect 395835 -22398 395921 -22342
rect 395977 -22398 396180 -22342
rect 396236 -22398 396322 -22342
rect 396378 -22398 396580 -22342
rect 396636 -22398 396722 -22342
rect 396778 -22398 396977 -22342
rect 397033 -22398 397119 -22342
rect 397175 -22398 397374 -22342
rect 397430 -22398 397516 -22342
rect 397572 -22398 397778 -22342
rect 397834 -22398 397920 -22342
rect 397976 -22398 398174 -22342
rect 398230 -22398 398316 -22342
rect 398372 -22398 398574 -22342
rect 398630 -22398 398716 -22342
rect 398772 -22398 398971 -22342
rect 399027 -22398 399113 -22342
rect 399169 -22398 399376 -22342
rect 399432 -22398 399518 -22342
rect 399574 -22398 399776 -22342
rect 399832 -22398 399918 -22342
rect 399974 -22398 400181 -22342
rect 400237 -22398 400323 -22342
rect 400379 -22368 400766 -22342
rect 400822 -22368 400890 -22312
rect 400946 -22368 401014 -22312
rect 401070 -22368 401138 -22312
rect 401194 -22368 401262 -22312
rect 401318 -22368 402640 -22312
rect 400379 -22398 402640 -22368
rect 387840 -22436 402640 -22398
rect 387840 -22492 387954 -22436
rect 388010 -22492 388078 -22436
rect 388134 -22492 388202 -22436
rect 388258 -22492 388326 -22436
rect 388382 -22492 388450 -22436
rect 388506 -22484 400766 -22436
rect 388506 -22492 388981 -22484
rect 387840 -22540 388981 -22492
rect 389037 -22540 389123 -22484
rect 389179 -22540 389382 -22484
rect 389438 -22540 389524 -22484
rect 389580 -22540 389782 -22484
rect 389838 -22540 389924 -22484
rect 389980 -22540 390179 -22484
rect 390235 -22540 390321 -22484
rect 390377 -22540 390576 -22484
rect 390632 -22540 390718 -22484
rect 390774 -22540 390980 -22484
rect 391036 -22540 391122 -22484
rect 391178 -22540 391376 -22484
rect 391432 -22540 391518 -22484
rect 391574 -22540 391776 -22484
rect 391832 -22540 391918 -22484
rect 391974 -22540 392173 -22484
rect 392229 -22540 392315 -22484
rect 392371 -22540 392578 -22484
rect 392634 -22540 392720 -22484
rect 392776 -22540 392978 -22484
rect 393034 -22540 393120 -22484
rect 393176 -22540 393383 -22484
rect 393439 -22540 393525 -22484
rect 393581 -22540 393780 -22484
rect 393836 -22540 393922 -22484
rect 393978 -22540 394177 -22484
rect 394233 -22540 394319 -22484
rect 394375 -22540 394580 -22484
rect 394636 -22540 394722 -22484
rect 394778 -22540 394982 -22484
rect 395038 -22540 395124 -22484
rect 395180 -22540 395385 -22484
rect 395441 -22540 395527 -22484
rect 395583 -22540 395779 -22484
rect 395835 -22540 395921 -22484
rect 395977 -22540 396180 -22484
rect 396236 -22540 396322 -22484
rect 396378 -22540 396580 -22484
rect 396636 -22540 396722 -22484
rect 396778 -22540 396977 -22484
rect 397033 -22540 397119 -22484
rect 397175 -22540 397374 -22484
rect 397430 -22540 397516 -22484
rect 397572 -22540 397778 -22484
rect 397834 -22540 397920 -22484
rect 397976 -22540 398174 -22484
rect 398230 -22540 398316 -22484
rect 398372 -22540 398574 -22484
rect 398630 -22540 398716 -22484
rect 398772 -22540 398971 -22484
rect 399027 -22540 399113 -22484
rect 399169 -22540 399376 -22484
rect 399432 -22540 399518 -22484
rect 399574 -22540 399776 -22484
rect 399832 -22540 399918 -22484
rect 399974 -22540 400181 -22484
rect 400237 -22540 400323 -22484
rect 400379 -22492 400766 -22484
rect 400822 -22492 400890 -22436
rect 400946 -22492 401014 -22436
rect 401070 -22492 401138 -22436
rect 401194 -22492 401262 -22436
rect 401318 -22492 402640 -22436
rect 400379 -22540 402640 -22492
rect 387840 -22560 402640 -22540
rect 387840 -22616 387954 -22560
rect 388010 -22616 388078 -22560
rect 388134 -22616 388202 -22560
rect 388258 -22616 388326 -22560
rect 388382 -22616 388450 -22560
rect 388506 -22616 400766 -22560
rect 400822 -22616 400890 -22560
rect 400946 -22616 401014 -22560
rect 401070 -22616 401138 -22560
rect 401194 -22616 401262 -22560
rect 401318 -22616 402640 -22560
rect 387840 -22626 402640 -22616
rect 387840 -22682 388981 -22626
rect 389037 -22682 389123 -22626
rect 389179 -22682 389382 -22626
rect 389438 -22682 389524 -22626
rect 389580 -22682 389782 -22626
rect 389838 -22682 389924 -22626
rect 389980 -22682 390179 -22626
rect 390235 -22682 390321 -22626
rect 390377 -22682 390576 -22626
rect 390632 -22682 390718 -22626
rect 390774 -22682 390980 -22626
rect 391036 -22682 391122 -22626
rect 391178 -22682 391376 -22626
rect 391432 -22682 391518 -22626
rect 391574 -22682 391776 -22626
rect 391832 -22682 391918 -22626
rect 391974 -22682 392173 -22626
rect 392229 -22682 392315 -22626
rect 392371 -22682 392578 -22626
rect 392634 -22682 392720 -22626
rect 392776 -22682 392978 -22626
rect 393034 -22682 393120 -22626
rect 393176 -22682 393383 -22626
rect 393439 -22682 393525 -22626
rect 393581 -22682 393780 -22626
rect 393836 -22682 393922 -22626
rect 393978 -22682 394177 -22626
rect 394233 -22682 394319 -22626
rect 394375 -22682 394580 -22626
rect 394636 -22682 394722 -22626
rect 394778 -22682 394982 -22626
rect 395038 -22682 395124 -22626
rect 395180 -22682 395385 -22626
rect 395441 -22682 395527 -22626
rect 395583 -22682 395779 -22626
rect 395835 -22682 395921 -22626
rect 395977 -22682 396180 -22626
rect 396236 -22682 396322 -22626
rect 396378 -22682 396580 -22626
rect 396636 -22682 396722 -22626
rect 396778 -22682 396977 -22626
rect 397033 -22682 397119 -22626
rect 397175 -22682 397374 -22626
rect 397430 -22682 397516 -22626
rect 397572 -22682 397778 -22626
rect 397834 -22682 397920 -22626
rect 397976 -22682 398174 -22626
rect 398230 -22682 398316 -22626
rect 398372 -22682 398574 -22626
rect 398630 -22682 398716 -22626
rect 398772 -22682 398971 -22626
rect 399027 -22682 399113 -22626
rect 399169 -22682 399376 -22626
rect 399432 -22682 399518 -22626
rect 399574 -22682 399776 -22626
rect 399832 -22682 399918 -22626
rect 399974 -22682 400181 -22626
rect 400237 -22682 400323 -22626
rect 400379 -22682 402640 -22626
rect 387840 -22684 402640 -22682
rect 387840 -22740 387954 -22684
rect 388010 -22740 388078 -22684
rect 388134 -22740 388202 -22684
rect 388258 -22740 388326 -22684
rect 388382 -22740 388450 -22684
rect 388506 -22740 400766 -22684
rect 400822 -22740 400890 -22684
rect 400946 -22740 401014 -22684
rect 401070 -22740 401138 -22684
rect 401194 -22740 401262 -22684
rect 401318 -22740 402640 -22684
rect 387840 -22768 402640 -22740
rect 387840 -22808 388981 -22768
rect 387840 -22864 387954 -22808
rect 388010 -22864 388078 -22808
rect 388134 -22864 388202 -22808
rect 388258 -22864 388326 -22808
rect 388382 -22864 388450 -22808
rect 388506 -22824 388981 -22808
rect 389037 -22824 389123 -22768
rect 389179 -22824 389382 -22768
rect 389438 -22824 389524 -22768
rect 389580 -22824 389782 -22768
rect 389838 -22824 389924 -22768
rect 389980 -22824 390179 -22768
rect 390235 -22824 390321 -22768
rect 390377 -22824 390576 -22768
rect 390632 -22824 390718 -22768
rect 390774 -22824 390980 -22768
rect 391036 -22824 391122 -22768
rect 391178 -22824 391376 -22768
rect 391432 -22824 391518 -22768
rect 391574 -22824 391776 -22768
rect 391832 -22824 391918 -22768
rect 391974 -22824 392173 -22768
rect 392229 -22824 392315 -22768
rect 392371 -22824 392578 -22768
rect 392634 -22824 392720 -22768
rect 392776 -22824 392978 -22768
rect 393034 -22824 393120 -22768
rect 393176 -22824 393383 -22768
rect 393439 -22824 393525 -22768
rect 393581 -22824 393780 -22768
rect 393836 -22824 393922 -22768
rect 393978 -22824 394177 -22768
rect 394233 -22824 394319 -22768
rect 394375 -22824 394580 -22768
rect 394636 -22824 394722 -22768
rect 394778 -22824 394982 -22768
rect 395038 -22824 395124 -22768
rect 395180 -22824 395385 -22768
rect 395441 -22824 395527 -22768
rect 395583 -22824 395779 -22768
rect 395835 -22824 395921 -22768
rect 395977 -22824 396180 -22768
rect 396236 -22824 396322 -22768
rect 396378 -22824 396580 -22768
rect 396636 -22824 396722 -22768
rect 396778 -22824 396977 -22768
rect 397033 -22824 397119 -22768
rect 397175 -22824 397374 -22768
rect 397430 -22824 397516 -22768
rect 397572 -22824 397778 -22768
rect 397834 -22824 397920 -22768
rect 397976 -22824 398174 -22768
rect 398230 -22824 398316 -22768
rect 398372 -22824 398574 -22768
rect 398630 -22824 398716 -22768
rect 398772 -22824 398971 -22768
rect 399027 -22824 399113 -22768
rect 399169 -22824 399376 -22768
rect 399432 -22824 399518 -22768
rect 399574 -22824 399776 -22768
rect 399832 -22824 399918 -22768
rect 399974 -22824 400181 -22768
rect 400237 -22824 400323 -22768
rect 400379 -22808 402640 -22768
rect 400379 -22824 400766 -22808
rect 388506 -22864 400766 -22824
rect 400822 -22864 400890 -22808
rect 400946 -22864 401014 -22808
rect 401070 -22864 401138 -22808
rect 401194 -22864 401262 -22808
rect 401318 -22864 402640 -22808
rect 387840 -22910 402640 -22864
rect 387840 -22932 388981 -22910
rect 387840 -22988 387954 -22932
rect 388010 -22988 388078 -22932
rect 388134 -22988 388202 -22932
rect 388258 -22988 388326 -22932
rect 388382 -22988 388450 -22932
rect 388506 -22966 388981 -22932
rect 389037 -22966 389123 -22910
rect 389179 -22966 389382 -22910
rect 389438 -22966 389524 -22910
rect 389580 -22966 389782 -22910
rect 389838 -22966 389924 -22910
rect 389980 -22966 390179 -22910
rect 390235 -22966 390321 -22910
rect 390377 -22966 390576 -22910
rect 390632 -22966 390718 -22910
rect 390774 -22966 390980 -22910
rect 391036 -22966 391122 -22910
rect 391178 -22966 391376 -22910
rect 391432 -22966 391518 -22910
rect 391574 -22966 391776 -22910
rect 391832 -22966 391918 -22910
rect 391974 -22966 392173 -22910
rect 392229 -22966 392315 -22910
rect 392371 -22966 392578 -22910
rect 392634 -22966 392720 -22910
rect 392776 -22966 392978 -22910
rect 393034 -22966 393120 -22910
rect 393176 -22966 393383 -22910
rect 393439 -22966 393525 -22910
rect 393581 -22966 393780 -22910
rect 393836 -22966 393922 -22910
rect 393978 -22966 394177 -22910
rect 394233 -22966 394319 -22910
rect 394375 -22966 394580 -22910
rect 394636 -22966 394722 -22910
rect 394778 -22966 394982 -22910
rect 395038 -22966 395124 -22910
rect 395180 -22966 395385 -22910
rect 395441 -22966 395527 -22910
rect 395583 -22966 395779 -22910
rect 395835 -22966 395921 -22910
rect 395977 -22966 396180 -22910
rect 396236 -22966 396322 -22910
rect 396378 -22966 396580 -22910
rect 396636 -22966 396722 -22910
rect 396778 -22966 396977 -22910
rect 397033 -22966 397119 -22910
rect 397175 -22966 397374 -22910
rect 397430 -22966 397516 -22910
rect 397572 -22966 397778 -22910
rect 397834 -22966 397920 -22910
rect 397976 -22966 398174 -22910
rect 398230 -22966 398316 -22910
rect 398372 -22966 398574 -22910
rect 398630 -22966 398716 -22910
rect 398772 -22966 398971 -22910
rect 399027 -22966 399113 -22910
rect 399169 -22966 399376 -22910
rect 399432 -22966 399518 -22910
rect 399574 -22966 399776 -22910
rect 399832 -22966 399918 -22910
rect 399974 -22966 400181 -22910
rect 400237 -22966 400323 -22910
rect 400379 -22932 402640 -22910
rect 400379 -22966 400766 -22932
rect 388506 -22988 400766 -22966
rect 400822 -22988 400890 -22932
rect 400946 -22988 401014 -22932
rect 401070 -22988 401138 -22932
rect 401194 -22988 401262 -22932
rect 401318 -22988 402640 -22932
rect 387840 -23052 402640 -22988
rect 387840 -23056 388981 -23052
rect 387840 -23112 387954 -23056
rect 388010 -23112 388078 -23056
rect 388134 -23112 388202 -23056
rect 388258 -23112 388326 -23056
rect 388382 -23112 388450 -23056
rect 388506 -23108 388981 -23056
rect 389037 -23108 389123 -23052
rect 389179 -23108 389382 -23052
rect 389438 -23108 389524 -23052
rect 389580 -23108 389782 -23052
rect 389838 -23108 389924 -23052
rect 389980 -23108 390179 -23052
rect 390235 -23108 390321 -23052
rect 390377 -23108 390576 -23052
rect 390632 -23108 390718 -23052
rect 390774 -23108 390980 -23052
rect 391036 -23108 391122 -23052
rect 391178 -23108 391376 -23052
rect 391432 -23108 391518 -23052
rect 391574 -23108 391776 -23052
rect 391832 -23108 391918 -23052
rect 391974 -23108 392173 -23052
rect 392229 -23108 392315 -23052
rect 392371 -23108 392578 -23052
rect 392634 -23108 392720 -23052
rect 392776 -23108 392978 -23052
rect 393034 -23108 393120 -23052
rect 393176 -23108 393383 -23052
rect 393439 -23108 393525 -23052
rect 393581 -23108 393780 -23052
rect 393836 -23108 393922 -23052
rect 393978 -23108 394177 -23052
rect 394233 -23108 394319 -23052
rect 394375 -23108 394580 -23052
rect 394636 -23108 394722 -23052
rect 394778 -23108 394982 -23052
rect 395038 -23108 395124 -23052
rect 395180 -23108 395385 -23052
rect 395441 -23108 395527 -23052
rect 395583 -23108 395779 -23052
rect 395835 -23108 395921 -23052
rect 395977 -23108 396180 -23052
rect 396236 -23108 396322 -23052
rect 396378 -23108 396580 -23052
rect 396636 -23108 396722 -23052
rect 396778 -23108 396977 -23052
rect 397033 -23108 397119 -23052
rect 397175 -23108 397374 -23052
rect 397430 -23108 397516 -23052
rect 397572 -23108 397778 -23052
rect 397834 -23108 397920 -23052
rect 397976 -23108 398174 -23052
rect 398230 -23108 398316 -23052
rect 398372 -23108 398574 -23052
rect 398630 -23108 398716 -23052
rect 398772 -23108 398971 -23052
rect 399027 -23108 399113 -23052
rect 399169 -23108 399376 -23052
rect 399432 -23108 399518 -23052
rect 399574 -23108 399776 -23052
rect 399832 -23108 399918 -23052
rect 399974 -23108 400181 -23052
rect 400237 -23108 400323 -23052
rect 400379 -23056 402640 -23052
rect 400379 -23108 400766 -23056
rect 388506 -23112 400766 -23108
rect 400822 -23112 400890 -23056
rect 400946 -23112 401014 -23056
rect 401070 -23112 401138 -23056
rect 401194 -23112 401262 -23056
rect 401318 -23112 402640 -23056
rect 387840 -23180 402640 -23112
rect 387840 -23236 387954 -23180
rect 388010 -23236 388078 -23180
rect 388134 -23236 388202 -23180
rect 388258 -23236 388326 -23180
rect 388382 -23236 388450 -23180
rect 388506 -23194 400766 -23180
rect 388506 -23236 388981 -23194
rect 387840 -23250 388981 -23236
rect 389037 -23250 389123 -23194
rect 389179 -23250 389382 -23194
rect 389438 -23250 389524 -23194
rect 389580 -23250 389782 -23194
rect 389838 -23250 389924 -23194
rect 389980 -23250 390179 -23194
rect 390235 -23250 390321 -23194
rect 390377 -23250 390576 -23194
rect 390632 -23250 390718 -23194
rect 390774 -23250 390980 -23194
rect 391036 -23250 391122 -23194
rect 391178 -23250 391376 -23194
rect 391432 -23250 391518 -23194
rect 391574 -23250 391776 -23194
rect 391832 -23250 391918 -23194
rect 391974 -23250 392173 -23194
rect 392229 -23250 392315 -23194
rect 392371 -23250 392578 -23194
rect 392634 -23250 392720 -23194
rect 392776 -23250 392978 -23194
rect 393034 -23250 393120 -23194
rect 393176 -23250 393383 -23194
rect 393439 -23250 393525 -23194
rect 393581 -23250 393780 -23194
rect 393836 -23250 393922 -23194
rect 393978 -23250 394177 -23194
rect 394233 -23250 394319 -23194
rect 394375 -23250 394580 -23194
rect 394636 -23250 394722 -23194
rect 394778 -23250 394982 -23194
rect 395038 -23250 395124 -23194
rect 395180 -23250 395385 -23194
rect 395441 -23250 395527 -23194
rect 395583 -23250 395779 -23194
rect 395835 -23250 395921 -23194
rect 395977 -23250 396180 -23194
rect 396236 -23250 396322 -23194
rect 396378 -23250 396580 -23194
rect 396636 -23250 396722 -23194
rect 396778 -23250 396977 -23194
rect 397033 -23250 397119 -23194
rect 397175 -23250 397374 -23194
rect 397430 -23250 397516 -23194
rect 397572 -23250 397778 -23194
rect 397834 -23250 397920 -23194
rect 397976 -23250 398174 -23194
rect 398230 -23250 398316 -23194
rect 398372 -23250 398574 -23194
rect 398630 -23250 398716 -23194
rect 398772 -23250 398971 -23194
rect 399027 -23250 399113 -23194
rect 399169 -23250 399376 -23194
rect 399432 -23250 399518 -23194
rect 399574 -23250 399776 -23194
rect 399832 -23250 399918 -23194
rect 399974 -23250 400181 -23194
rect 400237 -23250 400323 -23194
rect 400379 -23236 400766 -23194
rect 400822 -23236 400890 -23180
rect 400946 -23236 401014 -23180
rect 401070 -23236 401138 -23180
rect 401194 -23236 401262 -23180
rect 401318 -23236 402640 -23180
rect 400379 -23250 402640 -23236
rect 387840 -23304 402640 -23250
rect 387840 -23360 387954 -23304
rect 388010 -23360 388078 -23304
rect 388134 -23360 388202 -23304
rect 388258 -23360 388326 -23304
rect 388382 -23360 388450 -23304
rect 388506 -23336 400766 -23304
rect 388506 -23360 388981 -23336
rect 387840 -23392 388981 -23360
rect 389037 -23392 389123 -23336
rect 389179 -23392 389382 -23336
rect 389438 -23392 389524 -23336
rect 389580 -23392 389782 -23336
rect 389838 -23392 389924 -23336
rect 389980 -23392 390179 -23336
rect 390235 -23392 390321 -23336
rect 390377 -23392 390576 -23336
rect 390632 -23392 390718 -23336
rect 390774 -23392 390980 -23336
rect 391036 -23392 391122 -23336
rect 391178 -23392 391376 -23336
rect 391432 -23392 391518 -23336
rect 391574 -23392 391776 -23336
rect 391832 -23392 391918 -23336
rect 391974 -23392 392173 -23336
rect 392229 -23392 392315 -23336
rect 392371 -23392 392578 -23336
rect 392634 -23392 392720 -23336
rect 392776 -23392 392978 -23336
rect 393034 -23392 393120 -23336
rect 393176 -23392 393383 -23336
rect 393439 -23392 393525 -23336
rect 393581 -23392 393780 -23336
rect 393836 -23392 393922 -23336
rect 393978 -23392 394177 -23336
rect 394233 -23392 394319 -23336
rect 394375 -23392 394580 -23336
rect 394636 -23392 394722 -23336
rect 394778 -23392 394982 -23336
rect 395038 -23392 395124 -23336
rect 395180 -23392 395385 -23336
rect 395441 -23392 395527 -23336
rect 395583 -23392 395779 -23336
rect 395835 -23392 395921 -23336
rect 395977 -23392 396180 -23336
rect 396236 -23392 396322 -23336
rect 396378 -23392 396580 -23336
rect 396636 -23392 396722 -23336
rect 396778 -23392 396977 -23336
rect 397033 -23392 397119 -23336
rect 397175 -23392 397374 -23336
rect 397430 -23392 397516 -23336
rect 397572 -23392 397778 -23336
rect 397834 -23392 397920 -23336
rect 397976 -23392 398174 -23336
rect 398230 -23392 398316 -23336
rect 398372 -23392 398574 -23336
rect 398630 -23392 398716 -23336
rect 398772 -23392 398971 -23336
rect 399027 -23392 399113 -23336
rect 399169 -23392 399376 -23336
rect 399432 -23392 399518 -23336
rect 399574 -23392 399776 -23336
rect 399832 -23392 399918 -23336
rect 399974 -23392 400181 -23336
rect 400237 -23392 400323 -23336
rect 400379 -23360 400766 -23336
rect 400822 -23360 400890 -23304
rect 400946 -23360 401014 -23304
rect 401070 -23360 401138 -23304
rect 401194 -23360 401262 -23304
rect 401318 -23360 402640 -23304
rect 400379 -23392 402640 -23360
rect 387840 -23428 402640 -23392
rect 387840 -23484 387954 -23428
rect 388010 -23484 388078 -23428
rect 388134 -23484 388202 -23428
rect 388258 -23484 388326 -23428
rect 388382 -23484 388450 -23428
rect 388506 -23478 400766 -23428
rect 388506 -23484 388981 -23478
rect 387840 -23534 388981 -23484
rect 389037 -23534 389123 -23478
rect 389179 -23534 389382 -23478
rect 389438 -23534 389524 -23478
rect 389580 -23534 389782 -23478
rect 389838 -23534 389924 -23478
rect 389980 -23534 390179 -23478
rect 390235 -23534 390321 -23478
rect 390377 -23534 390576 -23478
rect 390632 -23534 390718 -23478
rect 390774 -23534 390980 -23478
rect 391036 -23534 391122 -23478
rect 391178 -23534 391376 -23478
rect 391432 -23534 391518 -23478
rect 391574 -23534 391776 -23478
rect 391832 -23534 391918 -23478
rect 391974 -23534 392173 -23478
rect 392229 -23534 392315 -23478
rect 392371 -23534 392578 -23478
rect 392634 -23534 392720 -23478
rect 392776 -23534 392978 -23478
rect 393034 -23534 393120 -23478
rect 393176 -23534 393383 -23478
rect 393439 -23534 393525 -23478
rect 393581 -23534 393780 -23478
rect 393836 -23534 393922 -23478
rect 393978 -23534 394177 -23478
rect 394233 -23534 394319 -23478
rect 394375 -23534 394580 -23478
rect 394636 -23534 394722 -23478
rect 394778 -23534 394982 -23478
rect 395038 -23534 395124 -23478
rect 395180 -23534 395385 -23478
rect 395441 -23534 395527 -23478
rect 395583 -23534 395779 -23478
rect 395835 -23534 395921 -23478
rect 395977 -23534 396180 -23478
rect 396236 -23534 396322 -23478
rect 396378 -23534 396580 -23478
rect 396636 -23534 396722 -23478
rect 396778 -23534 396977 -23478
rect 397033 -23534 397119 -23478
rect 397175 -23534 397374 -23478
rect 397430 -23534 397516 -23478
rect 397572 -23534 397778 -23478
rect 397834 -23534 397920 -23478
rect 397976 -23534 398174 -23478
rect 398230 -23534 398316 -23478
rect 398372 -23534 398574 -23478
rect 398630 -23534 398716 -23478
rect 398772 -23534 398971 -23478
rect 399027 -23534 399113 -23478
rect 399169 -23534 399376 -23478
rect 399432 -23534 399518 -23478
rect 399574 -23534 399776 -23478
rect 399832 -23534 399918 -23478
rect 399974 -23534 400181 -23478
rect 400237 -23534 400323 -23478
rect 400379 -23484 400766 -23478
rect 400822 -23484 400890 -23428
rect 400946 -23484 401014 -23428
rect 401070 -23484 401138 -23428
rect 401194 -23484 401262 -23428
rect 401318 -23484 402640 -23428
rect 400379 -23534 402640 -23484
rect 387840 -23552 402640 -23534
rect 387840 -23608 387954 -23552
rect 388010 -23608 388078 -23552
rect 388134 -23608 388202 -23552
rect 388258 -23608 388326 -23552
rect 388382 -23608 388450 -23552
rect 388506 -23608 400766 -23552
rect 400822 -23608 400890 -23552
rect 400946 -23608 401014 -23552
rect 401070 -23608 401138 -23552
rect 401194 -23608 401262 -23552
rect 401318 -23608 402640 -23552
rect 387840 -23620 402640 -23608
rect 387840 -23676 388981 -23620
rect 389037 -23676 389123 -23620
rect 389179 -23676 389382 -23620
rect 389438 -23676 389524 -23620
rect 389580 -23676 389782 -23620
rect 389838 -23676 389924 -23620
rect 389980 -23676 390179 -23620
rect 390235 -23676 390321 -23620
rect 390377 -23676 390576 -23620
rect 390632 -23676 390718 -23620
rect 390774 -23676 390980 -23620
rect 391036 -23676 391122 -23620
rect 391178 -23676 391376 -23620
rect 391432 -23676 391518 -23620
rect 391574 -23676 391776 -23620
rect 391832 -23676 391918 -23620
rect 391974 -23676 392173 -23620
rect 392229 -23676 392315 -23620
rect 392371 -23676 392578 -23620
rect 392634 -23676 392720 -23620
rect 392776 -23676 392978 -23620
rect 393034 -23676 393120 -23620
rect 393176 -23676 393383 -23620
rect 393439 -23676 393525 -23620
rect 393581 -23676 393780 -23620
rect 393836 -23676 393922 -23620
rect 393978 -23676 394177 -23620
rect 394233 -23676 394319 -23620
rect 394375 -23676 394580 -23620
rect 394636 -23676 394722 -23620
rect 394778 -23676 394982 -23620
rect 395038 -23676 395124 -23620
rect 395180 -23676 395385 -23620
rect 395441 -23676 395527 -23620
rect 395583 -23676 395779 -23620
rect 395835 -23676 395921 -23620
rect 395977 -23676 396180 -23620
rect 396236 -23676 396322 -23620
rect 396378 -23676 396580 -23620
rect 396636 -23676 396722 -23620
rect 396778 -23676 396977 -23620
rect 397033 -23676 397119 -23620
rect 397175 -23676 397374 -23620
rect 397430 -23676 397516 -23620
rect 397572 -23676 397778 -23620
rect 397834 -23676 397920 -23620
rect 397976 -23676 398174 -23620
rect 398230 -23676 398316 -23620
rect 398372 -23676 398574 -23620
rect 398630 -23676 398716 -23620
rect 398772 -23676 398971 -23620
rect 399027 -23676 399113 -23620
rect 399169 -23676 399376 -23620
rect 399432 -23676 399518 -23620
rect 399574 -23676 399776 -23620
rect 399832 -23676 399918 -23620
rect 399974 -23676 400181 -23620
rect 400237 -23676 400323 -23620
rect 400379 -23676 402640 -23620
rect 387840 -23732 387954 -23676
rect 388010 -23732 388078 -23676
rect 388134 -23732 388202 -23676
rect 388258 -23732 388326 -23676
rect 388382 -23732 388450 -23676
rect 388506 -23732 400766 -23676
rect 400822 -23732 400890 -23676
rect 400946 -23732 401014 -23676
rect 401070 -23732 401138 -23676
rect 401194 -23732 401262 -23676
rect 401318 -23732 402640 -23676
rect 387840 -23762 402640 -23732
rect 387840 -23800 388981 -23762
rect 387840 -23856 387954 -23800
rect 388010 -23856 388078 -23800
rect 388134 -23856 388202 -23800
rect 388258 -23856 388326 -23800
rect 388382 -23856 388450 -23800
rect 388506 -23818 388981 -23800
rect 389037 -23818 389123 -23762
rect 389179 -23818 389382 -23762
rect 389438 -23818 389524 -23762
rect 389580 -23818 389782 -23762
rect 389838 -23818 389924 -23762
rect 389980 -23818 390179 -23762
rect 390235 -23818 390321 -23762
rect 390377 -23818 390576 -23762
rect 390632 -23818 390718 -23762
rect 390774 -23818 390980 -23762
rect 391036 -23818 391122 -23762
rect 391178 -23818 391376 -23762
rect 391432 -23818 391518 -23762
rect 391574 -23818 391776 -23762
rect 391832 -23818 391918 -23762
rect 391974 -23818 392173 -23762
rect 392229 -23818 392315 -23762
rect 392371 -23818 392578 -23762
rect 392634 -23818 392720 -23762
rect 392776 -23818 392978 -23762
rect 393034 -23818 393120 -23762
rect 393176 -23818 393383 -23762
rect 393439 -23818 393525 -23762
rect 393581 -23818 393780 -23762
rect 393836 -23818 393922 -23762
rect 393978 -23818 394177 -23762
rect 394233 -23818 394319 -23762
rect 394375 -23818 394580 -23762
rect 394636 -23818 394722 -23762
rect 394778 -23818 394982 -23762
rect 395038 -23818 395124 -23762
rect 395180 -23818 395385 -23762
rect 395441 -23818 395527 -23762
rect 395583 -23818 395779 -23762
rect 395835 -23818 395921 -23762
rect 395977 -23818 396180 -23762
rect 396236 -23818 396322 -23762
rect 396378 -23818 396580 -23762
rect 396636 -23818 396722 -23762
rect 396778 -23818 396977 -23762
rect 397033 -23818 397119 -23762
rect 397175 -23818 397374 -23762
rect 397430 -23818 397516 -23762
rect 397572 -23818 397778 -23762
rect 397834 -23818 397920 -23762
rect 397976 -23818 398174 -23762
rect 398230 -23818 398316 -23762
rect 398372 -23818 398574 -23762
rect 398630 -23818 398716 -23762
rect 398772 -23818 398971 -23762
rect 399027 -23818 399113 -23762
rect 399169 -23818 399376 -23762
rect 399432 -23818 399518 -23762
rect 399574 -23818 399776 -23762
rect 399832 -23818 399918 -23762
rect 399974 -23818 400181 -23762
rect 400237 -23818 400323 -23762
rect 400379 -23800 402640 -23762
rect 400379 -23818 400766 -23800
rect 388506 -23856 400766 -23818
rect 400822 -23856 400890 -23800
rect 400946 -23856 401014 -23800
rect 401070 -23856 401138 -23800
rect 401194 -23856 401262 -23800
rect 401318 -23856 402640 -23800
rect 387840 -23904 402640 -23856
rect 387840 -23924 388981 -23904
rect 387840 -23980 387954 -23924
rect 388010 -23980 388078 -23924
rect 388134 -23980 388202 -23924
rect 388258 -23980 388326 -23924
rect 388382 -23980 388450 -23924
rect 388506 -23960 388981 -23924
rect 389037 -23960 389123 -23904
rect 389179 -23960 389382 -23904
rect 389438 -23960 389524 -23904
rect 389580 -23960 389782 -23904
rect 389838 -23960 389924 -23904
rect 389980 -23960 390179 -23904
rect 390235 -23960 390321 -23904
rect 390377 -23960 390576 -23904
rect 390632 -23960 390718 -23904
rect 390774 -23960 390980 -23904
rect 391036 -23960 391122 -23904
rect 391178 -23960 391376 -23904
rect 391432 -23960 391518 -23904
rect 391574 -23960 391776 -23904
rect 391832 -23960 391918 -23904
rect 391974 -23960 392173 -23904
rect 392229 -23960 392315 -23904
rect 392371 -23960 392578 -23904
rect 392634 -23960 392720 -23904
rect 392776 -23960 392978 -23904
rect 393034 -23960 393120 -23904
rect 393176 -23960 393383 -23904
rect 393439 -23960 393525 -23904
rect 393581 -23960 393780 -23904
rect 393836 -23960 393922 -23904
rect 393978 -23960 394177 -23904
rect 394233 -23960 394319 -23904
rect 394375 -23960 394580 -23904
rect 394636 -23960 394722 -23904
rect 394778 -23960 394982 -23904
rect 395038 -23960 395124 -23904
rect 395180 -23960 395385 -23904
rect 395441 -23960 395527 -23904
rect 395583 -23960 395779 -23904
rect 395835 -23960 395921 -23904
rect 395977 -23960 396180 -23904
rect 396236 -23960 396322 -23904
rect 396378 -23960 396580 -23904
rect 396636 -23960 396722 -23904
rect 396778 -23960 396977 -23904
rect 397033 -23960 397119 -23904
rect 397175 -23960 397374 -23904
rect 397430 -23960 397516 -23904
rect 397572 -23960 397778 -23904
rect 397834 -23960 397920 -23904
rect 397976 -23960 398174 -23904
rect 398230 -23960 398316 -23904
rect 398372 -23960 398574 -23904
rect 398630 -23960 398716 -23904
rect 398772 -23960 398971 -23904
rect 399027 -23960 399113 -23904
rect 399169 -23960 399376 -23904
rect 399432 -23960 399518 -23904
rect 399574 -23960 399776 -23904
rect 399832 -23960 399918 -23904
rect 399974 -23960 400181 -23904
rect 400237 -23960 400323 -23904
rect 400379 -23924 402640 -23904
rect 400379 -23960 400766 -23924
rect 388506 -23980 400766 -23960
rect 400822 -23980 400890 -23924
rect 400946 -23980 401014 -23924
rect 401070 -23980 401138 -23924
rect 401194 -23980 401262 -23924
rect 401318 -23980 402640 -23924
rect 387840 -24046 402640 -23980
rect 387840 -24048 388981 -24046
rect 387840 -24104 387954 -24048
rect 388010 -24104 388078 -24048
rect 388134 -24104 388202 -24048
rect 388258 -24104 388326 -24048
rect 388382 -24104 388450 -24048
rect 388506 -24102 388981 -24048
rect 389037 -24102 389123 -24046
rect 389179 -24102 389382 -24046
rect 389438 -24102 389524 -24046
rect 389580 -24102 389782 -24046
rect 389838 -24102 389924 -24046
rect 389980 -24102 390179 -24046
rect 390235 -24102 390321 -24046
rect 390377 -24102 390576 -24046
rect 390632 -24102 390718 -24046
rect 390774 -24102 390980 -24046
rect 391036 -24102 391122 -24046
rect 391178 -24102 391376 -24046
rect 391432 -24102 391518 -24046
rect 391574 -24102 391776 -24046
rect 391832 -24102 391918 -24046
rect 391974 -24102 392173 -24046
rect 392229 -24102 392315 -24046
rect 392371 -24102 392578 -24046
rect 392634 -24102 392720 -24046
rect 392776 -24102 392978 -24046
rect 393034 -24102 393120 -24046
rect 393176 -24102 393383 -24046
rect 393439 -24102 393525 -24046
rect 393581 -24102 393780 -24046
rect 393836 -24102 393922 -24046
rect 393978 -24102 394177 -24046
rect 394233 -24102 394319 -24046
rect 394375 -24102 394580 -24046
rect 394636 -24102 394722 -24046
rect 394778 -24102 394982 -24046
rect 395038 -24102 395124 -24046
rect 395180 -24102 395385 -24046
rect 395441 -24102 395527 -24046
rect 395583 -24102 395779 -24046
rect 395835 -24102 395921 -24046
rect 395977 -24102 396180 -24046
rect 396236 -24102 396322 -24046
rect 396378 -24102 396580 -24046
rect 396636 -24102 396722 -24046
rect 396778 -24102 396977 -24046
rect 397033 -24102 397119 -24046
rect 397175 -24102 397374 -24046
rect 397430 -24102 397516 -24046
rect 397572 -24102 397778 -24046
rect 397834 -24102 397920 -24046
rect 397976 -24102 398174 -24046
rect 398230 -24102 398316 -24046
rect 398372 -24102 398574 -24046
rect 398630 -24102 398716 -24046
rect 398772 -24102 398971 -24046
rect 399027 -24102 399113 -24046
rect 399169 -24102 399376 -24046
rect 399432 -24102 399518 -24046
rect 399574 -24102 399776 -24046
rect 399832 -24102 399918 -24046
rect 399974 -24102 400181 -24046
rect 400237 -24102 400323 -24046
rect 400379 -24048 402640 -24046
rect 400379 -24102 400766 -24048
rect 388506 -24104 400766 -24102
rect 400822 -24104 400890 -24048
rect 400946 -24104 401014 -24048
rect 401070 -24104 401138 -24048
rect 401194 -24104 401262 -24048
rect 401318 -24104 402640 -24048
rect 387840 -24172 402640 -24104
rect 387840 -24228 387954 -24172
rect 388010 -24228 388078 -24172
rect 388134 -24228 388202 -24172
rect 388258 -24228 388326 -24172
rect 388382 -24228 388450 -24172
rect 388506 -24188 400766 -24172
rect 388506 -24228 388981 -24188
rect 387840 -24244 388981 -24228
rect 389037 -24244 389123 -24188
rect 389179 -24244 389382 -24188
rect 389438 -24244 389524 -24188
rect 389580 -24244 389782 -24188
rect 389838 -24244 389924 -24188
rect 389980 -24244 390179 -24188
rect 390235 -24244 390321 -24188
rect 390377 -24244 390576 -24188
rect 390632 -24244 390718 -24188
rect 390774 -24244 390980 -24188
rect 391036 -24244 391122 -24188
rect 391178 -24244 391376 -24188
rect 391432 -24244 391518 -24188
rect 391574 -24244 391776 -24188
rect 391832 -24244 391918 -24188
rect 391974 -24244 392173 -24188
rect 392229 -24244 392315 -24188
rect 392371 -24244 392578 -24188
rect 392634 -24244 392720 -24188
rect 392776 -24244 392978 -24188
rect 393034 -24244 393120 -24188
rect 393176 -24244 393383 -24188
rect 393439 -24244 393525 -24188
rect 393581 -24244 393780 -24188
rect 393836 -24244 393922 -24188
rect 393978 -24244 394177 -24188
rect 394233 -24244 394319 -24188
rect 394375 -24244 394580 -24188
rect 394636 -24244 394722 -24188
rect 394778 -24244 394982 -24188
rect 395038 -24244 395124 -24188
rect 395180 -24244 395385 -24188
rect 395441 -24244 395527 -24188
rect 395583 -24244 395779 -24188
rect 395835 -24244 395921 -24188
rect 395977 -24244 396180 -24188
rect 396236 -24244 396322 -24188
rect 396378 -24244 396580 -24188
rect 396636 -24244 396722 -24188
rect 396778 -24244 396977 -24188
rect 397033 -24244 397119 -24188
rect 397175 -24244 397374 -24188
rect 397430 -24244 397516 -24188
rect 397572 -24244 397778 -24188
rect 397834 -24244 397920 -24188
rect 397976 -24244 398174 -24188
rect 398230 -24244 398316 -24188
rect 398372 -24244 398574 -24188
rect 398630 -24244 398716 -24188
rect 398772 -24244 398971 -24188
rect 399027 -24244 399113 -24188
rect 399169 -24244 399376 -24188
rect 399432 -24244 399518 -24188
rect 399574 -24244 399776 -24188
rect 399832 -24244 399918 -24188
rect 399974 -24244 400181 -24188
rect 400237 -24244 400323 -24188
rect 400379 -24228 400766 -24188
rect 400822 -24228 400890 -24172
rect 400946 -24228 401014 -24172
rect 401070 -24228 401138 -24172
rect 401194 -24228 401262 -24172
rect 401318 -24228 402640 -24172
rect 400379 -24244 402640 -24228
rect 387840 -24296 402640 -24244
rect 387840 -24352 387954 -24296
rect 388010 -24352 388078 -24296
rect 388134 -24352 388202 -24296
rect 388258 -24352 388326 -24296
rect 388382 -24352 388450 -24296
rect 388506 -24330 400766 -24296
rect 388506 -24352 388981 -24330
rect 387840 -24386 388981 -24352
rect 389037 -24386 389123 -24330
rect 389179 -24386 389382 -24330
rect 389438 -24386 389524 -24330
rect 389580 -24386 389782 -24330
rect 389838 -24386 389924 -24330
rect 389980 -24386 390179 -24330
rect 390235 -24386 390321 -24330
rect 390377 -24386 390576 -24330
rect 390632 -24386 390718 -24330
rect 390774 -24386 390980 -24330
rect 391036 -24386 391122 -24330
rect 391178 -24386 391376 -24330
rect 391432 -24386 391518 -24330
rect 391574 -24386 391776 -24330
rect 391832 -24386 391918 -24330
rect 391974 -24386 392173 -24330
rect 392229 -24386 392315 -24330
rect 392371 -24386 392578 -24330
rect 392634 -24386 392720 -24330
rect 392776 -24386 392978 -24330
rect 393034 -24386 393120 -24330
rect 393176 -24386 393383 -24330
rect 393439 -24386 393525 -24330
rect 393581 -24386 393780 -24330
rect 393836 -24386 393922 -24330
rect 393978 -24386 394177 -24330
rect 394233 -24386 394319 -24330
rect 394375 -24386 394580 -24330
rect 394636 -24386 394722 -24330
rect 394778 -24386 394982 -24330
rect 395038 -24386 395124 -24330
rect 395180 -24386 395385 -24330
rect 395441 -24386 395527 -24330
rect 395583 -24386 395779 -24330
rect 395835 -24386 395921 -24330
rect 395977 -24386 396180 -24330
rect 396236 -24386 396322 -24330
rect 396378 -24386 396580 -24330
rect 396636 -24386 396722 -24330
rect 396778 -24386 396977 -24330
rect 397033 -24386 397119 -24330
rect 397175 -24386 397374 -24330
rect 397430 -24386 397516 -24330
rect 397572 -24386 397778 -24330
rect 397834 -24386 397920 -24330
rect 397976 -24386 398174 -24330
rect 398230 -24386 398316 -24330
rect 398372 -24386 398574 -24330
rect 398630 -24386 398716 -24330
rect 398772 -24386 398971 -24330
rect 399027 -24386 399113 -24330
rect 399169 -24386 399376 -24330
rect 399432 -24386 399518 -24330
rect 399574 -24386 399776 -24330
rect 399832 -24386 399918 -24330
rect 399974 -24386 400181 -24330
rect 400237 -24386 400323 -24330
rect 400379 -24352 400766 -24330
rect 400822 -24352 400890 -24296
rect 400946 -24352 401014 -24296
rect 401070 -24352 401138 -24296
rect 401194 -24352 401262 -24296
rect 401318 -24352 402640 -24296
rect 400379 -24386 402640 -24352
rect 387840 -24420 402640 -24386
rect 387840 -24476 387954 -24420
rect 388010 -24476 388078 -24420
rect 388134 -24476 388202 -24420
rect 388258 -24476 388326 -24420
rect 388382 -24476 388450 -24420
rect 388506 -24472 400766 -24420
rect 388506 -24476 388981 -24472
rect 387840 -24528 388981 -24476
rect 389037 -24528 389123 -24472
rect 389179 -24528 389382 -24472
rect 389438 -24528 389524 -24472
rect 389580 -24528 389782 -24472
rect 389838 -24528 389924 -24472
rect 389980 -24528 390179 -24472
rect 390235 -24528 390321 -24472
rect 390377 -24528 390576 -24472
rect 390632 -24528 390718 -24472
rect 390774 -24528 390980 -24472
rect 391036 -24528 391122 -24472
rect 391178 -24528 391376 -24472
rect 391432 -24528 391518 -24472
rect 391574 -24528 391776 -24472
rect 391832 -24528 391918 -24472
rect 391974 -24528 392173 -24472
rect 392229 -24528 392315 -24472
rect 392371 -24528 392578 -24472
rect 392634 -24528 392720 -24472
rect 392776 -24528 392978 -24472
rect 393034 -24528 393120 -24472
rect 393176 -24528 393383 -24472
rect 393439 -24528 393525 -24472
rect 393581 -24528 393780 -24472
rect 393836 -24528 393922 -24472
rect 393978 -24528 394177 -24472
rect 394233 -24528 394319 -24472
rect 394375 -24528 394580 -24472
rect 394636 -24528 394722 -24472
rect 394778 -24528 394982 -24472
rect 395038 -24528 395124 -24472
rect 395180 -24528 395385 -24472
rect 395441 -24528 395527 -24472
rect 395583 -24528 395779 -24472
rect 395835 -24528 395921 -24472
rect 395977 -24528 396180 -24472
rect 396236 -24528 396322 -24472
rect 396378 -24528 396580 -24472
rect 396636 -24528 396722 -24472
rect 396778 -24528 396977 -24472
rect 397033 -24528 397119 -24472
rect 397175 -24528 397374 -24472
rect 397430 -24528 397516 -24472
rect 397572 -24528 397778 -24472
rect 397834 -24528 397920 -24472
rect 397976 -24528 398174 -24472
rect 398230 -24528 398316 -24472
rect 398372 -24528 398574 -24472
rect 398630 -24528 398716 -24472
rect 398772 -24528 398971 -24472
rect 399027 -24528 399113 -24472
rect 399169 -24528 399376 -24472
rect 399432 -24528 399518 -24472
rect 399574 -24528 399776 -24472
rect 399832 -24528 399918 -24472
rect 399974 -24528 400181 -24472
rect 400237 -24528 400323 -24472
rect 400379 -24476 400766 -24472
rect 400822 -24476 400890 -24420
rect 400946 -24476 401014 -24420
rect 401070 -24476 401138 -24420
rect 401194 -24476 401262 -24420
rect 401318 -24476 402640 -24420
rect 400379 -24528 402640 -24476
rect 387840 -24544 402640 -24528
rect 387840 -24600 387954 -24544
rect 388010 -24600 388078 -24544
rect 388134 -24600 388202 -24544
rect 388258 -24600 388326 -24544
rect 388382 -24600 388450 -24544
rect 388506 -24600 400766 -24544
rect 400822 -24600 400890 -24544
rect 400946 -24600 401014 -24544
rect 401070 -24600 401138 -24544
rect 401194 -24600 401262 -24544
rect 401318 -24600 402640 -24544
rect 387840 -24614 402640 -24600
rect 387840 -24668 388981 -24614
rect 387840 -24724 387954 -24668
rect 388010 -24724 388078 -24668
rect 388134 -24724 388202 -24668
rect 388258 -24724 388326 -24668
rect 388382 -24724 388450 -24668
rect 388506 -24670 388981 -24668
rect 389037 -24670 389123 -24614
rect 389179 -24670 389382 -24614
rect 389438 -24670 389524 -24614
rect 389580 -24670 389782 -24614
rect 389838 -24670 389924 -24614
rect 389980 -24670 390179 -24614
rect 390235 -24670 390321 -24614
rect 390377 -24670 390576 -24614
rect 390632 -24670 390718 -24614
rect 390774 -24670 390980 -24614
rect 391036 -24670 391122 -24614
rect 391178 -24670 391376 -24614
rect 391432 -24670 391518 -24614
rect 391574 -24670 391776 -24614
rect 391832 -24670 391918 -24614
rect 391974 -24670 392173 -24614
rect 392229 -24670 392315 -24614
rect 392371 -24670 392578 -24614
rect 392634 -24670 392720 -24614
rect 392776 -24670 392978 -24614
rect 393034 -24670 393120 -24614
rect 393176 -24670 393383 -24614
rect 393439 -24670 393525 -24614
rect 393581 -24670 393780 -24614
rect 393836 -24670 393922 -24614
rect 393978 -24670 394177 -24614
rect 394233 -24670 394319 -24614
rect 394375 -24670 394580 -24614
rect 394636 -24670 394722 -24614
rect 394778 -24670 394982 -24614
rect 395038 -24670 395124 -24614
rect 395180 -24670 395385 -24614
rect 395441 -24670 395527 -24614
rect 395583 -24670 395779 -24614
rect 395835 -24670 395921 -24614
rect 395977 -24670 396180 -24614
rect 396236 -24670 396322 -24614
rect 396378 -24670 396580 -24614
rect 396636 -24670 396722 -24614
rect 396778 -24670 396977 -24614
rect 397033 -24670 397119 -24614
rect 397175 -24670 397374 -24614
rect 397430 -24670 397516 -24614
rect 397572 -24670 397778 -24614
rect 397834 -24670 397920 -24614
rect 397976 -24670 398174 -24614
rect 398230 -24670 398316 -24614
rect 398372 -24670 398574 -24614
rect 398630 -24670 398716 -24614
rect 398772 -24670 398971 -24614
rect 399027 -24670 399113 -24614
rect 399169 -24670 399376 -24614
rect 399432 -24670 399518 -24614
rect 399574 -24670 399776 -24614
rect 399832 -24670 399918 -24614
rect 399974 -24670 400181 -24614
rect 400237 -24670 400323 -24614
rect 400379 -24668 402640 -24614
rect 400379 -24670 400766 -24668
rect 388506 -24724 400766 -24670
rect 400822 -24724 400890 -24668
rect 400946 -24724 401014 -24668
rect 401070 -24724 401138 -24668
rect 401194 -24724 401262 -24668
rect 401318 -24724 402640 -24668
rect 387840 -24756 402640 -24724
rect 387840 -24792 388981 -24756
rect 387840 -24848 387954 -24792
rect 388010 -24848 388078 -24792
rect 388134 -24848 388202 -24792
rect 388258 -24848 388326 -24792
rect 388382 -24848 388450 -24792
rect 388506 -24812 388981 -24792
rect 389037 -24812 389123 -24756
rect 389179 -24812 389382 -24756
rect 389438 -24812 389524 -24756
rect 389580 -24812 389782 -24756
rect 389838 -24812 389924 -24756
rect 389980 -24812 390179 -24756
rect 390235 -24812 390321 -24756
rect 390377 -24812 390576 -24756
rect 390632 -24812 390718 -24756
rect 390774 -24812 390980 -24756
rect 391036 -24812 391122 -24756
rect 391178 -24812 391376 -24756
rect 391432 -24812 391518 -24756
rect 391574 -24812 391776 -24756
rect 391832 -24812 391918 -24756
rect 391974 -24812 392173 -24756
rect 392229 -24812 392315 -24756
rect 392371 -24812 392578 -24756
rect 392634 -24812 392720 -24756
rect 392776 -24812 392978 -24756
rect 393034 -24812 393120 -24756
rect 393176 -24812 393383 -24756
rect 393439 -24812 393525 -24756
rect 393581 -24812 393780 -24756
rect 393836 -24812 393922 -24756
rect 393978 -24812 394177 -24756
rect 394233 -24812 394319 -24756
rect 394375 -24812 394580 -24756
rect 394636 -24812 394722 -24756
rect 394778 -24812 394982 -24756
rect 395038 -24812 395124 -24756
rect 395180 -24812 395385 -24756
rect 395441 -24812 395527 -24756
rect 395583 -24812 395779 -24756
rect 395835 -24812 395921 -24756
rect 395977 -24812 396180 -24756
rect 396236 -24812 396322 -24756
rect 396378 -24812 396580 -24756
rect 396636 -24812 396722 -24756
rect 396778 -24812 396977 -24756
rect 397033 -24812 397119 -24756
rect 397175 -24812 397374 -24756
rect 397430 -24812 397516 -24756
rect 397572 -24812 397778 -24756
rect 397834 -24812 397920 -24756
rect 397976 -24812 398174 -24756
rect 398230 -24812 398316 -24756
rect 398372 -24812 398574 -24756
rect 398630 -24812 398716 -24756
rect 398772 -24812 398971 -24756
rect 399027 -24812 399113 -24756
rect 399169 -24812 399376 -24756
rect 399432 -24812 399518 -24756
rect 399574 -24812 399776 -24756
rect 399832 -24812 399918 -24756
rect 399974 -24812 400181 -24756
rect 400237 -24812 400323 -24756
rect 400379 -24792 402640 -24756
rect 400379 -24812 400766 -24792
rect 388506 -24848 400766 -24812
rect 400822 -24848 400890 -24792
rect 400946 -24848 401014 -24792
rect 401070 -24848 401138 -24792
rect 401194 -24848 401262 -24792
rect 401318 -24848 402640 -24792
rect 387840 -24898 402640 -24848
rect 387840 -24916 388981 -24898
rect 387840 -24972 387954 -24916
rect 388010 -24972 388078 -24916
rect 388134 -24972 388202 -24916
rect 388258 -24972 388326 -24916
rect 388382 -24972 388450 -24916
rect 388506 -24954 388981 -24916
rect 389037 -24954 389123 -24898
rect 389179 -24954 389382 -24898
rect 389438 -24954 389524 -24898
rect 389580 -24954 389782 -24898
rect 389838 -24954 389924 -24898
rect 389980 -24954 390179 -24898
rect 390235 -24954 390321 -24898
rect 390377 -24954 390576 -24898
rect 390632 -24954 390718 -24898
rect 390774 -24954 390980 -24898
rect 391036 -24954 391122 -24898
rect 391178 -24954 391376 -24898
rect 391432 -24954 391518 -24898
rect 391574 -24954 391776 -24898
rect 391832 -24954 391918 -24898
rect 391974 -24954 392173 -24898
rect 392229 -24954 392315 -24898
rect 392371 -24954 392578 -24898
rect 392634 -24954 392720 -24898
rect 392776 -24954 392978 -24898
rect 393034 -24954 393120 -24898
rect 393176 -24954 393383 -24898
rect 393439 -24954 393525 -24898
rect 393581 -24954 393780 -24898
rect 393836 -24954 393922 -24898
rect 393978 -24954 394177 -24898
rect 394233 -24954 394319 -24898
rect 394375 -24954 394580 -24898
rect 394636 -24954 394722 -24898
rect 394778 -24954 394982 -24898
rect 395038 -24954 395124 -24898
rect 395180 -24954 395385 -24898
rect 395441 -24954 395527 -24898
rect 395583 -24954 395779 -24898
rect 395835 -24954 395921 -24898
rect 395977 -24954 396180 -24898
rect 396236 -24954 396322 -24898
rect 396378 -24954 396580 -24898
rect 396636 -24954 396722 -24898
rect 396778 -24954 396977 -24898
rect 397033 -24954 397119 -24898
rect 397175 -24954 397374 -24898
rect 397430 -24954 397516 -24898
rect 397572 -24954 397778 -24898
rect 397834 -24954 397920 -24898
rect 397976 -24954 398174 -24898
rect 398230 -24954 398316 -24898
rect 398372 -24954 398574 -24898
rect 398630 -24954 398716 -24898
rect 398772 -24954 398971 -24898
rect 399027 -24954 399113 -24898
rect 399169 -24954 399376 -24898
rect 399432 -24954 399518 -24898
rect 399574 -24954 399776 -24898
rect 399832 -24954 399918 -24898
rect 399974 -24954 400181 -24898
rect 400237 -24954 400323 -24898
rect 400379 -24916 402640 -24898
rect 400379 -24954 400766 -24916
rect 388506 -24972 400766 -24954
rect 400822 -24972 400890 -24916
rect 400946 -24972 401014 -24916
rect 401070 -24972 401138 -24916
rect 401194 -24972 401262 -24916
rect 401318 -24972 402640 -24916
rect 387840 -25040 402640 -24972
rect 387840 -25096 387954 -25040
rect 388010 -25096 388078 -25040
rect 388134 -25096 388202 -25040
rect 388258 -25096 388326 -25040
rect 388382 -25096 388450 -25040
rect 388506 -25096 388981 -25040
rect 389037 -25096 389123 -25040
rect 389179 -25096 389382 -25040
rect 389438 -25096 389524 -25040
rect 389580 -25096 389782 -25040
rect 389838 -25096 389924 -25040
rect 389980 -25096 390179 -25040
rect 390235 -25096 390321 -25040
rect 390377 -25096 390576 -25040
rect 390632 -25096 390718 -25040
rect 390774 -25096 390980 -25040
rect 391036 -25096 391122 -25040
rect 391178 -25096 391376 -25040
rect 391432 -25096 391518 -25040
rect 391574 -25096 391776 -25040
rect 391832 -25096 391918 -25040
rect 391974 -25096 392173 -25040
rect 392229 -25096 392315 -25040
rect 392371 -25096 392578 -25040
rect 392634 -25096 392720 -25040
rect 392776 -25096 392978 -25040
rect 393034 -25096 393120 -25040
rect 393176 -25096 393383 -25040
rect 393439 -25096 393525 -25040
rect 393581 -25096 393780 -25040
rect 393836 -25096 393922 -25040
rect 393978 -25096 394177 -25040
rect 394233 -25096 394319 -25040
rect 394375 -25096 394580 -25040
rect 394636 -25096 394722 -25040
rect 394778 -25096 394982 -25040
rect 395038 -25096 395124 -25040
rect 395180 -25096 395385 -25040
rect 395441 -25096 395527 -25040
rect 395583 -25096 395779 -25040
rect 395835 -25096 395921 -25040
rect 395977 -25096 396180 -25040
rect 396236 -25096 396322 -25040
rect 396378 -25096 396580 -25040
rect 396636 -25096 396722 -25040
rect 396778 -25096 396977 -25040
rect 397033 -25096 397119 -25040
rect 397175 -25096 397374 -25040
rect 397430 -25096 397516 -25040
rect 397572 -25096 397778 -25040
rect 397834 -25096 397920 -25040
rect 397976 -25096 398174 -25040
rect 398230 -25096 398316 -25040
rect 398372 -25096 398574 -25040
rect 398630 -25096 398716 -25040
rect 398772 -25096 398971 -25040
rect 399027 -25096 399113 -25040
rect 399169 -25096 399376 -25040
rect 399432 -25096 399518 -25040
rect 399574 -25096 399776 -25040
rect 399832 -25096 399918 -25040
rect 399974 -25096 400181 -25040
rect 400237 -25096 400323 -25040
rect 400379 -25096 400766 -25040
rect 400822 -25096 400890 -25040
rect 400946 -25096 401014 -25040
rect 401070 -25096 401138 -25040
rect 401194 -25096 401262 -25040
rect 401318 -25096 402640 -25040
rect 387840 -25164 402640 -25096
rect 387840 -25220 387954 -25164
rect 388010 -25220 388078 -25164
rect 388134 -25220 388202 -25164
rect 388258 -25220 388326 -25164
rect 388382 -25220 388450 -25164
rect 388506 -25182 400766 -25164
rect 388506 -25220 388981 -25182
rect 387840 -25238 388981 -25220
rect 389037 -25238 389123 -25182
rect 389179 -25238 389382 -25182
rect 389438 -25238 389524 -25182
rect 389580 -25238 389782 -25182
rect 389838 -25238 389924 -25182
rect 389980 -25238 390179 -25182
rect 390235 -25238 390321 -25182
rect 390377 -25238 390576 -25182
rect 390632 -25238 390718 -25182
rect 390774 -25238 390980 -25182
rect 391036 -25238 391122 -25182
rect 391178 -25238 391376 -25182
rect 391432 -25238 391518 -25182
rect 391574 -25238 391776 -25182
rect 391832 -25238 391918 -25182
rect 391974 -25238 392173 -25182
rect 392229 -25238 392315 -25182
rect 392371 -25238 392578 -25182
rect 392634 -25238 392720 -25182
rect 392776 -25238 392978 -25182
rect 393034 -25238 393120 -25182
rect 393176 -25238 393383 -25182
rect 393439 -25238 393525 -25182
rect 393581 -25238 393780 -25182
rect 393836 -25238 393922 -25182
rect 393978 -25238 394177 -25182
rect 394233 -25238 394319 -25182
rect 394375 -25238 394580 -25182
rect 394636 -25238 394722 -25182
rect 394778 -25238 394982 -25182
rect 395038 -25238 395124 -25182
rect 395180 -25238 395385 -25182
rect 395441 -25238 395527 -25182
rect 395583 -25238 395779 -25182
rect 395835 -25238 395921 -25182
rect 395977 -25238 396180 -25182
rect 396236 -25238 396322 -25182
rect 396378 -25238 396580 -25182
rect 396636 -25238 396722 -25182
rect 396778 -25238 396977 -25182
rect 397033 -25238 397119 -25182
rect 397175 -25238 397374 -25182
rect 397430 -25238 397516 -25182
rect 397572 -25238 397778 -25182
rect 397834 -25238 397920 -25182
rect 397976 -25238 398174 -25182
rect 398230 -25238 398316 -25182
rect 398372 -25238 398574 -25182
rect 398630 -25238 398716 -25182
rect 398772 -25238 398971 -25182
rect 399027 -25238 399113 -25182
rect 399169 -25238 399376 -25182
rect 399432 -25238 399518 -25182
rect 399574 -25238 399776 -25182
rect 399832 -25238 399918 -25182
rect 399974 -25238 400181 -25182
rect 400237 -25238 400323 -25182
rect 400379 -25220 400766 -25182
rect 400822 -25220 400890 -25164
rect 400946 -25220 401014 -25164
rect 401070 -25220 401138 -25164
rect 401194 -25220 401262 -25164
rect 401318 -25220 402640 -25164
rect 400379 -25238 402640 -25220
rect 387840 -25288 402640 -25238
rect 387840 -25344 387954 -25288
rect 388010 -25344 388078 -25288
rect 388134 -25344 388202 -25288
rect 388258 -25344 388326 -25288
rect 388382 -25344 388450 -25288
rect 388506 -25324 400766 -25288
rect 388506 -25344 388981 -25324
rect 387840 -25380 388981 -25344
rect 389037 -25380 389123 -25324
rect 389179 -25380 389382 -25324
rect 389438 -25380 389524 -25324
rect 389580 -25380 389782 -25324
rect 389838 -25380 389924 -25324
rect 389980 -25380 390179 -25324
rect 390235 -25380 390321 -25324
rect 390377 -25380 390576 -25324
rect 390632 -25380 390718 -25324
rect 390774 -25380 390980 -25324
rect 391036 -25380 391122 -25324
rect 391178 -25380 391376 -25324
rect 391432 -25380 391518 -25324
rect 391574 -25380 391776 -25324
rect 391832 -25380 391918 -25324
rect 391974 -25380 392173 -25324
rect 392229 -25380 392315 -25324
rect 392371 -25380 392578 -25324
rect 392634 -25380 392720 -25324
rect 392776 -25380 392978 -25324
rect 393034 -25380 393120 -25324
rect 393176 -25380 393383 -25324
rect 393439 -25380 393525 -25324
rect 393581 -25380 393780 -25324
rect 393836 -25380 393922 -25324
rect 393978 -25380 394177 -25324
rect 394233 -25380 394319 -25324
rect 394375 -25380 394580 -25324
rect 394636 -25380 394722 -25324
rect 394778 -25380 394982 -25324
rect 395038 -25380 395124 -25324
rect 395180 -25380 395385 -25324
rect 395441 -25380 395527 -25324
rect 395583 -25380 395779 -25324
rect 395835 -25380 395921 -25324
rect 395977 -25380 396180 -25324
rect 396236 -25380 396322 -25324
rect 396378 -25380 396580 -25324
rect 396636 -25380 396722 -25324
rect 396778 -25380 396977 -25324
rect 397033 -25380 397119 -25324
rect 397175 -25380 397374 -25324
rect 397430 -25380 397516 -25324
rect 397572 -25380 397778 -25324
rect 397834 -25380 397920 -25324
rect 397976 -25380 398174 -25324
rect 398230 -25380 398316 -25324
rect 398372 -25380 398574 -25324
rect 398630 -25380 398716 -25324
rect 398772 -25380 398971 -25324
rect 399027 -25380 399113 -25324
rect 399169 -25380 399376 -25324
rect 399432 -25380 399518 -25324
rect 399574 -25380 399776 -25324
rect 399832 -25380 399918 -25324
rect 399974 -25380 400181 -25324
rect 400237 -25380 400323 -25324
rect 400379 -25344 400766 -25324
rect 400822 -25344 400890 -25288
rect 400946 -25344 401014 -25288
rect 401070 -25344 401138 -25288
rect 401194 -25344 401262 -25288
rect 401318 -25344 402640 -25288
rect 400379 -25380 402640 -25344
rect 387840 -25412 402640 -25380
rect 387840 -25468 387954 -25412
rect 388010 -25468 388078 -25412
rect 388134 -25468 388202 -25412
rect 388258 -25468 388326 -25412
rect 388382 -25468 388450 -25412
rect 388506 -25466 400766 -25412
rect 388506 -25468 388981 -25466
rect 387840 -25522 388981 -25468
rect 389037 -25522 389123 -25466
rect 389179 -25522 389382 -25466
rect 389438 -25522 389524 -25466
rect 389580 -25522 389782 -25466
rect 389838 -25522 389924 -25466
rect 389980 -25522 390179 -25466
rect 390235 -25522 390321 -25466
rect 390377 -25522 390576 -25466
rect 390632 -25522 390718 -25466
rect 390774 -25522 390980 -25466
rect 391036 -25522 391122 -25466
rect 391178 -25522 391376 -25466
rect 391432 -25522 391518 -25466
rect 391574 -25522 391776 -25466
rect 391832 -25522 391918 -25466
rect 391974 -25522 392173 -25466
rect 392229 -25522 392315 -25466
rect 392371 -25522 392578 -25466
rect 392634 -25522 392720 -25466
rect 392776 -25522 392978 -25466
rect 393034 -25522 393120 -25466
rect 393176 -25522 393383 -25466
rect 393439 -25522 393525 -25466
rect 393581 -25522 393780 -25466
rect 393836 -25522 393922 -25466
rect 393978 -25522 394177 -25466
rect 394233 -25522 394319 -25466
rect 394375 -25522 394580 -25466
rect 394636 -25522 394722 -25466
rect 394778 -25522 394982 -25466
rect 395038 -25522 395124 -25466
rect 395180 -25522 395385 -25466
rect 395441 -25522 395527 -25466
rect 395583 -25522 395779 -25466
rect 395835 -25522 395921 -25466
rect 395977 -25522 396180 -25466
rect 396236 -25522 396322 -25466
rect 396378 -25522 396580 -25466
rect 396636 -25522 396722 -25466
rect 396778 -25522 396977 -25466
rect 397033 -25522 397119 -25466
rect 397175 -25522 397374 -25466
rect 397430 -25522 397516 -25466
rect 397572 -25522 397778 -25466
rect 397834 -25522 397920 -25466
rect 397976 -25522 398174 -25466
rect 398230 -25522 398316 -25466
rect 398372 -25522 398574 -25466
rect 398630 -25522 398716 -25466
rect 398772 -25522 398971 -25466
rect 399027 -25522 399113 -25466
rect 399169 -25522 399376 -25466
rect 399432 -25522 399518 -25466
rect 399574 -25522 399776 -25466
rect 399832 -25522 399918 -25466
rect 399974 -25522 400181 -25466
rect 400237 -25522 400323 -25466
rect 400379 -25468 400766 -25466
rect 400822 -25468 400890 -25412
rect 400946 -25468 401014 -25412
rect 401070 -25468 401138 -25412
rect 401194 -25468 401262 -25412
rect 401318 -25468 402640 -25412
rect 400379 -25522 402640 -25468
rect 387840 -25536 402640 -25522
rect 387840 -25592 387954 -25536
rect 388010 -25592 388078 -25536
rect 388134 -25592 388202 -25536
rect 388258 -25592 388326 -25536
rect 388382 -25592 388450 -25536
rect 388506 -25592 400766 -25536
rect 400822 -25592 400890 -25536
rect 400946 -25592 401014 -25536
rect 401070 -25592 401138 -25536
rect 401194 -25592 401262 -25536
rect 401318 -25590 402640 -25536
rect 401318 -25592 401440 -25590
rect 387840 -25660 401440 -25592
rect 387840 -25716 387954 -25660
rect 388010 -25716 388078 -25660
rect 388134 -25716 388202 -25660
rect 388258 -25716 388326 -25660
rect 388382 -25716 388450 -25660
rect 388506 -25688 400766 -25660
rect 388506 -25716 388655 -25688
rect 387840 -25744 388655 -25716
rect 388711 -25744 388797 -25688
rect 388853 -25744 388939 -25688
rect 388995 -25744 389081 -25688
rect 389137 -25744 389223 -25688
rect 389279 -25744 389365 -25688
rect 389421 -25744 389507 -25688
rect 389563 -25744 389649 -25688
rect 389705 -25744 389791 -25688
rect 389847 -25744 389933 -25688
rect 389989 -25744 390075 -25688
rect 390131 -25744 390217 -25688
rect 390273 -25744 390359 -25688
rect 390415 -25744 390501 -25688
rect 390557 -25744 390643 -25688
rect 390699 -25744 390785 -25688
rect 390841 -25744 390927 -25688
rect 390983 -25744 391069 -25688
rect 391125 -25744 391211 -25688
rect 391267 -25744 391353 -25688
rect 391409 -25744 391495 -25688
rect 391551 -25744 391637 -25688
rect 391693 -25744 391779 -25688
rect 391835 -25744 391921 -25688
rect 391977 -25744 392063 -25688
rect 392119 -25744 392205 -25688
rect 392261 -25744 392347 -25688
rect 392403 -25744 392489 -25688
rect 392545 -25744 392631 -25688
rect 392687 -25744 392773 -25688
rect 392829 -25744 392915 -25688
rect 392971 -25744 393057 -25688
rect 393113 -25744 393199 -25688
rect 393255 -25744 393341 -25688
rect 393397 -25744 393483 -25688
rect 393539 -25744 393625 -25688
rect 393681 -25744 393767 -25688
rect 393823 -25744 393909 -25688
rect 393965 -25744 394051 -25688
rect 394107 -25744 394193 -25688
rect 394249 -25744 394335 -25688
rect 394391 -25744 394477 -25688
rect 394533 -25744 394619 -25688
rect 394675 -25744 394761 -25688
rect 394817 -25744 394903 -25688
rect 394959 -25744 395045 -25688
rect 395101 -25744 395187 -25688
rect 395243 -25744 395329 -25688
rect 395385 -25744 395471 -25688
rect 395527 -25744 395613 -25688
rect 395669 -25744 395755 -25688
rect 395811 -25744 395897 -25688
rect 395953 -25744 396039 -25688
rect 396095 -25744 396181 -25688
rect 396237 -25744 396323 -25688
rect 396379 -25744 396465 -25688
rect 396521 -25744 396607 -25688
rect 396663 -25744 396749 -25688
rect 396805 -25744 396891 -25688
rect 396947 -25744 397033 -25688
rect 397089 -25744 397175 -25688
rect 397231 -25744 397317 -25688
rect 397373 -25744 397459 -25688
rect 397515 -25744 397601 -25688
rect 397657 -25744 397743 -25688
rect 397799 -25744 397885 -25688
rect 397941 -25744 398027 -25688
rect 398083 -25744 398169 -25688
rect 398225 -25744 398311 -25688
rect 398367 -25744 398453 -25688
rect 398509 -25744 398595 -25688
rect 398651 -25744 398737 -25688
rect 398793 -25744 398879 -25688
rect 398935 -25744 399021 -25688
rect 399077 -25744 399163 -25688
rect 399219 -25744 399305 -25688
rect 399361 -25744 399447 -25688
rect 399503 -25744 399589 -25688
rect 399645 -25744 399731 -25688
rect 399787 -25744 399873 -25688
rect 399929 -25744 400015 -25688
rect 400071 -25744 400157 -25688
rect 400213 -25744 400299 -25688
rect 400355 -25744 400441 -25688
rect 400497 -25744 400583 -25688
rect 400639 -25716 400766 -25688
rect 400822 -25716 400890 -25660
rect 400946 -25716 401014 -25660
rect 401070 -25716 401138 -25660
rect 401194 -25716 401262 -25660
rect 401318 -25716 401440 -25660
rect 400639 -25744 401440 -25716
rect 387840 -25784 401440 -25744
rect 387840 -25840 387954 -25784
rect 388010 -25840 388078 -25784
rect 388134 -25840 388202 -25784
rect 388258 -25840 388326 -25784
rect 388382 -25840 388450 -25784
rect 388506 -25830 400766 -25784
rect 388506 -25840 388655 -25830
rect 387840 -25886 388655 -25840
rect 388711 -25886 388797 -25830
rect 388853 -25886 388939 -25830
rect 388995 -25886 389081 -25830
rect 389137 -25886 389223 -25830
rect 389279 -25886 389365 -25830
rect 389421 -25886 389507 -25830
rect 389563 -25886 389649 -25830
rect 389705 -25886 389791 -25830
rect 389847 -25886 389933 -25830
rect 389989 -25886 390075 -25830
rect 390131 -25886 390217 -25830
rect 390273 -25886 390359 -25830
rect 390415 -25886 390501 -25830
rect 390557 -25886 390643 -25830
rect 390699 -25886 390785 -25830
rect 390841 -25886 390927 -25830
rect 390983 -25886 391069 -25830
rect 391125 -25886 391211 -25830
rect 391267 -25886 391353 -25830
rect 391409 -25886 391495 -25830
rect 391551 -25886 391637 -25830
rect 391693 -25886 391779 -25830
rect 391835 -25886 391921 -25830
rect 391977 -25886 392063 -25830
rect 392119 -25886 392205 -25830
rect 392261 -25886 392347 -25830
rect 392403 -25886 392489 -25830
rect 392545 -25886 392631 -25830
rect 392687 -25886 392773 -25830
rect 392829 -25886 392915 -25830
rect 392971 -25886 393057 -25830
rect 393113 -25886 393199 -25830
rect 393255 -25886 393341 -25830
rect 393397 -25886 393483 -25830
rect 393539 -25886 393625 -25830
rect 393681 -25886 393767 -25830
rect 393823 -25886 393909 -25830
rect 393965 -25886 394051 -25830
rect 394107 -25886 394193 -25830
rect 394249 -25886 394335 -25830
rect 394391 -25886 394477 -25830
rect 394533 -25886 394619 -25830
rect 394675 -25886 394761 -25830
rect 394817 -25886 394903 -25830
rect 394959 -25886 395045 -25830
rect 395101 -25886 395187 -25830
rect 395243 -25886 395329 -25830
rect 395385 -25886 395471 -25830
rect 395527 -25886 395613 -25830
rect 395669 -25886 395755 -25830
rect 395811 -25886 395897 -25830
rect 395953 -25886 396039 -25830
rect 396095 -25886 396181 -25830
rect 396237 -25886 396323 -25830
rect 396379 -25886 396465 -25830
rect 396521 -25886 396607 -25830
rect 396663 -25886 396749 -25830
rect 396805 -25886 396891 -25830
rect 396947 -25886 397033 -25830
rect 397089 -25886 397175 -25830
rect 397231 -25886 397317 -25830
rect 397373 -25886 397459 -25830
rect 397515 -25886 397601 -25830
rect 397657 -25886 397743 -25830
rect 397799 -25886 397885 -25830
rect 397941 -25886 398027 -25830
rect 398083 -25886 398169 -25830
rect 398225 -25886 398311 -25830
rect 398367 -25886 398453 -25830
rect 398509 -25886 398595 -25830
rect 398651 -25886 398737 -25830
rect 398793 -25886 398879 -25830
rect 398935 -25886 399021 -25830
rect 399077 -25886 399163 -25830
rect 399219 -25886 399305 -25830
rect 399361 -25886 399447 -25830
rect 399503 -25886 399589 -25830
rect 399645 -25886 399731 -25830
rect 399787 -25886 399873 -25830
rect 399929 -25886 400015 -25830
rect 400071 -25886 400157 -25830
rect 400213 -25886 400299 -25830
rect 400355 -25886 400441 -25830
rect 400497 -25886 400583 -25830
rect 400639 -25840 400766 -25830
rect 400822 -25840 400890 -25784
rect 400946 -25840 401014 -25784
rect 401070 -25840 401138 -25784
rect 401194 -25840 401262 -25784
rect 401318 -25840 401440 -25784
rect 400639 -25886 401440 -25840
rect 387840 -25990 401440 -25886
<< glass >>
rect 388640 -25590 400640 -13590
<< labels >>
flabel metal5 390640 -25590 402640 -13590 0 FreeSans 24000 0 0 0 flash_clk
port 2 nsew
flabel metal5 388640 -25590 400640 -13590 0 FreeSans 24000 0 0 0 flash_clk
port 2 nsew
rlabel metal5 s 392140 -21990 397140 -16990 4 PAD
port 7 nsew signal bidirectional
rlabel space 387140 -25590 387140 -25590 4 & Metric 1.00
rlabel space 387140 -25190 387140 -25190 4 & Version 2014q3v1
rlabel space 387140 -24790 387140 -24790 4 & Product GF018green_ipio_5p0c_75
rlabel space 387140 -24390 387140 -24390 4 & Vendor GLOBALFOUNDRIES
rlabel metal5 402140 -25590 402140 -25590 4 & Metric 1.00
rlabel metal5 402140 -25190 402140 -25190 4 & Version 2014q3v1
rlabel metal5 402140 -24790 402140 -24790 4 & Product GF018green_ipio_5p0c_75
rlabel metal5 402140 -24390 402140 -24390 4 & Vendor GLOBALFOUNDRIES
<< properties >>
string FIXED_BBOX 0 0 778000 1020000
<< end >>
